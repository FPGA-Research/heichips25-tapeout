* NGSPICE file created from NE_term.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

.subckt NE_term FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1END[0] N1END[1] N1END[2] N1END[3]
+ N2END[0] N2END[1] N2END[2] N2END[3] N2END[4] N2END[5] N2END[6] N2END[7] N2MID[0]
+ N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5] N2MID[6] N2MID[7] N4END[0] N4END[10]
+ N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2] N4END[3] N4END[4]
+ N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] S1BEG[0] S1BEG[1] S1BEG[2] S1BEG[3]
+ S2BEG[0] S2BEG[1] S2BEG[2] S2BEG[3] S2BEG[4] S2BEG[5] S2BEG[6] S2BEG[7] S2BEGb[0]
+ S2BEGb[1] S2BEGb[2] S2BEGb[3] S2BEGb[4] S2BEGb[5] S2BEGb[6] S2BEGb[7] S4BEG[0] S4BEG[10]
+ S4BEG[11] S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15] S4BEG[1] S4BEG[2] S4BEG[3] S4BEG[4]
+ S4BEG[5] S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9] UserCLK UserCLKo VGND VPWR
X_83_ N4END[4] S4BEG[11] VPWR VGND sg13g2_buf_1
XFILLER_3_67 VPWR VGND sg13g2_decap_8
XFILLER_9_126 VPWR VGND sg13g2_fill_2
XFILLER_8_192 VPWR VGND sg13g2_decap_8
XFILLER_10_147 VPWR VGND sg13g2_fill_1
X_66_ N2END[5] S2BEGb[2] VPWR VGND sg13g2_buf_1
XFILLER_5_151 VPWR VGND sg13g2_decap_8
XFILLER_0_35 VPWR VGND sg13g2_decap_8
XFILLER_9_77 VPWR VGND sg13g2_decap_8
X_49_ FrameStrobe[17] FrameStrobe_O[17] VPWR VGND sg13g2_buf_1
XFILLER_6_67 VPWR VGND sg13g2_decap_8
XFILLER_11_0 VPWR VGND sg13g2_decap_8
XFILLER_3_46 VPWR VGND sg13g2_decap_8
XFILLER_9_105 VPWR VGND sg13g2_decap_8
X_82_ N4END[5] S4BEG[10] VPWR VGND sg13g2_buf_1
XFILLER_8_182 VPWR VGND sg13g2_decap_4
X_65_ N2END[6] S2BEGb[1] VPWR VGND sg13g2_buf_1
XFILLER_5_130 VPWR VGND sg13g2_decap_8
XFILLER_5_185 VPWR VGND sg13g2_decap_8
XFILLER_0_14 VPWR VGND sg13g2_decap_8
XFILLER_9_56 VPWR VGND sg13g2_decap_8
X_48_ FrameStrobe[16] FrameStrobe_O[16] VPWR VGND sg13g2_buf_1
XFILLER_1_90 VPWR VGND sg13g2_fill_1
XFILLER_6_46 VPWR VGND sg13g2_decap_8
XFILLER_9_128 VPWR VGND sg13g2_fill_1
X_81_ N4END[6] S4BEG[9] VPWR VGND sg13g2_buf_1
XFILLER_3_25 VPWR VGND sg13g2_decap_8
XFILLER_8_161 VPWR VGND sg13g2_decap_8
XFILLER_6_109 VPWR VGND sg13g2_decap_8
XFILLER_10_116 VPWR VGND sg13g2_decap_8
XFILLER_10_127 VPWR VGND sg13g2_decap_8
XFILLER_10_138 VPWR VGND sg13g2_decap_8
X_64_ N2END[7] S2BEGb[0] VPWR VGND sg13g2_buf_1
XFILLER_2_134 VPWR VGND sg13g2_decap_8
XFILLER_9_35 VPWR VGND sg13g2_decap_8
X_47_ FrameStrobe[15] FrameStrobe_O[15] VPWR VGND sg13g2_buf_1
XFILLER_1_0 VPWR VGND sg13g2_decap_8
XFILLER_6_25 VPWR VGND sg13g2_decap_8
X_80_ N4END[7] S4BEG[8] VPWR VGND sg13g2_buf_1
XFILLER_8_140 VPWR VGND sg13g2_decap_8
XFILLER_5_165 VPWR VGND sg13g2_fill_2
X_63_ N2MID[0] S2BEG[7] VPWR VGND sg13g2_buf_1
XFILLER_0_49 VPWR VGND sg13g2_decap_8
XFILLER_2_113 VPWR VGND sg13g2_decap_8
XFILLER_2_157 VPWR VGND sg13g2_decap_8
XFILLER_2_179 VPWR VGND sg13g2_decap_8
X_46_ FrameStrobe[14] FrameStrobe_O[14] VPWR VGND sg13g2_buf_1
XFILLER_9_14 VPWR VGND sg13g2_decap_8
X_29_ FrameData[29] FrameData_O[29] VPWR VGND sg13g2_buf_1
XFILLER_9_119 VPWR VGND sg13g2_decap_8
XFILLER_5_144 VPWR VGND sg13g2_decap_8
X_62_ N2MID[1] S2BEG[6] VPWR VGND sg13g2_buf_1
XFILLER_5_199 VPWR VGND sg13g2_fill_1
XFILLER_4_81 VPWR VGND sg13g2_decap_8
XFILLER_0_28 VPWR VGND sg13g2_decap_8
X_45_ FrameStrobe[13] FrameStrobe_O[13] VPWR VGND sg13g2_buf_1
X_28_ FrameData[28] FrameData_O[28] VPWR VGND sg13g2_buf_1
XFILLER_7_81 VPWR VGND sg13g2_decap_8
XFILLER_3_39 VPWR VGND sg13g2_decap_8
XFILLER_8_175 VPWR VGND sg13g2_decap_8
XFILLER_8_186 VPWR VGND sg13g2_fill_2
X_61_ N2MID[2] S2BEG[5] VPWR VGND sg13g2_buf_1
XFILLER_5_123 VPWR VGND sg13g2_decap_8
XFILLER_5_178 VPWR VGND sg13g2_decap_8
XFILLER_4_60 VPWR VGND sg13g2_decap_8
XFILLER_9_49 VPWR VGND sg13g2_decap_8
X_44_ FrameStrobe[12] FrameStrobe_O[12] VPWR VGND sg13g2_buf_1
XFILLER_1_50 VPWR VGND sg13g2_fill_1
X_27_ FrameData[27] FrameData_O[27] VPWR VGND sg13g2_buf_1
XFILLER_6_39 VPWR VGND sg13g2_decap_8
XFILLER_7_60 VPWR VGND sg13g2_decap_8
XFILLER_3_18 VPWR VGND sg13g2_decap_8
XFILLER_8_154 VPWR VGND sg13g2_decap_8
X_60_ N2MID[3] S2BEG[4] VPWR VGND sg13g2_buf_1
XFILLER_5_102 VPWR VGND sg13g2_decap_8
XFILLER_2_127 VPWR VGND sg13g2_decap_8
XFILLER_9_28 VPWR VGND sg13g2_decap_8
X_43_ FrameStrobe[11] FrameStrobe_O[11] VPWR VGND sg13g2_buf_1
X_26_ FrameData[26] FrameData_O[26] VPWR VGND sg13g2_buf_1
XFILLER_1_40 VPWR VGND sg13g2_fill_1
XFILLER_6_18 VPWR VGND sg13g2_decap_8
XFILLER_10_60 VPWR VGND sg13g2_decap_8
X_09_ FrameData[9] FrameData_O[9] VPWR VGND sg13g2_buf_1
XFILLER_8_133 VPWR VGND sg13g2_decap_8
XFILLER_8_199 VPWR VGND sg13g2_fill_1
XFILLER_5_158 VPWR VGND sg13g2_fill_2
XFILLER_4_95 VPWR VGND sg13g2_decap_8
XFILLER_2_106 VPWR VGND sg13g2_decap_8
XFILLER_1_183 VPWR VGND sg13g2_fill_2
XFILLER_1_150 VPWR VGND sg13g2_fill_2
X_42_ FrameStrobe[10] FrameStrobe_O[10] VPWR VGND sg13g2_buf_1
X_25_ FrameData[25] FrameData_O[25] VPWR VGND sg13g2_buf_1
XFILLER_10_83 VPWR VGND sg13g2_fill_2
X_08_ FrameData[8] FrameData_O[8] VPWR VGND sg13g2_buf_1
XFILLER_11_7 VPWR VGND sg13g2_decap_8
XFILLER_7_95 VPWR VGND sg13g2_decap_8
XFILLER_8_112 VPWR VGND sg13g2_decap_8
XFILLER_5_137 VPWR VGND sg13g2_decap_8
XFILLER_4_74 VPWR VGND sg13g2_decap_8
X_41_ FrameStrobe[9] FrameStrobe_O[9] VPWR VGND sg13g2_buf_1
XFILLER_1_86 VPWR VGND sg13g2_decap_4
X_24_ FrameData[24] FrameData_O[24] VPWR VGND sg13g2_buf_1
XFILLER_10_51 VPWR VGND sg13g2_decap_4
XFILLER_10_73 VPWR VGND sg13g2_decap_4
X_07_ FrameData[7] FrameData_O[7] VPWR VGND sg13g2_buf_1
XFILLER_7_74 VPWR VGND sg13g2_decap_8
XFILLER_8_168 VPWR VGND sg13g2_decap_8
XFILLER_5_116 VPWR VGND sg13g2_decap_8
XFILLER_4_53 VPWR VGND sg13g2_decap_8
XFILLER_1_152 VPWR VGND sg13g2_fill_1
XFILLER_8_0 VPWR VGND sg13g2_decap_8
X_40_ FrameStrobe[8] FrameStrobe_O[8] VPWR VGND sg13g2_buf_1
X_23_ FrameData[23] FrameData_O[23] VPWR VGND sg13g2_buf_1
XFILLER_10_41 VPWR VGND sg13g2_decap_4
X_06_ FrameData[6] FrameData_O[6] VPWR VGND sg13g2_buf_1
XFILLER_7_53 VPWR VGND sg13g2_decap_8
XFILLER_8_147 VPWR VGND sg13g2_decap_8
XFILLER_4_32 VPWR VGND sg13g2_decap_8
XFILLER_4_172 VPWR VGND sg13g2_decap_8
XFILLER_1_120 VPWR VGND sg13g2_fill_1
XFILLER_1_197 VPWR VGND sg13g2_fill_2
XFILLER_1_99 VPWR VGND sg13g2_fill_1
XFILLER_1_55 VPWR VGND sg13g2_decap_4
X_22_ FrameData[22] FrameData_O[22] VPWR VGND sg13g2_buf_1
XFILLER_10_31 VPWR VGND sg13g2_decap_4
X_05_ FrameData[5] FrameData_O[5] VPWR VGND sg13g2_buf_1
XFILLER_7_32 VPWR VGND sg13g2_decap_8
XFILLER_8_126 VPWR VGND sg13g2_decap_8
XFILLER_4_11 VPWR VGND sg13g2_decap_8
XFILLER_4_88 VPWR VGND sg13g2_decap_8
XFILLER_4_151 VPWR VGND sg13g2_decap_8
XFILLER_4_195 VPWR VGND sg13g2_decap_4
XFILLER_1_176 VPWR VGND sg13g2_decap_8
XFILLER_1_143 VPWR VGND sg13g2_decap_8
X_21_ FrameData[21] FrameData_O[21] VPWR VGND sg13g2_buf_1
XFILLER_1_45 VPWR VGND sg13g2_fill_1
X_04_ FrameData[4] FrameData_O[4] VPWR VGND sg13g2_buf_1
XFILLER_7_88 VPWR VGND sg13g2_decap_8
XFILLER_8_105 VPWR VGND sg13g2_decap_8
XFILLER_4_67 VPWR VGND sg13g2_decap_8
XFILLER_4_130 VPWR VGND sg13g2_decap_8
XFILLER_1_199 VPWR VGND sg13g2_fill_1
XFILLER_6_0 VPWR VGND sg13g2_decap_8
XFILLER_1_79 VPWR VGND sg13g2_decap_8
X_20_ FrameData[20] FrameData_O[20] VPWR VGND sg13g2_buf_1
XFILLER_10_22 VPWR VGND sg13g2_fill_1
XFILLER_10_55 VPWR VGND sg13g2_fill_1
XFILLER_10_77 VPWR VGND sg13g2_fill_2
X_03_ FrameData[3] FrameData_O[3] VPWR VGND sg13g2_buf_1
XFILLER_7_67 VPWR VGND sg13g2_decap_8
XFILLER_7_172 VPWR VGND sg13g2_fill_2
XFILLER_5_109 VPWR VGND sg13g2_decap_8
XFILLER_4_46 VPWR VGND sg13g2_decap_8
X_79_ N4END[8] S4BEG[7] VPWR VGND sg13g2_buf_1
XFILLER_10_45 VPWR VGND sg13g2_fill_2
XFILLER_10_67 VPWR VGND sg13g2_fill_2
XFILLER_10_89 VPWR VGND sg13g2_decap_8
X_02_ FrameData[2] FrameData_O[2] VPWR VGND sg13g2_buf_1
XFILLER_7_46 VPWR VGND sg13g2_decap_8
XFILLER_7_151 VPWR VGND sg13g2_decap_8
XFILLER_4_25 VPWR VGND sg13g2_decap_8
XFILLER_4_165 VPWR VGND sg13g2_decap_8
XFILLER_1_157 VPWR VGND sg13g2_decap_8
X_78_ N4END[9] S4BEG[6] VPWR VGND sg13g2_buf_1
XFILLER_10_35 VPWR VGND sg13g2_fill_2
X_01_ FrameData[1] FrameData_O[1] VPWR VGND sg13g2_buf_1
XFILLER_7_25 VPWR VGND sg13g2_decap_8
XFILLER_8_119 VPWR VGND sg13g2_decap_8
XFILLER_7_130 VPWR VGND sg13g2_decap_8
XFILLER_7_185 VPWR VGND sg13g2_fill_2
XFILLER_7_196 VPWR VGND sg13g2_decap_4
XFILLER_4_144 VPWR VGND sg13g2_decap_8
XFILLER_4_199 VPWR VGND sg13g2_fill_1
XFILLER_1_38 VPWR VGND sg13g2_fill_2
X_77_ N4END[10] S4BEG[5] VPWR VGND sg13g2_buf_1
X_00_ FrameData[0] FrameData_O[0] VPWR VGND sg13g2_buf_1
XFILLER_4_0 VPWR VGND sg13g2_decap_8
XFILLER_2_92 VPWR VGND sg13g2_decap_8
XFILLER_11_182 VPWR VGND sg13g2_decap_8
XFILLER_8_91 VPWR VGND sg13g2_decap_8
XFILLER_4_123 VPWR VGND sg13g2_decap_8
XFILLER_1_137 VPWR VGND sg13g2_fill_2
XFILLER_8_7 VPWR VGND sg13g2_decap_8
XFILLER_5_81 VPWR VGND sg13g2_decap_8
X_76_ N4END[11] S4BEG[4] VPWR VGND sg13g2_buf_1
XFILLER_10_15 VPWR VGND sg13g2_decap_8
X_59_ N2MID[4] S2BEG[3] VPWR VGND sg13g2_buf_1
XFILLER_2_82 VPWR VGND sg13g2_decap_4
XFILLER_11_91 VPWR VGND sg13g2_decap_8
XFILLER_11_161 VPWR VGND sg13g2_decap_8
XFILLER_7_165 VPWR VGND sg13g2_decap_8
XFILLER_7_187 VPWR VGND sg13g2_fill_1
XFILLER_8_70 VPWR VGND sg13g2_decap_8
XFILLER_4_39 VPWR VGND sg13g2_decap_8
XFILLER_4_102 VPWR VGND sg13g2_decap_8
XFILLER_4_179 VPWR VGND sg13g2_decap_4
XFILLER_1_116 VPWR VGND sg13g2_decap_4
XFILLER_0_193 VPWR VGND sg13g2_decap_8
XFILLER_5_60 VPWR VGND sg13g2_decap_8
X_75_ N4END[12] S4BEG[3] VPWR VGND sg13g2_buf_1
XFILLER_2_61 VPWR VGND sg13g2_decap_8
X_58_ N2MID[5] S2BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_11_70 VPWR VGND sg13g2_decap_8
XFILLER_7_39 VPWR VGND sg13g2_decap_8
XFILLER_11_140 VPWR VGND sg13g2_decap_8
XFILLER_7_144 VPWR VGND sg13g2_decap_8
XFILLER_4_18 VPWR VGND sg13g2_decap_8
XFILLER_4_158 VPWR VGND sg13g2_decap_8
XFILLER_0_172 VPWR VGND sg13g2_decap_8
XFILLER_0_161 VPWR VGND sg13g2_decap_8
XFILLER_1_19 VPWR VGND sg13g2_decap_8
X_74_ N4END[13] S4BEG[2] VPWR VGND sg13g2_buf_1
X_57_ N2MID[6] S2BEG[1] VPWR VGND sg13g2_buf_1
XFILLER_2_0 VPWR VGND sg13g2_decap_8
XFILLER_7_18 VPWR VGND sg13g2_decap_8
XFILLER_11_196 VPWR VGND sg13g2_decap_4
XFILLER_7_123 VPWR VGND sg13g2_decap_8
XFILLER_7_178 VPWR VGND sg13g2_decap_8
XFILLER_4_137 VPWR VGND sg13g2_decap_8
XFILLER_3_192 VPWR VGND sg13g2_decap_8
XFILLER_0_140 VPWR VGND sg13g2_decap_8
XFILLER_5_95 VPWR VGND sg13g2_decap_8
X_73_ N4END[14] S4BEG[1] VPWR VGND sg13g2_buf_1
X_56_ N2MID[7] S2BEG[0] VPWR VGND sg13g2_buf_1
X_39_ FrameStrobe[7] FrameStrobe_O[7] VPWR VGND sg13g2_buf_1
XFILLER_11_175 VPWR VGND sg13g2_decap_8
XFILLER_7_102 VPWR VGND sg13g2_decap_8
XFILLER_8_84 VPWR VGND sg13g2_decap_8
XFILLER_4_116 VPWR VGND sg13g2_decap_8
XFILLER_5_74 VPWR VGND sg13g2_decap_8
XFILLER_10_0 VPWR VGND sg13g2_fill_2
X_72_ N4END[15] S4BEG[0] VPWR VGND sg13g2_buf_1
XFILLER_2_42 VPWR VGND sg13g2_decap_8
XFILLER_2_20 VPWR VGND sg13g2_decap_4
X_55_ N1END[0] S1BEG[3] VPWR VGND sg13g2_buf_1
XFILLER_2_75 VPWR VGND sg13g2_fill_2
XFILLER_2_86 VPWR VGND sg13g2_fill_2
XFILLER_11_84 VPWR VGND sg13g2_decap_8
X_38_ FrameStrobe[6] FrameStrobe_O[6] VPWR VGND sg13g2_buf_1
XFILLER_11_154 VPWR VGND sg13g2_decap_8
XFILLER_7_158 VPWR VGND sg13g2_decap_8
XFILLER_6_191 VPWR VGND sg13g2_decap_8
XFILLER_8_63 VPWR VGND sg13g2_decap_8
XFILLER_3_172 VPWR VGND sg13g2_decap_8
XFILLER_0_186 VPWR VGND sg13g2_decap_8
XFILLER_5_53 VPWR VGND sg13g2_decap_8
X_71_ N2END[0] S2BEGb[7] VPWR VGND sg13g2_buf_1
X_54_ N1END[1] S1BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_11_63 VPWR VGND sg13g2_decap_8
X_37_ FrameStrobe[5] FrameStrobe_O[5] VPWR VGND sg13g2_buf_1
XFILLER_11_133 VPWR VGND sg13g2_decap_8
XFILLER_0_0 VPWR VGND sg13g2_decap_8
XFILLER_7_137 VPWR VGND sg13g2_decap_8
XFILLER_8_42 VPWR VGND sg13g2_decap_8
XFILLER_3_151 VPWR VGND sg13g2_decap_8
XFILLER_0_154 VPWR VGND sg13g2_decap_8
XFILLER_5_32 VPWR VGND sg13g2_decap_8
XFILLER_10_2 VPWR VGND sg13g2_fill_1
X_70_ N2END[1] S2BEGb[6] VPWR VGND sg13g2_buf_1
XFILLER_2_11 VPWR VGND sg13g2_decap_4
X_53_ N1END[2] S1BEG[1] VPWR VGND sg13g2_buf_1
XFILLER_2_77 VPWR VGND sg13g2_fill_1
XFILLER_2_99 VPWR VGND sg13g2_decap_8
XFILLER_11_42 VPWR VGND sg13g2_decap_8
X_36_ FrameStrobe[4] FrameStrobe_O[4] VPWR VGND sg13g2_buf_1
XFILLER_11_189 VPWR VGND sg13g2_decap_8
XFILLER_11_112 VPWR VGND sg13g2_decap_8
XFILLER_7_116 VPWR VGND sg13g2_decap_8
XFILLER_8_21 VPWR VGND sg13g2_decap_8
XFILLER_8_98 VPWR VGND sg13g2_decap_8
X_19_ FrameData[19] FrameData_O[19] VPWR VGND sg13g2_buf_1
XFILLER_3_130 VPWR VGND sg13g2_decap_8
XFILLER_0_133 VPWR VGND sg13g2_decap_8
XFILLER_5_11 VPWR VGND sg13g2_decap_8
XFILLER_5_88 VPWR VGND sg13g2_decap_8
XFILLER_2_56 VPWR VGND sg13g2_fill_1
X_52_ N1END[3] S1BEG[0] VPWR VGND sg13g2_buf_1
XFILLER_11_98 VPWR VGND sg13g2_decap_8
XFILLER_11_21 VPWR VGND sg13g2_decap_8
X_35_ FrameStrobe[3] FrameStrobe_O[3] VPWR VGND sg13g2_buf_1
XFILLER_11_168 VPWR VGND sg13g2_decap_8
XFILLER_6_172 VPWR VGND sg13g2_decap_8
XFILLER_8_77 VPWR VGND sg13g2_decap_8
XFILLER_4_109 VPWR VGND sg13g2_decap_8
X_18_ FrameData[18] FrameData_O[18] VPWR VGND sg13g2_buf_1
XFILLER_3_186 VPWR VGND sg13g2_fill_2
XFILLER_0_112 VPWR VGND sg13g2_decap_8
XFILLER_5_67 VPWR VGND sg13g2_decap_8
X_51_ FrameStrobe[19] FrameStrobe_O[19] VPWR VGND sg13g2_buf_1
XFILLER_2_35 VPWR VGND sg13g2_decap_8
XFILLER_2_68 VPWR VGND sg13g2_decap_8
XFILLER_11_77 VPWR VGND sg13g2_decap_8
X_34_ FrameStrobe[2] FrameStrobe_O[2] VPWR VGND sg13g2_buf_1
XFILLER_11_147 VPWR VGND sg13g2_decap_8
XFILLER_8_56 VPWR VGND sg13g2_decap_8
XFILLER_6_151 VPWR VGND sg13g2_decap_8
X_17_ FrameData[17] FrameData_O[17] VPWR VGND sg13g2_buf_1
XFILLER_3_165 VPWR VGND sg13g2_decap_8
XFILLER_0_179 VPWR VGND sg13g2_decap_8
XFILLER_5_46 VPWR VGND sg13g2_decap_8
X_50_ FrameStrobe[18] FrameStrobe_O[18] VPWR VGND sg13g2_buf_1
XFILLER_9_0 VPWR VGND sg13g2_decap_8
XFILLER_11_56 VPWR VGND sg13g2_decap_8
X_33_ FrameStrobe[1] FrameStrobe_O[1] VPWR VGND sg13g2_buf_1
XFILLER_9_182 VPWR VGND sg13g2_decap_8
XFILLER_11_126 VPWR VGND sg13g2_decap_8
XFILLER_10_181 VPWR VGND sg13g2_decap_4
XFILLER_6_130 VPWR VGND sg13g2_decap_8
X_16_ FrameData[16] FrameData_O[16] VPWR VGND sg13g2_buf_1
XFILLER_8_35 VPWR VGND sg13g2_decap_8
XFILLER_3_144 VPWR VGND sg13g2_decap_8
XFILLER_3_199 VPWR VGND sg13g2_fill_1
XFILLER_0_91 VPWR VGND sg13g2_decap_8
XFILLER_0_147 VPWR VGND sg13g2_decap_8
XFILLER_5_25 VPWR VGND sg13g2_decap_8
XFILLER_2_15 VPWR VGND sg13g2_fill_1
XFILLER_11_35 VPWR VGND sg13g2_decap_8
XFILLER_9_161 VPWR VGND sg13g2_decap_8
X_32_ FrameStrobe[0] FrameStrobe_O[0] VPWR VGND sg13g2_buf_1
XFILLER_11_105 VPWR VGND sg13g2_decap_8
XFILLER_7_109 VPWR VGND sg13g2_decap_8
X_15_ FrameData[15] FrameData_O[15] VPWR VGND sg13g2_buf_1
XFILLER_6_186 VPWR VGND sg13g2_fill_1
XFILLER_8_14 VPWR VGND sg13g2_decap_8
XFILLER_3_123 VPWR VGND sg13g2_decap_8
XFILLER_0_70 VPWR VGND sg13g2_decap_8
XFILLER_0_126 VPWR VGND sg13g2_decap_8
XFILLER_2_49 VPWR VGND sg13g2_decap_8
XFILLER_11_14 VPWR VGND sg13g2_decap_8
X_31_ FrameData[31] FrameData_O[31] VPWR VGND sg13g2_buf_1
XFILLER_9_140 VPWR VGND sg13g2_decap_8
XFILLER_3_81 VPWR VGND sg13g2_decap_8
XFILLER_6_165 VPWR VGND sg13g2_decap_8
XFILLER_6_198 VPWR VGND sg13g2_fill_2
X_14_ FrameData[14] FrameData_O[14] VPWR VGND sg13g2_buf_1
XFILLER_3_102 VPWR VGND sg13g2_decap_8
XFILLER_3_179 VPWR VGND sg13g2_decap_8
XFILLER_0_105 VPWR VGND sg13g2_decap_8
XFILLER_9_91 VPWR VGND sg13g2_decap_8
XFILLER_6_81 VPWR VGND sg13g2_decap_8
XFILLER_2_28 VPWR VGND sg13g2_decap_8
XFILLER_7_0 VPWR VGND sg13g2_decap_4
X_30_ FrameData[30] FrameData_O[30] VPWR VGND sg13g2_buf_1
XFILLER_9_196 VPWR VGND sg13g2_decap_4
XFILLER_3_60 VPWR VGND sg13g2_decap_8
XFILLER_0_7 VPWR VGND sg13g2_decap_8
XFILLER_6_144 VPWR VGND sg13g2_decap_8
XFILLER_8_49 VPWR VGND sg13g2_decap_8
X_13_ FrameData[13] FrameData_O[13] VPWR VGND sg13g2_buf_1
XFILLER_3_158 VPWR VGND sg13g2_decap_8
XFILLER_9_70 VPWR VGND sg13g2_decap_8
XFILLER_5_39 VPWR VGND sg13g2_decap_8
XFILLER_6_60 VPWR VGND sg13g2_decap_8
XFILLER_11_49 VPWR VGND sg13g2_decap_8
XFILLER_11_119 VPWR VGND sg13g2_decap_8
XFILLER_9_175 VPWR VGND sg13g2_decap_8
XFILLER_8_28 VPWR VGND sg13g2_decap_8
XFILLER_10_152 VPWR VGND sg13g2_fill_2
X_12_ FrameData[12] FrameData_O[12] VPWR VGND sg13g2_buf_1
XFILLER_6_123 VPWR VGND sg13g2_decap_8
XFILLER_3_137 VPWR VGND sg13g2_decap_8
XFILLER_0_84 VPWR VGND sg13g2_decap_8
XFILLER_5_18 VPWR VGND sg13g2_decap_8
XFILLER_11_28 VPWR VGND sg13g2_decap_8
XFILLER_3_95 VPWR VGND sg13g2_decap_8
X_88_ UserCLK UserCLKo VPWR VGND sg13g2_buf_1
XFILLER_9_154 VPWR VGND sg13g2_decap_8
XFILLER_10_197 VPWR VGND sg13g2_fill_2
XFILLER_10_175 VPWR VGND sg13g2_fill_2
X_11_ FrameData[11] FrameData_O[11] VPWR VGND sg13g2_buf_1
XFILLER_6_102 VPWR VGND sg13g2_decap_8
XFILLER_6_179 VPWR VGND sg13g2_decap_8
XFILLER_3_116 VPWR VGND sg13g2_decap_8
XFILLER_0_63 VPWR VGND sg13g2_decap_8
XFILLER_2_193 VPWR VGND sg13g2_decap_8
XFILLER_0_119 VPWR VGND sg13g2_decap_8
XFILLER_6_95 VPWR VGND sg13g2_decap_8
XFILLER_3_74 VPWR VGND sg13g2_decap_8
XFILLER_9_133 VPWR VGND sg13g2_decap_8
X_87_ N4END[0] S4BEG[15] VPWR VGND sg13g2_buf_1
XFILLER_5_0 VPWR VGND sg13g2_decap_8
X_10_ FrameData[10] FrameData_O[10] VPWR VGND sg13g2_buf_1
XFILLER_6_158 VPWR VGND sg13g2_decap_8
XFILLER_10_154 VPWR VGND sg13g2_fill_1
XFILLER_0_42 VPWR VGND sg13g2_decap_8
XFILLER_2_172 VPWR VGND sg13g2_decap_8
XFILLER_9_84 VPWR VGND sg13g2_decap_8
XFILLER_6_74 VPWR VGND sg13g2_decap_8
XFILLER_9_7 VPWR VGND sg13g2_fill_2
XFILLER_9_189 VPWR VGND sg13g2_decap_8
XFILLER_7_4 VPWR VGND sg13g2_fill_2
XFILLER_9_112 VPWR VGND sg13g2_decap_8
X_86_ N4END[1] S4BEG[14] VPWR VGND sg13g2_buf_1
XFILLER_3_53 VPWR VGND sg13g2_decap_8
XFILLER_10_199 VPWR VGND sg13g2_fill_1
XFILLER_6_137 VPWR VGND sg13g2_decap_8
XFILLER_10_100 VPWR VGND sg13g2_decap_4
XFILLER_5_192 VPWR VGND sg13g2_decap_8
X_69_ N2END[2] S2BEGb[5] VPWR VGND sg13g2_buf_1
XFILLER_0_98 VPWR VGND sg13g2_decap_8
XFILLER_0_21 VPWR VGND sg13g2_decap_8
XFILLER_2_151 VPWR VGND sg13g2_fill_2
XFILLER_9_63 VPWR VGND sg13g2_decap_8
XFILLER_6_53 VPWR VGND sg13g2_decap_8
XFILLER_9_168 VPWR VGND sg13g2_decap_8
X_85_ N4END[2] S4BEG[13] VPWR VGND sg13g2_buf_1
XFILLER_3_32 VPWR VGND sg13g2_decap_8
XFILLER_10_167 VPWR VGND sg13g2_decap_4
XFILLER_6_116 VPWR VGND sg13g2_decap_8
XFILLER_10_145 VPWR VGND sg13g2_fill_2
XFILLER_5_160 VPWR VGND sg13g2_fill_1
XFILLER_5_171 VPWR VGND sg13g2_decap_8
X_68_ N2END[3] S2BEGb[4] VPWR VGND sg13g2_buf_1
XFILLER_2_141 VPWR VGND sg13g2_fill_2
XFILLER_0_77 VPWR VGND sg13g2_decap_8
XFILLER_9_42 VPWR VGND sg13g2_decap_8
XFILLER_6_32 VPWR VGND sg13g2_decap_8
XFILLER_9_9 VPWR VGND sg13g2_fill_1
X_84_ N4END[3] S4BEG[12] VPWR VGND sg13g2_buf_1
XFILLER_3_11 VPWR VGND sg13g2_decap_8
XFILLER_3_88 VPWR VGND sg13g2_decap_8
XFILLER_9_147 VPWR VGND sg13g2_decap_8
X_67_ N2END[4] S2BEGb[3] VPWR VGND sg13g2_buf_1
XFILLER_3_109 VPWR VGND sg13g2_decap_8
XFILLER_2_120 VPWR VGND sg13g2_decap_8
XFILLER_2_164 VPWR VGND sg13g2_decap_4
XFILLER_2_186 VPWR VGND sg13g2_decap_8
XFILLER_3_0 VPWR VGND sg13g2_decap_8
XFILLER_0_56 VPWR VGND sg13g2_decap_8
XFILLER_9_21 VPWR VGND sg13g2_decap_8
XFILLER_9_98 VPWR VGND sg13g2_decap_8
XFILLER_6_11 VPWR VGND sg13g2_decap_8
XFILLER_6_88 VPWR VGND sg13g2_decap_8
.ends

