magic
tech ihp-sg13g2
magscale 1 2
timestamp 1753389534
<< metal1 >>
rect 576 38576 89376 38600
rect 576 38536 4352 38576
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4720 38536 19472 38576
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19840 38536 34592 38576
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34960 38536 49712 38576
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 50080 38536 64832 38576
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 65200 38536 79952 38576
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 80320 38536 89376 38576
rect 576 38512 89376 38536
rect 576 37820 89376 37844
rect 576 37780 3112 37820
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3480 37780 18232 37820
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18600 37780 33352 37820
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33720 37780 48472 37820
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48840 37780 63592 37820
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63960 37780 78712 37820
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 79080 37780 89376 37820
rect 576 37756 89376 37780
rect 576 37064 89376 37088
rect 576 37024 4352 37064
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4720 37024 19472 37064
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19840 37024 34592 37064
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34960 37024 49712 37064
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 50080 37024 64832 37064
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 65200 37024 79952 37064
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 80320 37024 89376 37064
rect 576 37000 89376 37024
rect 576 36308 89376 36332
rect 576 36268 3112 36308
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3480 36268 18232 36308
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18600 36268 33352 36308
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33720 36268 48472 36308
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48840 36268 63592 36308
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63960 36268 78712 36308
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 79080 36268 89376 36308
rect 576 36244 89376 36268
rect 576 35552 89376 35576
rect 576 35512 4352 35552
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4720 35512 19472 35552
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19840 35512 34592 35552
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34960 35512 49712 35552
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 50080 35512 64832 35552
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 65200 35512 79952 35552
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 80320 35512 89376 35552
rect 576 35488 89376 35512
rect 643 35132 701 35133
rect 643 35092 652 35132
rect 692 35092 701 35132
rect 643 35091 701 35092
rect 843 34964 885 34973
rect 843 34924 844 34964
rect 884 34924 885 34964
rect 843 34915 885 34924
rect 576 34796 89376 34820
rect 576 34756 3112 34796
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3480 34756 18232 34796
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18600 34756 33352 34796
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33720 34756 48472 34796
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48840 34756 63592 34796
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63960 34756 78712 34796
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 79080 34756 89376 34796
rect 576 34732 89376 34756
rect 643 34460 701 34461
rect 643 34420 652 34460
rect 692 34420 701 34460
rect 643 34419 701 34420
rect 843 34208 885 34217
rect 843 34168 844 34208
rect 884 34168 885 34208
rect 843 34159 885 34168
rect 576 34040 89376 34064
rect 576 34000 4352 34040
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4720 34000 19472 34040
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19840 34000 34592 34040
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34960 34000 49712 34040
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 50080 34000 64832 34040
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 65200 34000 79952 34040
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 80320 34000 89376 34040
rect 576 33976 89376 34000
rect 643 33620 701 33621
rect 643 33580 652 33620
rect 692 33580 701 33620
rect 643 33579 701 33580
rect 843 33452 885 33461
rect 843 33412 844 33452
rect 884 33412 885 33452
rect 843 33403 885 33412
rect 576 33284 89376 33308
rect 576 33244 3112 33284
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3480 33244 18232 33284
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18600 33244 33352 33284
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33720 33244 48472 33284
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48840 33244 63592 33284
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63960 33244 78712 33284
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 79080 33244 89376 33284
rect 576 33220 89376 33244
rect 643 32948 701 32949
rect 643 32908 652 32948
rect 692 32908 701 32948
rect 643 32907 701 32908
rect 4291 32864 4349 32865
rect 4291 32824 4300 32864
rect 4340 32824 4349 32864
rect 4291 32823 4349 32824
rect 4387 32864 4445 32865
rect 4387 32824 4396 32864
rect 4436 32824 4445 32864
rect 4387 32823 4445 32824
rect 843 32696 885 32705
rect 843 32656 844 32696
rect 884 32656 885 32696
rect 843 32647 885 32656
rect 4587 32696 4629 32705
rect 4587 32656 4588 32696
rect 4628 32656 4629 32696
rect 4587 32647 4629 32656
rect 576 32528 89376 32552
rect 576 32488 4352 32528
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4720 32488 19472 32528
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19840 32488 34592 32528
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34960 32488 49712 32528
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 50080 32488 64832 32528
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 65200 32488 79952 32528
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 80320 32488 89376 32528
rect 576 32464 89376 32488
rect 4387 32192 4445 32193
rect 4387 32152 4396 32192
rect 4436 32152 4445 32192
rect 4387 32151 4445 32152
rect 4491 32192 4533 32201
rect 4491 32152 4492 32192
rect 4532 32152 4533 32192
rect 4491 32143 4533 32152
rect 643 32108 701 32109
rect 643 32068 652 32108
rect 692 32068 701 32108
rect 643 32067 701 32068
rect 843 31940 885 31949
rect 843 31900 844 31940
rect 884 31900 885 31940
rect 843 31891 885 31900
rect 4203 31940 4245 31949
rect 4203 31900 4204 31940
rect 4244 31900 4245 31940
rect 4203 31891 4245 31900
rect 576 31772 89376 31796
rect 576 31732 3112 31772
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3480 31732 18232 31772
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18600 31732 33352 31772
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33720 31732 48472 31772
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48840 31732 63592 31772
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63960 31732 78712 31772
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 79080 31732 89376 31772
rect 576 31708 89376 31732
rect 643 31436 701 31437
rect 643 31396 652 31436
rect 692 31396 701 31436
rect 643 31395 701 31396
rect 843 31184 885 31193
rect 843 31144 844 31184
rect 884 31144 885 31184
rect 843 31135 885 31144
rect 576 31016 89376 31040
rect 576 30976 4352 31016
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4720 30976 19472 31016
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19840 30976 34592 31016
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34960 30976 49712 31016
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 50080 30976 64832 31016
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 65200 30976 79952 31016
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 80320 30976 89376 31016
rect 576 30952 89376 30976
rect 3811 30848 3869 30849
rect 3811 30808 3820 30848
rect 3860 30808 3869 30848
rect 3811 30807 3869 30808
rect 2667 30680 2709 30689
rect 2667 30640 2668 30680
rect 2708 30640 2709 30680
rect 2667 30631 2709 30640
rect 2859 30680 2901 30689
rect 2859 30640 2860 30680
rect 2900 30640 2901 30680
rect 2859 30631 2901 30640
rect 3051 30680 3093 30689
rect 3051 30640 3052 30680
rect 3092 30640 3093 30680
rect 3051 30631 3093 30640
rect 3235 30680 3293 30681
rect 3235 30640 3244 30680
rect 3284 30640 3293 30680
rect 3235 30639 3293 30640
rect 3531 30680 3573 30689
rect 3531 30640 3532 30680
rect 3572 30640 3573 30680
rect 3531 30631 3573 30640
rect 3627 30680 3669 30689
rect 3627 30640 3628 30680
rect 3668 30640 3669 30680
rect 3627 30631 3669 30640
rect 3723 30680 3765 30689
rect 3723 30640 3724 30680
rect 3764 30640 3765 30680
rect 3723 30631 3765 30640
rect 643 30596 701 30597
rect 643 30556 652 30596
rect 692 30556 701 30596
rect 643 30555 701 30556
rect 3147 30512 3189 30521
rect 3147 30472 3148 30512
rect 3188 30472 3189 30512
rect 3147 30463 3189 30472
rect 843 30428 885 30437
rect 843 30388 844 30428
rect 884 30388 885 30428
rect 843 30379 885 30388
rect 2859 30428 2901 30437
rect 2859 30388 2860 30428
rect 2900 30388 2901 30428
rect 2859 30379 2901 30388
rect 576 30260 89376 30284
rect 576 30220 3112 30260
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3480 30220 18232 30260
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18600 30220 33352 30260
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33720 30220 48472 30260
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48840 30220 63592 30260
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63960 30220 78712 30260
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 79080 30220 89376 30260
rect 576 30196 89376 30220
rect 643 29924 701 29925
rect 643 29884 652 29924
rect 692 29884 701 29924
rect 643 29883 701 29884
rect 2275 29840 2333 29841
rect 2275 29800 2284 29840
rect 2324 29800 2333 29840
rect 2275 29799 2333 29800
rect 2563 29840 2621 29841
rect 2563 29800 2572 29840
rect 2612 29800 2621 29840
rect 2563 29799 2621 29800
rect 3235 29840 3293 29841
rect 3235 29800 3244 29840
rect 3284 29800 3293 29840
rect 3235 29799 3293 29800
rect 3331 29840 3389 29841
rect 3331 29800 3340 29840
rect 3380 29800 3389 29840
rect 3331 29799 3389 29800
rect 2755 29756 2813 29757
rect 2755 29716 2764 29756
rect 2804 29716 2813 29756
rect 2755 29715 2813 29716
rect 843 29672 885 29681
rect 843 29632 844 29672
rect 884 29632 885 29672
rect 843 29623 885 29632
rect 3051 29672 3093 29681
rect 3051 29632 3052 29672
rect 3092 29632 3093 29672
rect 3051 29623 3093 29632
rect 576 29504 89376 29528
rect 576 29464 4352 29504
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4720 29464 19472 29504
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19840 29464 34592 29504
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34960 29464 49712 29504
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 50080 29464 64832 29504
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 65200 29464 79952 29504
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 80320 29464 89376 29504
rect 576 29440 89376 29464
rect 576 28748 89376 28772
rect 576 28708 3112 28748
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3480 28708 18232 28748
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18600 28708 33352 28748
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33720 28708 48472 28748
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48840 28708 63592 28748
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63960 28708 78712 28748
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 79080 28708 89376 28748
rect 576 28684 89376 28708
rect 843 28580 885 28589
rect 843 28540 844 28580
rect 884 28540 885 28580
rect 843 28531 885 28540
rect 643 28412 701 28413
rect 643 28372 652 28412
rect 692 28372 701 28412
rect 643 28371 701 28372
rect 576 27992 89376 28016
rect 576 27952 4352 27992
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4720 27952 19472 27992
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19840 27952 34592 27992
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34960 27952 49712 27992
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 50080 27952 64832 27992
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 65200 27952 79952 27992
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 80320 27952 89376 27992
rect 576 27928 89376 27952
rect 843 27824 885 27833
rect 843 27784 844 27824
rect 884 27784 885 27824
rect 843 27775 885 27784
rect 11395 27824 11453 27825
rect 11395 27784 11404 27824
rect 11444 27784 11453 27824
rect 11395 27783 11453 27784
rect 11299 27656 11357 27657
rect 11299 27616 11308 27656
rect 11348 27616 11357 27656
rect 11299 27615 11357 27616
rect 643 27572 701 27573
rect 643 27532 652 27572
rect 692 27532 701 27572
rect 643 27531 701 27532
rect 11107 27404 11165 27405
rect 11107 27364 11116 27404
rect 11156 27364 11165 27404
rect 11107 27363 11165 27364
rect 576 27236 89376 27260
rect 576 27196 3112 27236
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3480 27196 18232 27236
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18600 27196 33352 27236
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33720 27196 48472 27236
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48840 27196 63592 27236
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63960 27196 78712 27236
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 79080 27196 89376 27236
rect 576 27172 89376 27196
rect 3819 27068 3861 27077
rect 3819 27028 3820 27068
rect 3860 27028 3861 27068
rect 3819 27019 3861 27028
rect 843 26984 885 26993
rect 843 26944 844 26984
rect 884 26944 885 26984
rect 843 26935 885 26944
rect 10827 26984 10869 26993
rect 10827 26944 10828 26984
rect 10868 26944 10869 26984
rect 10827 26935 10869 26944
rect 643 26900 701 26901
rect 643 26860 652 26900
rect 692 26860 701 26900
rect 643 26859 701 26860
rect 3435 26816 3477 26825
rect 3435 26776 3436 26816
rect 3476 26776 3477 26816
rect 3435 26767 3477 26776
rect 3627 26816 3669 26825
rect 3627 26776 3628 26816
rect 3668 26776 3669 26816
rect 3627 26767 3669 26776
rect 3811 26816 3869 26817
rect 3811 26776 3820 26816
rect 3860 26776 3869 26816
rect 3811 26775 3869 26776
rect 3907 26816 3965 26817
rect 3907 26776 3916 26816
rect 3956 26776 3965 26816
rect 3907 26775 3965 26776
rect 4107 26816 4149 26825
rect 4107 26776 4108 26816
rect 4148 26776 4149 26816
rect 4107 26767 4149 26776
rect 4203 26816 4245 26825
rect 4203 26776 4204 26816
rect 4244 26776 4245 26816
rect 4203 26767 4245 26776
rect 4296 26816 4354 26817
rect 4296 26776 4305 26816
rect 4345 26776 4354 26816
rect 4296 26775 4354 26776
rect 4779 26816 4821 26825
rect 4779 26776 4780 26816
rect 4820 26776 4821 26816
rect 4779 26767 4821 26776
rect 4867 26816 4925 26817
rect 4867 26776 4876 26816
rect 4916 26776 4925 26816
rect 4867 26775 4925 26776
rect 10827 26816 10869 26825
rect 10827 26776 10828 26816
rect 10868 26776 10869 26816
rect 10827 26767 10869 26776
rect 11203 26816 11261 26817
rect 11203 26776 11212 26816
rect 11252 26776 11261 26816
rect 11203 26775 11261 26776
rect 11491 26816 11549 26817
rect 11491 26776 11500 26816
rect 11540 26776 11549 26816
rect 11491 26775 11549 26776
rect 3531 26648 3573 26657
rect 3531 26608 3532 26648
rect 3572 26608 3573 26648
rect 3531 26599 3573 26608
rect 5163 26648 5205 26657
rect 5163 26608 5164 26648
rect 5204 26608 5205 26648
rect 5163 26599 5205 26608
rect 11019 26648 11061 26657
rect 11019 26608 11020 26648
rect 11060 26608 11061 26648
rect 11019 26599 11061 26608
rect 11691 26648 11733 26657
rect 11691 26608 11692 26648
rect 11732 26608 11733 26648
rect 11691 26599 11733 26608
rect 576 26480 89376 26504
rect 576 26440 4352 26480
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4720 26440 19472 26480
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19840 26440 34592 26480
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34960 26440 49712 26480
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 50080 26440 64832 26480
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 65200 26440 79952 26480
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 80320 26440 89376 26480
rect 576 26416 89376 26440
rect 5259 26312 5301 26321
rect 5259 26272 5260 26312
rect 5300 26272 5301 26312
rect 5259 26263 5301 26272
rect 3435 26144 3477 26153
rect 3435 26104 3436 26144
rect 3476 26104 3477 26144
rect 3435 26095 3477 26104
rect 3627 26144 3669 26153
rect 3627 26104 3628 26144
rect 3668 26104 3669 26144
rect 3627 26095 3669 26104
rect 5163 26144 5205 26153
rect 5163 26104 5164 26144
rect 5204 26104 5205 26144
rect 5163 26095 5205 26104
rect 5355 26144 5397 26153
rect 5355 26104 5356 26144
rect 5396 26104 5397 26144
rect 5355 26095 5397 26104
rect 11115 26144 11157 26153
rect 11115 26104 11116 26144
rect 11156 26104 11157 26144
rect 11115 26095 11157 26104
rect 11307 26144 11349 26153
rect 11307 26104 11308 26144
rect 11348 26104 11349 26144
rect 11307 26095 11349 26104
rect 11395 26144 11453 26145
rect 11395 26104 11404 26144
rect 11444 26104 11453 26144
rect 11395 26103 11453 26104
rect 643 26060 701 26061
rect 643 26020 652 26060
rect 692 26020 701 26060
rect 643 26019 701 26020
rect 3627 25976 3669 25985
rect 3627 25936 3628 25976
rect 3668 25936 3669 25976
rect 3627 25927 3669 25936
rect 843 25892 885 25901
rect 843 25852 844 25892
rect 884 25852 885 25892
rect 843 25843 885 25852
rect 11115 25892 11157 25901
rect 11115 25852 11116 25892
rect 11156 25852 11157 25892
rect 11115 25843 11157 25852
rect 576 25724 89376 25748
rect 576 25684 3112 25724
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3480 25684 18232 25724
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18600 25684 33352 25724
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33720 25684 48472 25724
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48840 25684 63592 25724
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63960 25684 78712 25724
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 79080 25684 89376 25724
rect 576 25660 89376 25684
rect 843 25556 885 25565
rect 843 25516 844 25556
rect 884 25516 885 25556
rect 843 25507 885 25516
rect 643 25388 701 25389
rect 643 25348 652 25388
rect 692 25348 701 25388
rect 643 25347 701 25348
rect 12355 25388 12413 25389
rect 12355 25348 12364 25388
rect 12404 25348 12413 25388
rect 12355 25347 12413 25348
rect 12547 25304 12605 25305
rect 12547 25264 12556 25304
rect 12596 25264 12605 25304
rect 12547 25263 12605 25264
rect 12643 25304 12701 25305
rect 12643 25264 12652 25304
rect 12692 25264 12701 25304
rect 12643 25263 12701 25264
rect 576 24968 89376 24992
rect 576 24928 4352 24968
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4720 24928 19472 24968
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19840 24928 34592 24968
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34960 24928 49712 24968
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 50080 24928 64832 24968
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 65200 24928 79952 24968
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 80320 24928 89376 24968
rect 576 24904 89376 24928
rect 10819 24800 10877 24801
rect 10819 24760 10828 24800
rect 10868 24760 10877 24800
rect 10819 24759 10877 24760
rect 12075 24800 12117 24809
rect 12075 24760 12076 24800
rect 12116 24760 12117 24800
rect 12075 24751 12117 24760
rect 4779 24716 4821 24725
rect 4779 24676 4780 24716
rect 4820 24676 4821 24716
rect 4779 24667 4821 24676
rect 9771 24716 9813 24725
rect 9771 24676 9772 24716
rect 9812 24676 9813 24716
rect 9771 24667 9813 24676
rect 4107 24632 4149 24641
rect 4107 24592 4108 24632
rect 4148 24592 4149 24632
rect 4107 24583 4149 24592
rect 4203 24632 4245 24641
rect 4203 24592 4204 24632
rect 4244 24592 4245 24632
rect 4203 24583 4245 24592
rect 4291 24632 4349 24633
rect 4291 24592 4300 24632
rect 4340 24592 4349 24632
rect 4291 24591 4349 24592
rect 4675 24632 4733 24633
rect 4675 24592 4684 24632
rect 4724 24592 4733 24632
rect 4675 24591 4733 24592
rect 5443 24632 5501 24633
rect 5443 24592 5452 24632
rect 5492 24592 5501 24632
rect 5443 24591 5501 24592
rect 5539 24632 5597 24633
rect 5539 24592 5548 24632
rect 5588 24592 5597 24632
rect 5539 24591 5597 24592
rect 6499 24632 6557 24633
rect 6499 24592 6508 24632
rect 6548 24592 6557 24632
rect 6499 24591 6557 24592
rect 6595 24632 6653 24633
rect 6595 24592 6604 24632
rect 6644 24592 6653 24632
rect 6595 24591 6653 24592
rect 9867 24632 9909 24641
rect 9867 24592 9868 24632
rect 9908 24592 9909 24632
rect 9867 24583 9909 24592
rect 9963 24632 10005 24641
rect 9963 24592 9964 24632
rect 10004 24592 10005 24632
rect 9963 24583 10005 24592
rect 10059 24632 10101 24641
rect 10059 24592 10060 24632
rect 10100 24592 10101 24632
rect 10059 24583 10101 24592
rect 11019 24632 11061 24641
rect 11019 24592 11020 24632
rect 11060 24592 11061 24632
rect 11019 24583 11061 24592
rect 11115 24632 11157 24641
rect 11115 24592 11116 24632
rect 11156 24592 11157 24632
rect 11115 24583 11157 24592
rect 11979 24632 12021 24641
rect 11979 24592 11980 24632
rect 12020 24592 12021 24632
rect 11979 24583 12021 24592
rect 12171 24632 12213 24641
rect 12171 24592 12172 24632
rect 12212 24592 12213 24632
rect 12171 24583 12213 24592
rect 643 24548 701 24549
rect 643 24508 652 24548
rect 692 24508 701 24548
rect 643 24507 701 24508
rect 843 24380 885 24389
rect 843 24340 844 24380
rect 884 24340 885 24380
rect 843 24331 885 24340
rect 5355 24380 5397 24389
rect 5355 24340 5356 24380
rect 5396 24340 5397 24380
rect 5355 24331 5397 24340
rect 6411 24380 6453 24389
rect 6411 24340 6412 24380
rect 6452 24340 6453 24380
rect 6411 24331 6453 24340
rect 576 24212 89376 24236
rect 576 24172 3112 24212
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3480 24172 18232 24212
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18600 24172 33352 24212
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33720 24172 48472 24212
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48840 24172 63592 24212
rect 63632 24172 63674 24212
rect 63714 24172 63756 24212
rect 63796 24172 63838 24212
rect 63878 24172 63920 24212
rect 63960 24172 78712 24212
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 79080 24172 89376 24212
rect 576 24148 89376 24172
rect 1899 24044 1941 24053
rect 1899 24004 1900 24044
rect 1940 24004 1941 24044
rect 1899 23995 1941 24004
rect 4203 24044 4245 24053
rect 4203 24004 4204 24044
rect 4244 24004 4245 24044
rect 4203 23995 4245 24004
rect 11403 24044 11445 24053
rect 11403 24004 11404 24044
rect 11444 24004 11445 24044
rect 11403 23995 11445 24004
rect 643 23876 701 23877
rect 643 23836 652 23876
rect 692 23836 701 23876
rect 643 23835 701 23836
rect 1803 23792 1845 23801
rect 1803 23752 1804 23792
rect 1844 23752 1845 23792
rect 1803 23743 1845 23752
rect 1987 23792 2045 23793
rect 1987 23752 1996 23792
rect 2036 23752 2045 23792
rect 1987 23751 2045 23752
rect 2179 23792 2237 23793
rect 2179 23752 2188 23792
rect 2228 23752 2237 23792
rect 2179 23751 2237 23752
rect 2467 23792 2525 23793
rect 2467 23752 2476 23792
rect 2516 23752 2525 23792
rect 2467 23751 2525 23752
rect 4099 23792 4157 23793
rect 4099 23752 4108 23792
rect 4148 23752 4157 23792
rect 4099 23751 4157 23752
rect 4299 23792 4341 23801
rect 4299 23752 4300 23792
rect 4340 23752 4341 23792
rect 4299 23743 4341 23752
rect 11211 23792 11253 23801
rect 11211 23752 11212 23792
rect 11252 23752 11253 23792
rect 11211 23743 11253 23752
rect 11403 23792 11445 23801
rect 11403 23752 11404 23792
rect 11444 23752 11445 23792
rect 11403 23743 11445 23752
rect 2659 23708 2717 23709
rect 2659 23668 2668 23708
rect 2708 23668 2717 23708
rect 2659 23667 2717 23668
rect 843 23624 885 23633
rect 843 23584 844 23624
rect 884 23584 885 23624
rect 843 23575 885 23584
rect 576 23456 89376 23480
rect 576 23416 4352 23456
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4720 23416 19472 23456
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19840 23416 34592 23456
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34960 23416 49712 23456
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 50080 23416 64832 23456
rect 64872 23416 64914 23456
rect 64954 23416 64996 23456
rect 65036 23416 65078 23456
rect 65118 23416 65160 23456
rect 65200 23416 79952 23456
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 80320 23416 89376 23456
rect 576 23392 89376 23416
rect 12067 23288 12125 23289
rect 12067 23248 12076 23288
rect 12116 23248 12125 23288
rect 12067 23247 12125 23248
rect 12355 23288 12413 23289
rect 12355 23248 12364 23288
rect 12404 23248 12413 23288
rect 12355 23247 12413 23248
rect 12259 23120 12317 23121
rect 12259 23080 12268 23120
rect 12308 23080 12317 23120
rect 12259 23079 12317 23080
rect 643 23036 701 23037
rect 643 22996 652 23036
rect 692 22996 701 23036
rect 643 22995 701 22996
rect 843 22868 885 22877
rect 843 22828 844 22868
rect 884 22828 885 22868
rect 843 22819 885 22828
rect 576 22700 89376 22724
rect 576 22660 3112 22700
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3480 22660 18232 22700
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18600 22660 33352 22700
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33720 22660 48472 22700
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48840 22660 63592 22700
rect 63632 22660 63674 22700
rect 63714 22660 63756 22700
rect 63796 22660 63838 22700
rect 63878 22660 63920 22700
rect 63960 22660 78712 22700
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 79080 22660 89376 22700
rect 576 22636 89376 22660
rect 11875 22364 11933 22365
rect 11875 22324 11884 22364
rect 11924 22324 11933 22364
rect 11875 22323 11933 22324
rect 11299 22280 11357 22281
rect 11299 22240 11308 22280
rect 11348 22240 11357 22280
rect 11299 22239 11357 22240
rect 11587 22280 11645 22281
rect 11587 22240 11596 22280
rect 11636 22240 11645 22280
rect 11587 22239 11645 22240
rect 12067 22280 12125 22281
rect 12067 22240 12076 22280
rect 12116 22240 12125 22280
rect 12067 22239 12125 22240
rect 12163 22280 12221 22281
rect 12163 22240 12172 22280
rect 12212 22240 12221 22280
rect 12163 22239 12221 22240
rect 643 22112 701 22113
rect 643 22072 652 22112
rect 692 22072 701 22112
rect 643 22071 701 22072
rect 11115 22112 11157 22121
rect 11115 22072 11116 22112
rect 11156 22072 11157 22112
rect 11115 22063 11157 22072
rect 576 21944 89376 21968
rect 576 21904 4352 21944
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4720 21904 19472 21944
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19840 21904 34592 21944
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34960 21904 49712 21944
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 50080 21904 64832 21944
rect 64872 21904 64914 21944
rect 64954 21904 64996 21944
rect 65036 21904 65078 21944
rect 65118 21904 65160 21944
rect 65200 21904 79952 21944
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 80320 21904 89376 21944
rect 576 21880 89376 21904
rect 576 21188 89376 21212
rect 576 21148 3112 21188
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3480 21148 18232 21188
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18600 21148 33352 21188
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33720 21148 48472 21188
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48840 21148 63592 21188
rect 63632 21148 63674 21188
rect 63714 21148 63756 21188
rect 63796 21148 63838 21188
rect 63878 21148 63920 21188
rect 63960 21148 78712 21188
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 79080 21148 89376 21188
rect 576 21124 89376 21148
rect 8811 20936 8853 20945
rect 8811 20896 8812 20936
rect 8852 20896 8853 20936
rect 8811 20887 8853 20896
rect 3427 20768 3485 20769
rect 3427 20728 3436 20768
rect 3476 20728 3485 20768
rect 3427 20727 3485 20728
rect 3811 20768 3869 20769
rect 3811 20728 3820 20768
rect 3860 20728 3869 20768
rect 3811 20727 3869 20728
rect 4099 20768 4157 20769
rect 4099 20728 4108 20768
rect 4148 20728 4157 20768
rect 4099 20727 4157 20728
rect 8323 20768 8381 20769
rect 8323 20728 8332 20768
rect 8372 20728 8381 20768
rect 8323 20727 8381 20728
rect 8515 20768 8573 20769
rect 8515 20728 8524 20768
rect 8564 20728 8573 20768
rect 8515 20727 8573 20728
rect 8907 20768 8949 20777
rect 8907 20728 8908 20768
rect 8948 20728 8949 20768
rect 8907 20719 8949 20728
rect 4291 20684 4349 20685
rect 4291 20644 4300 20684
rect 4340 20644 4349 20684
rect 4291 20643 4349 20644
rect 643 20600 701 20601
rect 643 20560 652 20600
rect 692 20560 701 20600
rect 643 20559 701 20560
rect 3339 20600 3381 20609
rect 3339 20560 3340 20600
rect 3380 20560 3381 20600
rect 3339 20551 3381 20560
rect 4003 20600 4061 20601
rect 4003 20560 4012 20600
rect 4052 20560 4061 20600
rect 4003 20559 4061 20560
rect 576 20432 89376 20456
rect 576 20392 4352 20432
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4720 20392 19472 20432
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19840 20392 34592 20432
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34960 20392 49712 20432
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 50080 20392 64832 20432
rect 64872 20392 64914 20432
rect 64954 20392 64996 20432
rect 65036 20392 65078 20432
rect 65118 20392 65160 20432
rect 65200 20392 79952 20432
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 80320 20392 89376 20432
rect 576 20368 89376 20392
rect 643 20264 701 20265
rect 643 20224 652 20264
rect 692 20224 701 20264
rect 643 20223 701 20224
rect 8619 20264 8661 20273
rect 8619 20224 8620 20264
rect 8660 20224 8661 20264
rect 8619 20215 8661 20224
rect 7843 20180 7901 20181
rect 7843 20140 7852 20180
rect 7892 20140 7901 20180
rect 7843 20139 7901 20140
rect 8035 20096 8093 20097
rect 8035 20056 8044 20096
rect 8084 20056 8093 20096
rect 8035 20055 8093 20056
rect 8323 20096 8381 20097
rect 8323 20056 8332 20096
rect 8372 20056 8381 20096
rect 8323 20055 8381 20056
rect 8707 20096 8765 20097
rect 8707 20056 8716 20096
rect 8756 20056 8765 20096
rect 8707 20055 8765 20056
rect 9091 20096 9149 20097
rect 9091 20056 9100 20096
rect 9140 20056 9149 20096
rect 9091 20055 9149 20056
rect 576 19676 89376 19700
rect 576 19636 3112 19676
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3480 19636 18232 19676
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18600 19636 33352 19676
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33720 19636 48472 19676
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48840 19636 63592 19676
rect 63632 19636 63674 19676
rect 63714 19636 63756 19676
rect 63796 19636 63838 19676
rect 63878 19636 63920 19676
rect 63960 19636 78712 19676
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 79080 19636 89376 19676
rect 576 19612 89376 19636
rect 8323 19508 8381 19509
rect 8323 19468 8332 19508
rect 8372 19468 8381 19508
rect 8323 19467 8381 19468
rect 8131 19256 8189 19257
rect 8131 19216 8140 19256
rect 8180 19216 8189 19256
rect 8131 19215 8189 19216
rect 643 19088 701 19089
rect 643 19048 652 19088
rect 692 19048 701 19088
rect 643 19047 701 19048
rect 8035 19088 8093 19089
rect 8035 19048 8044 19088
rect 8084 19048 8093 19088
rect 8035 19047 8093 19048
rect 576 18920 89376 18944
rect 576 18880 4352 18920
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4720 18880 19472 18920
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19840 18880 34592 18920
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34960 18880 49712 18920
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 50080 18880 64832 18920
rect 64872 18880 64914 18920
rect 64954 18880 64996 18920
rect 65036 18880 65078 18920
rect 65118 18880 65160 18920
rect 65200 18880 79952 18920
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 80320 18880 89376 18920
rect 576 18856 89376 18880
rect 643 18752 701 18753
rect 643 18712 652 18752
rect 692 18712 701 18752
rect 643 18711 701 18712
rect 576 18164 89376 18188
rect 576 18124 3112 18164
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3480 18124 18232 18164
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18600 18124 33352 18164
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33720 18124 48472 18164
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48840 18124 63592 18164
rect 63632 18124 63674 18164
rect 63714 18124 63756 18164
rect 63796 18124 63838 18164
rect 63878 18124 63920 18164
rect 63960 18124 78712 18164
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 79080 18124 89376 18164
rect 576 18100 89376 18124
rect 643 17576 701 17577
rect 643 17536 652 17576
rect 692 17536 701 17576
rect 643 17535 701 17536
rect 576 17408 89376 17432
rect 576 17368 4352 17408
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4720 17368 19472 17408
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19840 17368 34592 17408
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34960 17368 49712 17408
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 50080 17368 64832 17408
rect 64872 17368 64914 17408
rect 64954 17368 64996 17408
rect 65036 17368 65078 17408
rect 65118 17368 65160 17408
rect 65200 17368 79952 17408
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 80320 17368 89376 17408
rect 576 17344 89376 17368
rect 643 17240 701 17241
rect 643 17200 652 17240
rect 692 17200 701 17240
rect 643 17199 701 17200
rect 576 16652 89376 16676
rect 576 16612 3112 16652
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3480 16612 18232 16652
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18600 16612 33352 16652
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33720 16612 48472 16652
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48840 16612 63592 16652
rect 63632 16612 63674 16652
rect 63714 16612 63756 16652
rect 63796 16612 63838 16652
rect 63878 16612 63920 16652
rect 63960 16612 78712 16652
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 79080 16612 89376 16652
rect 576 16588 89376 16612
rect 643 16064 701 16065
rect 643 16024 652 16064
rect 692 16024 701 16064
rect 643 16023 701 16024
rect 576 15896 89376 15920
rect 576 15856 4352 15896
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4720 15856 19472 15896
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19840 15856 34592 15896
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34960 15856 49712 15896
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 50080 15856 64832 15896
rect 64872 15856 64914 15896
rect 64954 15856 64996 15896
rect 65036 15856 65078 15896
rect 65118 15856 65160 15896
rect 65200 15856 79952 15896
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 80320 15856 89376 15896
rect 576 15832 89376 15856
rect 643 15728 701 15729
rect 643 15688 652 15728
rect 692 15688 701 15728
rect 643 15687 701 15688
rect 576 15140 89376 15164
rect 576 15100 3112 15140
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3480 15100 18232 15140
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18600 15100 33352 15140
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 33720 15100 48472 15140
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48840 15100 63592 15140
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63960 15100 78712 15140
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 79080 15100 89376 15140
rect 576 15076 89376 15100
rect 643 14552 701 14553
rect 643 14512 652 14552
rect 692 14512 701 14552
rect 643 14511 701 14512
rect 576 14384 89376 14408
rect 576 14344 4352 14384
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4720 14344 19472 14384
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19840 14344 34592 14384
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34960 14344 49712 14384
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 50080 14344 64832 14384
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 65200 14344 79952 14384
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 80320 14344 89376 14384
rect 576 14320 89376 14344
rect 576 13628 89376 13652
rect 576 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 18232 13628
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18600 13588 33352 13628
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33720 13588 48472 13628
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48840 13588 63592 13628
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63960 13588 78712 13628
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 79080 13588 89376 13628
rect 576 13564 89376 13588
rect 643 13040 701 13041
rect 643 13000 652 13040
rect 692 13000 701 13040
rect 643 12999 701 13000
rect 576 12872 89376 12896
rect 576 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 19472 12872
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19840 12832 34592 12872
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34960 12832 49712 12872
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 50080 12832 64832 12872
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 65200 12832 79952 12872
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 80320 12832 89376 12872
rect 576 12808 89376 12832
rect 643 12704 701 12705
rect 643 12664 652 12704
rect 692 12664 701 12704
rect 643 12663 701 12664
rect 576 12116 89376 12140
rect 576 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 18232 12116
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18600 12076 33352 12116
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33720 12076 48472 12116
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48840 12076 63592 12116
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63960 12076 78712 12116
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 79080 12076 89376 12116
rect 576 12052 89376 12076
rect 643 11528 701 11529
rect 643 11488 652 11528
rect 692 11488 701 11528
rect 643 11487 701 11488
rect 576 11360 89376 11384
rect 576 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 19472 11360
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19840 11320 34592 11360
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34960 11320 49712 11360
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 50080 11320 64832 11360
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 65200 11320 79952 11360
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 80320 11320 89376 11360
rect 576 11296 89376 11320
rect 643 11192 701 11193
rect 643 11152 652 11192
rect 692 11152 701 11192
rect 643 11151 701 11152
rect 576 10604 89376 10628
rect 576 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 18232 10604
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18600 10564 33352 10604
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33720 10564 48472 10604
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48840 10564 63592 10604
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63960 10564 78712 10604
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 79080 10564 89376 10604
rect 576 10540 89376 10564
rect 643 10016 701 10017
rect 643 9976 652 10016
rect 692 9976 701 10016
rect 643 9975 701 9976
rect 576 9848 89376 9872
rect 576 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 19472 9848
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19840 9808 34592 9848
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34960 9808 49712 9848
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 50080 9808 64832 9848
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 65200 9808 79952 9848
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 80320 9808 89376 9848
rect 576 9784 89376 9808
rect 643 9680 701 9681
rect 643 9640 652 9680
rect 692 9640 701 9680
rect 643 9639 701 9640
rect 576 9092 89376 9116
rect 576 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 18232 9092
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18600 9052 33352 9092
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33720 9052 48472 9092
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48840 9052 63592 9092
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63960 9052 78712 9092
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 79080 9052 89376 9092
rect 576 9028 89376 9052
rect 835 8756 893 8757
rect 835 8716 844 8756
rect 884 8716 893 8756
rect 835 8715 893 8716
rect 651 8504 693 8513
rect 651 8464 652 8504
rect 692 8464 693 8504
rect 651 8455 693 8464
rect 576 8336 89376 8360
rect 576 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 19472 8336
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19840 8296 34592 8336
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34960 8296 49712 8336
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 50080 8296 64832 8336
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 65200 8296 79952 8336
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 80320 8296 89376 8336
rect 576 8272 89376 8296
rect 835 7916 893 7917
rect 835 7876 844 7916
rect 884 7876 893 7916
rect 835 7875 893 7876
rect 651 7748 693 7757
rect 651 7708 652 7748
rect 692 7708 693 7748
rect 651 7699 693 7708
rect 576 7580 89376 7604
rect 576 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 18232 7580
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18600 7540 33352 7580
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33720 7540 48472 7580
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48840 7540 63592 7580
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63960 7540 78712 7580
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 79080 7540 89376 7580
rect 576 7516 89376 7540
rect 835 7244 893 7245
rect 835 7204 844 7244
rect 884 7204 893 7244
rect 835 7203 893 7204
rect 651 6992 693 7001
rect 651 6952 652 6992
rect 692 6952 693 6992
rect 651 6943 693 6952
rect 576 6824 89376 6848
rect 576 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 19472 6824
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19840 6784 34592 6824
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34960 6784 49712 6824
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 50080 6784 64832 6824
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 65200 6784 79952 6824
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 80320 6784 89376 6824
rect 576 6760 89376 6784
rect 576 6068 89376 6092
rect 576 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 18232 6068
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18600 6028 33352 6068
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33720 6028 48472 6068
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48840 6028 63592 6068
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63960 6028 78712 6068
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 79080 6028 89376 6068
rect 576 6004 89376 6028
rect 835 5732 893 5733
rect 835 5692 844 5732
rect 884 5692 893 5732
rect 835 5691 893 5692
rect 651 5480 693 5489
rect 651 5440 652 5480
rect 692 5440 693 5480
rect 651 5431 693 5440
rect 576 5312 89376 5336
rect 576 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 19472 5312
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19840 5272 34592 5312
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34960 5272 49712 5312
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 50080 5272 64832 5312
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 65200 5272 79952 5312
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 80320 5272 89376 5312
rect 576 5248 89376 5272
rect 835 4892 893 4893
rect 835 4852 844 4892
rect 884 4852 893 4892
rect 835 4851 893 4852
rect 651 4808 693 4817
rect 651 4768 652 4808
rect 692 4768 693 4808
rect 651 4759 693 4768
rect 576 4556 89376 4580
rect 576 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 18232 4556
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18600 4516 33352 4556
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33720 4516 48472 4556
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48840 4516 63592 4556
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63960 4516 78712 4556
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 79080 4516 89376 4556
rect 576 4492 89376 4516
rect 835 4220 893 4221
rect 835 4180 844 4220
rect 884 4180 893 4220
rect 835 4179 893 4180
rect 651 3968 693 3977
rect 651 3928 652 3968
rect 692 3928 693 3968
rect 651 3919 693 3928
rect 576 3800 89376 3824
rect 576 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 19472 3800
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19840 3760 34592 3800
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34960 3760 49712 3800
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 50080 3760 64832 3800
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 65200 3760 79952 3800
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 80320 3760 89376 3800
rect 576 3736 89376 3760
rect 835 3380 893 3381
rect 835 3340 844 3380
rect 884 3340 893 3380
rect 835 3339 893 3340
rect 651 3212 693 3221
rect 651 3172 652 3212
rect 692 3172 693 3212
rect 651 3163 693 3172
rect 576 3044 89376 3068
rect 576 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 18232 3044
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18600 3004 33352 3044
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33720 3004 48472 3044
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48840 3004 63592 3044
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63960 3004 78712 3044
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 79080 3004 89376 3044
rect 576 2980 89376 3004
rect 835 2708 893 2709
rect 835 2668 844 2708
rect 884 2668 893 2708
rect 835 2667 893 2668
rect 651 2456 693 2465
rect 651 2416 652 2456
rect 692 2416 693 2456
rect 651 2407 693 2416
rect 576 2288 89376 2312
rect 576 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 19472 2288
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19840 2248 34592 2288
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34960 2248 49712 2288
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 50080 2248 64832 2288
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 65200 2248 79952 2288
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 80320 2248 89376 2288
rect 576 2224 89376 2248
rect 576 1532 89376 1556
rect 576 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 18232 1532
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18600 1492 33352 1532
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33720 1492 48472 1532
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48840 1492 63592 1532
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63960 1492 78712 1532
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 79080 1492 89376 1532
rect 576 1468 89376 1492
rect 576 776 89376 800
rect 576 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 19472 776
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19840 736 34592 776
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34960 736 49712 776
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 50080 736 64832 776
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 65200 736 79952 776
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 80320 736 89376 776
rect 576 712 89376 736
<< via1 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 652 35092 692 35132
rect 844 34924 884 34964
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 652 34420 692 34460
rect 844 34168 884 34208
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 652 33580 692 33620
rect 844 33412 884 33452
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 652 32908 692 32948
rect 4300 32824 4340 32864
rect 4396 32824 4436 32864
rect 844 32656 884 32696
rect 4588 32656 4628 32696
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 4396 32152 4436 32192
rect 4492 32152 4532 32192
rect 652 32068 692 32108
rect 844 31900 884 31940
rect 4204 31900 4244 31940
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 652 31396 692 31436
rect 844 31144 884 31184
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 3820 30808 3860 30848
rect 2668 30640 2708 30680
rect 2860 30640 2900 30680
rect 3052 30640 3092 30680
rect 3244 30640 3284 30680
rect 3532 30640 3572 30680
rect 3628 30640 3668 30680
rect 3724 30640 3764 30680
rect 652 30556 692 30596
rect 3148 30472 3188 30512
rect 844 30388 884 30428
rect 2860 30388 2900 30428
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 652 29884 692 29924
rect 2284 29800 2324 29840
rect 2572 29800 2612 29840
rect 3244 29800 3284 29840
rect 3340 29800 3380 29840
rect 2764 29716 2804 29756
rect 844 29632 884 29672
rect 3052 29632 3092 29672
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 844 28540 884 28580
rect 652 28372 692 28412
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 844 27784 884 27824
rect 11404 27784 11444 27824
rect 11308 27616 11348 27656
rect 652 27532 692 27572
rect 11116 27364 11156 27404
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 3820 27028 3860 27068
rect 844 26944 884 26984
rect 10828 26944 10868 26984
rect 652 26860 692 26900
rect 3436 26776 3476 26816
rect 3628 26776 3668 26816
rect 3820 26776 3860 26816
rect 3916 26776 3956 26816
rect 4108 26776 4148 26816
rect 4204 26776 4244 26816
rect 4305 26776 4345 26816
rect 4780 26776 4820 26816
rect 4876 26776 4916 26816
rect 10828 26776 10868 26816
rect 11212 26776 11252 26816
rect 11500 26776 11540 26816
rect 3532 26608 3572 26648
rect 5164 26608 5204 26648
rect 11020 26608 11060 26648
rect 11692 26608 11732 26648
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 5260 26272 5300 26312
rect 3436 26104 3476 26144
rect 3628 26104 3668 26144
rect 5164 26104 5204 26144
rect 5356 26104 5396 26144
rect 11116 26104 11156 26144
rect 11308 26104 11348 26144
rect 11404 26104 11444 26144
rect 652 26020 692 26060
rect 3628 25936 3668 25976
rect 844 25852 884 25892
rect 11116 25852 11156 25892
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 844 25516 884 25556
rect 652 25348 692 25388
rect 12364 25348 12404 25388
rect 12556 25264 12596 25304
rect 12652 25264 12692 25304
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 10828 24760 10868 24800
rect 12076 24760 12116 24800
rect 4780 24676 4820 24716
rect 9772 24676 9812 24716
rect 4108 24592 4148 24632
rect 4204 24592 4244 24632
rect 4300 24592 4340 24632
rect 4684 24592 4724 24632
rect 5452 24592 5492 24632
rect 5548 24592 5588 24632
rect 6508 24592 6548 24632
rect 6604 24592 6644 24632
rect 9868 24592 9908 24632
rect 9964 24592 10004 24632
rect 10060 24592 10100 24632
rect 11020 24592 11060 24632
rect 11116 24592 11156 24632
rect 11980 24592 12020 24632
rect 12172 24592 12212 24632
rect 652 24508 692 24548
rect 844 24340 884 24380
rect 5356 24340 5396 24380
rect 6412 24340 6452 24380
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 63592 24172 63632 24212
rect 63674 24172 63714 24212
rect 63756 24172 63796 24212
rect 63838 24172 63878 24212
rect 63920 24172 63960 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 1900 24004 1940 24044
rect 4204 24004 4244 24044
rect 11404 24004 11444 24044
rect 652 23836 692 23876
rect 1804 23752 1844 23792
rect 1996 23752 2036 23792
rect 2188 23752 2228 23792
rect 2476 23752 2516 23792
rect 4108 23752 4148 23792
rect 4300 23752 4340 23792
rect 11212 23752 11252 23792
rect 11404 23752 11444 23792
rect 2668 23668 2708 23708
rect 844 23584 884 23624
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 64832 23416 64872 23456
rect 64914 23416 64954 23456
rect 64996 23416 65036 23456
rect 65078 23416 65118 23456
rect 65160 23416 65200 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 12076 23248 12116 23288
rect 12364 23248 12404 23288
rect 12268 23080 12308 23120
rect 652 22996 692 23036
rect 844 22828 884 22868
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 63592 22660 63632 22700
rect 63674 22660 63714 22700
rect 63756 22660 63796 22700
rect 63838 22660 63878 22700
rect 63920 22660 63960 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 11884 22324 11924 22364
rect 11308 22240 11348 22280
rect 11596 22240 11636 22280
rect 12076 22240 12116 22280
rect 12172 22240 12212 22280
rect 652 22072 692 22112
rect 11116 22072 11156 22112
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 64832 21904 64872 21944
rect 64914 21904 64954 21944
rect 64996 21904 65036 21944
rect 65078 21904 65118 21944
rect 65160 21904 65200 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 63592 21148 63632 21188
rect 63674 21148 63714 21188
rect 63756 21148 63796 21188
rect 63838 21148 63878 21188
rect 63920 21148 63960 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 8812 20896 8852 20936
rect 3436 20728 3476 20768
rect 3820 20728 3860 20768
rect 4108 20728 4148 20768
rect 8332 20728 8372 20768
rect 8524 20728 8564 20768
rect 8908 20728 8948 20768
rect 4300 20644 4340 20684
rect 652 20560 692 20600
rect 3340 20560 3380 20600
rect 4012 20560 4052 20600
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 64832 20392 64872 20432
rect 64914 20392 64954 20432
rect 64996 20392 65036 20432
rect 65078 20392 65118 20432
rect 65160 20392 65200 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 652 20224 692 20264
rect 8620 20224 8660 20264
rect 7852 20140 7892 20180
rect 8044 20056 8084 20096
rect 8332 20056 8372 20096
rect 8716 20056 8756 20096
rect 9100 20056 9140 20096
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 63592 19636 63632 19676
rect 63674 19636 63714 19676
rect 63756 19636 63796 19676
rect 63838 19636 63878 19676
rect 63920 19636 63960 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 8332 19468 8372 19508
rect 8140 19216 8180 19256
rect 652 19048 692 19088
rect 8044 19048 8084 19088
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 64832 18880 64872 18920
rect 64914 18880 64954 18920
rect 64996 18880 65036 18920
rect 65078 18880 65118 18920
rect 65160 18880 65200 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 652 18712 692 18752
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 63592 18124 63632 18164
rect 63674 18124 63714 18164
rect 63756 18124 63796 18164
rect 63838 18124 63878 18164
rect 63920 18124 63960 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 652 17536 692 17576
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 64832 17368 64872 17408
rect 64914 17368 64954 17408
rect 64996 17368 65036 17408
rect 65078 17368 65118 17408
rect 65160 17368 65200 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 652 17200 692 17240
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 63592 16612 63632 16652
rect 63674 16612 63714 16652
rect 63756 16612 63796 16652
rect 63838 16612 63878 16652
rect 63920 16612 63960 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 652 16024 692 16064
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 64832 15856 64872 15896
rect 64914 15856 64954 15896
rect 64996 15856 65036 15896
rect 65078 15856 65118 15896
rect 65160 15856 65200 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 652 15688 692 15728
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 652 14512 692 14552
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 652 13000 692 13040
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 652 12664 692 12704
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 652 11488 692 11528
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 652 11152 692 11192
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 652 9976 692 10016
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 652 9640 692 9680
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 844 8716 884 8756
rect 652 8464 692 8504
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 844 7876 884 7916
rect 652 7708 692 7748
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 844 7204 884 7244
rect 652 6952 692 6992
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 844 5692 884 5732
rect 652 5440 692 5480
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 844 4852 884 4892
rect 652 4768 692 4808
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 844 4180 884 4220
rect 652 3928 692 3968
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 844 3340 884 3380
rect 652 3172 692 3212
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 844 2668 884 2708
rect 652 2416 692 2456
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
<< metal2 >>
rect 4352 38576 4720 38585
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4352 38527 4720 38536
rect 19472 38576 19840 38585
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19472 38527 19840 38536
rect 34592 38576 34960 38585
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34592 38527 34960 38536
rect 49712 38576 50080 38585
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 49712 38527 50080 38536
rect 64832 38576 65200 38585
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 64832 38527 65200 38536
rect 79952 38576 80320 38585
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 79952 38527 80320 38536
rect 3112 37820 3480 37829
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3112 37771 3480 37780
rect 18232 37820 18600 37829
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18232 37771 18600 37780
rect 33352 37820 33720 37829
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33352 37771 33720 37780
rect 48472 37820 48840 37829
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48472 37771 48840 37780
rect 63592 37820 63960 37829
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63592 37771 63960 37780
rect 78712 37820 79080 37829
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 78712 37771 79080 37780
rect 4352 37064 4720 37073
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4352 37015 4720 37024
rect 19472 37064 19840 37073
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19472 37015 19840 37024
rect 34592 37064 34960 37073
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34592 37015 34960 37024
rect 49712 37064 50080 37073
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 49712 37015 50080 37024
rect 64832 37064 65200 37073
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 64832 37015 65200 37024
rect 79952 37064 80320 37073
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 79952 37015 80320 37024
rect 3112 36308 3480 36317
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3112 36259 3480 36268
rect 18232 36308 18600 36317
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18232 36259 18600 36268
rect 33352 36308 33720 36317
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33352 36259 33720 36268
rect 48472 36308 48840 36317
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48472 36259 48840 36268
rect 63592 36308 63960 36317
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63592 36259 63960 36268
rect 78712 36308 79080 36317
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 78712 36259 79080 36268
rect 4352 35552 4720 35561
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4352 35503 4720 35512
rect 19472 35552 19840 35561
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19472 35503 19840 35512
rect 34592 35552 34960 35561
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34592 35503 34960 35512
rect 49712 35552 50080 35561
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 49712 35503 50080 35512
rect 64832 35552 65200 35561
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 64832 35503 65200 35512
rect 79952 35552 80320 35561
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 79952 35503 80320 35512
rect 651 35132 693 35141
rect 651 35092 652 35132
rect 692 35092 693 35132
rect 651 35083 693 35092
rect 652 34998 692 35083
rect 844 34964 884 34973
rect 748 34924 844 34964
rect 652 34460 692 34469
rect 652 34217 692 34420
rect 651 34208 693 34217
rect 651 34168 652 34208
rect 692 34168 693 34208
rect 651 34159 693 34168
rect 748 33629 788 34924
rect 844 34915 884 34924
rect 3112 34796 3480 34805
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3112 34747 3480 34756
rect 18232 34796 18600 34805
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18232 34747 18600 34756
rect 33352 34796 33720 34805
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33352 34747 33720 34756
rect 48472 34796 48840 34805
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48472 34747 48840 34756
rect 63592 34796 63960 34805
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63592 34747 63960 34756
rect 78712 34796 79080 34805
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 78712 34747 79080 34756
rect 844 34208 884 34217
rect 884 34168 1076 34208
rect 844 34159 884 34168
rect 652 33620 692 33629
rect 652 33377 692 33580
rect 747 33620 789 33629
rect 747 33580 748 33620
rect 788 33580 789 33620
rect 747 33571 789 33580
rect 844 33452 884 33461
rect 748 33412 844 33452
rect 651 33368 693 33377
rect 651 33328 652 33368
rect 692 33328 693 33368
rect 651 33319 693 33328
rect 748 33116 788 33412
rect 844 33403 884 33412
rect 460 33076 788 33116
rect 363 31520 405 31529
rect 363 31480 364 31520
rect 404 31480 405 31520
rect 363 31471 405 31480
rect 364 26732 404 31471
rect 460 26909 500 33076
rect 652 32948 692 32957
rect 652 32537 692 32908
rect 844 32696 884 32705
rect 748 32656 844 32696
rect 651 32528 693 32537
rect 651 32488 652 32528
rect 692 32488 693 32528
rect 651 32479 693 32488
rect 652 32108 692 32117
rect 555 31940 597 31949
rect 555 31900 556 31940
rect 596 31900 597 31940
rect 555 31891 597 31900
rect 556 26993 596 31891
rect 652 31697 692 32068
rect 651 31688 693 31697
rect 651 31648 652 31688
rect 692 31648 693 31688
rect 651 31639 693 31648
rect 652 31436 692 31445
rect 652 30857 692 31396
rect 651 30848 693 30857
rect 651 30808 652 30848
rect 692 30808 693 30848
rect 651 30799 693 30808
rect 652 30596 692 30605
rect 652 30101 692 30556
rect 651 30092 693 30101
rect 651 30052 652 30092
rect 692 30052 693 30092
rect 651 30043 693 30052
rect 652 29924 692 29933
rect 652 29177 692 29884
rect 748 29504 788 32656
rect 844 32647 884 32656
rect 843 31940 885 31949
rect 843 31900 844 31940
rect 884 31900 885 31940
rect 843 31891 885 31900
rect 844 31806 884 31891
rect 844 31184 884 31193
rect 884 31144 980 31184
rect 844 31135 884 31144
rect 844 30428 884 30437
rect 844 29933 884 30388
rect 843 29924 885 29933
rect 843 29884 844 29924
rect 884 29884 885 29924
rect 843 29875 885 29884
rect 844 29681 884 29766
rect 843 29672 885 29681
rect 843 29632 844 29672
rect 884 29632 885 29672
rect 843 29623 885 29632
rect 940 29588 980 31144
rect 1036 30689 1076 34168
rect 4352 34040 4720 34049
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4352 33991 4720 34000
rect 19472 34040 19840 34049
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19472 33991 19840 34000
rect 34592 34040 34960 34049
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34592 33991 34960 34000
rect 49712 34040 50080 34049
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 49712 33991 50080 34000
rect 64832 34040 65200 34049
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 64832 33991 65200 34000
rect 79952 34040 80320 34049
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 79952 33991 80320 34000
rect 4395 33620 4437 33629
rect 4395 33580 4396 33620
rect 4436 33580 4437 33620
rect 4395 33571 4437 33580
rect 3112 33284 3480 33293
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3112 33235 3480 33244
rect 4300 32864 4340 32873
rect 4300 32780 4340 32824
rect 4396 32864 4436 33571
rect 18232 33284 18600 33293
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18232 33235 18600 33244
rect 33352 33284 33720 33293
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33352 33235 33720 33244
rect 48472 33284 48840 33293
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48472 33235 48840 33244
rect 63592 33284 63960 33293
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63592 33235 63960 33244
rect 78712 33284 79080 33293
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 78712 33235 79080 33244
rect 4396 32815 4436 32824
rect 4108 32740 4340 32780
rect 3819 32192 3861 32201
rect 3819 32152 3820 32192
rect 3860 32152 3861 32192
rect 3819 32143 3861 32152
rect 3112 31772 3480 31781
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3112 31723 3480 31732
rect 3820 30848 3860 32143
rect 3820 30799 3860 30808
rect 3244 30689 3284 30774
rect 1035 30680 1077 30689
rect 1035 30640 1036 30680
rect 1076 30640 1077 30680
rect 1035 30631 1077 30640
rect 2571 30680 2613 30689
rect 2571 30640 2572 30680
rect 2612 30640 2613 30680
rect 2571 30631 2613 30640
rect 2668 30680 2708 30689
rect 2283 29840 2325 29849
rect 2283 29800 2284 29840
rect 2324 29800 2325 29840
rect 2283 29791 2325 29800
rect 2572 29840 2612 30631
rect 2668 30605 2708 30640
rect 2859 30680 2901 30689
rect 2859 30640 2860 30680
rect 2900 30640 2901 30680
rect 2859 30631 2901 30640
rect 3051 30680 3093 30689
rect 3051 30640 3052 30680
rect 3092 30640 3093 30680
rect 3051 30631 3093 30640
rect 3243 30680 3285 30689
rect 3243 30640 3244 30680
rect 3284 30640 3285 30680
rect 3243 30631 3285 30640
rect 3532 30680 3572 30689
rect 2667 30596 2709 30605
rect 2667 30556 2668 30596
rect 2708 30556 2709 30596
rect 2667 30547 2709 30556
rect 2668 29849 2708 30547
rect 2860 30546 2900 30631
rect 3052 30546 3092 30631
rect 3148 30521 3188 30606
rect 3147 30512 3189 30521
rect 3147 30472 3148 30512
rect 3188 30472 3189 30512
rect 3147 30463 3189 30472
rect 2859 30428 2901 30437
rect 2859 30388 2860 30428
rect 2900 30388 2901 30428
rect 2859 30379 2901 30388
rect 2860 30294 2900 30379
rect 3112 30260 3480 30269
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3112 30211 3480 30220
rect 3532 29849 3572 30640
rect 3628 30680 3668 30689
rect 3628 30437 3668 30640
rect 3724 30680 3764 30689
rect 3724 30521 3764 30640
rect 3723 30512 3765 30521
rect 3723 30472 3724 30512
rect 3764 30472 3765 30512
rect 3723 30463 3765 30472
rect 3627 30428 3669 30437
rect 3627 30388 3628 30428
rect 3668 30388 3669 30428
rect 3627 30379 3669 30388
rect 2572 29791 2612 29800
rect 2667 29840 2709 29849
rect 3244 29840 3284 29849
rect 2667 29800 2668 29840
rect 2708 29800 2709 29840
rect 2667 29791 2709 29800
rect 2764 29800 3244 29840
rect 1227 29672 1269 29681
rect 1227 29632 1228 29672
rect 1268 29632 1269 29672
rect 1227 29623 1269 29632
rect 2091 29672 2133 29681
rect 2091 29632 2092 29672
rect 2132 29632 2133 29672
rect 2091 29623 2133 29632
rect 940 29548 1076 29588
rect 748 29464 980 29504
rect 747 29336 789 29345
rect 747 29296 748 29336
rect 788 29296 789 29336
rect 747 29287 789 29296
rect 651 29168 693 29177
rect 651 29128 652 29168
rect 692 29128 693 29168
rect 651 29119 693 29128
rect 651 28412 693 28421
rect 651 28372 652 28412
rect 692 28372 693 28412
rect 651 28363 693 28372
rect 652 28278 692 28363
rect 748 27824 788 29287
rect 843 29000 885 29009
rect 843 28960 844 29000
rect 884 28960 885 29000
rect 843 28951 885 28960
rect 844 28580 884 28951
rect 844 28531 884 28540
rect 844 27824 884 27833
rect 748 27784 844 27824
rect 844 27775 884 27784
rect 651 27572 693 27581
rect 651 27532 652 27572
rect 692 27532 693 27572
rect 651 27523 693 27532
rect 652 27438 692 27523
rect 555 26984 597 26993
rect 555 26944 556 26984
rect 596 26944 597 26984
rect 555 26935 597 26944
rect 844 26984 884 26993
rect 459 26900 501 26909
rect 459 26860 460 26900
rect 500 26860 501 26900
rect 459 26851 501 26860
rect 652 26900 692 26909
rect 364 26692 596 26732
rect 459 25220 501 25229
rect 459 25180 460 25220
rect 500 25180 501 25220
rect 459 25171 501 25180
rect 363 20096 405 20105
rect 363 20056 364 20096
rect 404 20056 405 20096
rect 363 20047 405 20056
rect 364 11360 404 20047
rect 460 15821 500 25171
rect 556 16232 596 26692
rect 652 26657 692 26860
rect 844 26825 884 26944
rect 940 26900 980 29464
rect 1036 27077 1076 29548
rect 1131 27152 1173 27161
rect 1131 27112 1132 27152
rect 1172 27112 1173 27152
rect 1131 27103 1173 27112
rect 1035 27068 1077 27077
rect 1035 27028 1036 27068
rect 1076 27028 1077 27068
rect 1035 27019 1077 27028
rect 940 26860 1076 26900
rect 843 26816 885 26825
rect 843 26776 844 26816
rect 884 26776 885 26816
rect 843 26767 885 26776
rect 651 26648 693 26657
rect 651 26608 652 26648
rect 692 26608 693 26648
rect 651 26599 693 26608
rect 652 26060 692 26069
rect 652 25817 692 26020
rect 844 25892 884 25901
rect 748 25852 844 25892
rect 651 25808 693 25817
rect 651 25768 652 25808
rect 692 25768 693 25808
rect 651 25759 693 25768
rect 652 25388 692 25397
rect 652 24977 692 25348
rect 651 24968 693 24977
rect 651 24928 652 24968
rect 692 24928 693 24968
rect 651 24919 693 24928
rect 652 24548 692 24557
rect 652 24137 692 24508
rect 651 24128 693 24137
rect 651 24088 652 24128
rect 692 24088 693 24128
rect 651 24079 693 24088
rect 652 23876 692 23885
rect 652 23297 692 23836
rect 748 23801 788 25852
rect 844 25843 884 25852
rect 843 25556 885 25565
rect 843 25516 844 25556
rect 884 25516 885 25556
rect 843 25507 885 25516
rect 844 25422 884 25507
rect 843 24380 885 24389
rect 843 24340 844 24380
rect 884 24340 885 24380
rect 843 24331 885 24340
rect 844 24246 884 24331
rect 1036 23885 1076 26860
rect 1132 25565 1172 27103
rect 1131 25556 1173 25565
rect 1131 25516 1132 25556
rect 1172 25516 1173 25556
rect 1131 25507 1173 25516
rect 1131 24128 1173 24137
rect 1131 24088 1132 24128
rect 1172 24088 1173 24128
rect 1131 24079 1173 24088
rect 1035 23876 1077 23885
rect 1035 23836 1036 23876
rect 1076 23836 1077 23876
rect 1035 23827 1077 23836
rect 747 23792 789 23801
rect 747 23752 748 23792
rect 788 23752 789 23792
rect 747 23743 789 23752
rect 844 23624 884 23633
rect 884 23584 980 23624
rect 844 23575 884 23584
rect 651 23288 693 23297
rect 651 23248 652 23288
rect 692 23248 693 23288
rect 651 23239 693 23248
rect 652 23036 692 23045
rect 652 22457 692 22996
rect 844 22868 884 22877
rect 651 22448 693 22457
rect 651 22408 652 22448
rect 692 22408 693 22448
rect 651 22399 693 22408
rect 652 22112 692 22121
rect 652 21617 692 22072
rect 651 21608 693 21617
rect 651 21568 652 21608
rect 692 21568 693 21608
rect 651 21559 693 21568
rect 844 20777 884 22828
rect 651 20768 693 20777
rect 651 20728 652 20768
rect 692 20728 693 20768
rect 651 20719 693 20728
rect 843 20768 885 20777
rect 843 20728 844 20768
rect 884 20728 885 20768
rect 843 20719 885 20728
rect 652 20600 692 20719
rect 652 20551 692 20560
rect 652 20264 692 20273
rect 652 19937 692 20224
rect 651 19928 693 19937
rect 651 19888 652 19928
rect 692 19888 693 19928
rect 651 19879 693 19888
rect 940 19097 980 23584
rect 1035 22112 1077 22121
rect 1035 22072 1036 22112
rect 1076 22072 1077 22112
rect 1035 22063 1077 22072
rect 651 19088 693 19097
rect 651 19048 652 19088
rect 692 19048 693 19088
rect 651 19039 693 19048
rect 939 19088 981 19097
rect 939 19048 940 19088
rect 980 19048 981 19088
rect 939 19039 981 19048
rect 652 18954 692 19039
rect 652 18752 692 18761
rect 652 18257 692 18712
rect 651 18248 693 18257
rect 651 18208 652 18248
rect 692 18208 693 18248
rect 651 18199 693 18208
rect 652 17576 692 17585
rect 652 17417 692 17536
rect 651 17408 693 17417
rect 651 17368 652 17408
rect 692 17368 693 17408
rect 651 17359 693 17368
rect 652 17240 692 17249
rect 652 16577 692 17200
rect 651 16568 693 16577
rect 651 16528 652 16568
rect 692 16528 693 16568
rect 651 16519 693 16528
rect 556 16192 788 16232
rect 652 16064 692 16073
rect 556 16024 652 16064
rect 459 15812 501 15821
rect 459 15772 460 15812
rect 500 15772 501 15812
rect 459 15763 501 15772
rect 556 15737 596 16024
rect 652 16015 692 16024
rect 555 15728 597 15737
rect 555 15688 556 15728
rect 596 15688 597 15728
rect 555 15679 597 15688
rect 652 15728 692 15737
rect 652 14897 692 15688
rect 651 14888 693 14897
rect 651 14848 652 14888
rect 692 14848 693 14888
rect 651 14839 693 14848
rect 652 14552 692 14561
rect 652 14057 692 14512
rect 651 14048 693 14057
rect 651 14008 652 14048
rect 692 14008 693 14048
rect 651 13999 693 14008
rect 651 13208 693 13217
rect 651 13168 652 13208
rect 692 13168 693 13208
rect 651 13159 693 13168
rect 652 13040 692 13159
rect 652 12991 692 13000
rect 652 12704 692 12713
rect 652 12377 692 12664
rect 651 12368 693 12377
rect 651 12328 652 12368
rect 692 12328 693 12368
rect 651 12319 693 12328
rect 651 11528 693 11537
rect 651 11488 652 11528
rect 692 11488 693 11528
rect 651 11479 693 11488
rect 652 11394 692 11479
rect 748 11360 788 16192
rect 939 15812 981 15821
rect 939 15772 940 15812
rect 980 15772 981 15812
rect 939 15763 981 15772
rect 364 11320 596 11360
rect 748 11320 884 11360
rect 556 6320 596 11320
rect 652 11192 692 11201
rect 652 10697 692 11152
rect 651 10688 693 10697
rect 651 10648 652 10688
rect 692 10648 693 10688
rect 651 10639 693 10648
rect 652 10016 692 10025
rect 652 9857 692 9976
rect 651 9848 693 9857
rect 651 9808 652 9848
rect 692 9808 693 9848
rect 651 9799 693 9808
rect 652 9680 692 9689
rect 652 9017 692 9640
rect 651 9008 693 9017
rect 651 8968 652 9008
rect 692 8968 693 9008
rect 651 8959 693 8968
rect 844 8756 884 11320
rect 844 8707 884 8716
rect 652 8504 692 8513
rect 652 8177 692 8464
rect 651 8168 693 8177
rect 651 8128 652 8168
rect 692 8128 693 8168
rect 651 8119 693 8128
rect 843 7916 885 7925
rect 843 7876 844 7916
rect 884 7876 885 7916
rect 843 7867 885 7876
rect 844 7782 884 7867
rect 652 7748 692 7757
rect 652 7337 692 7708
rect 651 7328 693 7337
rect 651 7288 652 7328
rect 692 7288 693 7328
rect 651 7279 693 7288
rect 843 7244 885 7253
rect 843 7204 844 7244
rect 884 7204 885 7244
rect 843 7195 885 7204
rect 844 7110 884 7195
rect 652 6992 692 7001
rect 652 6497 692 6952
rect 651 6488 693 6497
rect 651 6448 652 6488
rect 692 6448 693 6488
rect 651 6439 693 6448
rect 556 6280 788 6320
rect 651 5648 693 5657
rect 651 5608 652 5648
rect 692 5608 693 5648
rect 651 5599 693 5608
rect 652 5480 692 5599
rect 652 5431 692 5440
rect 651 4808 693 4817
rect 651 4768 652 4808
rect 692 4768 693 4808
rect 651 4759 693 4768
rect 652 4674 692 4759
rect 651 3968 693 3977
rect 651 3928 652 3968
rect 692 3928 693 3968
rect 651 3919 693 3928
rect 652 3834 692 3919
rect 748 3380 788 6280
rect 843 5732 885 5741
rect 843 5692 844 5732
rect 884 5692 885 5732
rect 843 5683 885 5692
rect 844 5598 884 5683
rect 844 4892 884 4901
rect 940 4892 980 15763
rect 884 4852 980 4892
rect 844 4843 884 4852
rect 844 4220 884 4229
rect 1036 4220 1076 22063
rect 1132 7253 1172 24079
rect 1228 20861 1268 29623
rect 1900 24053 1940 24138
rect 1899 24044 1941 24053
rect 1899 24004 1900 24044
rect 1940 24004 1941 24044
rect 1899 23995 1941 24004
rect 1803 23876 1845 23885
rect 1803 23836 1804 23876
rect 1844 23836 1845 23876
rect 1803 23827 1845 23836
rect 1804 23792 1844 23827
rect 1804 23741 1844 23752
rect 1995 23792 2037 23801
rect 1995 23752 1996 23792
rect 2036 23752 2037 23792
rect 1995 23743 2037 23752
rect 1996 23658 2036 23743
rect 1227 20852 1269 20861
rect 1227 20812 1228 20852
rect 1268 20812 1269 20852
rect 1227 20803 1269 20812
rect 1227 19844 1269 19853
rect 1227 19804 1228 19844
rect 1268 19804 1269 19844
rect 1227 19795 1269 19804
rect 1131 7244 1173 7253
rect 1131 7204 1132 7244
rect 1172 7204 1173 7244
rect 1131 7195 1173 7204
rect 884 4180 1076 4220
rect 844 4171 884 4180
rect 844 3380 884 3389
rect 748 3340 844 3380
rect 844 3331 884 3340
rect 651 3212 693 3221
rect 651 3172 652 3212
rect 692 3172 693 3212
rect 651 3163 693 3172
rect 652 3078 692 3163
rect 844 2708 884 2717
rect 1228 2708 1268 19795
rect 2092 7925 2132 29623
rect 2284 29345 2324 29791
rect 2764 29756 2804 29800
rect 3244 29791 3284 29800
rect 3339 29840 3381 29849
rect 3339 29800 3340 29840
rect 3380 29800 3381 29840
rect 3339 29791 3381 29800
rect 3531 29840 3573 29849
rect 3531 29800 3532 29840
rect 3572 29800 3573 29840
rect 3531 29791 3573 29800
rect 3819 29840 3861 29849
rect 3819 29800 3820 29840
rect 3860 29800 3861 29840
rect 3819 29791 3861 29800
rect 2764 29707 2804 29716
rect 3340 29706 3380 29791
rect 3051 29672 3093 29681
rect 3051 29632 3052 29672
rect 3092 29632 3093 29672
rect 3051 29623 3093 29632
rect 3052 29538 3092 29623
rect 2283 29336 2325 29345
rect 2283 29296 2284 29336
rect 2324 29296 2325 29336
rect 2283 29287 2325 29296
rect 3112 28748 3480 28757
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3112 28699 3480 28708
rect 3112 27236 3480 27245
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3112 27187 3480 27196
rect 3820 27068 3860 29791
rect 4108 29009 4148 32740
rect 4588 32696 4628 32705
rect 4628 32656 4820 32696
rect 4588 32647 4628 32656
rect 4352 32528 4720 32537
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4352 32479 4720 32488
rect 4395 32192 4437 32201
rect 4395 32152 4396 32192
rect 4436 32152 4437 32192
rect 4395 32143 4437 32152
rect 4492 32192 4532 32201
rect 4780 32192 4820 32656
rect 19472 32528 19840 32537
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19472 32479 19840 32488
rect 34592 32528 34960 32537
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34592 32479 34960 32488
rect 49712 32528 50080 32537
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 49712 32479 50080 32488
rect 64832 32528 65200 32537
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 64832 32479 65200 32488
rect 79952 32528 80320 32537
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 79952 32479 80320 32488
rect 4532 32152 4820 32192
rect 4492 32143 4532 32152
rect 4396 32058 4436 32143
rect 4204 31940 4244 31949
rect 4204 31529 4244 31900
rect 18232 31772 18600 31781
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18232 31723 18600 31732
rect 33352 31772 33720 31781
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33352 31723 33720 31732
rect 48472 31772 48840 31781
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48472 31723 48840 31732
rect 63592 31772 63960 31781
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63592 31723 63960 31732
rect 78712 31772 79080 31781
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 78712 31723 79080 31732
rect 4203 31520 4245 31529
rect 4203 31480 4204 31520
rect 4244 31480 4245 31520
rect 4203 31471 4245 31480
rect 4352 31016 4720 31025
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4352 30967 4720 30976
rect 19472 31016 19840 31025
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19472 30967 19840 30976
rect 34592 31016 34960 31025
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34592 30967 34960 30976
rect 49712 31016 50080 31025
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 49712 30967 50080 30976
rect 64832 31016 65200 31025
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 64832 30967 65200 30976
rect 79952 31016 80320 31025
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 79952 30967 80320 30976
rect 18232 30260 18600 30269
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18232 30211 18600 30220
rect 33352 30260 33720 30269
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33352 30211 33720 30220
rect 48472 30260 48840 30269
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48472 30211 48840 30220
rect 63592 30260 63960 30269
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63592 30211 63960 30220
rect 78712 30260 79080 30269
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 78712 30211 79080 30220
rect 8715 29924 8757 29933
rect 8715 29884 8716 29924
rect 8756 29884 8757 29924
rect 8715 29875 8757 29884
rect 4352 29504 4720 29513
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4352 29455 4720 29464
rect 4107 29000 4149 29009
rect 4107 28960 4108 29000
rect 4148 28960 4149 29000
rect 4107 28951 4149 28960
rect 4352 27992 4720 28001
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4352 27943 4720 27952
rect 3820 27019 3860 27028
rect 3627 26900 3669 26909
rect 3627 26860 3628 26900
rect 3668 26860 3669 26900
rect 3627 26851 3669 26860
rect 4304 26900 4346 26909
rect 4304 26860 4305 26900
rect 4345 26860 4346 26900
rect 4304 26851 4346 26860
rect 4779 26900 4821 26909
rect 4779 26860 4780 26900
rect 4820 26860 4821 26900
rect 4779 26851 4821 26860
rect 3435 26816 3477 26825
rect 3435 26776 3436 26816
rect 3476 26776 3477 26816
rect 3435 26767 3477 26776
rect 3628 26816 3668 26851
rect 3820 26816 3860 26825
rect 3436 26682 3476 26767
rect 3628 26765 3668 26776
rect 3724 26776 3820 26816
rect 3532 26648 3572 26657
rect 3572 26608 3668 26648
rect 3532 26599 3572 26608
rect 3436 26144 3476 26153
rect 3628 26144 3668 26608
rect 3476 26104 3572 26144
rect 3436 26095 3476 26104
rect 3112 25724 3480 25733
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3112 25675 3480 25684
rect 3112 24212 3480 24221
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3112 24163 3480 24172
rect 3532 24053 3572 26104
rect 3628 26095 3668 26104
rect 3628 25976 3668 25985
rect 3724 25976 3764 26776
rect 3820 26767 3860 26776
rect 3915 26816 3957 26825
rect 4108 26816 4148 26825
rect 3915 26776 3916 26816
rect 3956 26776 3957 26816
rect 3915 26767 3957 26776
rect 4012 26776 4108 26816
rect 3916 26682 3956 26767
rect 3668 25936 3764 25976
rect 3628 25927 3668 25936
rect 4012 24557 4052 26776
rect 4108 26767 4148 26776
rect 4204 26816 4244 26827
rect 4204 26741 4244 26776
rect 4305 26816 4345 26851
rect 4305 26765 4345 26776
rect 4780 26816 4820 26851
rect 4780 26765 4820 26776
rect 4876 26816 4916 26827
rect 4876 26741 4916 26776
rect 5259 26816 5301 26825
rect 5259 26776 5260 26816
rect 5300 26776 5301 26816
rect 5259 26767 5301 26776
rect 4203 26732 4245 26741
rect 4203 26692 4204 26732
rect 4244 26692 4245 26732
rect 4203 26683 4245 26692
rect 4875 26732 4917 26741
rect 4875 26692 4876 26732
rect 4916 26692 4917 26732
rect 4875 26683 4917 26692
rect 5164 26648 5204 26657
rect 4352 26480 4720 26489
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4352 26431 4720 26440
rect 5164 26153 5204 26608
rect 5260 26312 5300 26767
rect 5260 26263 5300 26272
rect 5163 26144 5205 26153
rect 5163 26104 5164 26144
rect 5204 26104 5205 26144
rect 5163 26095 5205 26104
rect 5356 26144 5396 26153
rect 5164 26010 5204 26095
rect 4352 24968 4720 24977
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4352 24919 4720 24928
rect 5356 24725 5396 26104
rect 5547 26144 5589 26153
rect 5547 26104 5548 26144
rect 5588 26104 5589 26144
rect 5547 26095 5589 26104
rect 4779 24716 4821 24725
rect 4779 24676 4780 24716
rect 4820 24676 4821 24716
rect 4779 24667 4821 24676
rect 5355 24716 5397 24725
rect 5355 24676 5356 24716
rect 5396 24676 5397 24716
rect 5355 24667 5397 24676
rect 4108 24632 4148 24641
rect 4011 24548 4053 24557
rect 4011 24508 4012 24548
rect 4052 24508 4053 24548
rect 4011 24499 4053 24508
rect 3531 24044 3573 24053
rect 3531 24004 3532 24044
rect 3572 24004 3573 24044
rect 3531 23995 3573 24004
rect 4012 23960 4052 24499
rect 4108 24044 4148 24592
rect 4203 24632 4245 24641
rect 4203 24592 4204 24632
rect 4244 24592 4245 24632
rect 4203 24583 4245 24592
rect 4300 24632 4340 24641
rect 4204 24498 4244 24583
rect 4300 24053 4340 24592
rect 4684 24632 4724 24641
rect 4204 24044 4244 24053
rect 4108 24004 4204 24044
rect 4204 23995 4244 24004
rect 4299 24044 4341 24053
rect 4299 24004 4300 24044
rect 4340 24004 4341 24044
rect 4299 23995 4341 24004
rect 4012 23920 4148 23960
rect 2475 23876 2517 23885
rect 2475 23836 2476 23876
rect 2516 23836 2517 23876
rect 2475 23827 2517 23836
rect 2187 23792 2229 23801
rect 2187 23752 2188 23792
rect 2228 23752 2229 23792
rect 2187 23743 2229 23752
rect 2476 23792 2516 23827
rect 2188 23658 2228 23743
rect 2476 23741 2516 23752
rect 4108 23792 4148 23920
rect 4108 23743 4148 23752
rect 4300 23792 4340 23803
rect 4300 23717 4340 23752
rect 4684 23717 4724 24592
rect 4780 24582 4820 24667
rect 5451 24632 5493 24641
rect 5451 24592 5452 24632
rect 5492 24592 5493 24632
rect 5451 24583 5493 24592
rect 5548 24632 5588 26095
rect 6603 24716 6645 24725
rect 6603 24676 6604 24716
rect 6644 24676 6645 24716
rect 6603 24667 6645 24676
rect 5548 24583 5588 24592
rect 6507 24632 6549 24641
rect 6507 24592 6508 24632
rect 6548 24592 6549 24632
rect 6507 24583 6549 24592
rect 6604 24632 6644 24667
rect 5452 24498 5492 24583
rect 6508 24498 6548 24583
rect 6604 24557 6644 24592
rect 6603 24548 6645 24557
rect 6603 24508 6604 24548
rect 6644 24508 6645 24548
rect 6603 24499 6645 24508
rect 6604 24468 6644 24499
rect 5356 24380 5396 24389
rect 5356 24137 5396 24340
rect 6412 24380 6452 24389
rect 5355 24128 5397 24137
rect 5355 24088 5356 24128
rect 5396 24088 5397 24128
rect 5355 24079 5397 24088
rect 2667 23708 2709 23717
rect 2667 23668 2668 23708
rect 2708 23668 2709 23708
rect 2667 23659 2709 23668
rect 4299 23708 4341 23717
rect 4299 23668 4300 23708
rect 4340 23668 4341 23708
rect 4299 23659 4341 23668
rect 4683 23708 4725 23717
rect 4683 23668 4684 23708
rect 4724 23668 4725 23708
rect 4683 23659 4725 23668
rect 2668 23574 2708 23659
rect 4352 23456 4720 23465
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4352 23407 4720 23416
rect 3112 22700 3480 22709
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3112 22651 3480 22660
rect 4352 21944 4720 21953
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4352 21895 4720 21904
rect 3112 21188 3480 21197
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3112 21139 3480 21148
rect 3435 20852 3477 20861
rect 3435 20812 3436 20852
rect 3476 20812 3477 20852
rect 3435 20803 3477 20812
rect 4107 20852 4149 20861
rect 4107 20812 4108 20852
rect 4148 20812 4149 20852
rect 4107 20803 4149 20812
rect 3436 20768 3476 20803
rect 3436 20717 3476 20728
rect 3819 20768 3861 20777
rect 3819 20728 3820 20768
rect 3860 20728 3861 20768
rect 3819 20719 3861 20728
rect 4011 20768 4053 20777
rect 4011 20728 4012 20768
rect 4052 20728 4053 20768
rect 4011 20719 4053 20728
rect 4108 20768 4148 20803
rect 3820 20634 3860 20719
rect 3340 20600 3380 20609
rect 3340 19853 3380 20560
rect 4012 20600 4052 20719
rect 4108 20717 4148 20728
rect 4299 20684 4341 20693
rect 4299 20644 4300 20684
rect 4340 20644 4341 20684
rect 4299 20635 4341 20644
rect 4012 20551 4052 20560
rect 4300 20550 4340 20635
rect 4352 20432 4720 20441
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4352 20383 4720 20392
rect 3339 19844 3381 19853
rect 3339 19804 3340 19844
rect 3380 19804 3381 19844
rect 3339 19795 3381 19804
rect 3112 19676 3480 19685
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3112 19627 3480 19636
rect 4352 18920 4720 18929
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4352 18871 4720 18880
rect 3112 18164 3480 18173
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3112 18115 3480 18124
rect 4352 17408 4720 17417
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4352 17359 4720 17368
rect 3112 16652 3480 16661
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3112 16603 3480 16612
rect 4352 15896 4720 15905
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4352 15847 4720 15856
rect 3112 15140 3480 15149
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3112 15091 3480 15100
rect 4352 14384 4720 14393
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4352 14335 4720 14344
rect 3112 13628 3480 13637
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3112 13579 3480 13588
rect 4352 12872 4720 12881
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4352 12823 4720 12832
rect 3112 12116 3480 12125
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3112 12067 3480 12076
rect 4352 11360 4720 11369
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4352 11311 4720 11320
rect 3112 10604 3480 10613
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3112 10555 3480 10564
rect 4352 9848 4720 9857
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4352 9799 4720 9808
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 2091 7916 2133 7925
rect 2091 7876 2092 7916
rect 2132 7876 2133 7916
rect 2091 7867 2133 7876
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 6412 5741 6452 24340
rect 8332 20768 8372 20777
rect 8332 20273 8372 20728
rect 8524 20768 8564 20779
rect 8524 20693 8564 20728
rect 8523 20684 8565 20693
rect 8523 20644 8524 20684
rect 8564 20644 8565 20684
rect 8523 20635 8565 20644
rect 8043 20264 8085 20273
rect 8043 20224 8044 20264
rect 8084 20224 8085 20264
rect 8043 20215 8085 20224
rect 8331 20264 8373 20273
rect 8331 20224 8332 20264
rect 8372 20224 8373 20264
rect 8331 20215 8373 20224
rect 7851 20180 7893 20189
rect 7851 20140 7852 20180
rect 7892 20140 7893 20180
rect 7851 20131 7893 20140
rect 7852 20046 7892 20131
rect 8044 20096 8084 20215
rect 8044 20047 8084 20056
rect 8235 20096 8277 20105
rect 8235 20056 8236 20096
rect 8276 20056 8277 20096
rect 8235 20047 8277 20056
rect 8332 20096 8372 20105
rect 8524 20096 8564 20635
rect 8620 20273 8660 20358
rect 8619 20264 8661 20273
rect 8619 20224 8620 20264
rect 8660 20224 8661 20264
rect 8619 20215 8661 20224
rect 8716 20096 8756 29875
rect 19472 29504 19840 29513
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19472 29455 19840 29464
rect 34592 29504 34960 29513
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34592 29455 34960 29464
rect 49712 29504 50080 29513
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 49712 29455 50080 29464
rect 64832 29504 65200 29513
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 64832 29455 65200 29464
rect 79952 29504 80320 29513
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 79952 29455 80320 29464
rect 18232 28748 18600 28757
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18232 28699 18600 28708
rect 33352 28748 33720 28757
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33352 28699 33720 28708
rect 48472 28748 48840 28757
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48472 28699 48840 28708
rect 63592 28748 63960 28757
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63592 28699 63960 28708
rect 78712 28748 79080 28757
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 78712 28699 79080 28708
rect 19472 27992 19840 28001
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19472 27943 19840 27952
rect 34592 27992 34960 28001
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34592 27943 34960 27952
rect 49712 27992 50080 28001
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 49712 27943 50080 27952
rect 64832 27992 65200 28001
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 64832 27943 65200 27952
rect 79952 27992 80320 28001
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 79952 27943 80320 27952
rect 11404 27824 11444 27833
rect 11308 27656 11348 27665
rect 11116 27404 11156 27413
rect 10731 27152 10773 27161
rect 10731 27112 10732 27152
rect 10772 27112 10773 27152
rect 10731 27103 10773 27112
rect 10732 26816 10772 27103
rect 10828 26993 10868 27078
rect 10827 26984 10869 26993
rect 10827 26944 10828 26984
rect 10868 26944 10869 26984
rect 10827 26935 10869 26944
rect 10827 26816 10869 26825
rect 10732 26776 10828 26816
rect 10868 26776 10869 26816
rect 10827 26767 10869 26776
rect 10828 26682 10868 26767
rect 11019 26648 11061 26657
rect 11019 26608 11020 26648
rect 11060 26608 11061 26648
rect 11019 26599 11061 26608
rect 11020 26514 11060 26599
rect 11116 26144 11156 27364
rect 11308 26993 11348 27616
rect 11307 26984 11349 26993
rect 11307 26944 11308 26984
rect 11348 26944 11349 26984
rect 11307 26935 11349 26944
rect 11404 26825 11444 27784
rect 18232 27236 18600 27245
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18232 27187 18600 27196
rect 33352 27236 33720 27245
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33352 27187 33720 27196
rect 48472 27236 48840 27245
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48472 27187 48840 27196
rect 63592 27236 63960 27245
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63592 27187 63960 27196
rect 78712 27236 79080 27245
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 78712 27187 79080 27196
rect 12267 27068 12309 27077
rect 12267 27028 12268 27068
rect 12308 27028 12309 27068
rect 12267 27019 12309 27028
rect 11499 26984 11541 26993
rect 11499 26944 11500 26984
rect 11540 26944 11541 26984
rect 11499 26935 11541 26944
rect 11211 26816 11253 26825
rect 11211 26776 11212 26816
rect 11252 26776 11253 26816
rect 11211 26767 11253 26776
rect 11403 26816 11445 26825
rect 11403 26776 11404 26816
rect 11444 26776 11445 26816
rect 11403 26767 11445 26776
rect 11500 26816 11540 26935
rect 11500 26767 11540 26776
rect 11212 26682 11252 26767
rect 11403 26648 11445 26657
rect 11403 26608 11404 26648
rect 11444 26608 11445 26648
rect 11403 26599 11445 26608
rect 11692 26648 11732 26657
rect 11116 26095 11156 26104
rect 11307 26144 11349 26153
rect 11307 26104 11308 26144
rect 11348 26104 11349 26144
rect 11307 26095 11349 26104
rect 11404 26144 11444 26599
rect 11404 26095 11444 26104
rect 11308 26010 11348 26095
rect 9867 25892 9909 25901
rect 9867 25852 9868 25892
rect 9908 25852 9909 25892
rect 9867 25843 9909 25852
rect 11115 25892 11157 25901
rect 11115 25852 11116 25892
rect 11156 25852 11157 25892
rect 11115 25843 11157 25852
rect 9771 24716 9813 24725
rect 9771 24676 9772 24716
rect 9812 24676 9813 24716
rect 9771 24667 9813 24676
rect 9772 24582 9812 24667
rect 9868 24632 9908 25843
rect 11116 25758 11156 25843
rect 11692 25397 11732 26608
rect 11979 26144 12021 26153
rect 11979 26104 11980 26144
rect 12020 26104 12021 26144
rect 11979 26095 12021 26104
rect 11019 25388 11061 25397
rect 11019 25348 11020 25388
rect 11060 25348 11061 25388
rect 11019 25339 11061 25348
rect 11691 25388 11733 25397
rect 11691 25348 11692 25388
rect 11732 25348 11733 25388
rect 11691 25339 11733 25348
rect 9963 24800 10005 24809
rect 9963 24760 9964 24800
rect 10004 24760 10005 24800
rect 9963 24751 10005 24760
rect 10827 24800 10869 24809
rect 10827 24760 10828 24800
rect 10868 24760 10869 24800
rect 10827 24751 10869 24760
rect 9868 24583 9908 24592
rect 9964 24632 10004 24751
rect 10828 24666 10868 24751
rect 9964 24583 10004 24592
rect 10060 24632 10100 24641
rect 10060 22289 10100 24592
rect 11020 24632 11060 25339
rect 11020 24583 11060 24592
rect 11116 24632 11156 24641
rect 11116 23960 11156 24592
rect 11980 24632 12020 26095
rect 12075 25304 12117 25313
rect 12075 25264 12076 25304
rect 12116 25264 12117 25304
rect 12075 25255 12117 25264
rect 12076 24800 12116 25255
rect 12076 24751 12116 24760
rect 11404 24053 11444 24138
rect 11403 24044 11445 24053
rect 11403 24004 11404 24044
rect 11444 24004 11445 24044
rect 11403 23995 11445 24004
rect 11116 23920 11348 23960
rect 11212 23792 11252 23801
rect 11308 23792 11348 23920
rect 11404 23792 11444 23801
rect 11308 23752 11404 23792
rect 11212 22289 11252 23752
rect 11307 22364 11349 22373
rect 11404 22364 11444 23752
rect 11980 23288 12020 24592
rect 12172 24632 12212 24641
rect 12172 24053 12212 24592
rect 12171 24044 12213 24053
rect 12171 24004 12172 24044
rect 12212 24004 12213 24044
rect 12171 23995 12213 24004
rect 12076 23288 12116 23297
rect 11980 23248 12076 23288
rect 12076 23239 12116 23248
rect 12268 23120 12308 27019
rect 19472 26480 19840 26489
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19472 26431 19840 26440
rect 34592 26480 34960 26489
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34592 26431 34960 26440
rect 49712 26480 50080 26489
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 49712 26431 50080 26440
rect 64832 26480 65200 26489
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 64832 26431 65200 26440
rect 79952 26480 80320 26489
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 79952 26431 80320 26440
rect 18232 25724 18600 25733
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18232 25675 18600 25684
rect 33352 25724 33720 25733
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33352 25675 33720 25684
rect 48472 25724 48840 25733
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48472 25675 48840 25684
rect 63592 25724 63960 25733
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63592 25675 63960 25684
rect 78712 25724 79080 25733
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 78712 25675 79080 25684
rect 12364 25388 12404 25397
rect 12364 25229 12404 25348
rect 12651 25388 12693 25397
rect 12651 25348 12652 25388
rect 12692 25348 12693 25388
rect 12651 25339 12693 25348
rect 12555 25304 12597 25313
rect 12555 25264 12556 25304
rect 12596 25264 12597 25304
rect 12555 25255 12597 25264
rect 12652 25304 12692 25339
rect 12363 25220 12405 25229
rect 12363 25180 12364 25220
rect 12404 25180 12405 25220
rect 12363 25171 12405 25180
rect 12556 25170 12596 25255
rect 12652 25253 12692 25264
rect 19472 24968 19840 24977
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19472 24919 19840 24928
rect 34592 24968 34960 24977
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34592 24919 34960 24928
rect 49712 24968 50080 24977
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 49712 24919 50080 24928
rect 64832 24968 65200 24977
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 64832 24919 65200 24928
rect 79952 24968 80320 24977
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 79952 24919 80320 24928
rect 12363 24380 12405 24389
rect 12363 24340 12364 24380
rect 12404 24340 12405 24380
rect 12363 24331 12405 24340
rect 12076 23080 12268 23120
rect 11307 22324 11308 22364
rect 11348 22324 11444 22364
rect 11883 22364 11925 22373
rect 11883 22324 11884 22364
rect 11924 22324 11925 22364
rect 11307 22315 11349 22324
rect 11883 22315 11925 22324
rect 8811 22280 8853 22289
rect 8811 22240 8812 22280
rect 8852 22240 8853 22280
rect 8811 22231 8853 22240
rect 10059 22280 10101 22289
rect 10059 22240 10060 22280
rect 10100 22240 10101 22280
rect 10059 22231 10101 22240
rect 11211 22280 11253 22289
rect 11211 22240 11212 22280
rect 11252 22240 11253 22280
rect 11211 22231 11253 22240
rect 11308 22280 11348 22315
rect 8812 20936 8852 22231
rect 11308 22229 11348 22240
rect 11595 22280 11637 22289
rect 11595 22240 11596 22280
rect 11636 22240 11637 22280
rect 11595 22231 11637 22240
rect 11596 22146 11636 22231
rect 11884 22230 11924 22315
rect 12076 22280 12116 23080
rect 12268 23071 12308 23080
rect 12364 23288 12404 24331
rect 18232 24212 18600 24221
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18232 24163 18600 24172
rect 33352 24212 33720 24221
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33352 24163 33720 24172
rect 48472 24212 48840 24221
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48472 24163 48840 24172
rect 63592 24212 63960 24221
rect 63632 24172 63674 24212
rect 63714 24172 63756 24212
rect 63796 24172 63838 24212
rect 63878 24172 63920 24212
rect 63592 24163 63960 24172
rect 78712 24212 79080 24221
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 78712 24163 79080 24172
rect 19472 23456 19840 23465
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19472 23407 19840 23416
rect 34592 23456 34960 23465
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34592 23407 34960 23416
rect 49712 23456 50080 23465
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 49712 23407 50080 23416
rect 64832 23456 65200 23465
rect 64872 23416 64914 23456
rect 64954 23416 64996 23456
rect 65036 23416 65078 23456
rect 65118 23416 65160 23456
rect 64832 23407 65200 23416
rect 79952 23456 80320 23465
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 79952 23407 80320 23416
rect 12076 22231 12116 22240
rect 12172 22280 12212 22289
rect 12364 22280 12404 23248
rect 18232 22700 18600 22709
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18232 22651 18600 22660
rect 33352 22700 33720 22709
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33352 22651 33720 22660
rect 48472 22700 48840 22709
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48472 22651 48840 22660
rect 63592 22700 63960 22709
rect 63632 22660 63674 22700
rect 63714 22660 63756 22700
rect 63796 22660 63838 22700
rect 63878 22660 63920 22700
rect 63592 22651 63960 22660
rect 78712 22700 79080 22709
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 78712 22651 79080 22660
rect 12212 22240 12404 22280
rect 12172 22231 12212 22240
rect 11115 22112 11157 22121
rect 11115 22072 11116 22112
rect 11156 22072 11157 22112
rect 11115 22063 11157 22072
rect 11116 21978 11156 22063
rect 19472 21944 19840 21953
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19472 21895 19840 21904
rect 34592 21944 34960 21953
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34592 21895 34960 21904
rect 49712 21944 50080 21953
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 49712 21895 50080 21904
rect 64832 21944 65200 21953
rect 64872 21904 64914 21944
rect 64954 21904 64996 21944
rect 65036 21904 65078 21944
rect 65118 21904 65160 21944
rect 64832 21895 65200 21904
rect 79952 21944 80320 21953
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 79952 21895 80320 21904
rect 18232 21188 18600 21197
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18232 21139 18600 21148
rect 33352 21188 33720 21197
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33352 21139 33720 21148
rect 48472 21188 48840 21197
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48472 21139 48840 21148
rect 63592 21188 63960 21197
rect 63632 21148 63674 21188
rect 63714 21148 63756 21188
rect 63796 21148 63838 21188
rect 63878 21148 63920 21188
rect 63592 21139 63960 21148
rect 78712 21188 79080 21197
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 78712 21139 79080 21148
rect 8812 20887 8852 20896
rect 8908 20768 8948 20777
rect 8908 20189 8948 20728
rect 19472 20432 19840 20441
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19472 20383 19840 20392
rect 34592 20432 34960 20441
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34592 20383 34960 20392
rect 49712 20432 50080 20441
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 49712 20383 50080 20392
rect 64832 20432 65200 20441
rect 64872 20392 64914 20432
rect 64954 20392 64996 20432
rect 65036 20392 65078 20432
rect 65118 20392 65160 20432
rect 64832 20383 65200 20392
rect 79952 20432 80320 20441
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 79952 20383 80320 20392
rect 8907 20180 8949 20189
rect 8907 20140 8908 20180
rect 8948 20140 8949 20180
rect 8907 20131 8949 20140
rect 8372 20056 8564 20096
rect 8620 20056 8716 20096
rect 8332 20047 8372 20056
rect 8236 19508 8276 20047
rect 8332 19508 8372 19517
rect 8236 19468 8332 19508
rect 8332 19459 8372 19468
rect 8140 19256 8180 19265
rect 8620 19256 8660 20056
rect 8716 20047 8756 20056
rect 9100 20096 9140 20105
rect 8180 19216 8660 19256
rect 8140 19207 8180 19216
rect 9100 19097 9140 20056
rect 18232 19676 18600 19685
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18232 19627 18600 19636
rect 33352 19676 33720 19685
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33352 19627 33720 19636
rect 48472 19676 48840 19685
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48472 19627 48840 19636
rect 63592 19676 63960 19685
rect 63632 19636 63674 19676
rect 63714 19636 63756 19676
rect 63796 19636 63838 19676
rect 63878 19636 63920 19676
rect 63592 19627 63960 19636
rect 78712 19676 79080 19685
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 78712 19627 79080 19636
rect 8043 19088 8085 19097
rect 8043 19048 8044 19088
rect 8084 19048 8085 19088
rect 8043 19039 8085 19048
rect 9099 19088 9141 19097
rect 9099 19048 9100 19088
rect 9140 19048 9141 19088
rect 9099 19039 9141 19048
rect 8044 18954 8084 19039
rect 19472 18920 19840 18929
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19472 18871 19840 18880
rect 34592 18920 34960 18929
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34592 18871 34960 18880
rect 49712 18920 50080 18929
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 49712 18871 50080 18880
rect 64832 18920 65200 18929
rect 64872 18880 64914 18920
rect 64954 18880 64996 18920
rect 65036 18880 65078 18920
rect 65118 18880 65160 18920
rect 64832 18871 65200 18880
rect 79952 18920 80320 18929
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 79952 18871 80320 18880
rect 18232 18164 18600 18173
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18232 18115 18600 18124
rect 33352 18164 33720 18173
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33352 18115 33720 18124
rect 48472 18164 48840 18173
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48472 18115 48840 18124
rect 63592 18164 63960 18173
rect 63632 18124 63674 18164
rect 63714 18124 63756 18164
rect 63796 18124 63838 18164
rect 63878 18124 63920 18164
rect 63592 18115 63960 18124
rect 78712 18164 79080 18173
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 78712 18115 79080 18124
rect 19472 17408 19840 17417
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19472 17359 19840 17368
rect 34592 17408 34960 17417
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34592 17359 34960 17368
rect 49712 17408 50080 17417
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 49712 17359 50080 17368
rect 64832 17408 65200 17417
rect 64872 17368 64914 17408
rect 64954 17368 64996 17408
rect 65036 17368 65078 17408
rect 65118 17368 65160 17408
rect 64832 17359 65200 17368
rect 79952 17408 80320 17417
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 79952 17359 80320 17368
rect 18232 16652 18600 16661
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18232 16603 18600 16612
rect 33352 16652 33720 16661
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33352 16603 33720 16612
rect 48472 16652 48840 16661
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48472 16603 48840 16612
rect 63592 16652 63960 16661
rect 63632 16612 63674 16652
rect 63714 16612 63756 16652
rect 63796 16612 63838 16652
rect 63878 16612 63920 16652
rect 63592 16603 63960 16612
rect 78712 16652 79080 16661
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 78712 16603 79080 16612
rect 19472 15896 19840 15905
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19472 15847 19840 15856
rect 34592 15896 34960 15905
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34592 15847 34960 15856
rect 49712 15896 50080 15905
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 49712 15847 50080 15856
rect 64832 15896 65200 15905
rect 64872 15856 64914 15896
rect 64954 15856 64996 15896
rect 65036 15856 65078 15896
rect 65118 15856 65160 15896
rect 64832 15847 65200 15856
rect 79952 15896 80320 15905
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 79952 15847 80320 15856
rect 18232 15140 18600 15149
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18232 15091 18600 15100
rect 33352 15140 33720 15149
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 33352 15091 33720 15100
rect 48472 15140 48840 15149
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48472 15091 48840 15100
rect 63592 15140 63960 15149
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63592 15091 63960 15100
rect 78712 15140 79080 15149
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 78712 15091 79080 15100
rect 19472 14384 19840 14393
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19472 14335 19840 14344
rect 34592 14384 34960 14393
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34592 14335 34960 14344
rect 49712 14384 50080 14393
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 49712 14335 50080 14344
rect 64832 14384 65200 14393
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 64832 14335 65200 14344
rect 79952 14384 80320 14393
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 79952 14335 80320 14344
rect 18232 13628 18600 13637
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18232 13579 18600 13588
rect 33352 13628 33720 13637
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33352 13579 33720 13588
rect 48472 13628 48840 13637
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48472 13579 48840 13588
rect 63592 13628 63960 13637
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63592 13579 63960 13588
rect 78712 13628 79080 13637
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 78712 13579 79080 13588
rect 19472 12872 19840 12881
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19472 12823 19840 12832
rect 34592 12872 34960 12881
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34592 12823 34960 12832
rect 49712 12872 50080 12881
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 49712 12823 50080 12832
rect 64832 12872 65200 12881
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 64832 12823 65200 12832
rect 79952 12872 80320 12881
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 79952 12823 80320 12832
rect 18232 12116 18600 12125
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18232 12067 18600 12076
rect 33352 12116 33720 12125
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33352 12067 33720 12076
rect 48472 12116 48840 12125
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48472 12067 48840 12076
rect 63592 12116 63960 12125
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63592 12067 63960 12076
rect 78712 12116 79080 12125
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 78712 12067 79080 12076
rect 19472 11360 19840 11369
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19472 11311 19840 11320
rect 34592 11360 34960 11369
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34592 11311 34960 11320
rect 49712 11360 50080 11369
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 49712 11311 50080 11320
rect 64832 11360 65200 11369
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 64832 11311 65200 11320
rect 79952 11360 80320 11369
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 79952 11311 80320 11320
rect 18232 10604 18600 10613
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18232 10555 18600 10564
rect 33352 10604 33720 10613
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33352 10555 33720 10564
rect 48472 10604 48840 10613
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48472 10555 48840 10564
rect 63592 10604 63960 10613
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63592 10555 63960 10564
rect 78712 10604 79080 10613
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 78712 10555 79080 10564
rect 19472 9848 19840 9857
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19472 9799 19840 9808
rect 34592 9848 34960 9857
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34592 9799 34960 9808
rect 49712 9848 50080 9857
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 49712 9799 50080 9808
rect 64832 9848 65200 9857
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 64832 9799 65200 9808
rect 79952 9848 80320 9857
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 79952 9799 80320 9808
rect 18232 9092 18600 9101
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18232 9043 18600 9052
rect 33352 9092 33720 9101
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33352 9043 33720 9052
rect 48472 9092 48840 9101
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48472 9043 48840 9052
rect 63592 9092 63960 9101
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63592 9043 63960 9052
rect 78712 9092 79080 9101
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 78712 9043 79080 9052
rect 19472 8336 19840 8345
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19472 8287 19840 8296
rect 34592 8336 34960 8345
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34592 8287 34960 8296
rect 49712 8336 50080 8345
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 49712 8287 50080 8296
rect 64832 8336 65200 8345
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 64832 8287 65200 8296
rect 79952 8336 80320 8345
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 79952 8287 80320 8296
rect 18232 7580 18600 7589
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18232 7531 18600 7540
rect 33352 7580 33720 7589
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33352 7531 33720 7540
rect 48472 7580 48840 7589
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48472 7531 48840 7540
rect 63592 7580 63960 7589
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63592 7531 63960 7540
rect 78712 7580 79080 7589
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 78712 7531 79080 7540
rect 19472 6824 19840 6833
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19472 6775 19840 6784
rect 34592 6824 34960 6833
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34592 6775 34960 6784
rect 49712 6824 50080 6833
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 49712 6775 50080 6784
rect 64832 6824 65200 6833
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 64832 6775 65200 6784
rect 79952 6824 80320 6833
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 79952 6775 80320 6784
rect 18232 6068 18600 6077
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18232 6019 18600 6028
rect 33352 6068 33720 6077
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33352 6019 33720 6028
rect 48472 6068 48840 6077
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48472 6019 48840 6028
rect 63592 6068 63960 6077
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63592 6019 63960 6028
rect 78712 6068 79080 6077
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 78712 6019 79080 6028
rect 6411 5732 6453 5741
rect 6411 5692 6412 5732
rect 6452 5692 6453 5732
rect 6411 5683 6453 5692
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 19472 5312 19840 5321
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19472 5263 19840 5272
rect 34592 5312 34960 5321
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34592 5263 34960 5272
rect 49712 5312 50080 5321
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 49712 5263 50080 5272
rect 64832 5312 65200 5321
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 64832 5263 65200 5272
rect 79952 5312 80320 5321
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 79952 5263 80320 5272
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 18232 4556 18600 4565
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18232 4507 18600 4516
rect 33352 4556 33720 4565
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33352 4507 33720 4516
rect 48472 4556 48840 4565
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48472 4507 48840 4516
rect 63592 4556 63960 4565
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63592 4507 63960 4516
rect 78712 4556 79080 4565
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 78712 4507 79080 4516
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 19472 3800 19840 3809
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19472 3751 19840 3760
rect 34592 3800 34960 3809
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34592 3751 34960 3760
rect 49712 3800 50080 3809
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 49712 3751 50080 3760
rect 64832 3800 65200 3809
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 64832 3751 65200 3760
rect 79952 3800 80320 3809
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 79952 3751 80320 3760
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 18232 3044 18600 3053
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18232 2995 18600 3004
rect 33352 3044 33720 3053
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33352 2995 33720 3004
rect 48472 3044 48840 3053
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48472 2995 48840 3004
rect 63592 3044 63960 3053
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63592 2995 63960 3004
rect 78712 3044 79080 3053
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 78712 2995 79080 3004
rect 884 2668 1268 2708
rect 844 2659 884 2668
rect 652 2456 692 2465
rect 652 2297 692 2416
rect 651 2288 693 2297
rect 651 2248 652 2288
rect 692 2248 693 2288
rect 651 2239 693 2248
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 19472 2288 19840 2297
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19472 2239 19840 2248
rect 34592 2288 34960 2297
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34592 2239 34960 2248
rect 49712 2288 50080 2297
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 49712 2239 50080 2248
rect 64832 2288 65200 2297
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 64832 2239 65200 2248
rect 79952 2288 80320 2297
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 79952 2239 80320 2248
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 18232 1532 18600 1541
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18232 1483 18600 1492
rect 33352 1532 33720 1541
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33352 1483 33720 1492
rect 48472 1532 48840 1541
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48472 1483 48840 1492
rect 63592 1532 63960 1541
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63592 1483 63960 1492
rect 78712 1532 79080 1541
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 78712 1483 79080 1492
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
rect 19472 776 19840 785
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19472 727 19840 736
rect 34592 776 34960 785
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34592 727 34960 736
rect 49712 776 50080 785
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 49712 727 50080 736
rect 64832 776 65200 785
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 64832 727 65200 736
rect 79952 776 80320 785
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 79952 727 80320 736
<< via2 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 652 35092 692 35132
rect 652 34168 692 34208
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 748 33580 788 33620
rect 652 33328 692 33368
rect 364 31480 404 31520
rect 652 32488 692 32528
rect 556 31900 596 31940
rect 652 31648 692 31688
rect 652 30808 692 30848
rect 652 30052 692 30092
rect 844 31900 884 31940
rect 844 29884 884 29924
rect 844 29632 884 29672
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 4396 33580 4436 33620
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 3820 32152 3860 32192
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 1036 30640 1076 30680
rect 2572 30640 2612 30680
rect 2284 29800 2324 29840
rect 2860 30640 2900 30680
rect 3052 30640 3092 30680
rect 3244 30640 3284 30680
rect 2668 30556 2708 30596
rect 3148 30472 3188 30512
rect 2860 30388 2900 30428
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 3724 30472 3764 30512
rect 3628 30388 3668 30428
rect 2668 29800 2708 29840
rect 1228 29632 1268 29672
rect 2092 29632 2132 29672
rect 748 29296 788 29336
rect 652 29128 692 29168
rect 652 28372 692 28412
rect 844 28960 884 29000
rect 652 27532 692 27572
rect 556 26944 596 26984
rect 460 26860 500 26900
rect 460 25180 500 25220
rect 364 20056 404 20096
rect 1132 27112 1172 27152
rect 1036 27028 1076 27068
rect 844 26776 884 26816
rect 652 26608 692 26648
rect 652 25768 692 25808
rect 652 24928 692 24968
rect 652 24088 692 24128
rect 844 25516 884 25556
rect 844 24340 884 24380
rect 1132 25516 1172 25556
rect 1132 24088 1172 24128
rect 1036 23836 1076 23876
rect 748 23752 788 23792
rect 652 23248 692 23288
rect 652 22408 692 22448
rect 652 21568 692 21608
rect 652 20728 692 20768
rect 844 20728 884 20768
rect 652 19888 692 19928
rect 1036 22072 1076 22112
rect 652 19048 692 19088
rect 940 19048 980 19088
rect 652 18208 692 18248
rect 652 17368 692 17408
rect 652 16528 692 16568
rect 460 15772 500 15812
rect 556 15688 596 15728
rect 652 14848 692 14888
rect 652 14008 692 14048
rect 652 13168 692 13208
rect 652 12328 692 12368
rect 652 11488 692 11528
rect 940 15772 980 15812
rect 652 10648 692 10688
rect 652 9808 692 9848
rect 652 8968 692 9008
rect 652 8128 692 8168
rect 844 7876 884 7916
rect 652 7288 692 7328
rect 844 7204 884 7244
rect 652 6448 692 6488
rect 652 5608 692 5648
rect 652 4768 692 4808
rect 652 3928 692 3968
rect 844 5692 884 5732
rect 1900 24004 1940 24044
rect 1804 23836 1844 23876
rect 1996 23752 2036 23792
rect 1228 20812 1268 20852
rect 1228 19804 1268 19844
rect 1132 7204 1172 7244
rect 652 3172 692 3212
rect 3340 29800 3380 29840
rect 3532 29800 3572 29840
rect 3820 29800 3860 29840
rect 3052 29632 3092 29672
rect 2284 29296 2324 29336
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 4396 32152 4436 32192
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 4204 31480 4244 31520
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 8716 29884 8756 29924
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 4108 28960 4148 29000
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 3628 26860 3668 26900
rect 4305 26860 4345 26900
rect 4780 26860 4820 26900
rect 3436 26776 3476 26816
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 3916 26776 3956 26816
rect 5260 26776 5300 26816
rect 4204 26692 4244 26732
rect 4876 26692 4916 26732
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 5164 26104 5204 26144
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 5548 26104 5588 26144
rect 4780 24676 4820 24716
rect 5356 24676 5396 24716
rect 4012 24508 4052 24548
rect 3532 24004 3572 24044
rect 4204 24592 4244 24632
rect 4300 24004 4340 24044
rect 2476 23836 2516 23876
rect 2188 23752 2228 23792
rect 5452 24592 5492 24632
rect 6604 24676 6644 24716
rect 6508 24592 6548 24632
rect 6604 24508 6644 24548
rect 5356 24088 5396 24128
rect 2668 23668 2708 23708
rect 4300 23668 4340 23708
rect 4684 23668 4724 23708
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 3436 20812 3476 20852
rect 4108 20812 4148 20852
rect 3820 20728 3860 20768
rect 4012 20728 4052 20768
rect 4300 20644 4340 20684
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 3340 19804 3380 19844
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 2092 7876 2132 7916
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 8524 20644 8564 20684
rect 8044 20224 8084 20264
rect 8332 20224 8372 20264
rect 7852 20140 7892 20180
rect 8236 20056 8276 20096
rect 8620 20224 8660 20264
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 10732 27112 10772 27152
rect 10828 26944 10868 26984
rect 10828 26776 10868 26816
rect 11020 26608 11060 26648
rect 11308 26944 11348 26984
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 12268 27028 12308 27068
rect 11500 26944 11540 26984
rect 11212 26776 11252 26816
rect 11404 26776 11444 26816
rect 11404 26608 11444 26648
rect 11308 26104 11348 26144
rect 9868 25852 9908 25892
rect 11116 25852 11156 25892
rect 9772 24676 9812 24716
rect 11980 26104 12020 26144
rect 11020 25348 11060 25388
rect 11692 25348 11732 25388
rect 9964 24760 10004 24800
rect 10828 24760 10868 24800
rect 12076 25264 12116 25304
rect 11404 24004 11444 24044
rect 12172 24004 12212 24044
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 12652 25348 12692 25388
rect 12556 25264 12596 25304
rect 12364 25180 12404 25220
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 12364 24340 12404 24380
rect 11308 22324 11348 22364
rect 11884 22324 11924 22364
rect 8812 22240 8852 22280
rect 10060 22240 10100 22280
rect 11212 22240 11252 22280
rect 11596 22240 11636 22280
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 63592 24172 63632 24212
rect 63674 24172 63714 24212
rect 63756 24172 63796 24212
rect 63838 24172 63878 24212
rect 63920 24172 63960 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 64832 23416 64872 23456
rect 64914 23416 64954 23456
rect 64996 23416 65036 23456
rect 65078 23416 65118 23456
rect 65160 23416 65200 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 63592 22660 63632 22700
rect 63674 22660 63714 22700
rect 63756 22660 63796 22700
rect 63838 22660 63878 22700
rect 63920 22660 63960 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 11116 22072 11156 22112
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 64832 21904 64872 21944
rect 64914 21904 64954 21944
rect 64996 21904 65036 21944
rect 65078 21904 65118 21944
rect 65160 21904 65200 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 63592 21148 63632 21188
rect 63674 21148 63714 21188
rect 63756 21148 63796 21188
rect 63838 21148 63878 21188
rect 63920 21148 63960 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 64832 20392 64872 20432
rect 64914 20392 64954 20432
rect 64996 20392 65036 20432
rect 65078 20392 65118 20432
rect 65160 20392 65200 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 8908 20140 8948 20180
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 63592 19636 63632 19676
rect 63674 19636 63714 19676
rect 63756 19636 63796 19676
rect 63838 19636 63878 19676
rect 63920 19636 63960 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 8044 19048 8084 19088
rect 9100 19048 9140 19088
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 64832 18880 64872 18920
rect 64914 18880 64954 18920
rect 64996 18880 65036 18920
rect 65078 18880 65118 18920
rect 65160 18880 65200 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 63592 18124 63632 18164
rect 63674 18124 63714 18164
rect 63756 18124 63796 18164
rect 63838 18124 63878 18164
rect 63920 18124 63960 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 64832 17368 64872 17408
rect 64914 17368 64954 17408
rect 64996 17368 65036 17408
rect 65078 17368 65118 17408
rect 65160 17368 65200 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 63592 16612 63632 16652
rect 63674 16612 63714 16652
rect 63756 16612 63796 16652
rect 63838 16612 63878 16652
rect 63920 16612 63960 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 64832 15856 64872 15896
rect 64914 15856 64954 15896
rect 64996 15856 65036 15896
rect 65078 15856 65118 15896
rect 65160 15856 65200 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 6412 5692 6452 5732
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 652 2248 692 2288
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
<< metal3 >>
rect 4343 38536 4352 38576
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4720 38536 4729 38576
rect 19463 38536 19472 38576
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19840 38536 19849 38576
rect 34583 38536 34592 38576
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34960 38536 34969 38576
rect 49703 38536 49712 38576
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 50080 38536 50089 38576
rect 64823 38536 64832 38576
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 65200 38536 65209 38576
rect 79943 38536 79952 38576
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 80320 38536 80329 38576
rect 3103 37780 3112 37820
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3480 37780 3489 37820
rect 18223 37780 18232 37820
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18600 37780 18609 37820
rect 33343 37780 33352 37820
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33720 37780 33729 37820
rect 48463 37780 48472 37820
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48840 37780 48849 37820
rect 63583 37780 63592 37820
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63960 37780 63969 37820
rect 78703 37780 78712 37820
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 79080 37780 79089 37820
rect 0 37508 80 37588
rect 4343 37024 4352 37064
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4720 37024 4729 37064
rect 19463 37024 19472 37064
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19840 37024 19849 37064
rect 34583 37024 34592 37064
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34960 37024 34969 37064
rect 49703 37024 49712 37064
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 50080 37024 50089 37064
rect 64823 37024 64832 37064
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 65200 37024 65209 37064
rect 79943 37024 79952 37064
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 80320 37024 80329 37064
rect 0 36668 80 36748
rect 3103 36268 3112 36308
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3480 36268 3489 36308
rect 18223 36268 18232 36308
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18600 36268 18609 36308
rect 33343 36268 33352 36308
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33720 36268 33729 36308
rect 48463 36268 48472 36308
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48840 36268 48849 36308
rect 63583 36268 63592 36308
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63960 36268 63969 36308
rect 78703 36268 78712 36308
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 79080 36268 79089 36308
rect 0 35828 80 35908
rect 4343 35512 4352 35552
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4720 35512 4729 35552
rect 19463 35512 19472 35552
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19840 35512 19849 35552
rect 34583 35512 34592 35552
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34960 35512 34969 35552
rect 49703 35512 49712 35552
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 50080 35512 50089 35552
rect 64823 35512 64832 35552
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 65200 35512 65209 35552
rect 79943 35512 79952 35552
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 80320 35512 80329 35552
rect 643 35092 652 35132
rect 692 35092 701 35132
rect 0 35048 80 35068
rect 652 35048 692 35092
rect 0 35008 692 35048
rect 0 34988 80 35008
rect 3103 34756 3112 34796
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3480 34756 3489 34796
rect 18223 34756 18232 34796
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18600 34756 18609 34796
rect 33343 34756 33352 34796
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33720 34756 33729 34796
rect 48463 34756 48472 34796
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48840 34756 48849 34796
rect 63583 34756 63592 34796
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63960 34756 63969 34796
rect 78703 34756 78712 34796
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 79080 34756 79089 34796
rect 0 34208 80 34228
rect 0 34168 652 34208
rect 692 34168 701 34208
rect 0 34148 80 34168
rect 4343 34000 4352 34040
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4720 34000 4729 34040
rect 19463 34000 19472 34040
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19840 34000 19849 34040
rect 34583 34000 34592 34040
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34960 34000 34969 34040
rect 49703 34000 49712 34040
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 50080 34000 50089 34040
rect 64823 34000 64832 34040
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 65200 34000 65209 34040
rect 79943 34000 79952 34040
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 80320 34000 80329 34040
rect 739 33580 748 33620
rect 788 33580 4396 33620
rect 4436 33580 4445 33620
rect 0 33368 80 33388
rect 0 33328 652 33368
rect 692 33328 701 33368
rect 0 33308 80 33328
rect 3103 33244 3112 33284
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3480 33244 3489 33284
rect 18223 33244 18232 33284
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18600 33244 18609 33284
rect 33343 33244 33352 33284
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33720 33244 33729 33284
rect 48463 33244 48472 33284
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48840 33244 48849 33284
rect 63583 33244 63592 33284
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63960 33244 63969 33284
rect 78703 33244 78712 33284
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 79080 33244 79089 33284
rect 0 32528 80 32548
rect 0 32488 652 32528
rect 692 32488 701 32528
rect 4343 32488 4352 32528
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4720 32488 4729 32528
rect 19463 32488 19472 32528
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19840 32488 19849 32528
rect 34583 32488 34592 32528
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34960 32488 34969 32528
rect 49703 32488 49712 32528
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 50080 32488 50089 32528
rect 64823 32488 64832 32528
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 65200 32488 65209 32528
rect 79943 32488 79952 32528
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 80320 32488 80329 32528
rect 0 32468 80 32488
rect 3811 32152 3820 32192
rect 3860 32152 4396 32192
rect 4436 32152 4445 32192
rect 547 31900 556 31940
rect 596 31900 844 31940
rect 884 31900 893 31940
rect 3103 31732 3112 31772
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3480 31732 3489 31772
rect 18223 31732 18232 31772
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18600 31732 18609 31772
rect 33343 31732 33352 31772
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33720 31732 33729 31772
rect 48463 31732 48472 31772
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48840 31732 48849 31772
rect 63583 31732 63592 31772
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63960 31732 63969 31772
rect 78703 31732 78712 31772
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 79080 31732 79089 31772
rect 0 31688 80 31708
rect 0 31648 652 31688
rect 692 31648 701 31688
rect 0 31628 80 31648
rect 355 31480 364 31520
rect 404 31480 4204 31520
rect 4244 31480 4253 31520
rect 4343 30976 4352 31016
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4720 30976 4729 31016
rect 19463 30976 19472 31016
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19840 30976 19849 31016
rect 34583 30976 34592 31016
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34960 30976 34969 31016
rect 49703 30976 49712 31016
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 50080 30976 50089 31016
rect 64823 30976 64832 31016
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 65200 30976 65209 31016
rect 79943 30976 79952 31016
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 80320 30976 80329 31016
rect 0 30848 80 30868
rect 0 30808 652 30848
rect 692 30808 701 30848
rect 0 30788 80 30808
rect 1027 30640 1036 30680
rect 1076 30640 2572 30680
rect 2612 30640 2860 30680
rect 2900 30640 3052 30680
rect 3092 30640 3101 30680
rect 3235 30640 3244 30680
rect 3284 30640 3293 30680
rect 3244 30596 3284 30640
rect 2659 30556 2668 30596
rect 2708 30556 3284 30596
rect 3139 30472 3148 30512
rect 3188 30472 3724 30512
rect 3764 30472 3773 30512
rect 2851 30388 2860 30428
rect 2900 30388 3628 30428
rect 3668 30388 3677 30428
rect 3103 30220 3112 30260
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3480 30220 3489 30260
rect 18223 30220 18232 30260
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18600 30220 18609 30260
rect 33343 30220 33352 30260
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33720 30220 33729 30260
rect 48463 30220 48472 30260
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48840 30220 48849 30260
rect 63583 30220 63592 30260
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63960 30220 63969 30260
rect 78703 30220 78712 30260
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 79080 30220 79089 30260
rect 643 30052 652 30092
rect 692 30052 701 30092
rect 0 30008 80 30028
rect 652 30008 692 30052
rect 0 29968 692 30008
rect 0 29948 80 29968
rect 835 29884 844 29924
rect 884 29884 8716 29924
rect 8756 29884 8765 29924
rect 2275 29800 2284 29840
rect 2324 29800 2668 29840
rect 2708 29800 2717 29840
rect 3331 29800 3340 29840
rect 3380 29800 3532 29840
rect 3572 29800 3820 29840
rect 3860 29800 3869 29840
rect 835 29632 844 29672
rect 884 29632 1228 29672
rect 1268 29632 1277 29672
rect 2083 29632 2092 29672
rect 2132 29632 3052 29672
rect 3092 29632 3101 29672
rect 4343 29464 4352 29504
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4720 29464 4729 29504
rect 19463 29464 19472 29504
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19840 29464 19849 29504
rect 34583 29464 34592 29504
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34960 29464 34969 29504
rect 49703 29464 49712 29504
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 50080 29464 50089 29504
rect 64823 29464 64832 29504
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 65200 29464 65209 29504
rect 79943 29464 79952 29504
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 80320 29464 80329 29504
rect 739 29296 748 29336
rect 788 29296 2284 29336
rect 2324 29296 2333 29336
rect 0 29168 80 29188
rect 0 29128 652 29168
rect 692 29128 701 29168
rect 0 29108 80 29128
rect 835 28960 844 29000
rect 884 28960 4108 29000
rect 4148 28960 4157 29000
rect 3103 28708 3112 28748
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3480 28708 3489 28748
rect 18223 28708 18232 28748
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18600 28708 18609 28748
rect 33343 28708 33352 28748
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33720 28708 33729 28748
rect 48463 28708 48472 28748
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48840 28708 48849 28748
rect 63583 28708 63592 28748
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63960 28708 63969 28748
rect 78703 28708 78712 28748
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 79080 28708 79089 28748
rect 643 28372 652 28412
rect 692 28372 701 28412
rect 0 28328 80 28348
rect 652 28328 692 28372
rect 0 28288 692 28328
rect 0 28268 80 28288
rect 4343 27952 4352 27992
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4720 27952 4729 27992
rect 19463 27952 19472 27992
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19840 27952 19849 27992
rect 34583 27952 34592 27992
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34960 27952 34969 27992
rect 49703 27952 49712 27992
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 50080 27952 50089 27992
rect 64823 27952 64832 27992
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 65200 27952 65209 27992
rect 79943 27952 79952 27992
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 80320 27952 80329 27992
rect 643 27532 652 27572
rect 692 27532 701 27572
rect 0 27488 80 27508
rect 652 27488 692 27532
rect 0 27448 692 27488
rect 0 27428 80 27448
rect 3103 27196 3112 27236
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3480 27196 3489 27236
rect 18223 27196 18232 27236
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18600 27196 18609 27236
rect 33343 27196 33352 27236
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33720 27196 33729 27236
rect 48463 27196 48472 27236
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48840 27196 48849 27236
rect 63583 27196 63592 27236
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63960 27196 63969 27236
rect 78703 27196 78712 27236
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 79080 27196 79089 27236
rect 1123 27112 1132 27152
rect 1172 27112 10732 27152
rect 10772 27112 10781 27152
rect 1027 27028 1036 27068
rect 1076 27028 12268 27068
rect 12308 27028 12317 27068
rect 547 26944 556 26984
rect 596 26944 10828 26984
rect 10868 26944 11308 26984
rect 11348 26944 11500 26984
rect 11540 26944 11549 26984
rect 451 26860 460 26900
rect 500 26860 3628 26900
rect 3668 26860 4305 26900
rect 4345 26860 4780 26900
rect 4820 26860 4829 26900
rect 835 26776 844 26816
rect 884 26776 3436 26816
rect 3476 26776 3485 26816
rect 3907 26776 3916 26816
rect 3956 26776 5260 26816
rect 5300 26776 5309 26816
rect 10819 26776 10828 26816
rect 10868 26776 11212 26816
rect 11252 26776 11404 26816
rect 11444 26776 11453 26816
rect 3436 26732 3476 26776
rect 3436 26692 4204 26732
rect 4244 26692 4876 26732
rect 4916 26692 4925 26732
rect 0 26648 80 26668
rect 0 26608 652 26648
rect 692 26608 701 26648
rect 11011 26608 11020 26648
rect 11060 26608 11404 26648
rect 11444 26608 11453 26648
rect 0 26588 80 26608
rect 4343 26440 4352 26480
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4720 26440 4729 26480
rect 19463 26440 19472 26480
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19840 26440 19849 26480
rect 34583 26440 34592 26480
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34960 26440 34969 26480
rect 49703 26440 49712 26480
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 50080 26440 50089 26480
rect 64823 26440 64832 26480
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 65200 26440 65209 26480
rect 79943 26440 79952 26480
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 80320 26440 80329 26480
rect 5155 26104 5164 26144
rect 5204 26104 5548 26144
rect 5588 26104 5597 26144
rect 11299 26104 11308 26144
rect 11348 26104 11980 26144
rect 12020 26104 12029 26144
rect 9859 25852 9868 25892
rect 9908 25852 11116 25892
rect 11156 25852 11165 25892
rect 0 25808 80 25828
rect 0 25768 652 25808
rect 692 25768 701 25808
rect 0 25748 80 25768
rect 3103 25684 3112 25724
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3480 25684 3489 25724
rect 18223 25684 18232 25724
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18600 25684 18609 25724
rect 33343 25684 33352 25724
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33720 25684 33729 25724
rect 48463 25684 48472 25724
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48840 25684 48849 25724
rect 63583 25684 63592 25724
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63960 25684 63969 25724
rect 78703 25684 78712 25724
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 79080 25684 79089 25724
rect 835 25516 844 25556
rect 884 25516 1132 25556
rect 1172 25516 1181 25556
rect 11011 25348 11020 25388
rect 11060 25348 11692 25388
rect 11732 25348 12652 25388
rect 12692 25348 12701 25388
rect 12067 25264 12076 25304
rect 12116 25264 12556 25304
rect 12596 25264 12605 25304
rect 451 25180 460 25220
rect 500 25180 12364 25220
rect 12404 25180 12413 25220
rect 0 24968 80 24988
rect 0 24928 652 24968
rect 692 24928 701 24968
rect 4343 24928 4352 24968
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4720 24928 4729 24968
rect 19463 24928 19472 24968
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19840 24928 19849 24968
rect 34583 24928 34592 24968
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34960 24928 34969 24968
rect 49703 24928 49712 24968
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 50080 24928 50089 24968
rect 64823 24928 64832 24968
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 65200 24928 65209 24968
rect 79943 24928 79952 24968
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 80320 24928 80329 24968
rect 0 24908 80 24928
rect 9955 24760 9964 24800
rect 10004 24760 10828 24800
rect 10868 24760 10877 24800
rect 4771 24676 4780 24716
rect 4820 24676 5356 24716
rect 5396 24676 6320 24716
rect 6595 24676 6604 24716
rect 6644 24676 9772 24716
rect 9812 24676 9821 24716
rect 6280 24632 6320 24676
rect 4195 24592 4204 24632
rect 4244 24592 5452 24632
rect 5492 24592 5501 24632
rect 6280 24592 6508 24632
rect 6548 24592 6557 24632
rect 4003 24508 4012 24548
rect 4052 24508 6604 24548
rect 6644 24508 6653 24548
rect 835 24340 844 24380
rect 884 24340 12364 24380
rect 12404 24340 12413 24380
rect 3103 24172 3112 24212
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3480 24172 3489 24212
rect 18223 24172 18232 24212
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18600 24172 18609 24212
rect 33343 24172 33352 24212
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33720 24172 33729 24212
rect 48463 24172 48472 24212
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48840 24172 48849 24212
rect 63583 24172 63592 24212
rect 63632 24172 63674 24212
rect 63714 24172 63756 24212
rect 63796 24172 63838 24212
rect 63878 24172 63920 24212
rect 63960 24172 63969 24212
rect 78703 24172 78712 24212
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 79080 24172 79089 24212
rect 0 24128 80 24148
rect 0 24088 652 24128
rect 692 24088 701 24128
rect 1123 24088 1132 24128
rect 1172 24088 5356 24128
rect 5396 24088 5405 24128
rect 0 24068 80 24088
rect 1891 24004 1900 24044
rect 1940 24004 3532 24044
rect 3572 24004 4300 24044
rect 4340 24004 4349 24044
rect 11395 24004 11404 24044
rect 11444 24004 12172 24044
rect 12212 24004 12221 24044
rect 1027 23836 1036 23876
rect 1076 23836 1804 23876
rect 1844 23836 2476 23876
rect 2516 23836 2525 23876
rect 739 23752 748 23792
rect 788 23752 1996 23792
rect 2036 23752 2188 23792
rect 2228 23752 2237 23792
rect 2659 23668 2668 23708
rect 2708 23668 4300 23708
rect 4340 23668 4684 23708
rect 4724 23668 4733 23708
rect 4343 23416 4352 23456
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4720 23416 4729 23456
rect 19463 23416 19472 23456
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19840 23416 19849 23456
rect 34583 23416 34592 23456
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34960 23416 34969 23456
rect 49703 23416 49712 23456
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 50080 23416 50089 23456
rect 64823 23416 64832 23456
rect 64872 23416 64914 23456
rect 64954 23416 64996 23456
rect 65036 23416 65078 23456
rect 65118 23416 65160 23456
rect 65200 23416 65209 23456
rect 79943 23416 79952 23456
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 80320 23416 80329 23456
rect 0 23288 80 23308
rect 0 23248 652 23288
rect 692 23248 701 23288
rect 0 23228 80 23248
rect 3103 22660 3112 22700
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3480 22660 3489 22700
rect 18223 22660 18232 22700
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18600 22660 18609 22700
rect 33343 22660 33352 22700
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33720 22660 33729 22700
rect 48463 22660 48472 22700
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48840 22660 48849 22700
rect 63583 22660 63592 22700
rect 63632 22660 63674 22700
rect 63714 22660 63756 22700
rect 63796 22660 63838 22700
rect 63878 22660 63920 22700
rect 63960 22660 63969 22700
rect 78703 22660 78712 22700
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 79080 22660 79089 22700
rect 0 22448 80 22468
rect 0 22408 652 22448
rect 692 22408 701 22448
rect 0 22388 80 22408
rect 11299 22324 11308 22364
rect 11348 22324 11884 22364
rect 11924 22324 11933 22364
rect 8803 22240 8812 22280
rect 8852 22240 10060 22280
rect 10100 22240 11212 22280
rect 11252 22240 11596 22280
rect 11636 22240 11645 22280
rect 1027 22072 1036 22112
rect 1076 22072 11116 22112
rect 11156 22072 11165 22112
rect 4343 21904 4352 21944
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4720 21904 4729 21944
rect 19463 21904 19472 21944
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19840 21904 19849 21944
rect 34583 21904 34592 21944
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34960 21904 34969 21944
rect 49703 21904 49712 21944
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 50080 21904 50089 21944
rect 64823 21904 64832 21944
rect 64872 21904 64914 21944
rect 64954 21904 64996 21944
rect 65036 21904 65078 21944
rect 65118 21904 65160 21944
rect 65200 21904 65209 21944
rect 79943 21904 79952 21944
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 80320 21904 80329 21944
rect 0 21608 80 21628
rect 0 21568 652 21608
rect 692 21568 701 21608
rect 0 21548 80 21568
rect 3103 21148 3112 21188
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3480 21148 3489 21188
rect 18223 21148 18232 21188
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18600 21148 18609 21188
rect 33343 21148 33352 21188
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33720 21148 33729 21188
rect 48463 21148 48472 21188
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48840 21148 48849 21188
rect 63583 21148 63592 21188
rect 63632 21148 63674 21188
rect 63714 21148 63756 21188
rect 63796 21148 63838 21188
rect 63878 21148 63920 21188
rect 63960 21148 63969 21188
rect 78703 21148 78712 21188
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 79080 21148 79089 21188
rect 1219 20812 1228 20852
rect 1268 20812 3436 20852
rect 3476 20812 4108 20852
rect 4148 20812 4157 20852
rect 0 20768 80 20788
rect 0 20728 652 20768
rect 692 20728 701 20768
rect 835 20728 844 20768
rect 884 20728 3820 20768
rect 3860 20728 4012 20768
rect 4052 20728 4061 20768
rect 0 20708 80 20728
rect 4291 20644 4300 20684
rect 4340 20644 8524 20684
rect 8564 20644 8573 20684
rect 4343 20392 4352 20432
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4720 20392 4729 20432
rect 19463 20392 19472 20432
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19840 20392 19849 20432
rect 34583 20392 34592 20432
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34960 20392 34969 20432
rect 49703 20392 49712 20432
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 50080 20392 50089 20432
rect 64823 20392 64832 20432
rect 64872 20392 64914 20432
rect 64954 20392 64996 20432
rect 65036 20392 65078 20432
rect 65118 20392 65160 20432
rect 65200 20392 65209 20432
rect 79943 20392 79952 20432
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 80320 20392 80329 20432
rect 8035 20224 8044 20264
rect 8084 20224 8332 20264
rect 8372 20224 8620 20264
rect 8660 20224 8669 20264
rect 2500 20140 7852 20180
rect 7892 20140 7901 20180
rect 8236 20140 8908 20180
rect 8948 20140 8957 20180
rect 2500 20096 2540 20140
rect 8236 20096 8276 20140
rect 355 20056 364 20096
rect 404 20056 2540 20096
rect 8227 20056 8236 20096
rect 8276 20056 8285 20096
rect 0 19928 80 19948
rect 0 19888 652 19928
rect 692 19888 701 19928
rect 0 19868 80 19888
rect 1219 19804 1228 19844
rect 1268 19804 3340 19844
rect 3380 19804 3389 19844
rect 3103 19636 3112 19676
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3480 19636 3489 19676
rect 18223 19636 18232 19676
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18600 19636 18609 19676
rect 33343 19636 33352 19676
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33720 19636 33729 19676
rect 48463 19636 48472 19676
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48840 19636 48849 19676
rect 63583 19636 63592 19676
rect 63632 19636 63674 19676
rect 63714 19636 63756 19676
rect 63796 19636 63838 19676
rect 63878 19636 63920 19676
rect 63960 19636 63969 19676
rect 78703 19636 78712 19676
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 79080 19636 79089 19676
rect 0 19088 80 19108
rect 0 19048 652 19088
rect 692 19048 701 19088
rect 931 19048 940 19088
rect 980 19048 8044 19088
rect 8084 19048 9100 19088
rect 9140 19048 9149 19088
rect 0 19028 80 19048
rect 4343 18880 4352 18920
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4720 18880 4729 18920
rect 19463 18880 19472 18920
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19840 18880 19849 18920
rect 34583 18880 34592 18920
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34960 18880 34969 18920
rect 49703 18880 49712 18920
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 50080 18880 50089 18920
rect 64823 18880 64832 18920
rect 64872 18880 64914 18920
rect 64954 18880 64996 18920
rect 65036 18880 65078 18920
rect 65118 18880 65160 18920
rect 65200 18880 65209 18920
rect 79943 18880 79952 18920
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 80320 18880 80329 18920
rect 0 18248 80 18268
rect 0 18208 652 18248
rect 692 18208 701 18248
rect 0 18188 80 18208
rect 3103 18124 3112 18164
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3480 18124 3489 18164
rect 18223 18124 18232 18164
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18600 18124 18609 18164
rect 33343 18124 33352 18164
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33720 18124 33729 18164
rect 48463 18124 48472 18164
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48840 18124 48849 18164
rect 63583 18124 63592 18164
rect 63632 18124 63674 18164
rect 63714 18124 63756 18164
rect 63796 18124 63838 18164
rect 63878 18124 63920 18164
rect 63960 18124 63969 18164
rect 78703 18124 78712 18164
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 79080 18124 79089 18164
rect 0 17408 80 17428
rect 0 17368 652 17408
rect 692 17368 701 17408
rect 4343 17368 4352 17408
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4720 17368 4729 17408
rect 19463 17368 19472 17408
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19840 17368 19849 17408
rect 34583 17368 34592 17408
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34960 17368 34969 17408
rect 49703 17368 49712 17408
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 50080 17368 50089 17408
rect 64823 17368 64832 17408
rect 64872 17368 64914 17408
rect 64954 17368 64996 17408
rect 65036 17368 65078 17408
rect 65118 17368 65160 17408
rect 65200 17368 65209 17408
rect 79943 17368 79952 17408
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 80320 17368 80329 17408
rect 0 17348 80 17368
rect 3103 16612 3112 16652
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3480 16612 3489 16652
rect 18223 16612 18232 16652
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18600 16612 18609 16652
rect 33343 16612 33352 16652
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33720 16612 33729 16652
rect 48463 16612 48472 16652
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48840 16612 48849 16652
rect 63583 16612 63592 16652
rect 63632 16612 63674 16652
rect 63714 16612 63756 16652
rect 63796 16612 63838 16652
rect 63878 16612 63920 16652
rect 63960 16612 63969 16652
rect 78703 16612 78712 16652
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 79080 16612 79089 16652
rect 0 16568 80 16588
rect 0 16528 652 16568
rect 692 16528 701 16568
rect 0 16508 80 16528
rect 4343 15856 4352 15896
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4720 15856 4729 15896
rect 19463 15856 19472 15896
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19840 15856 19849 15896
rect 34583 15856 34592 15896
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34960 15856 34969 15896
rect 49703 15856 49712 15896
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 50080 15856 50089 15896
rect 64823 15856 64832 15896
rect 64872 15856 64914 15896
rect 64954 15856 64996 15896
rect 65036 15856 65078 15896
rect 65118 15856 65160 15896
rect 65200 15856 65209 15896
rect 79943 15856 79952 15896
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 80320 15856 80329 15896
rect 451 15772 460 15812
rect 500 15772 940 15812
rect 980 15772 989 15812
rect 0 15728 80 15748
rect 0 15688 556 15728
rect 596 15688 605 15728
rect 0 15668 80 15688
rect 3103 15100 3112 15140
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3480 15100 3489 15140
rect 18223 15100 18232 15140
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18600 15100 18609 15140
rect 33343 15100 33352 15140
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 33720 15100 33729 15140
rect 48463 15100 48472 15140
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48840 15100 48849 15140
rect 63583 15100 63592 15140
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63960 15100 63969 15140
rect 78703 15100 78712 15140
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 79080 15100 79089 15140
rect 0 14888 80 14908
rect 0 14848 652 14888
rect 692 14848 701 14888
rect 0 14828 80 14848
rect 4343 14344 4352 14384
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4720 14344 4729 14384
rect 19463 14344 19472 14384
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19840 14344 19849 14384
rect 34583 14344 34592 14384
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34960 14344 34969 14384
rect 49703 14344 49712 14384
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 50080 14344 50089 14384
rect 64823 14344 64832 14384
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 65200 14344 65209 14384
rect 79943 14344 79952 14384
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 80320 14344 80329 14384
rect 0 14048 80 14068
rect 0 14008 652 14048
rect 692 14008 701 14048
rect 0 13988 80 14008
rect 3103 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 3489 13628
rect 18223 13588 18232 13628
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18600 13588 18609 13628
rect 33343 13588 33352 13628
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33720 13588 33729 13628
rect 48463 13588 48472 13628
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48840 13588 48849 13628
rect 63583 13588 63592 13628
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63960 13588 63969 13628
rect 78703 13588 78712 13628
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 79080 13588 79089 13628
rect 0 13208 80 13228
rect 0 13168 652 13208
rect 692 13168 701 13208
rect 0 13148 80 13168
rect 4343 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 4729 12872
rect 19463 12832 19472 12872
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19840 12832 19849 12872
rect 34583 12832 34592 12872
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34960 12832 34969 12872
rect 49703 12832 49712 12872
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 50080 12832 50089 12872
rect 64823 12832 64832 12872
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 65200 12832 65209 12872
rect 79943 12832 79952 12872
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 80320 12832 80329 12872
rect 0 12368 80 12388
rect 0 12328 652 12368
rect 692 12328 701 12368
rect 0 12308 80 12328
rect 3103 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 3489 12116
rect 18223 12076 18232 12116
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18600 12076 18609 12116
rect 33343 12076 33352 12116
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33720 12076 33729 12116
rect 48463 12076 48472 12116
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48840 12076 48849 12116
rect 63583 12076 63592 12116
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63960 12076 63969 12116
rect 78703 12076 78712 12116
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 79080 12076 79089 12116
rect 0 11528 80 11548
rect 0 11488 652 11528
rect 692 11488 701 11528
rect 0 11468 80 11488
rect 4343 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 4729 11360
rect 19463 11320 19472 11360
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19840 11320 19849 11360
rect 34583 11320 34592 11360
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34960 11320 34969 11360
rect 49703 11320 49712 11360
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 50080 11320 50089 11360
rect 64823 11320 64832 11360
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 65200 11320 65209 11360
rect 79943 11320 79952 11360
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 80320 11320 80329 11360
rect 0 10688 80 10708
rect 0 10648 652 10688
rect 692 10648 701 10688
rect 0 10628 80 10648
rect 3103 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 3489 10604
rect 18223 10564 18232 10604
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18600 10564 18609 10604
rect 33343 10564 33352 10604
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33720 10564 33729 10604
rect 48463 10564 48472 10604
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48840 10564 48849 10604
rect 63583 10564 63592 10604
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63960 10564 63969 10604
rect 78703 10564 78712 10604
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 79080 10564 79089 10604
rect 0 9848 80 9868
rect 0 9808 652 9848
rect 692 9808 701 9848
rect 4343 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 4729 9848
rect 19463 9808 19472 9848
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19840 9808 19849 9848
rect 34583 9808 34592 9848
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34960 9808 34969 9848
rect 49703 9808 49712 9848
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 50080 9808 50089 9848
rect 64823 9808 64832 9848
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 65200 9808 65209 9848
rect 79943 9808 79952 9848
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 80320 9808 80329 9848
rect 0 9788 80 9808
rect 3103 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 3489 9092
rect 18223 9052 18232 9092
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18600 9052 18609 9092
rect 33343 9052 33352 9092
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33720 9052 33729 9092
rect 48463 9052 48472 9092
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48840 9052 48849 9092
rect 63583 9052 63592 9092
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63960 9052 63969 9092
rect 78703 9052 78712 9092
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 79080 9052 79089 9092
rect 0 9008 80 9028
rect 0 8968 652 9008
rect 692 8968 701 9008
rect 0 8948 80 8968
rect 4343 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 4729 8336
rect 19463 8296 19472 8336
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19840 8296 19849 8336
rect 34583 8296 34592 8336
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34960 8296 34969 8336
rect 49703 8296 49712 8336
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 50080 8296 50089 8336
rect 64823 8296 64832 8336
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 65200 8296 65209 8336
rect 79943 8296 79952 8336
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 80320 8296 80329 8336
rect 0 8168 80 8188
rect 0 8128 652 8168
rect 692 8128 701 8168
rect 0 8108 80 8128
rect 835 7876 844 7916
rect 884 7876 2092 7916
rect 2132 7876 2141 7916
rect 3103 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 3489 7580
rect 18223 7540 18232 7580
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18600 7540 18609 7580
rect 33343 7540 33352 7580
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33720 7540 33729 7580
rect 48463 7540 48472 7580
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48840 7540 48849 7580
rect 63583 7540 63592 7580
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63960 7540 63969 7580
rect 78703 7540 78712 7580
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 79080 7540 79089 7580
rect 0 7328 80 7348
rect 0 7288 652 7328
rect 692 7288 701 7328
rect 0 7268 80 7288
rect 835 7204 844 7244
rect 884 7204 1132 7244
rect 1172 7204 1181 7244
rect 4343 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 4729 6824
rect 19463 6784 19472 6824
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19840 6784 19849 6824
rect 34583 6784 34592 6824
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34960 6784 34969 6824
rect 49703 6784 49712 6824
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 50080 6784 50089 6824
rect 64823 6784 64832 6824
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 65200 6784 65209 6824
rect 79943 6784 79952 6824
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 80320 6784 80329 6824
rect 0 6488 80 6508
rect 0 6448 652 6488
rect 692 6448 701 6488
rect 0 6428 80 6448
rect 3103 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 3489 6068
rect 18223 6028 18232 6068
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18600 6028 18609 6068
rect 33343 6028 33352 6068
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33720 6028 33729 6068
rect 48463 6028 48472 6068
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48840 6028 48849 6068
rect 63583 6028 63592 6068
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63960 6028 63969 6068
rect 78703 6028 78712 6068
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 79080 6028 79089 6068
rect 835 5692 844 5732
rect 884 5692 6412 5732
rect 6452 5692 6461 5732
rect 0 5648 80 5668
rect 0 5608 652 5648
rect 692 5608 701 5648
rect 0 5588 80 5608
rect 4343 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 4729 5312
rect 19463 5272 19472 5312
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19840 5272 19849 5312
rect 34583 5272 34592 5312
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34960 5272 34969 5312
rect 49703 5272 49712 5312
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 50080 5272 50089 5312
rect 64823 5272 64832 5312
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 65200 5272 65209 5312
rect 79943 5272 79952 5312
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 80320 5272 80329 5312
rect 0 4808 80 4828
rect 0 4768 652 4808
rect 692 4768 701 4808
rect 0 4748 80 4768
rect 3103 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 3489 4556
rect 18223 4516 18232 4556
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18600 4516 18609 4556
rect 33343 4516 33352 4556
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33720 4516 33729 4556
rect 48463 4516 48472 4556
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48840 4516 48849 4556
rect 63583 4516 63592 4556
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63960 4516 63969 4556
rect 78703 4516 78712 4556
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 79080 4516 79089 4556
rect 0 3968 80 3988
rect 0 3928 652 3968
rect 692 3928 701 3968
rect 0 3908 80 3928
rect 4343 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 4729 3800
rect 19463 3760 19472 3800
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19840 3760 19849 3800
rect 34583 3760 34592 3800
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34960 3760 34969 3800
rect 49703 3760 49712 3800
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 50080 3760 50089 3800
rect 64823 3760 64832 3800
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 65200 3760 65209 3800
rect 79943 3760 79952 3800
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 80320 3760 80329 3800
rect 643 3172 652 3212
rect 692 3172 701 3212
rect 0 3128 80 3148
rect 652 3128 692 3172
rect 0 3088 692 3128
rect 0 3068 80 3088
rect 3103 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 3489 3044
rect 18223 3004 18232 3044
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18600 3004 18609 3044
rect 33343 3004 33352 3044
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33720 3004 33729 3044
rect 48463 3004 48472 3044
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48840 3004 48849 3044
rect 63583 3004 63592 3044
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63960 3004 63969 3044
rect 78703 3004 78712 3044
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 79080 3004 79089 3044
rect 0 2288 80 2308
rect 0 2248 652 2288
rect 692 2248 701 2288
rect 4343 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 4729 2288
rect 19463 2248 19472 2288
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19840 2248 19849 2288
rect 34583 2248 34592 2288
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34960 2248 34969 2288
rect 49703 2248 49712 2288
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 50080 2248 50089 2288
rect 64823 2248 64832 2288
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 65200 2248 65209 2288
rect 79943 2248 79952 2288
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 80320 2248 80329 2288
rect 0 2228 80 2248
rect 3103 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 3489 1532
rect 18223 1492 18232 1532
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18600 1492 18609 1532
rect 33343 1492 33352 1532
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33720 1492 33729 1532
rect 48463 1492 48472 1532
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48840 1492 48849 1532
rect 63583 1492 63592 1532
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63960 1492 63969 1532
rect 78703 1492 78712 1532
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 79080 1492 79089 1532
rect 4343 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 4729 776
rect 19463 736 19472 776
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19840 736 19849 776
rect 34583 736 34592 776
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34960 736 34969 776
rect 49703 736 49712 776
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 50080 736 50089 776
rect 64823 736 64832 776
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 65200 736 65209 776
rect 79943 736 79952 776
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 80320 736 80329 776
<< via3 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 63592 24172 63632 24212
rect 63674 24172 63714 24212
rect 63756 24172 63796 24212
rect 63838 24172 63878 24212
rect 63920 24172 63960 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 64832 23416 64872 23456
rect 64914 23416 64954 23456
rect 64996 23416 65036 23456
rect 65078 23416 65118 23456
rect 65160 23416 65200 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 63592 22660 63632 22700
rect 63674 22660 63714 22700
rect 63756 22660 63796 22700
rect 63838 22660 63878 22700
rect 63920 22660 63960 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 64832 21904 64872 21944
rect 64914 21904 64954 21944
rect 64996 21904 65036 21944
rect 65078 21904 65118 21944
rect 65160 21904 65200 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 63592 21148 63632 21188
rect 63674 21148 63714 21188
rect 63756 21148 63796 21188
rect 63838 21148 63878 21188
rect 63920 21148 63960 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 64832 20392 64872 20432
rect 64914 20392 64954 20432
rect 64996 20392 65036 20432
rect 65078 20392 65118 20432
rect 65160 20392 65200 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 63592 19636 63632 19676
rect 63674 19636 63714 19676
rect 63756 19636 63796 19676
rect 63838 19636 63878 19676
rect 63920 19636 63960 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 64832 18880 64872 18920
rect 64914 18880 64954 18920
rect 64996 18880 65036 18920
rect 65078 18880 65118 18920
rect 65160 18880 65200 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 63592 18124 63632 18164
rect 63674 18124 63714 18164
rect 63756 18124 63796 18164
rect 63838 18124 63878 18164
rect 63920 18124 63960 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 64832 17368 64872 17408
rect 64914 17368 64954 17408
rect 64996 17368 65036 17408
rect 65078 17368 65118 17408
rect 65160 17368 65200 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 63592 16612 63632 16652
rect 63674 16612 63714 16652
rect 63756 16612 63796 16652
rect 63838 16612 63878 16652
rect 63920 16612 63960 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 64832 15856 64872 15896
rect 64914 15856 64954 15896
rect 64996 15856 65036 15896
rect 65078 15856 65118 15896
rect 65160 15856 65200 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
<< metal4 >>
rect 4352 38576 4720 38585
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4352 38527 4720 38536
rect 19472 38576 19840 38585
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19472 38527 19840 38536
rect 34592 38576 34960 38585
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34592 38527 34960 38536
rect 49712 38576 50080 38585
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 49712 38527 50080 38536
rect 64832 38576 65200 38585
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 64832 38527 65200 38536
rect 79952 38576 80320 38585
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 79952 38527 80320 38536
rect 3112 37820 3480 37829
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3112 37771 3480 37780
rect 18232 37820 18600 37829
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18232 37771 18600 37780
rect 33352 37820 33720 37829
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33352 37771 33720 37780
rect 48472 37820 48840 37829
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48472 37771 48840 37780
rect 63592 37820 63960 37829
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63592 37771 63960 37780
rect 78712 37820 79080 37829
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 78712 37771 79080 37780
rect 4352 37064 4720 37073
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4352 37015 4720 37024
rect 19472 37064 19840 37073
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19472 37015 19840 37024
rect 34592 37064 34960 37073
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34592 37015 34960 37024
rect 49712 37064 50080 37073
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 49712 37015 50080 37024
rect 64832 37064 65200 37073
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 64832 37015 65200 37024
rect 79952 37064 80320 37073
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 79952 37015 80320 37024
rect 3112 36308 3480 36317
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3112 36259 3480 36268
rect 18232 36308 18600 36317
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18232 36259 18600 36268
rect 33352 36308 33720 36317
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33352 36259 33720 36268
rect 48472 36308 48840 36317
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48472 36259 48840 36268
rect 63592 36308 63960 36317
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63592 36259 63960 36268
rect 78712 36308 79080 36317
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 78712 36259 79080 36268
rect 4352 35552 4720 35561
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4352 35503 4720 35512
rect 19472 35552 19840 35561
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19472 35503 19840 35512
rect 34592 35552 34960 35561
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34592 35503 34960 35512
rect 49712 35552 50080 35561
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 49712 35503 50080 35512
rect 64832 35552 65200 35561
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 64832 35503 65200 35512
rect 79952 35552 80320 35561
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 79952 35503 80320 35512
rect 3112 34796 3480 34805
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3112 34747 3480 34756
rect 18232 34796 18600 34805
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18232 34747 18600 34756
rect 33352 34796 33720 34805
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33352 34747 33720 34756
rect 48472 34796 48840 34805
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48472 34747 48840 34756
rect 63592 34796 63960 34805
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63592 34747 63960 34756
rect 78712 34796 79080 34805
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 78712 34747 79080 34756
rect 4352 34040 4720 34049
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4352 33991 4720 34000
rect 19472 34040 19840 34049
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19472 33991 19840 34000
rect 34592 34040 34960 34049
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34592 33991 34960 34000
rect 49712 34040 50080 34049
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 49712 33991 50080 34000
rect 64832 34040 65200 34049
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 64832 33991 65200 34000
rect 79952 34040 80320 34049
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 79952 33991 80320 34000
rect 3112 33284 3480 33293
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3112 33235 3480 33244
rect 18232 33284 18600 33293
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18232 33235 18600 33244
rect 33352 33284 33720 33293
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33352 33235 33720 33244
rect 48472 33284 48840 33293
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48472 33235 48840 33244
rect 63592 33284 63960 33293
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63592 33235 63960 33244
rect 78712 33284 79080 33293
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 78712 33235 79080 33244
rect 4352 32528 4720 32537
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4352 32479 4720 32488
rect 19472 32528 19840 32537
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19472 32479 19840 32488
rect 34592 32528 34960 32537
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34592 32479 34960 32488
rect 49712 32528 50080 32537
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 49712 32479 50080 32488
rect 64832 32528 65200 32537
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 64832 32479 65200 32488
rect 79952 32528 80320 32537
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 79952 32479 80320 32488
rect 3112 31772 3480 31781
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3112 31723 3480 31732
rect 18232 31772 18600 31781
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18232 31723 18600 31732
rect 33352 31772 33720 31781
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33352 31723 33720 31732
rect 48472 31772 48840 31781
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48472 31723 48840 31732
rect 63592 31772 63960 31781
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63592 31723 63960 31732
rect 78712 31772 79080 31781
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 78712 31723 79080 31732
rect 4352 31016 4720 31025
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4352 30967 4720 30976
rect 19472 31016 19840 31025
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19472 30967 19840 30976
rect 34592 31016 34960 31025
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34592 30967 34960 30976
rect 49712 31016 50080 31025
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 49712 30967 50080 30976
rect 64832 31016 65200 31025
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 64832 30967 65200 30976
rect 79952 31016 80320 31025
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 79952 30967 80320 30976
rect 3112 30260 3480 30269
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3112 30211 3480 30220
rect 18232 30260 18600 30269
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18232 30211 18600 30220
rect 33352 30260 33720 30269
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33352 30211 33720 30220
rect 48472 30260 48840 30269
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48472 30211 48840 30220
rect 63592 30260 63960 30269
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63592 30211 63960 30220
rect 78712 30260 79080 30269
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 78712 30211 79080 30220
rect 4352 29504 4720 29513
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4352 29455 4720 29464
rect 19472 29504 19840 29513
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19472 29455 19840 29464
rect 34592 29504 34960 29513
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34592 29455 34960 29464
rect 49712 29504 50080 29513
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 49712 29455 50080 29464
rect 64832 29504 65200 29513
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 64832 29455 65200 29464
rect 79952 29504 80320 29513
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 79952 29455 80320 29464
rect 3112 28748 3480 28757
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3112 28699 3480 28708
rect 18232 28748 18600 28757
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18232 28699 18600 28708
rect 33352 28748 33720 28757
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33352 28699 33720 28708
rect 48472 28748 48840 28757
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48472 28699 48840 28708
rect 63592 28748 63960 28757
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63592 28699 63960 28708
rect 78712 28748 79080 28757
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 78712 28699 79080 28708
rect 4352 27992 4720 28001
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4352 27943 4720 27952
rect 19472 27992 19840 28001
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19472 27943 19840 27952
rect 34592 27992 34960 28001
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34592 27943 34960 27952
rect 49712 27992 50080 28001
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 49712 27943 50080 27952
rect 64832 27992 65200 28001
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 64832 27943 65200 27952
rect 79952 27992 80320 28001
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 79952 27943 80320 27952
rect 3112 27236 3480 27245
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3112 27187 3480 27196
rect 18232 27236 18600 27245
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18232 27187 18600 27196
rect 33352 27236 33720 27245
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33352 27187 33720 27196
rect 48472 27236 48840 27245
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48472 27187 48840 27196
rect 63592 27236 63960 27245
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63592 27187 63960 27196
rect 78712 27236 79080 27245
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 78712 27187 79080 27196
rect 4352 26480 4720 26489
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4352 26431 4720 26440
rect 19472 26480 19840 26489
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19472 26431 19840 26440
rect 34592 26480 34960 26489
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34592 26431 34960 26440
rect 49712 26480 50080 26489
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 49712 26431 50080 26440
rect 64832 26480 65200 26489
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 64832 26431 65200 26440
rect 79952 26480 80320 26489
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 79952 26431 80320 26440
rect 3112 25724 3480 25733
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3112 25675 3480 25684
rect 18232 25724 18600 25733
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18232 25675 18600 25684
rect 33352 25724 33720 25733
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33352 25675 33720 25684
rect 48472 25724 48840 25733
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48472 25675 48840 25684
rect 63592 25724 63960 25733
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63592 25675 63960 25684
rect 78712 25724 79080 25733
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 78712 25675 79080 25684
rect 4352 24968 4720 24977
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4352 24919 4720 24928
rect 19472 24968 19840 24977
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19472 24919 19840 24928
rect 34592 24968 34960 24977
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34592 24919 34960 24928
rect 49712 24968 50080 24977
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 49712 24919 50080 24928
rect 64832 24968 65200 24977
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 64832 24919 65200 24928
rect 79952 24968 80320 24977
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 79952 24919 80320 24928
rect 3112 24212 3480 24221
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3112 24163 3480 24172
rect 18232 24212 18600 24221
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18232 24163 18600 24172
rect 33352 24212 33720 24221
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33352 24163 33720 24172
rect 48472 24212 48840 24221
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48472 24163 48840 24172
rect 63592 24212 63960 24221
rect 63632 24172 63674 24212
rect 63714 24172 63756 24212
rect 63796 24172 63838 24212
rect 63878 24172 63920 24212
rect 63592 24163 63960 24172
rect 78712 24212 79080 24221
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 78712 24163 79080 24172
rect 4352 23456 4720 23465
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4352 23407 4720 23416
rect 19472 23456 19840 23465
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19472 23407 19840 23416
rect 34592 23456 34960 23465
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34592 23407 34960 23416
rect 49712 23456 50080 23465
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 49712 23407 50080 23416
rect 64832 23456 65200 23465
rect 64872 23416 64914 23456
rect 64954 23416 64996 23456
rect 65036 23416 65078 23456
rect 65118 23416 65160 23456
rect 64832 23407 65200 23416
rect 79952 23456 80320 23465
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 79952 23407 80320 23416
rect 3112 22700 3480 22709
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3112 22651 3480 22660
rect 18232 22700 18600 22709
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18232 22651 18600 22660
rect 33352 22700 33720 22709
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33352 22651 33720 22660
rect 48472 22700 48840 22709
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48472 22651 48840 22660
rect 63592 22700 63960 22709
rect 63632 22660 63674 22700
rect 63714 22660 63756 22700
rect 63796 22660 63838 22700
rect 63878 22660 63920 22700
rect 63592 22651 63960 22660
rect 78712 22700 79080 22709
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 78712 22651 79080 22660
rect 4352 21944 4720 21953
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4352 21895 4720 21904
rect 19472 21944 19840 21953
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19472 21895 19840 21904
rect 34592 21944 34960 21953
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34592 21895 34960 21904
rect 49712 21944 50080 21953
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 49712 21895 50080 21904
rect 64832 21944 65200 21953
rect 64872 21904 64914 21944
rect 64954 21904 64996 21944
rect 65036 21904 65078 21944
rect 65118 21904 65160 21944
rect 64832 21895 65200 21904
rect 79952 21944 80320 21953
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 79952 21895 80320 21904
rect 3112 21188 3480 21197
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3112 21139 3480 21148
rect 18232 21188 18600 21197
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18232 21139 18600 21148
rect 33352 21188 33720 21197
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33352 21139 33720 21148
rect 48472 21188 48840 21197
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48472 21139 48840 21148
rect 63592 21188 63960 21197
rect 63632 21148 63674 21188
rect 63714 21148 63756 21188
rect 63796 21148 63838 21188
rect 63878 21148 63920 21188
rect 63592 21139 63960 21148
rect 78712 21188 79080 21197
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 78712 21139 79080 21148
rect 4352 20432 4720 20441
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4352 20383 4720 20392
rect 19472 20432 19840 20441
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19472 20383 19840 20392
rect 34592 20432 34960 20441
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34592 20383 34960 20392
rect 49712 20432 50080 20441
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 49712 20383 50080 20392
rect 64832 20432 65200 20441
rect 64872 20392 64914 20432
rect 64954 20392 64996 20432
rect 65036 20392 65078 20432
rect 65118 20392 65160 20432
rect 64832 20383 65200 20392
rect 79952 20432 80320 20441
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 79952 20383 80320 20392
rect 3112 19676 3480 19685
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3112 19627 3480 19636
rect 18232 19676 18600 19685
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18232 19627 18600 19636
rect 33352 19676 33720 19685
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33352 19627 33720 19636
rect 48472 19676 48840 19685
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48472 19627 48840 19636
rect 63592 19676 63960 19685
rect 63632 19636 63674 19676
rect 63714 19636 63756 19676
rect 63796 19636 63838 19676
rect 63878 19636 63920 19676
rect 63592 19627 63960 19636
rect 78712 19676 79080 19685
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 78712 19627 79080 19636
rect 4352 18920 4720 18929
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4352 18871 4720 18880
rect 19472 18920 19840 18929
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19472 18871 19840 18880
rect 34592 18920 34960 18929
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34592 18871 34960 18880
rect 49712 18920 50080 18929
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 49712 18871 50080 18880
rect 64832 18920 65200 18929
rect 64872 18880 64914 18920
rect 64954 18880 64996 18920
rect 65036 18880 65078 18920
rect 65118 18880 65160 18920
rect 64832 18871 65200 18880
rect 79952 18920 80320 18929
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 79952 18871 80320 18880
rect 3112 18164 3480 18173
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3112 18115 3480 18124
rect 18232 18164 18600 18173
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18232 18115 18600 18124
rect 33352 18164 33720 18173
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33352 18115 33720 18124
rect 48472 18164 48840 18173
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48472 18115 48840 18124
rect 63592 18164 63960 18173
rect 63632 18124 63674 18164
rect 63714 18124 63756 18164
rect 63796 18124 63838 18164
rect 63878 18124 63920 18164
rect 63592 18115 63960 18124
rect 78712 18164 79080 18173
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 78712 18115 79080 18124
rect 4352 17408 4720 17417
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4352 17359 4720 17368
rect 19472 17408 19840 17417
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19472 17359 19840 17368
rect 34592 17408 34960 17417
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34592 17359 34960 17368
rect 49712 17408 50080 17417
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 49712 17359 50080 17368
rect 64832 17408 65200 17417
rect 64872 17368 64914 17408
rect 64954 17368 64996 17408
rect 65036 17368 65078 17408
rect 65118 17368 65160 17408
rect 64832 17359 65200 17368
rect 79952 17408 80320 17417
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 79952 17359 80320 17368
rect 3112 16652 3480 16661
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3112 16603 3480 16612
rect 18232 16652 18600 16661
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18232 16603 18600 16612
rect 33352 16652 33720 16661
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33352 16603 33720 16612
rect 48472 16652 48840 16661
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48472 16603 48840 16612
rect 63592 16652 63960 16661
rect 63632 16612 63674 16652
rect 63714 16612 63756 16652
rect 63796 16612 63838 16652
rect 63878 16612 63920 16652
rect 63592 16603 63960 16612
rect 78712 16652 79080 16661
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 78712 16603 79080 16612
rect 4352 15896 4720 15905
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4352 15847 4720 15856
rect 19472 15896 19840 15905
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19472 15847 19840 15856
rect 34592 15896 34960 15905
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34592 15847 34960 15856
rect 49712 15896 50080 15905
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 49712 15847 50080 15856
rect 64832 15896 65200 15905
rect 64872 15856 64914 15896
rect 64954 15856 64996 15896
rect 65036 15856 65078 15896
rect 65118 15856 65160 15896
rect 64832 15847 65200 15856
rect 79952 15896 80320 15905
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 79952 15847 80320 15856
rect 3112 15140 3480 15149
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3112 15091 3480 15100
rect 18232 15140 18600 15149
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18232 15091 18600 15100
rect 33352 15140 33720 15149
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 33352 15091 33720 15100
rect 48472 15140 48840 15149
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48472 15091 48840 15100
rect 63592 15140 63960 15149
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63592 15091 63960 15100
rect 78712 15140 79080 15149
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 78712 15091 79080 15100
rect 4352 14384 4720 14393
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4352 14335 4720 14344
rect 19472 14384 19840 14393
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19472 14335 19840 14344
rect 34592 14384 34960 14393
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34592 14335 34960 14344
rect 49712 14384 50080 14393
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 49712 14335 50080 14344
rect 64832 14384 65200 14393
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 64832 14335 65200 14344
rect 79952 14384 80320 14393
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 79952 14335 80320 14344
rect 3112 13628 3480 13637
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3112 13579 3480 13588
rect 18232 13628 18600 13637
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18232 13579 18600 13588
rect 33352 13628 33720 13637
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33352 13579 33720 13588
rect 48472 13628 48840 13637
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48472 13579 48840 13588
rect 63592 13628 63960 13637
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63592 13579 63960 13588
rect 78712 13628 79080 13637
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 78712 13579 79080 13588
rect 4352 12872 4720 12881
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4352 12823 4720 12832
rect 19472 12872 19840 12881
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19472 12823 19840 12832
rect 34592 12872 34960 12881
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34592 12823 34960 12832
rect 49712 12872 50080 12881
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 49712 12823 50080 12832
rect 64832 12872 65200 12881
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 64832 12823 65200 12832
rect 79952 12872 80320 12881
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 79952 12823 80320 12832
rect 3112 12116 3480 12125
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3112 12067 3480 12076
rect 18232 12116 18600 12125
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18232 12067 18600 12076
rect 33352 12116 33720 12125
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33352 12067 33720 12076
rect 48472 12116 48840 12125
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48472 12067 48840 12076
rect 63592 12116 63960 12125
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63592 12067 63960 12076
rect 78712 12116 79080 12125
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 78712 12067 79080 12076
rect 4352 11360 4720 11369
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4352 11311 4720 11320
rect 19472 11360 19840 11369
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19472 11311 19840 11320
rect 34592 11360 34960 11369
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34592 11311 34960 11320
rect 49712 11360 50080 11369
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 49712 11311 50080 11320
rect 64832 11360 65200 11369
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 64832 11311 65200 11320
rect 79952 11360 80320 11369
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 79952 11311 80320 11320
rect 3112 10604 3480 10613
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3112 10555 3480 10564
rect 18232 10604 18600 10613
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18232 10555 18600 10564
rect 33352 10604 33720 10613
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33352 10555 33720 10564
rect 48472 10604 48840 10613
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48472 10555 48840 10564
rect 63592 10604 63960 10613
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63592 10555 63960 10564
rect 78712 10604 79080 10613
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 78712 10555 79080 10564
rect 4352 9848 4720 9857
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4352 9799 4720 9808
rect 19472 9848 19840 9857
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19472 9799 19840 9808
rect 34592 9848 34960 9857
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34592 9799 34960 9808
rect 49712 9848 50080 9857
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 49712 9799 50080 9808
rect 64832 9848 65200 9857
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 64832 9799 65200 9808
rect 79952 9848 80320 9857
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 79952 9799 80320 9808
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 18232 9092 18600 9101
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18232 9043 18600 9052
rect 33352 9092 33720 9101
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33352 9043 33720 9052
rect 48472 9092 48840 9101
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48472 9043 48840 9052
rect 63592 9092 63960 9101
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63592 9043 63960 9052
rect 78712 9092 79080 9101
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 78712 9043 79080 9052
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 19472 8336 19840 8345
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19472 8287 19840 8296
rect 34592 8336 34960 8345
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34592 8287 34960 8296
rect 49712 8336 50080 8345
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 49712 8287 50080 8296
rect 64832 8336 65200 8345
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 64832 8287 65200 8296
rect 79952 8336 80320 8345
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 79952 8287 80320 8296
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 18232 7580 18600 7589
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18232 7531 18600 7540
rect 33352 7580 33720 7589
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33352 7531 33720 7540
rect 48472 7580 48840 7589
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48472 7531 48840 7540
rect 63592 7580 63960 7589
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63592 7531 63960 7540
rect 78712 7580 79080 7589
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 78712 7531 79080 7540
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 19472 6824 19840 6833
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19472 6775 19840 6784
rect 34592 6824 34960 6833
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34592 6775 34960 6784
rect 49712 6824 50080 6833
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 49712 6775 50080 6784
rect 64832 6824 65200 6833
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 64832 6775 65200 6784
rect 79952 6824 80320 6833
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 79952 6775 80320 6784
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 18232 6068 18600 6077
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18232 6019 18600 6028
rect 33352 6068 33720 6077
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33352 6019 33720 6028
rect 48472 6068 48840 6077
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48472 6019 48840 6028
rect 63592 6068 63960 6077
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63592 6019 63960 6028
rect 78712 6068 79080 6077
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 78712 6019 79080 6028
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 19472 5312 19840 5321
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19472 5263 19840 5272
rect 34592 5312 34960 5321
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34592 5263 34960 5272
rect 49712 5312 50080 5321
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 49712 5263 50080 5272
rect 64832 5312 65200 5321
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 64832 5263 65200 5272
rect 79952 5312 80320 5321
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 79952 5263 80320 5272
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 18232 4556 18600 4565
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18232 4507 18600 4516
rect 33352 4556 33720 4565
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33352 4507 33720 4516
rect 48472 4556 48840 4565
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48472 4507 48840 4516
rect 63592 4556 63960 4565
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63592 4507 63960 4516
rect 78712 4556 79080 4565
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 78712 4507 79080 4516
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 19472 3800 19840 3809
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19472 3751 19840 3760
rect 34592 3800 34960 3809
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34592 3751 34960 3760
rect 49712 3800 50080 3809
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 49712 3751 50080 3760
rect 64832 3800 65200 3809
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 64832 3751 65200 3760
rect 79952 3800 80320 3809
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 79952 3751 80320 3760
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 18232 3044 18600 3053
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18232 2995 18600 3004
rect 33352 3044 33720 3053
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33352 2995 33720 3004
rect 48472 3044 48840 3053
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48472 2995 48840 3004
rect 63592 3044 63960 3053
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63592 2995 63960 3004
rect 78712 3044 79080 3053
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 78712 2995 79080 3004
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 19472 2288 19840 2297
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19472 2239 19840 2248
rect 34592 2288 34960 2297
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34592 2239 34960 2248
rect 49712 2288 50080 2297
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 49712 2239 50080 2248
rect 64832 2288 65200 2297
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 64832 2239 65200 2248
rect 79952 2288 80320 2297
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 79952 2239 80320 2248
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 18232 1532 18600 1541
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18232 1483 18600 1492
rect 33352 1532 33720 1541
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33352 1483 33720 1492
rect 48472 1532 48840 1541
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48472 1483 48840 1492
rect 63592 1532 63960 1541
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63592 1483 63960 1492
rect 78712 1532 79080 1541
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 78712 1483 79080 1492
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
rect 19472 776 19840 785
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19472 727 19840 736
rect 34592 776 34960 785
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34592 727 34960 736
rect 49712 776 50080 785
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 49712 727 50080 736
rect 64832 776 65200 785
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 64832 727 65200 736
rect 79952 776 80320 785
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 79952 727 80320 736
<< via4 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 63592 24172 63632 24212
rect 63674 24172 63714 24212
rect 63756 24172 63796 24212
rect 63838 24172 63878 24212
rect 63920 24172 63960 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 64832 23416 64872 23456
rect 64914 23416 64954 23456
rect 64996 23416 65036 23456
rect 65078 23416 65118 23456
rect 65160 23416 65200 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 63592 22660 63632 22700
rect 63674 22660 63714 22700
rect 63756 22660 63796 22700
rect 63838 22660 63878 22700
rect 63920 22660 63960 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 64832 21904 64872 21944
rect 64914 21904 64954 21944
rect 64996 21904 65036 21944
rect 65078 21904 65118 21944
rect 65160 21904 65200 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 63592 21148 63632 21188
rect 63674 21148 63714 21188
rect 63756 21148 63796 21188
rect 63838 21148 63878 21188
rect 63920 21148 63960 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 64832 20392 64872 20432
rect 64914 20392 64954 20432
rect 64996 20392 65036 20432
rect 65078 20392 65118 20432
rect 65160 20392 65200 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 63592 19636 63632 19676
rect 63674 19636 63714 19676
rect 63756 19636 63796 19676
rect 63838 19636 63878 19676
rect 63920 19636 63960 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 64832 18880 64872 18920
rect 64914 18880 64954 18920
rect 64996 18880 65036 18920
rect 65078 18880 65118 18920
rect 65160 18880 65200 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 63592 18124 63632 18164
rect 63674 18124 63714 18164
rect 63756 18124 63796 18164
rect 63838 18124 63878 18164
rect 63920 18124 63960 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 64832 17368 64872 17408
rect 64914 17368 64954 17408
rect 64996 17368 65036 17408
rect 65078 17368 65118 17408
rect 65160 17368 65200 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 63592 16612 63632 16652
rect 63674 16612 63714 16652
rect 63756 16612 63796 16652
rect 63838 16612 63878 16652
rect 63920 16612 63960 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 64832 15856 64872 15896
rect 64914 15856 64954 15896
rect 64996 15856 65036 15896
rect 65078 15856 65118 15896
rect 65160 15856 65200 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
<< metal5 >>
rect 4343 38599 4729 38618
rect 4343 38576 4409 38599
rect 4495 38576 4577 38599
rect 4663 38576 4729 38599
rect 4343 38536 4352 38576
rect 4392 38536 4409 38576
rect 4495 38536 4516 38576
rect 4556 38536 4577 38576
rect 4663 38536 4680 38576
rect 4720 38536 4729 38576
rect 4343 38513 4409 38536
rect 4495 38513 4577 38536
rect 4663 38513 4729 38536
rect 4343 38494 4729 38513
rect 19463 38599 19849 38618
rect 19463 38576 19529 38599
rect 19615 38576 19697 38599
rect 19783 38576 19849 38599
rect 19463 38536 19472 38576
rect 19512 38536 19529 38576
rect 19615 38536 19636 38576
rect 19676 38536 19697 38576
rect 19783 38536 19800 38576
rect 19840 38536 19849 38576
rect 19463 38513 19529 38536
rect 19615 38513 19697 38536
rect 19783 38513 19849 38536
rect 19463 38494 19849 38513
rect 34583 38599 34969 38618
rect 34583 38576 34649 38599
rect 34735 38576 34817 38599
rect 34903 38576 34969 38599
rect 34583 38536 34592 38576
rect 34632 38536 34649 38576
rect 34735 38536 34756 38576
rect 34796 38536 34817 38576
rect 34903 38536 34920 38576
rect 34960 38536 34969 38576
rect 34583 38513 34649 38536
rect 34735 38513 34817 38536
rect 34903 38513 34969 38536
rect 34583 38494 34969 38513
rect 49703 38599 50089 38618
rect 49703 38576 49769 38599
rect 49855 38576 49937 38599
rect 50023 38576 50089 38599
rect 49703 38536 49712 38576
rect 49752 38536 49769 38576
rect 49855 38536 49876 38576
rect 49916 38536 49937 38576
rect 50023 38536 50040 38576
rect 50080 38536 50089 38576
rect 49703 38513 49769 38536
rect 49855 38513 49937 38536
rect 50023 38513 50089 38536
rect 49703 38494 50089 38513
rect 64823 38599 65209 38618
rect 64823 38576 64889 38599
rect 64975 38576 65057 38599
rect 65143 38576 65209 38599
rect 64823 38536 64832 38576
rect 64872 38536 64889 38576
rect 64975 38536 64996 38576
rect 65036 38536 65057 38576
rect 65143 38536 65160 38576
rect 65200 38536 65209 38576
rect 64823 38513 64889 38536
rect 64975 38513 65057 38536
rect 65143 38513 65209 38536
rect 64823 38494 65209 38513
rect 79943 38599 80329 38618
rect 79943 38576 80009 38599
rect 80095 38576 80177 38599
rect 80263 38576 80329 38599
rect 79943 38536 79952 38576
rect 79992 38536 80009 38576
rect 80095 38536 80116 38576
rect 80156 38536 80177 38576
rect 80263 38536 80280 38576
rect 80320 38536 80329 38576
rect 79943 38513 80009 38536
rect 80095 38513 80177 38536
rect 80263 38513 80329 38536
rect 79943 38494 80329 38513
rect 3103 37843 3489 37862
rect 3103 37820 3169 37843
rect 3255 37820 3337 37843
rect 3423 37820 3489 37843
rect 3103 37780 3112 37820
rect 3152 37780 3169 37820
rect 3255 37780 3276 37820
rect 3316 37780 3337 37820
rect 3423 37780 3440 37820
rect 3480 37780 3489 37820
rect 3103 37757 3169 37780
rect 3255 37757 3337 37780
rect 3423 37757 3489 37780
rect 3103 37738 3489 37757
rect 18223 37843 18609 37862
rect 18223 37820 18289 37843
rect 18375 37820 18457 37843
rect 18543 37820 18609 37843
rect 18223 37780 18232 37820
rect 18272 37780 18289 37820
rect 18375 37780 18396 37820
rect 18436 37780 18457 37820
rect 18543 37780 18560 37820
rect 18600 37780 18609 37820
rect 18223 37757 18289 37780
rect 18375 37757 18457 37780
rect 18543 37757 18609 37780
rect 18223 37738 18609 37757
rect 33343 37843 33729 37862
rect 33343 37820 33409 37843
rect 33495 37820 33577 37843
rect 33663 37820 33729 37843
rect 33343 37780 33352 37820
rect 33392 37780 33409 37820
rect 33495 37780 33516 37820
rect 33556 37780 33577 37820
rect 33663 37780 33680 37820
rect 33720 37780 33729 37820
rect 33343 37757 33409 37780
rect 33495 37757 33577 37780
rect 33663 37757 33729 37780
rect 33343 37738 33729 37757
rect 48463 37843 48849 37862
rect 48463 37820 48529 37843
rect 48615 37820 48697 37843
rect 48783 37820 48849 37843
rect 48463 37780 48472 37820
rect 48512 37780 48529 37820
rect 48615 37780 48636 37820
rect 48676 37780 48697 37820
rect 48783 37780 48800 37820
rect 48840 37780 48849 37820
rect 48463 37757 48529 37780
rect 48615 37757 48697 37780
rect 48783 37757 48849 37780
rect 48463 37738 48849 37757
rect 63583 37843 63969 37862
rect 63583 37820 63649 37843
rect 63735 37820 63817 37843
rect 63903 37820 63969 37843
rect 63583 37780 63592 37820
rect 63632 37780 63649 37820
rect 63735 37780 63756 37820
rect 63796 37780 63817 37820
rect 63903 37780 63920 37820
rect 63960 37780 63969 37820
rect 63583 37757 63649 37780
rect 63735 37757 63817 37780
rect 63903 37757 63969 37780
rect 63583 37738 63969 37757
rect 78703 37843 79089 37862
rect 78703 37820 78769 37843
rect 78855 37820 78937 37843
rect 79023 37820 79089 37843
rect 78703 37780 78712 37820
rect 78752 37780 78769 37820
rect 78855 37780 78876 37820
rect 78916 37780 78937 37820
rect 79023 37780 79040 37820
rect 79080 37780 79089 37820
rect 78703 37757 78769 37780
rect 78855 37757 78937 37780
rect 79023 37757 79089 37780
rect 78703 37738 79089 37757
rect 4343 37087 4729 37106
rect 4343 37064 4409 37087
rect 4495 37064 4577 37087
rect 4663 37064 4729 37087
rect 4343 37024 4352 37064
rect 4392 37024 4409 37064
rect 4495 37024 4516 37064
rect 4556 37024 4577 37064
rect 4663 37024 4680 37064
rect 4720 37024 4729 37064
rect 4343 37001 4409 37024
rect 4495 37001 4577 37024
rect 4663 37001 4729 37024
rect 4343 36982 4729 37001
rect 19463 37087 19849 37106
rect 19463 37064 19529 37087
rect 19615 37064 19697 37087
rect 19783 37064 19849 37087
rect 19463 37024 19472 37064
rect 19512 37024 19529 37064
rect 19615 37024 19636 37064
rect 19676 37024 19697 37064
rect 19783 37024 19800 37064
rect 19840 37024 19849 37064
rect 19463 37001 19529 37024
rect 19615 37001 19697 37024
rect 19783 37001 19849 37024
rect 19463 36982 19849 37001
rect 34583 37087 34969 37106
rect 34583 37064 34649 37087
rect 34735 37064 34817 37087
rect 34903 37064 34969 37087
rect 34583 37024 34592 37064
rect 34632 37024 34649 37064
rect 34735 37024 34756 37064
rect 34796 37024 34817 37064
rect 34903 37024 34920 37064
rect 34960 37024 34969 37064
rect 34583 37001 34649 37024
rect 34735 37001 34817 37024
rect 34903 37001 34969 37024
rect 34583 36982 34969 37001
rect 49703 37087 50089 37106
rect 49703 37064 49769 37087
rect 49855 37064 49937 37087
rect 50023 37064 50089 37087
rect 49703 37024 49712 37064
rect 49752 37024 49769 37064
rect 49855 37024 49876 37064
rect 49916 37024 49937 37064
rect 50023 37024 50040 37064
rect 50080 37024 50089 37064
rect 49703 37001 49769 37024
rect 49855 37001 49937 37024
rect 50023 37001 50089 37024
rect 49703 36982 50089 37001
rect 64823 37087 65209 37106
rect 64823 37064 64889 37087
rect 64975 37064 65057 37087
rect 65143 37064 65209 37087
rect 64823 37024 64832 37064
rect 64872 37024 64889 37064
rect 64975 37024 64996 37064
rect 65036 37024 65057 37064
rect 65143 37024 65160 37064
rect 65200 37024 65209 37064
rect 64823 37001 64889 37024
rect 64975 37001 65057 37024
rect 65143 37001 65209 37024
rect 64823 36982 65209 37001
rect 79943 37087 80329 37106
rect 79943 37064 80009 37087
rect 80095 37064 80177 37087
rect 80263 37064 80329 37087
rect 79943 37024 79952 37064
rect 79992 37024 80009 37064
rect 80095 37024 80116 37064
rect 80156 37024 80177 37064
rect 80263 37024 80280 37064
rect 80320 37024 80329 37064
rect 79943 37001 80009 37024
rect 80095 37001 80177 37024
rect 80263 37001 80329 37024
rect 79943 36982 80329 37001
rect 3103 36331 3489 36350
rect 3103 36308 3169 36331
rect 3255 36308 3337 36331
rect 3423 36308 3489 36331
rect 3103 36268 3112 36308
rect 3152 36268 3169 36308
rect 3255 36268 3276 36308
rect 3316 36268 3337 36308
rect 3423 36268 3440 36308
rect 3480 36268 3489 36308
rect 3103 36245 3169 36268
rect 3255 36245 3337 36268
rect 3423 36245 3489 36268
rect 3103 36226 3489 36245
rect 18223 36331 18609 36350
rect 18223 36308 18289 36331
rect 18375 36308 18457 36331
rect 18543 36308 18609 36331
rect 18223 36268 18232 36308
rect 18272 36268 18289 36308
rect 18375 36268 18396 36308
rect 18436 36268 18457 36308
rect 18543 36268 18560 36308
rect 18600 36268 18609 36308
rect 18223 36245 18289 36268
rect 18375 36245 18457 36268
rect 18543 36245 18609 36268
rect 18223 36226 18609 36245
rect 33343 36331 33729 36350
rect 33343 36308 33409 36331
rect 33495 36308 33577 36331
rect 33663 36308 33729 36331
rect 33343 36268 33352 36308
rect 33392 36268 33409 36308
rect 33495 36268 33516 36308
rect 33556 36268 33577 36308
rect 33663 36268 33680 36308
rect 33720 36268 33729 36308
rect 33343 36245 33409 36268
rect 33495 36245 33577 36268
rect 33663 36245 33729 36268
rect 33343 36226 33729 36245
rect 48463 36331 48849 36350
rect 48463 36308 48529 36331
rect 48615 36308 48697 36331
rect 48783 36308 48849 36331
rect 48463 36268 48472 36308
rect 48512 36268 48529 36308
rect 48615 36268 48636 36308
rect 48676 36268 48697 36308
rect 48783 36268 48800 36308
rect 48840 36268 48849 36308
rect 48463 36245 48529 36268
rect 48615 36245 48697 36268
rect 48783 36245 48849 36268
rect 48463 36226 48849 36245
rect 63583 36331 63969 36350
rect 63583 36308 63649 36331
rect 63735 36308 63817 36331
rect 63903 36308 63969 36331
rect 63583 36268 63592 36308
rect 63632 36268 63649 36308
rect 63735 36268 63756 36308
rect 63796 36268 63817 36308
rect 63903 36268 63920 36308
rect 63960 36268 63969 36308
rect 63583 36245 63649 36268
rect 63735 36245 63817 36268
rect 63903 36245 63969 36268
rect 63583 36226 63969 36245
rect 78703 36331 79089 36350
rect 78703 36308 78769 36331
rect 78855 36308 78937 36331
rect 79023 36308 79089 36331
rect 78703 36268 78712 36308
rect 78752 36268 78769 36308
rect 78855 36268 78876 36308
rect 78916 36268 78937 36308
rect 79023 36268 79040 36308
rect 79080 36268 79089 36308
rect 78703 36245 78769 36268
rect 78855 36245 78937 36268
rect 79023 36245 79089 36268
rect 78703 36226 79089 36245
rect 4343 35575 4729 35594
rect 4343 35552 4409 35575
rect 4495 35552 4577 35575
rect 4663 35552 4729 35575
rect 4343 35512 4352 35552
rect 4392 35512 4409 35552
rect 4495 35512 4516 35552
rect 4556 35512 4577 35552
rect 4663 35512 4680 35552
rect 4720 35512 4729 35552
rect 4343 35489 4409 35512
rect 4495 35489 4577 35512
rect 4663 35489 4729 35512
rect 4343 35470 4729 35489
rect 19463 35575 19849 35594
rect 19463 35552 19529 35575
rect 19615 35552 19697 35575
rect 19783 35552 19849 35575
rect 19463 35512 19472 35552
rect 19512 35512 19529 35552
rect 19615 35512 19636 35552
rect 19676 35512 19697 35552
rect 19783 35512 19800 35552
rect 19840 35512 19849 35552
rect 19463 35489 19529 35512
rect 19615 35489 19697 35512
rect 19783 35489 19849 35512
rect 19463 35470 19849 35489
rect 34583 35575 34969 35594
rect 34583 35552 34649 35575
rect 34735 35552 34817 35575
rect 34903 35552 34969 35575
rect 34583 35512 34592 35552
rect 34632 35512 34649 35552
rect 34735 35512 34756 35552
rect 34796 35512 34817 35552
rect 34903 35512 34920 35552
rect 34960 35512 34969 35552
rect 34583 35489 34649 35512
rect 34735 35489 34817 35512
rect 34903 35489 34969 35512
rect 34583 35470 34969 35489
rect 49703 35575 50089 35594
rect 49703 35552 49769 35575
rect 49855 35552 49937 35575
rect 50023 35552 50089 35575
rect 49703 35512 49712 35552
rect 49752 35512 49769 35552
rect 49855 35512 49876 35552
rect 49916 35512 49937 35552
rect 50023 35512 50040 35552
rect 50080 35512 50089 35552
rect 49703 35489 49769 35512
rect 49855 35489 49937 35512
rect 50023 35489 50089 35512
rect 49703 35470 50089 35489
rect 64823 35575 65209 35594
rect 64823 35552 64889 35575
rect 64975 35552 65057 35575
rect 65143 35552 65209 35575
rect 64823 35512 64832 35552
rect 64872 35512 64889 35552
rect 64975 35512 64996 35552
rect 65036 35512 65057 35552
rect 65143 35512 65160 35552
rect 65200 35512 65209 35552
rect 64823 35489 64889 35512
rect 64975 35489 65057 35512
rect 65143 35489 65209 35512
rect 64823 35470 65209 35489
rect 79943 35575 80329 35594
rect 79943 35552 80009 35575
rect 80095 35552 80177 35575
rect 80263 35552 80329 35575
rect 79943 35512 79952 35552
rect 79992 35512 80009 35552
rect 80095 35512 80116 35552
rect 80156 35512 80177 35552
rect 80263 35512 80280 35552
rect 80320 35512 80329 35552
rect 79943 35489 80009 35512
rect 80095 35489 80177 35512
rect 80263 35489 80329 35512
rect 79943 35470 80329 35489
rect 3103 34819 3489 34838
rect 3103 34796 3169 34819
rect 3255 34796 3337 34819
rect 3423 34796 3489 34819
rect 3103 34756 3112 34796
rect 3152 34756 3169 34796
rect 3255 34756 3276 34796
rect 3316 34756 3337 34796
rect 3423 34756 3440 34796
rect 3480 34756 3489 34796
rect 3103 34733 3169 34756
rect 3255 34733 3337 34756
rect 3423 34733 3489 34756
rect 3103 34714 3489 34733
rect 18223 34819 18609 34838
rect 18223 34796 18289 34819
rect 18375 34796 18457 34819
rect 18543 34796 18609 34819
rect 18223 34756 18232 34796
rect 18272 34756 18289 34796
rect 18375 34756 18396 34796
rect 18436 34756 18457 34796
rect 18543 34756 18560 34796
rect 18600 34756 18609 34796
rect 18223 34733 18289 34756
rect 18375 34733 18457 34756
rect 18543 34733 18609 34756
rect 18223 34714 18609 34733
rect 33343 34819 33729 34838
rect 33343 34796 33409 34819
rect 33495 34796 33577 34819
rect 33663 34796 33729 34819
rect 33343 34756 33352 34796
rect 33392 34756 33409 34796
rect 33495 34756 33516 34796
rect 33556 34756 33577 34796
rect 33663 34756 33680 34796
rect 33720 34756 33729 34796
rect 33343 34733 33409 34756
rect 33495 34733 33577 34756
rect 33663 34733 33729 34756
rect 33343 34714 33729 34733
rect 48463 34819 48849 34838
rect 48463 34796 48529 34819
rect 48615 34796 48697 34819
rect 48783 34796 48849 34819
rect 48463 34756 48472 34796
rect 48512 34756 48529 34796
rect 48615 34756 48636 34796
rect 48676 34756 48697 34796
rect 48783 34756 48800 34796
rect 48840 34756 48849 34796
rect 48463 34733 48529 34756
rect 48615 34733 48697 34756
rect 48783 34733 48849 34756
rect 48463 34714 48849 34733
rect 63583 34819 63969 34838
rect 63583 34796 63649 34819
rect 63735 34796 63817 34819
rect 63903 34796 63969 34819
rect 63583 34756 63592 34796
rect 63632 34756 63649 34796
rect 63735 34756 63756 34796
rect 63796 34756 63817 34796
rect 63903 34756 63920 34796
rect 63960 34756 63969 34796
rect 63583 34733 63649 34756
rect 63735 34733 63817 34756
rect 63903 34733 63969 34756
rect 63583 34714 63969 34733
rect 78703 34819 79089 34838
rect 78703 34796 78769 34819
rect 78855 34796 78937 34819
rect 79023 34796 79089 34819
rect 78703 34756 78712 34796
rect 78752 34756 78769 34796
rect 78855 34756 78876 34796
rect 78916 34756 78937 34796
rect 79023 34756 79040 34796
rect 79080 34756 79089 34796
rect 78703 34733 78769 34756
rect 78855 34733 78937 34756
rect 79023 34733 79089 34756
rect 78703 34714 79089 34733
rect 4343 34063 4729 34082
rect 4343 34040 4409 34063
rect 4495 34040 4577 34063
rect 4663 34040 4729 34063
rect 4343 34000 4352 34040
rect 4392 34000 4409 34040
rect 4495 34000 4516 34040
rect 4556 34000 4577 34040
rect 4663 34000 4680 34040
rect 4720 34000 4729 34040
rect 4343 33977 4409 34000
rect 4495 33977 4577 34000
rect 4663 33977 4729 34000
rect 4343 33958 4729 33977
rect 19463 34063 19849 34082
rect 19463 34040 19529 34063
rect 19615 34040 19697 34063
rect 19783 34040 19849 34063
rect 19463 34000 19472 34040
rect 19512 34000 19529 34040
rect 19615 34000 19636 34040
rect 19676 34000 19697 34040
rect 19783 34000 19800 34040
rect 19840 34000 19849 34040
rect 19463 33977 19529 34000
rect 19615 33977 19697 34000
rect 19783 33977 19849 34000
rect 19463 33958 19849 33977
rect 34583 34063 34969 34082
rect 34583 34040 34649 34063
rect 34735 34040 34817 34063
rect 34903 34040 34969 34063
rect 34583 34000 34592 34040
rect 34632 34000 34649 34040
rect 34735 34000 34756 34040
rect 34796 34000 34817 34040
rect 34903 34000 34920 34040
rect 34960 34000 34969 34040
rect 34583 33977 34649 34000
rect 34735 33977 34817 34000
rect 34903 33977 34969 34000
rect 34583 33958 34969 33977
rect 49703 34063 50089 34082
rect 49703 34040 49769 34063
rect 49855 34040 49937 34063
rect 50023 34040 50089 34063
rect 49703 34000 49712 34040
rect 49752 34000 49769 34040
rect 49855 34000 49876 34040
rect 49916 34000 49937 34040
rect 50023 34000 50040 34040
rect 50080 34000 50089 34040
rect 49703 33977 49769 34000
rect 49855 33977 49937 34000
rect 50023 33977 50089 34000
rect 49703 33958 50089 33977
rect 64823 34063 65209 34082
rect 64823 34040 64889 34063
rect 64975 34040 65057 34063
rect 65143 34040 65209 34063
rect 64823 34000 64832 34040
rect 64872 34000 64889 34040
rect 64975 34000 64996 34040
rect 65036 34000 65057 34040
rect 65143 34000 65160 34040
rect 65200 34000 65209 34040
rect 64823 33977 64889 34000
rect 64975 33977 65057 34000
rect 65143 33977 65209 34000
rect 64823 33958 65209 33977
rect 79943 34063 80329 34082
rect 79943 34040 80009 34063
rect 80095 34040 80177 34063
rect 80263 34040 80329 34063
rect 79943 34000 79952 34040
rect 79992 34000 80009 34040
rect 80095 34000 80116 34040
rect 80156 34000 80177 34040
rect 80263 34000 80280 34040
rect 80320 34000 80329 34040
rect 79943 33977 80009 34000
rect 80095 33977 80177 34000
rect 80263 33977 80329 34000
rect 79943 33958 80329 33977
rect 3103 33307 3489 33326
rect 3103 33284 3169 33307
rect 3255 33284 3337 33307
rect 3423 33284 3489 33307
rect 3103 33244 3112 33284
rect 3152 33244 3169 33284
rect 3255 33244 3276 33284
rect 3316 33244 3337 33284
rect 3423 33244 3440 33284
rect 3480 33244 3489 33284
rect 3103 33221 3169 33244
rect 3255 33221 3337 33244
rect 3423 33221 3489 33244
rect 3103 33202 3489 33221
rect 18223 33307 18609 33326
rect 18223 33284 18289 33307
rect 18375 33284 18457 33307
rect 18543 33284 18609 33307
rect 18223 33244 18232 33284
rect 18272 33244 18289 33284
rect 18375 33244 18396 33284
rect 18436 33244 18457 33284
rect 18543 33244 18560 33284
rect 18600 33244 18609 33284
rect 18223 33221 18289 33244
rect 18375 33221 18457 33244
rect 18543 33221 18609 33244
rect 18223 33202 18609 33221
rect 33343 33307 33729 33326
rect 33343 33284 33409 33307
rect 33495 33284 33577 33307
rect 33663 33284 33729 33307
rect 33343 33244 33352 33284
rect 33392 33244 33409 33284
rect 33495 33244 33516 33284
rect 33556 33244 33577 33284
rect 33663 33244 33680 33284
rect 33720 33244 33729 33284
rect 33343 33221 33409 33244
rect 33495 33221 33577 33244
rect 33663 33221 33729 33244
rect 33343 33202 33729 33221
rect 48463 33307 48849 33326
rect 48463 33284 48529 33307
rect 48615 33284 48697 33307
rect 48783 33284 48849 33307
rect 48463 33244 48472 33284
rect 48512 33244 48529 33284
rect 48615 33244 48636 33284
rect 48676 33244 48697 33284
rect 48783 33244 48800 33284
rect 48840 33244 48849 33284
rect 48463 33221 48529 33244
rect 48615 33221 48697 33244
rect 48783 33221 48849 33244
rect 48463 33202 48849 33221
rect 63583 33307 63969 33326
rect 63583 33284 63649 33307
rect 63735 33284 63817 33307
rect 63903 33284 63969 33307
rect 63583 33244 63592 33284
rect 63632 33244 63649 33284
rect 63735 33244 63756 33284
rect 63796 33244 63817 33284
rect 63903 33244 63920 33284
rect 63960 33244 63969 33284
rect 63583 33221 63649 33244
rect 63735 33221 63817 33244
rect 63903 33221 63969 33244
rect 63583 33202 63969 33221
rect 78703 33307 79089 33326
rect 78703 33284 78769 33307
rect 78855 33284 78937 33307
rect 79023 33284 79089 33307
rect 78703 33244 78712 33284
rect 78752 33244 78769 33284
rect 78855 33244 78876 33284
rect 78916 33244 78937 33284
rect 79023 33244 79040 33284
rect 79080 33244 79089 33284
rect 78703 33221 78769 33244
rect 78855 33221 78937 33244
rect 79023 33221 79089 33244
rect 78703 33202 79089 33221
rect 4343 32551 4729 32570
rect 4343 32528 4409 32551
rect 4495 32528 4577 32551
rect 4663 32528 4729 32551
rect 4343 32488 4352 32528
rect 4392 32488 4409 32528
rect 4495 32488 4516 32528
rect 4556 32488 4577 32528
rect 4663 32488 4680 32528
rect 4720 32488 4729 32528
rect 4343 32465 4409 32488
rect 4495 32465 4577 32488
rect 4663 32465 4729 32488
rect 4343 32446 4729 32465
rect 19463 32551 19849 32570
rect 19463 32528 19529 32551
rect 19615 32528 19697 32551
rect 19783 32528 19849 32551
rect 19463 32488 19472 32528
rect 19512 32488 19529 32528
rect 19615 32488 19636 32528
rect 19676 32488 19697 32528
rect 19783 32488 19800 32528
rect 19840 32488 19849 32528
rect 19463 32465 19529 32488
rect 19615 32465 19697 32488
rect 19783 32465 19849 32488
rect 19463 32446 19849 32465
rect 34583 32551 34969 32570
rect 34583 32528 34649 32551
rect 34735 32528 34817 32551
rect 34903 32528 34969 32551
rect 34583 32488 34592 32528
rect 34632 32488 34649 32528
rect 34735 32488 34756 32528
rect 34796 32488 34817 32528
rect 34903 32488 34920 32528
rect 34960 32488 34969 32528
rect 34583 32465 34649 32488
rect 34735 32465 34817 32488
rect 34903 32465 34969 32488
rect 34583 32446 34969 32465
rect 49703 32551 50089 32570
rect 49703 32528 49769 32551
rect 49855 32528 49937 32551
rect 50023 32528 50089 32551
rect 49703 32488 49712 32528
rect 49752 32488 49769 32528
rect 49855 32488 49876 32528
rect 49916 32488 49937 32528
rect 50023 32488 50040 32528
rect 50080 32488 50089 32528
rect 49703 32465 49769 32488
rect 49855 32465 49937 32488
rect 50023 32465 50089 32488
rect 49703 32446 50089 32465
rect 64823 32551 65209 32570
rect 64823 32528 64889 32551
rect 64975 32528 65057 32551
rect 65143 32528 65209 32551
rect 64823 32488 64832 32528
rect 64872 32488 64889 32528
rect 64975 32488 64996 32528
rect 65036 32488 65057 32528
rect 65143 32488 65160 32528
rect 65200 32488 65209 32528
rect 64823 32465 64889 32488
rect 64975 32465 65057 32488
rect 65143 32465 65209 32488
rect 64823 32446 65209 32465
rect 79943 32551 80329 32570
rect 79943 32528 80009 32551
rect 80095 32528 80177 32551
rect 80263 32528 80329 32551
rect 79943 32488 79952 32528
rect 79992 32488 80009 32528
rect 80095 32488 80116 32528
rect 80156 32488 80177 32528
rect 80263 32488 80280 32528
rect 80320 32488 80329 32528
rect 79943 32465 80009 32488
rect 80095 32465 80177 32488
rect 80263 32465 80329 32488
rect 79943 32446 80329 32465
rect 3103 31795 3489 31814
rect 3103 31772 3169 31795
rect 3255 31772 3337 31795
rect 3423 31772 3489 31795
rect 3103 31732 3112 31772
rect 3152 31732 3169 31772
rect 3255 31732 3276 31772
rect 3316 31732 3337 31772
rect 3423 31732 3440 31772
rect 3480 31732 3489 31772
rect 3103 31709 3169 31732
rect 3255 31709 3337 31732
rect 3423 31709 3489 31732
rect 3103 31690 3489 31709
rect 18223 31795 18609 31814
rect 18223 31772 18289 31795
rect 18375 31772 18457 31795
rect 18543 31772 18609 31795
rect 18223 31732 18232 31772
rect 18272 31732 18289 31772
rect 18375 31732 18396 31772
rect 18436 31732 18457 31772
rect 18543 31732 18560 31772
rect 18600 31732 18609 31772
rect 18223 31709 18289 31732
rect 18375 31709 18457 31732
rect 18543 31709 18609 31732
rect 18223 31690 18609 31709
rect 33343 31795 33729 31814
rect 33343 31772 33409 31795
rect 33495 31772 33577 31795
rect 33663 31772 33729 31795
rect 33343 31732 33352 31772
rect 33392 31732 33409 31772
rect 33495 31732 33516 31772
rect 33556 31732 33577 31772
rect 33663 31732 33680 31772
rect 33720 31732 33729 31772
rect 33343 31709 33409 31732
rect 33495 31709 33577 31732
rect 33663 31709 33729 31732
rect 33343 31690 33729 31709
rect 48463 31795 48849 31814
rect 48463 31772 48529 31795
rect 48615 31772 48697 31795
rect 48783 31772 48849 31795
rect 48463 31732 48472 31772
rect 48512 31732 48529 31772
rect 48615 31732 48636 31772
rect 48676 31732 48697 31772
rect 48783 31732 48800 31772
rect 48840 31732 48849 31772
rect 48463 31709 48529 31732
rect 48615 31709 48697 31732
rect 48783 31709 48849 31732
rect 48463 31690 48849 31709
rect 63583 31795 63969 31814
rect 63583 31772 63649 31795
rect 63735 31772 63817 31795
rect 63903 31772 63969 31795
rect 63583 31732 63592 31772
rect 63632 31732 63649 31772
rect 63735 31732 63756 31772
rect 63796 31732 63817 31772
rect 63903 31732 63920 31772
rect 63960 31732 63969 31772
rect 63583 31709 63649 31732
rect 63735 31709 63817 31732
rect 63903 31709 63969 31732
rect 63583 31690 63969 31709
rect 78703 31795 79089 31814
rect 78703 31772 78769 31795
rect 78855 31772 78937 31795
rect 79023 31772 79089 31795
rect 78703 31732 78712 31772
rect 78752 31732 78769 31772
rect 78855 31732 78876 31772
rect 78916 31732 78937 31772
rect 79023 31732 79040 31772
rect 79080 31732 79089 31772
rect 78703 31709 78769 31732
rect 78855 31709 78937 31732
rect 79023 31709 79089 31732
rect 78703 31690 79089 31709
rect 4343 31039 4729 31058
rect 4343 31016 4409 31039
rect 4495 31016 4577 31039
rect 4663 31016 4729 31039
rect 4343 30976 4352 31016
rect 4392 30976 4409 31016
rect 4495 30976 4516 31016
rect 4556 30976 4577 31016
rect 4663 30976 4680 31016
rect 4720 30976 4729 31016
rect 4343 30953 4409 30976
rect 4495 30953 4577 30976
rect 4663 30953 4729 30976
rect 4343 30934 4729 30953
rect 19463 31039 19849 31058
rect 19463 31016 19529 31039
rect 19615 31016 19697 31039
rect 19783 31016 19849 31039
rect 19463 30976 19472 31016
rect 19512 30976 19529 31016
rect 19615 30976 19636 31016
rect 19676 30976 19697 31016
rect 19783 30976 19800 31016
rect 19840 30976 19849 31016
rect 19463 30953 19529 30976
rect 19615 30953 19697 30976
rect 19783 30953 19849 30976
rect 19463 30934 19849 30953
rect 34583 31039 34969 31058
rect 34583 31016 34649 31039
rect 34735 31016 34817 31039
rect 34903 31016 34969 31039
rect 34583 30976 34592 31016
rect 34632 30976 34649 31016
rect 34735 30976 34756 31016
rect 34796 30976 34817 31016
rect 34903 30976 34920 31016
rect 34960 30976 34969 31016
rect 34583 30953 34649 30976
rect 34735 30953 34817 30976
rect 34903 30953 34969 30976
rect 34583 30934 34969 30953
rect 49703 31039 50089 31058
rect 49703 31016 49769 31039
rect 49855 31016 49937 31039
rect 50023 31016 50089 31039
rect 49703 30976 49712 31016
rect 49752 30976 49769 31016
rect 49855 30976 49876 31016
rect 49916 30976 49937 31016
rect 50023 30976 50040 31016
rect 50080 30976 50089 31016
rect 49703 30953 49769 30976
rect 49855 30953 49937 30976
rect 50023 30953 50089 30976
rect 49703 30934 50089 30953
rect 64823 31039 65209 31058
rect 64823 31016 64889 31039
rect 64975 31016 65057 31039
rect 65143 31016 65209 31039
rect 64823 30976 64832 31016
rect 64872 30976 64889 31016
rect 64975 30976 64996 31016
rect 65036 30976 65057 31016
rect 65143 30976 65160 31016
rect 65200 30976 65209 31016
rect 64823 30953 64889 30976
rect 64975 30953 65057 30976
rect 65143 30953 65209 30976
rect 64823 30934 65209 30953
rect 79943 31039 80329 31058
rect 79943 31016 80009 31039
rect 80095 31016 80177 31039
rect 80263 31016 80329 31039
rect 79943 30976 79952 31016
rect 79992 30976 80009 31016
rect 80095 30976 80116 31016
rect 80156 30976 80177 31016
rect 80263 30976 80280 31016
rect 80320 30976 80329 31016
rect 79943 30953 80009 30976
rect 80095 30953 80177 30976
rect 80263 30953 80329 30976
rect 79943 30934 80329 30953
rect 3103 30283 3489 30302
rect 3103 30260 3169 30283
rect 3255 30260 3337 30283
rect 3423 30260 3489 30283
rect 3103 30220 3112 30260
rect 3152 30220 3169 30260
rect 3255 30220 3276 30260
rect 3316 30220 3337 30260
rect 3423 30220 3440 30260
rect 3480 30220 3489 30260
rect 3103 30197 3169 30220
rect 3255 30197 3337 30220
rect 3423 30197 3489 30220
rect 3103 30178 3489 30197
rect 18223 30283 18609 30302
rect 18223 30260 18289 30283
rect 18375 30260 18457 30283
rect 18543 30260 18609 30283
rect 18223 30220 18232 30260
rect 18272 30220 18289 30260
rect 18375 30220 18396 30260
rect 18436 30220 18457 30260
rect 18543 30220 18560 30260
rect 18600 30220 18609 30260
rect 18223 30197 18289 30220
rect 18375 30197 18457 30220
rect 18543 30197 18609 30220
rect 18223 30178 18609 30197
rect 33343 30283 33729 30302
rect 33343 30260 33409 30283
rect 33495 30260 33577 30283
rect 33663 30260 33729 30283
rect 33343 30220 33352 30260
rect 33392 30220 33409 30260
rect 33495 30220 33516 30260
rect 33556 30220 33577 30260
rect 33663 30220 33680 30260
rect 33720 30220 33729 30260
rect 33343 30197 33409 30220
rect 33495 30197 33577 30220
rect 33663 30197 33729 30220
rect 33343 30178 33729 30197
rect 48463 30283 48849 30302
rect 48463 30260 48529 30283
rect 48615 30260 48697 30283
rect 48783 30260 48849 30283
rect 48463 30220 48472 30260
rect 48512 30220 48529 30260
rect 48615 30220 48636 30260
rect 48676 30220 48697 30260
rect 48783 30220 48800 30260
rect 48840 30220 48849 30260
rect 48463 30197 48529 30220
rect 48615 30197 48697 30220
rect 48783 30197 48849 30220
rect 48463 30178 48849 30197
rect 63583 30283 63969 30302
rect 63583 30260 63649 30283
rect 63735 30260 63817 30283
rect 63903 30260 63969 30283
rect 63583 30220 63592 30260
rect 63632 30220 63649 30260
rect 63735 30220 63756 30260
rect 63796 30220 63817 30260
rect 63903 30220 63920 30260
rect 63960 30220 63969 30260
rect 63583 30197 63649 30220
rect 63735 30197 63817 30220
rect 63903 30197 63969 30220
rect 63583 30178 63969 30197
rect 78703 30283 79089 30302
rect 78703 30260 78769 30283
rect 78855 30260 78937 30283
rect 79023 30260 79089 30283
rect 78703 30220 78712 30260
rect 78752 30220 78769 30260
rect 78855 30220 78876 30260
rect 78916 30220 78937 30260
rect 79023 30220 79040 30260
rect 79080 30220 79089 30260
rect 78703 30197 78769 30220
rect 78855 30197 78937 30220
rect 79023 30197 79089 30220
rect 78703 30178 79089 30197
rect 4343 29527 4729 29546
rect 4343 29504 4409 29527
rect 4495 29504 4577 29527
rect 4663 29504 4729 29527
rect 4343 29464 4352 29504
rect 4392 29464 4409 29504
rect 4495 29464 4516 29504
rect 4556 29464 4577 29504
rect 4663 29464 4680 29504
rect 4720 29464 4729 29504
rect 4343 29441 4409 29464
rect 4495 29441 4577 29464
rect 4663 29441 4729 29464
rect 4343 29422 4729 29441
rect 19463 29527 19849 29546
rect 19463 29504 19529 29527
rect 19615 29504 19697 29527
rect 19783 29504 19849 29527
rect 19463 29464 19472 29504
rect 19512 29464 19529 29504
rect 19615 29464 19636 29504
rect 19676 29464 19697 29504
rect 19783 29464 19800 29504
rect 19840 29464 19849 29504
rect 19463 29441 19529 29464
rect 19615 29441 19697 29464
rect 19783 29441 19849 29464
rect 19463 29422 19849 29441
rect 34583 29527 34969 29546
rect 34583 29504 34649 29527
rect 34735 29504 34817 29527
rect 34903 29504 34969 29527
rect 34583 29464 34592 29504
rect 34632 29464 34649 29504
rect 34735 29464 34756 29504
rect 34796 29464 34817 29504
rect 34903 29464 34920 29504
rect 34960 29464 34969 29504
rect 34583 29441 34649 29464
rect 34735 29441 34817 29464
rect 34903 29441 34969 29464
rect 34583 29422 34969 29441
rect 49703 29527 50089 29546
rect 49703 29504 49769 29527
rect 49855 29504 49937 29527
rect 50023 29504 50089 29527
rect 49703 29464 49712 29504
rect 49752 29464 49769 29504
rect 49855 29464 49876 29504
rect 49916 29464 49937 29504
rect 50023 29464 50040 29504
rect 50080 29464 50089 29504
rect 49703 29441 49769 29464
rect 49855 29441 49937 29464
rect 50023 29441 50089 29464
rect 49703 29422 50089 29441
rect 64823 29527 65209 29546
rect 64823 29504 64889 29527
rect 64975 29504 65057 29527
rect 65143 29504 65209 29527
rect 64823 29464 64832 29504
rect 64872 29464 64889 29504
rect 64975 29464 64996 29504
rect 65036 29464 65057 29504
rect 65143 29464 65160 29504
rect 65200 29464 65209 29504
rect 64823 29441 64889 29464
rect 64975 29441 65057 29464
rect 65143 29441 65209 29464
rect 64823 29422 65209 29441
rect 79943 29527 80329 29546
rect 79943 29504 80009 29527
rect 80095 29504 80177 29527
rect 80263 29504 80329 29527
rect 79943 29464 79952 29504
rect 79992 29464 80009 29504
rect 80095 29464 80116 29504
rect 80156 29464 80177 29504
rect 80263 29464 80280 29504
rect 80320 29464 80329 29504
rect 79943 29441 80009 29464
rect 80095 29441 80177 29464
rect 80263 29441 80329 29464
rect 79943 29422 80329 29441
rect 3103 28771 3489 28790
rect 3103 28748 3169 28771
rect 3255 28748 3337 28771
rect 3423 28748 3489 28771
rect 3103 28708 3112 28748
rect 3152 28708 3169 28748
rect 3255 28708 3276 28748
rect 3316 28708 3337 28748
rect 3423 28708 3440 28748
rect 3480 28708 3489 28748
rect 3103 28685 3169 28708
rect 3255 28685 3337 28708
rect 3423 28685 3489 28708
rect 3103 28666 3489 28685
rect 18223 28771 18609 28790
rect 18223 28748 18289 28771
rect 18375 28748 18457 28771
rect 18543 28748 18609 28771
rect 18223 28708 18232 28748
rect 18272 28708 18289 28748
rect 18375 28708 18396 28748
rect 18436 28708 18457 28748
rect 18543 28708 18560 28748
rect 18600 28708 18609 28748
rect 18223 28685 18289 28708
rect 18375 28685 18457 28708
rect 18543 28685 18609 28708
rect 18223 28666 18609 28685
rect 33343 28771 33729 28790
rect 33343 28748 33409 28771
rect 33495 28748 33577 28771
rect 33663 28748 33729 28771
rect 33343 28708 33352 28748
rect 33392 28708 33409 28748
rect 33495 28708 33516 28748
rect 33556 28708 33577 28748
rect 33663 28708 33680 28748
rect 33720 28708 33729 28748
rect 33343 28685 33409 28708
rect 33495 28685 33577 28708
rect 33663 28685 33729 28708
rect 33343 28666 33729 28685
rect 48463 28771 48849 28790
rect 48463 28748 48529 28771
rect 48615 28748 48697 28771
rect 48783 28748 48849 28771
rect 48463 28708 48472 28748
rect 48512 28708 48529 28748
rect 48615 28708 48636 28748
rect 48676 28708 48697 28748
rect 48783 28708 48800 28748
rect 48840 28708 48849 28748
rect 48463 28685 48529 28708
rect 48615 28685 48697 28708
rect 48783 28685 48849 28708
rect 48463 28666 48849 28685
rect 63583 28771 63969 28790
rect 63583 28748 63649 28771
rect 63735 28748 63817 28771
rect 63903 28748 63969 28771
rect 63583 28708 63592 28748
rect 63632 28708 63649 28748
rect 63735 28708 63756 28748
rect 63796 28708 63817 28748
rect 63903 28708 63920 28748
rect 63960 28708 63969 28748
rect 63583 28685 63649 28708
rect 63735 28685 63817 28708
rect 63903 28685 63969 28708
rect 63583 28666 63969 28685
rect 78703 28771 79089 28790
rect 78703 28748 78769 28771
rect 78855 28748 78937 28771
rect 79023 28748 79089 28771
rect 78703 28708 78712 28748
rect 78752 28708 78769 28748
rect 78855 28708 78876 28748
rect 78916 28708 78937 28748
rect 79023 28708 79040 28748
rect 79080 28708 79089 28748
rect 78703 28685 78769 28708
rect 78855 28685 78937 28708
rect 79023 28685 79089 28708
rect 78703 28666 79089 28685
rect 4343 28015 4729 28034
rect 4343 27992 4409 28015
rect 4495 27992 4577 28015
rect 4663 27992 4729 28015
rect 4343 27952 4352 27992
rect 4392 27952 4409 27992
rect 4495 27952 4516 27992
rect 4556 27952 4577 27992
rect 4663 27952 4680 27992
rect 4720 27952 4729 27992
rect 4343 27929 4409 27952
rect 4495 27929 4577 27952
rect 4663 27929 4729 27952
rect 4343 27910 4729 27929
rect 19463 28015 19849 28034
rect 19463 27992 19529 28015
rect 19615 27992 19697 28015
rect 19783 27992 19849 28015
rect 19463 27952 19472 27992
rect 19512 27952 19529 27992
rect 19615 27952 19636 27992
rect 19676 27952 19697 27992
rect 19783 27952 19800 27992
rect 19840 27952 19849 27992
rect 19463 27929 19529 27952
rect 19615 27929 19697 27952
rect 19783 27929 19849 27952
rect 19463 27910 19849 27929
rect 34583 28015 34969 28034
rect 34583 27992 34649 28015
rect 34735 27992 34817 28015
rect 34903 27992 34969 28015
rect 34583 27952 34592 27992
rect 34632 27952 34649 27992
rect 34735 27952 34756 27992
rect 34796 27952 34817 27992
rect 34903 27952 34920 27992
rect 34960 27952 34969 27992
rect 34583 27929 34649 27952
rect 34735 27929 34817 27952
rect 34903 27929 34969 27952
rect 34583 27910 34969 27929
rect 49703 28015 50089 28034
rect 49703 27992 49769 28015
rect 49855 27992 49937 28015
rect 50023 27992 50089 28015
rect 49703 27952 49712 27992
rect 49752 27952 49769 27992
rect 49855 27952 49876 27992
rect 49916 27952 49937 27992
rect 50023 27952 50040 27992
rect 50080 27952 50089 27992
rect 49703 27929 49769 27952
rect 49855 27929 49937 27952
rect 50023 27929 50089 27952
rect 49703 27910 50089 27929
rect 64823 28015 65209 28034
rect 64823 27992 64889 28015
rect 64975 27992 65057 28015
rect 65143 27992 65209 28015
rect 64823 27952 64832 27992
rect 64872 27952 64889 27992
rect 64975 27952 64996 27992
rect 65036 27952 65057 27992
rect 65143 27952 65160 27992
rect 65200 27952 65209 27992
rect 64823 27929 64889 27952
rect 64975 27929 65057 27952
rect 65143 27929 65209 27952
rect 64823 27910 65209 27929
rect 79943 28015 80329 28034
rect 79943 27992 80009 28015
rect 80095 27992 80177 28015
rect 80263 27992 80329 28015
rect 79943 27952 79952 27992
rect 79992 27952 80009 27992
rect 80095 27952 80116 27992
rect 80156 27952 80177 27992
rect 80263 27952 80280 27992
rect 80320 27952 80329 27992
rect 79943 27929 80009 27952
rect 80095 27929 80177 27952
rect 80263 27929 80329 27952
rect 79943 27910 80329 27929
rect 3103 27259 3489 27278
rect 3103 27236 3169 27259
rect 3255 27236 3337 27259
rect 3423 27236 3489 27259
rect 3103 27196 3112 27236
rect 3152 27196 3169 27236
rect 3255 27196 3276 27236
rect 3316 27196 3337 27236
rect 3423 27196 3440 27236
rect 3480 27196 3489 27236
rect 3103 27173 3169 27196
rect 3255 27173 3337 27196
rect 3423 27173 3489 27196
rect 3103 27154 3489 27173
rect 18223 27259 18609 27278
rect 18223 27236 18289 27259
rect 18375 27236 18457 27259
rect 18543 27236 18609 27259
rect 18223 27196 18232 27236
rect 18272 27196 18289 27236
rect 18375 27196 18396 27236
rect 18436 27196 18457 27236
rect 18543 27196 18560 27236
rect 18600 27196 18609 27236
rect 18223 27173 18289 27196
rect 18375 27173 18457 27196
rect 18543 27173 18609 27196
rect 18223 27154 18609 27173
rect 33343 27259 33729 27278
rect 33343 27236 33409 27259
rect 33495 27236 33577 27259
rect 33663 27236 33729 27259
rect 33343 27196 33352 27236
rect 33392 27196 33409 27236
rect 33495 27196 33516 27236
rect 33556 27196 33577 27236
rect 33663 27196 33680 27236
rect 33720 27196 33729 27236
rect 33343 27173 33409 27196
rect 33495 27173 33577 27196
rect 33663 27173 33729 27196
rect 33343 27154 33729 27173
rect 48463 27259 48849 27278
rect 48463 27236 48529 27259
rect 48615 27236 48697 27259
rect 48783 27236 48849 27259
rect 48463 27196 48472 27236
rect 48512 27196 48529 27236
rect 48615 27196 48636 27236
rect 48676 27196 48697 27236
rect 48783 27196 48800 27236
rect 48840 27196 48849 27236
rect 48463 27173 48529 27196
rect 48615 27173 48697 27196
rect 48783 27173 48849 27196
rect 48463 27154 48849 27173
rect 63583 27259 63969 27278
rect 63583 27236 63649 27259
rect 63735 27236 63817 27259
rect 63903 27236 63969 27259
rect 63583 27196 63592 27236
rect 63632 27196 63649 27236
rect 63735 27196 63756 27236
rect 63796 27196 63817 27236
rect 63903 27196 63920 27236
rect 63960 27196 63969 27236
rect 63583 27173 63649 27196
rect 63735 27173 63817 27196
rect 63903 27173 63969 27196
rect 63583 27154 63969 27173
rect 78703 27259 79089 27278
rect 78703 27236 78769 27259
rect 78855 27236 78937 27259
rect 79023 27236 79089 27259
rect 78703 27196 78712 27236
rect 78752 27196 78769 27236
rect 78855 27196 78876 27236
rect 78916 27196 78937 27236
rect 79023 27196 79040 27236
rect 79080 27196 79089 27236
rect 78703 27173 78769 27196
rect 78855 27173 78937 27196
rect 79023 27173 79089 27196
rect 78703 27154 79089 27173
rect 4343 26503 4729 26522
rect 4343 26480 4409 26503
rect 4495 26480 4577 26503
rect 4663 26480 4729 26503
rect 4343 26440 4352 26480
rect 4392 26440 4409 26480
rect 4495 26440 4516 26480
rect 4556 26440 4577 26480
rect 4663 26440 4680 26480
rect 4720 26440 4729 26480
rect 4343 26417 4409 26440
rect 4495 26417 4577 26440
rect 4663 26417 4729 26440
rect 4343 26398 4729 26417
rect 19463 26503 19849 26522
rect 19463 26480 19529 26503
rect 19615 26480 19697 26503
rect 19783 26480 19849 26503
rect 19463 26440 19472 26480
rect 19512 26440 19529 26480
rect 19615 26440 19636 26480
rect 19676 26440 19697 26480
rect 19783 26440 19800 26480
rect 19840 26440 19849 26480
rect 19463 26417 19529 26440
rect 19615 26417 19697 26440
rect 19783 26417 19849 26440
rect 19463 26398 19849 26417
rect 34583 26503 34969 26522
rect 34583 26480 34649 26503
rect 34735 26480 34817 26503
rect 34903 26480 34969 26503
rect 34583 26440 34592 26480
rect 34632 26440 34649 26480
rect 34735 26440 34756 26480
rect 34796 26440 34817 26480
rect 34903 26440 34920 26480
rect 34960 26440 34969 26480
rect 34583 26417 34649 26440
rect 34735 26417 34817 26440
rect 34903 26417 34969 26440
rect 34583 26398 34969 26417
rect 49703 26503 50089 26522
rect 49703 26480 49769 26503
rect 49855 26480 49937 26503
rect 50023 26480 50089 26503
rect 49703 26440 49712 26480
rect 49752 26440 49769 26480
rect 49855 26440 49876 26480
rect 49916 26440 49937 26480
rect 50023 26440 50040 26480
rect 50080 26440 50089 26480
rect 49703 26417 49769 26440
rect 49855 26417 49937 26440
rect 50023 26417 50089 26440
rect 49703 26398 50089 26417
rect 64823 26503 65209 26522
rect 64823 26480 64889 26503
rect 64975 26480 65057 26503
rect 65143 26480 65209 26503
rect 64823 26440 64832 26480
rect 64872 26440 64889 26480
rect 64975 26440 64996 26480
rect 65036 26440 65057 26480
rect 65143 26440 65160 26480
rect 65200 26440 65209 26480
rect 64823 26417 64889 26440
rect 64975 26417 65057 26440
rect 65143 26417 65209 26440
rect 64823 26398 65209 26417
rect 79943 26503 80329 26522
rect 79943 26480 80009 26503
rect 80095 26480 80177 26503
rect 80263 26480 80329 26503
rect 79943 26440 79952 26480
rect 79992 26440 80009 26480
rect 80095 26440 80116 26480
rect 80156 26440 80177 26480
rect 80263 26440 80280 26480
rect 80320 26440 80329 26480
rect 79943 26417 80009 26440
rect 80095 26417 80177 26440
rect 80263 26417 80329 26440
rect 79943 26398 80329 26417
rect 3103 25747 3489 25766
rect 3103 25724 3169 25747
rect 3255 25724 3337 25747
rect 3423 25724 3489 25747
rect 3103 25684 3112 25724
rect 3152 25684 3169 25724
rect 3255 25684 3276 25724
rect 3316 25684 3337 25724
rect 3423 25684 3440 25724
rect 3480 25684 3489 25724
rect 3103 25661 3169 25684
rect 3255 25661 3337 25684
rect 3423 25661 3489 25684
rect 3103 25642 3489 25661
rect 18223 25747 18609 25766
rect 18223 25724 18289 25747
rect 18375 25724 18457 25747
rect 18543 25724 18609 25747
rect 18223 25684 18232 25724
rect 18272 25684 18289 25724
rect 18375 25684 18396 25724
rect 18436 25684 18457 25724
rect 18543 25684 18560 25724
rect 18600 25684 18609 25724
rect 18223 25661 18289 25684
rect 18375 25661 18457 25684
rect 18543 25661 18609 25684
rect 18223 25642 18609 25661
rect 33343 25747 33729 25766
rect 33343 25724 33409 25747
rect 33495 25724 33577 25747
rect 33663 25724 33729 25747
rect 33343 25684 33352 25724
rect 33392 25684 33409 25724
rect 33495 25684 33516 25724
rect 33556 25684 33577 25724
rect 33663 25684 33680 25724
rect 33720 25684 33729 25724
rect 33343 25661 33409 25684
rect 33495 25661 33577 25684
rect 33663 25661 33729 25684
rect 33343 25642 33729 25661
rect 48463 25747 48849 25766
rect 48463 25724 48529 25747
rect 48615 25724 48697 25747
rect 48783 25724 48849 25747
rect 48463 25684 48472 25724
rect 48512 25684 48529 25724
rect 48615 25684 48636 25724
rect 48676 25684 48697 25724
rect 48783 25684 48800 25724
rect 48840 25684 48849 25724
rect 48463 25661 48529 25684
rect 48615 25661 48697 25684
rect 48783 25661 48849 25684
rect 48463 25642 48849 25661
rect 63583 25747 63969 25766
rect 63583 25724 63649 25747
rect 63735 25724 63817 25747
rect 63903 25724 63969 25747
rect 63583 25684 63592 25724
rect 63632 25684 63649 25724
rect 63735 25684 63756 25724
rect 63796 25684 63817 25724
rect 63903 25684 63920 25724
rect 63960 25684 63969 25724
rect 63583 25661 63649 25684
rect 63735 25661 63817 25684
rect 63903 25661 63969 25684
rect 63583 25642 63969 25661
rect 78703 25747 79089 25766
rect 78703 25724 78769 25747
rect 78855 25724 78937 25747
rect 79023 25724 79089 25747
rect 78703 25684 78712 25724
rect 78752 25684 78769 25724
rect 78855 25684 78876 25724
rect 78916 25684 78937 25724
rect 79023 25684 79040 25724
rect 79080 25684 79089 25724
rect 78703 25661 78769 25684
rect 78855 25661 78937 25684
rect 79023 25661 79089 25684
rect 78703 25642 79089 25661
rect 4343 24991 4729 25010
rect 4343 24968 4409 24991
rect 4495 24968 4577 24991
rect 4663 24968 4729 24991
rect 4343 24928 4352 24968
rect 4392 24928 4409 24968
rect 4495 24928 4516 24968
rect 4556 24928 4577 24968
rect 4663 24928 4680 24968
rect 4720 24928 4729 24968
rect 4343 24905 4409 24928
rect 4495 24905 4577 24928
rect 4663 24905 4729 24928
rect 4343 24886 4729 24905
rect 19463 24991 19849 25010
rect 19463 24968 19529 24991
rect 19615 24968 19697 24991
rect 19783 24968 19849 24991
rect 19463 24928 19472 24968
rect 19512 24928 19529 24968
rect 19615 24928 19636 24968
rect 19676 24928 19697 24968
rect 19783 24928 19800 24968
rect 19840 24928 19849 24968
rect 19463 24905 19529 24928
rect 19615 24905 19697 24928
rect 19783 24905 19849 24928
rect 19463 24886 19849 24905
rect 34583 24991 34969 25010
rect 34583 24968 34649 24991
rect 34735 24968 34817 24991
rect 34903 24968 34969 24991
rect 34583 24928 34592 24968
rect 34632 24928 34649 24968
rect 34735 24928 34756 24968
rect 34796 24928 34817 24968
rect 34903 24928 34920 24968
rect 34960 24928 34969 24968
rect 34583 24905 34649 24928
rect 34735 24905 34817 24928
rect 34903 24905 34969 24928
rect 34583 24886 34969 24905
rect 49703 24991 50089 25010
rect 49703 24968 49769 24991
rect 49855 24968 49937 24991
rect 50023 24968 50089 24991
rect 49703 24928 49712 24968
rect 49752 24928 49769 24968
rect 49855 24928 49876 24968
rect 49916 24928 49937 24968
rect 50023 24928 50040 24968
rect 50080 24928 50089 24968
rect 49703 24905 49769 24928
rect 49855 24905 49937 24928
rect 50023 24905 50089 24928
rect 49703 24886 50089 24905
rect 64823 24991 65209 25010
rect 64823 24968 64889 24991
rect 64975 24968 65057 24991
rect 65143 24968 65209 24991
rect 64823 24928 64832 24968
rect 64872 24928 64889 24968
rect 64975 24928 64996 24968
rect 65036 24928 65057 24968
rect 65143 24928 65160 24968
rect 65200 24928 65209 24968
rect 64823 24905 64889 24928
rect 64975 24905 65057 24928
rect 65143 24905 65209 24928
rect 64823 24886 65209 24905
rect 79943 24991 80329 25010
rect 79943 24968 80009 24991
rect 80095 24968 80177 24991
rect 80263 24968 80329 24991
rect 79943 24928 79952 24968
rect 79992 24928 80009 24968
rect 80095 24928 80116 24968
rect 80156 24928 80177 24968
rect 80263 24928 80280 24968
rect 80320 24928 80329 24968
rect 79943 24905 80009 24928
rect 80095 24905 80177 24928
rect 80263 24905 80329 24928
rect 79943 24886 80329 24905
rect 3103 24235 3489 24254
rect 3103 24212 3169 24235
rect 3255 24212 3337 24235
rect 3423 24212 3489 24235
rect 3103 24172 3112 24212
rect 3152 24172 3169 24212
rect 3255 24172 3276 24212
rect 3316 24172 3337 24212
rect 3423 24172 3440 24212
rect 3480 24172 3489 24212
rect 3103 24149 3169 24172
rect 3255 24149 3337 24172
rect 3423 24149 3489 24172
rect 3103 24130 3489 24149
rect 18223 24235 18609 24254
rect 18223 24212 18289 24235
rect 18375 24212 18457 24235
rect 18543 24212 18609 24235
rect 18223 24172 18232 24212
rect 18272 24172 18289 24212
rect 18375 24172 18396 24212
rect 18436 24172 18457 24212
rect 18543 24172 18560 24212
rect 18600 24172 18609 24212
rect 18223 24149 18289 24172
rect 18375 24149 18457 24172
rect 18543 24149 18609 24172
rect 18223 24130 18609 24149
rect 33343 24235 33729 24254
rect 33343 24212 33409 24235
rect 33495 24212 33577 24235
rect 33663 24212 33729 24235
rect 33343 24172 33352 24212
rect 33392 24172 33409 24212
rect 33495 24172 33516 24212
rect 33556 24172 33577 24212
rect 33663 24172 33680 24212
rect 33720 24172 33729 24212
rect 33343 24149 33409 24172
rect 33495 24149 33577 24172
rect 33663 24149 33729 24172
rect 33343 24130 33729 24149
rect 48463 24235 48849 24254
rect 48463 24212 48529 24235
rect 48615 24212 48697 24235
rect 48783 24212 48849 24235
rect 48463 24172 48472 24212
rect 48512 24172 48529 24212
rect 48615 24172 48636 24212
rect 48676 24172 48697 24212
rect 48783 24172 48800 24212
rect 48840 24172 48849 24212
rect 48463 24149 48529 24172
rect 48615 24149 48697 24172
rect 48783 24149 48849 24172
rect 48463 24130 48849 24149
rect 63583 24235 63969 24254
rect 63583 24212 63649 24235
rect 63735 24212 63817 24235
rect 63903 24212 63969 24235
rect 63583 24172 63592 24212
rect 63632 24172 63649 24212
rect 63735 24172 63756 24212
rect 63796 24172 63817 24212
rect 63903 24172 63920 24212
rect 63960 24172 63969 24212
rect 63583 24149 63649 24172
rect 63735 24149 63817 24172
rect 63903 24149 63969 24172
rect 63583 24130 63969 24149
rect 78703 24235 79089 24254
rect 78703 24212 78769 24235
rect 78855 24212 78937 24235
rect 79023 24212 79089 24235
rect 78703 24172 78712 24212
rect 78752 24172 78769 24212
rect 78855 24172 78876 24212
rect 78916 24172 78937 24212
rect 79023 24172 79040 24212
rect 79080 24172 79089 24212
rect 78703 24149 78769 24172
rect 78855 24149 78937 24172
rect 79023 24149 79089 24172
rect 78703 24130 79089 24149
rect 4343 23479 4729 23498
rect 4343 23456 4409 23479
rect 4495 23456 4577 23479
rect 4663 23456 4729 23479
rect 4343 23416 4352 23456
rect 4392 23416 4409 23456
rect 4495 23416 4516 23456
rect 4556 23416 4577 23456
rect 4663 23416 4680 23456
rect 4720 23416 4729 23456
rect 4343 23393 4409 23416
rect 4495 23393 4577 23416
rect 4663 23393 4729 23416
rect 4343 23374 4729 23393
rect 19463 23479 19849 23498
rect 19463 23456 19529 23479
rect 19615 23456 19697 23479
rect 19783 23456 19849 23479
rect 19463 23416 19472 23456
rect 19512 23416 19529 23456
rect 19615 23416 19636 23456
rect 19676 23416 19697 23456
rect 19783 23416 19800 23456
rect 19840 23416 19849 23456
rect 19463 23393 19529 23416
rect 19615 23393 19697 23416
rect 19783 23393 19849 23416
rect 19463 23374 19849 23393
rect 34583 23479 34969 23498
rect 34583 23456 34649 23479
rect 34735 23456 34817 23479
rect 34903 23456 34969 23479
rect 34583 23416 34592 23456
rect 34632 23416 34649 23456
rect 34735 23416 34756 23456
rect 34796 23416 34817 23456
rect 34903 23416 34920 23456
rect 34960 23416 34969 23456
rect 34583 23393 34649 23416
rect 34735 23393 34817 23416
rect 34903 23393 34969 23416
rect 34583 23374 34969 23393
rect 49703 23479 50089 23498
rect 49703 23456 49769 23479
rect 49855 23456 49937 23479
rect 50023 23456 50089 23479
rect 49703 23416 49712 23456
rect 49752 23416 49769 23456
rect 49855 23416 49876 23456
rect 49916 23416 49937 23456
rect 50023 23416 50040 23456
rect 50080 23416 50089 23456
rect 49703 23393 49769 23416
rect 49855 23393 49937 23416
rect 50023 23393 50089 23416
rect 49703 23374 50089 23393
rect 64823 23479 65209 23498
rect 64823 23456 64889 23479
rect 64975 23456 65057 23479
rect 65143 23456 65209 23479
rect 64823 23416 64832 23456
rect 64872 23416 64889 23456
rect 64975 23416 64996 23456
rect 65036 23416 65057 23456
rect 65143 23416 65160 23456
rect 65200 23416 65209 23456
rect 64823 23393 64889 23416
rect 64975 23393 65057 23416
rect 65143 23393 65209 23416
rect 64823 23374 65209 23393
rect 79943 23479 80329 23498
rect 79943 23456 80009 23479
rect 80095 23456 80177 23479
rect 80263 23456 80329 23479
rect 79943 23416 79952 23456
rect 79992 23416 80009 23456
rect 80095 23416 80116 23456
rect 80156 23416 80177 23456
rect 80263 23416 80280 23456
rect 80320 23416 80329 23456
rect 79943 23393 80009 23416
rect 80095 23393 80177 23416
rect 80263 23393 80329 23416
rect 79943 23374 80329 23393
rect 3103 22723 3489 22742
rect 3103 22700 3169 22723
rect 3255 22700 3337 22723
rect 3423 22700 3489 22723
rect 3103 22660 3112 22700
rect 3152 22660 3169 22700
rect 3255 22660 3276 22700
rect 3316 22660 3337 22700
rect 3423 22660 3440 22700
rect 3480 22660 3489 22700
rect 3103 22637 3169 22660
rect 3255 22637 3337 22660
rect 3423 22637 3489 22660
rect 3103 22618 3489 22637
rect 18223 22723 18609 22742
rect 18223 22700 18289 22723
rect 18375 22700 18457 22723
rect 18543 22700 18609 22723
rect 18223 22660 18232 22700
rect 18272 22660 18289 22700
rect 18375 22660 18396 22700
rect 18436 22660 18457 22700
rect 18543 22660 18560 22700
rect 18600 22660 18609 22700
rect 18223 22637 18289 22660
rect 18375 22637 18457 22660
rect 18543 22637 18609 22660
rect 18223 22618 18609 22637
rect 33343 22723 33729 22742
rect 33343 22700 33409 22723
rect 33495 22700 33577 22723
rect 33663 22700 33729 22723
rect 33343 22660 33352 22700
rect 33392 22660 33409 22700
rect 33495 22660 33516 22700
rect 33556 22660 33577 22700
rect 33663 22660 33680 22700
rect 33720 22660 33729 22700
rect 33343 22637 33409 22660
rect 33495 22637 33577 22660
rect 33663 22637 33729 22660
rect 33343 22618 33729 22637
rect 48463 22723 48849 22742
rect 48463 22700 48529 22723
rect 48615 22700 48697 22723
rect 48783 22700 48849 22723
rect 48463 22660 48472 22700
rect 48512 22660 48529 22700
rect 48615 22660 48636 22700
rect 48676 22660 48697 22700
rect 48783 22660 48800 22700
rect 48840 22660 48849 22700
rect 48463 22637 48529 22660
rect 48615 22637 48697 22660
rect 48783 22637 48849 22660
rect 48463 22618 48849 22637
rect 63583 22723 63969 22742
rect 63583 22700 63649 22723
rect 63735 22700 63817 22723
rect 63903 22700 63969 22723
rect 63583 22660 63592 22700
rect 63632 22660 63649 22700
rect 63735 22660 63756 22700
rect 63796 22660 63817 22700
rect 63903 22660 63920 22700
rect 63960 22660 63969 22700
rect 63583 22637 63649 22660
rect 63735 22637 63817 22660
rect 63903 22637 63969 22660
rect 63583 22618 63969 22637
rect 78703 22723 79089 22742
rect 78703 22700 78769 22723
rect 78855 22700 78937 22723
rect 79023 22700 79089 22723
rect 78703 22660 78712 22700
rect 78752 22660 78769 22700
rect 78855 22660 78876 22700
rect 78916 22660 78937 22700
rect 79023 22660 79040 22700
rect 79080 22660 79089 22700
rect 78703 22637 78769 22660
rect 78855 22637 78937 22660
rect 79023 22637 79089 22660
rect 78703 22618 79089 22637
rect 4343 21967 4729 21986
rect 4343 21944 4409 21967
rect 4495 21944 4577 21967
rect 4663 21944 4729 21967
rect 4343 21904 4352 21944
rect 4392 21904 4409 21944
rect 4495 21904 4516 21944
rect 4556 21904 4577 21944
rect 4663 21904 4680 21944
rect 4720 21904 4729 21944
rect 4343 21881 4409 21904
rect 4495 21881 4577 21904
rect 4663 21881 4729 21904
rect 4343 21862 4729 21881
rect 19463 21967 19849 21986
rect 19463 21944 19529 21967
rect 19615 21944 19697 21967
rect 19783 21944 19849 21967
rect 19463 21904 19472 21944
rect 19512 21904 19529 21944
rect 19615 21904 19636 21944
rect 19676 21904 19697 21944
rect 19783 21904 19800 21944
rect 19840 21904 19849 21944
rect 19463 21881 19529 21904
rect 19615 21881 19697 21904
rect 19783 21881 19849 21904
rect 19463 21862 19849 21881
rect 34583 21967 34969 21986
rect 34583 21944 34649 21967
rect 34735 21944 34817 21967
rect 34903 21944 34969 21967
rect 34583 21904 34592 21944
rect 34632 21904 34649 21944
rect 34735 21904 34756 21944
rect 34796 21904 34817 21944
rect 34903 21904 34920 21944
rect 34960 21904 34969 21944
rect 34583 21881 34649 21904
rect 34735 21881 34817 21904
rect 34903 21881 34969 21904
rect 34583 21862 34969 21881
rect 49703 21967 50089 21986
rect 49703 21944 49769 21967
rect 49855 21944 49937 21967
rect 50023 21944 50089 21967
rect 49703 21904 49712 21944
rect 49752 21904 49769 21944
rect 49855 21904 49876 21944
rect 49916 21904 49937 21944
rect 50023 21904 50040 21944
rect 50080 21904 50089 21944
rect 49703 21881 49769 21904
rect 49855 21881 49937 21904
rect 50023 21881 50089 21904
rect 49703 21862 50089 21881
rect 64823 21967 65209 21986
rect 64823 21944 64889 21967
rect 64975 21944 65057 21967
rect 65143 21944 65209 21967
rect 64823 21904 64832 21944
rect 64872 21904 64889 21944
rect 64975 21904 64996 21944
rect 65036 21904 65057 21944
rect 65143 21904 65160 21944
rect 65200 21904 65209 21944
rect 64823 21881 64889 21904
rect 64975 21881 65057 21904
rect 65143 21881 65209 21904
rect 64823 21862 65209 21881
rect 79943 21967 80329 21986
rect 79943 21944 80009 21967
rect 80095 21944 80177 21967
rect 80263 21944 80329 21967
rect 79943 21904 79952 21944
rect 79992 21904 80009 21944
rect 80095 21904 80116 21944
rect 80156 21904 80177 21944
rect 80263 21904 80280 21944
rect 80320 21904 80329 21944
rect 79943 21881 80009 21904
rect 80095 21881 80177 21904
rect 80263 21881 80329 21904
rect 79943 21862 80329 21881
rect 3103 21211 3489 21230
rect 3103 21188 3169 21211
rect 3255 21188 3337 21211
rect 3423 21188 3489 21211
rect 3103 21148 3112 21188
rect 3152 21148 3169 21188
rect 3255 21148 3276 21188
rect 3316 21148 3337 21188
rect 3423 21148 3440 21188
rect 3480 21148 3489 21188
rect 3103 21125 3169 21148
rect 3255 21125 3337 21148
rect 3423 21125 3489 21148
rect 3103 21106 3489 21125
rect 18223 21211 18609 21230
rect 18223 21188 18289 21211
rect 18375 21188 18457 21211
rect 18543 21188 18609 21211
rect 18223 21148 18232 21188
rect 18272 21148 18289 21188
rect 18375 21148 18396 21188
rect 18436 21148 18457 21188
rect 18543 21148 18560 21188
rect 18600 21148 18609 21188
rect 18223 21125 18289 21148
rect 18375 21125 18457 21148
rect 18543 21125 18609 21148
rect 18223 21106 18609 21125
rect 33343 21211 33729 21230
rect 33343 21188 33409 21211
rect 33495 21188 33577 21211
rect 33663 21188 33729 21211
rect 33343 21148 33352 21188
rect 33392 21148 33409 21188
rect 33495 21148 33516 21188
rect 33556 21148 33577 21188
rect 33663 21148 33680 21188
rect 33720 21148 33729 21188
rect 33343 21125 33409 21148
rect 33495 21125 33577 21148
rect 33663 21125 33729 21148
rect 33343 21106 33729 21125
rect 48463 21211 48849 21230
rect 48463 21188 48529 21211
rect 48615 21188 48697 21211
rect 48783 21188 48849 21211
rect 48463 21148 48472 21188
rect 48512 21148 48529 21188
rect 48615 21148 48636 21188
rect 48676 21148 48697 21188
rect 48783 21148 48800 21188
rect 48840 21148 48849 21188
rect 48463 21125 48529 21148
rect 48615 21125 48697 21148
rect 48783 21125 48849 21148
rect 48463 21106 48849 21125
rect 63583 21211 63969 21230
rect 63583 21188 63649 21211
rect 63735 21188 63817 21211
rect 63903 21188 63969 21211
rect 63583 21148 63592 21188
rect 63632 21148 63649 21188
rect 63735 21148 63756 21188
rect 63796 21148 63817 21188
rect 63903 21148 63920 21188
rect 63960 21148 63969 21188
rect 63583 21125 63649 21148
rect 63735 21125 63817 21148
rect 63903 21125 63969 21148
rect 63583 21106 63969 21125
rect 78703 21211 79089 21230
rect 78703 21188 78769 21211
rect 78855 21188 78937 21211
rect 79023 21188 79089 21211
rect 78703 21148 78712 21188
rect 78752 21148 78769 21188
rect 78855 21148 78876 21188
rect 78916 21148 78937 21188
rect 79023 21148 79040 21188
rect 79080 21148 79089 21188
rect 78703 21125 78769 21148
rect 78855 21125 78937 21148
rect 79023 21125 79089 21148
rect 78703 21106 79089 21125
rect 4343 20455 4729 20474
rect 4343 20432 4409 20455
rect 4495 20432 4577 20455
rect 4663 20432 4729 20455
rect 4343 20392 4352 20432
rect 4392 20392 4409 20432
rect 4495 20392 4516 20432
rect 4556 20392 4577 20432
rect 4663 20392 4680 20432
rect 4720 20392 4729 20432
rect 4343 20369 4409 20392
rect 4495 20369 4577 20392
rect 4663 20369 4729 20392
rect 4343 20350 4729 20369
rect 19463 20455 19849 20474
rect 19463 20432 19529 20455
rect 19615 20432 19697 20455
rect 19783 20432 19849 20455
rect 19463 20392 19472 20432
rect 19512 20392 19529 20432
rect 19615 20392 19636 20432
rect 19676 20392 19697 20432
rect 19783 20392 19800 20432
rect 19840 20392 19849 20432
rect 19463 20369 19529 20392
rect 19615 20369 19697 20392
rect 19783 20369 19849 20392
rect 19463 20350 19849 20369
rect 34583 20455 34969 20474
rect 34583 20432 34649 20455
rect 34735 20432 34817 20455
rect 34903 20432 34969 20455
rect 34583 20392 34592 20432
rect 34632 20392 34649 20432
rect 34735 20392 34756 20432
rect 34796 20392 34817 20432
rect 34903 20392 34920 20432
rect 34960 20392 34969 20432
rect 34583 20369 34649 20392
rect 34735 20369 34817 20392
rect 34903 20369 34969 20392
rect 34583 20350 34969 20369
rect 49703 20455 50089 20474
rect 49703 20432 49769 20455
rect 49855 20432 49937 20455
rect 50023 20432 50089 20455
rect 49703 20392 49712 20432
rect 49752 20392 49769 20432
rect 49855 20392 49876 20432
rect 49916 20392 49937 20432
rect 50023 20392 50040 20432
rect 50080 20392 50089 20432
rect 49703 20369 49769 20392
rect 49855 20369 49937 20392
rect 50023 20369 50089 20392
rect 49703 20350 50089 20369
rect 64823 20455 65209 20474
rect 64823 20432 64889 20455
rect 64975 20432 65057 20455
rect 65143 20432 65209 20455
rect 64823 20392 64832 20432
rect 64872 20392 64889 20432
rect 64975 20392 64996 20432
rect 65036 20392 65057 20432
rect 65143 20392 65160 20432
rect 65200 20392 65209 20432
rect 64823 20369 64889 20392
rect 64975 20369 65057 20392
rect 65143 20369 65209 20392
rect 64823 20350 65209 20369
rect 79943 20455 80329 20474
rect 79943 20432 80009 20455
rect 80095 20432 80177 20455
rect 80263 20432 80329 20455
rect 79943 20392 79952 20432
rect 79992 20392 80009 20432
rect 80095 20392 80116 20432
rect 80156 20392 80177 20432
rect 80263 20392 80280 20432
rect 80320 20392 80329 20432
rect 79943 20369 80009 20392
rect 80095 20369 80177 20392
rect 80263 20369 80329 20392
rect 79943 20350 80329 20369
rect 3103 19699 3489 19718
rect 3103 19676 3169 19699
rect 3255 19676 3337 19699
rect 3423 19676 3489 19699
rect 3103 19636 3112 19676
rect 3152 19636 3169 19676
rect 3255 19636 3276 19676
rect 3316 19636 3337 19676
rect 3423 19636 3440 19676
rect 3480 19636 3489 19676
rect 3103 19613 3169 19636
rect 3255 19613 3337 19636
rect 3423 19613 3489 19636
rect 3103 19594 3489 19613
rect 18223 19699 18609 19718
rect 18223 19676 18289 19699
rect 18375 19676 18457 19699
rect 18543 19676 18609 19699
rect 18223 19636 18232 19676
rect 18272 19636 18289 19676
rect 18375 19636 18396 19676
rect 18436 19636 18457 19676
rect 18543 19636 18560 19676
rect 18600 19636 18609 19676
rect 18223 19613 18289 19636
rect 18375 19613 18457 19636
rect 18543 19613 18609 19636
rect 18223 19594 18609 19613
rect 33343 19699 33729 19718
rect 33343 19676 33409 19699
rect 33495 19676 33577 19699
rect 33663 19676 33729 19699
rect 33343 19636 33352 19676
rect 33392 19636 33409 19676
rect 33495 19636 33516 19676
rect 33556 19636 33577 19676
rect 33663 19636 33680 19676
rect 33720 19636 33729 19676
rect 33343 19613 33409 19636
rect 33495 19613 33577 19636
rect 33663 19613 33729 19636
rect 33343 19594 33729 19613
rect 48463 19699 48849 19718
rect 48463 19676 48529 19699
rect 48615 19676 48697 19699
rect 48783 19676 48849 19699
rect 48463 19636 48472 19676
rect 48512 19636 48529 19676
rect 48615 19636 48636 19676
rect 48676 19636 48697 19676
rect 48783 19636 48800 19676
rect 48840 19636 48849 19676
rect 48463 19613 48529 19636
rect 48615 19613 48697 19636
rect 48783 19613 48849 19636
rect 48463 19594 48849 19613
rect 63583 19699 63969 19718
rect 63583 19676 63649 19699
rect 63735 19676 63817 19699
rect 63903 19676 63969 19699
rect 63583 19636 63592 19676
rect 63632 19636 63649 19676
rect 63735 19636 63756 19676
rect 63796 19636 63817 19676
rect 63903 19636 63920 19676
rect 63960 19636 63969 19676
rect 63583 19613 63649 19636
rect 63735 19613 63817 19636
rect 63903 19613 63969 19636
rect 63583 19594 63969 19613
rect 78703 19699 79089 19718
rect 78703 19676 78769 19699
rect 78855 19676 78937 19699
rect 79023 19676 79089 19699
rect 78703 19636 78712 19676
rect 78752 19636 78769 19676
rect 78855 19636 78876 19676
rect 78916 19636 78937 19676
rect 79023 19636 79040 19676
rect 79080 19636 79089 19676
rect 78703 19613 78769 19636
rect 78855 19613 78937 19636
rect 79023 19613 79089 19636
rect 78703 19594 79089 19613
rect 4343 18943 4729 18962
rect 4343 18920 4409 18943
rect 4495 18920 4577 18943
rect 4663 18920 4729 18943
rect 4343 18880 4352 18920
rect 4392 18880 4409 18920
rect 4495 18880 4516 18920
rect 4556 18880 4577 18920
rect 4663 18880 4680 18920
rect 4720 18880 4729 18920
rect 4343 18857 4409 18880
rect 4495 18857 4577 18880
rect 4663 18857 4729 18880
rect 4343 18838 4729 18857
rect 19463 18943 19849 18962
rect 19463 18920 19529 18943
rect 19615 18920 19697 18943
rect 19783 18920 19849 18943
rect 19463 18880 19472 18920
rect 19512 18880 19529 18920
rect 19615 18880 19636 18920
rect 19676 18880 19697 18920
rect 19783 18880 19800 18920
rect 19840 18880 19849 18920
rect 19463 18857 19529 18880
rect 19615 18857 19697 18880
rect 19783 18857 19849 18880
rect 19463 18838 19849 18857
rect 34583 18943 34969 18962
rect 34583 18920 34649 18943
rect 34735 18920 34817 18943
rect 34903 18920 34969 18943
rect 34583 18880 34592 18920
rect 34632 18880 34649 18920
rect 34735 18880 34756 18920
rect 34796 18880 34817 18920
rect 34903 18880 34920 18920
rect 34960 18880 34969 18920
rect 34583 18857 34649 18880
rect 34735 18857 34817 18880
rect 34903 18857 34969 18880
rect 34583 18838 34969 18857
rect 49703 18943 50089 18962
rect 49703 18920 49769 18943
rect 49855 18920 49937 18943
rect 50023 18920 50089 18943
rect 49703 18880 49712 18920
rect 49752 18880 49769 18920
rect 49855 18880 49876 18920
rect 49916 18880 49937 18920
rect 50023 18880 50040 18920
rect 50080 18880 50089 18920
rect 49703 18857 49769 18880
rect 49855 18857 49937 18880
rect 50023 18857 50089 18880
rect 49703 18838 50089 18857
rect 64823 18943 65209 18962
rect 64823 18920 64889 18943
rect 64975 18920 65057 18943
rect 65143 18920 65209 18943
rect 64823 18880 64832 18920
rect 64872 18880 64889 18920
rect 64975 18880 64996 18920
rect 65036 18880 65057 18920
rect 65143 18880 65160 18920
rect 65200 18880 65209 18920
rect 64823 18857 64889 18880
rect 64975 18857 65057 18880
rect 65143 18857 65209 18880
rect 64823 18838 65209 18857
rect 79943 18943 80329 18962
rect 79943 18920 80009 18943
rect 80095 18920 80177 18943
rect 80263 18920 80329 18943
rect 79943 18880 79952 18920
rect 79992 18880 80009 18920
rect 80095 18880 80116 18920
rect 80156 18880 80177 18920
rect 80263 18880 80280 18920
rect 80320 18880 80329 18920
rect 79943 18857 80009 18880
rect 80095 18857 80177 18880
rect 80263 18857 80329 18880
rect 79943 18838 80329 18857
rect 3103 18187 3489 18206
rect 3103 18164 3169 18187
rect 3255 18164 3337 18187
rect 3423 18164 3489 18187
rect 3103 18124 3112 18164
rect 3152 18124 3169 18164
rect 3255 18124 3276 18164
rect 3316 18124 3337 18164
rect 3423 18124 3440 18164
rect 3480 18124 3489 18164
rect 3103 18101 3169 18124
rect 3255 18101 3337 18124
rect 3423 18101 3489 18124
rect 3103 18082 3489 18101
rect 18223 18187 18609 18206
rect 18223 18164 18289 18187
rect 18375 18164 18457 18187
rect 18543 18164 18609 18187
rect 18223 18124 18232 18164
rect 18272 18124 18289 18164
rect 18375 18124 18396 18164
rect 18436 18124 18457 18164
rect 18543 18124 18560 18164
rect 18600 18124 18609 18164
rect 18223 18101 18289 18124
rect 18375 18101 18457 18124
rect 18543 18101 18609 18124
rect 18223 18082 18609 18101
rect 33343 18187 33729 18206
rect 33343 18164 33409 18187
rect 33495 18164 33577 18187
rect 33663 18164 33729 18187
rect 33343 18124 33352 18164
rect 33392 18124 33409 18164
rect 33495 18124 33516 18164
rect 33556 18124 33577 18164
rect 33663 18124 33680 18164
rect 33720 18124 33729 18164
rect 33343 18101 33409 18124
rect 33495 18101 33577 18124
rect 33663 18101 33729 18124
rect 33343 18082 33729 18101
rect 48463 18187 48849 18206
rect 48463 18164 48529 18187
rect 48615 18164 48697 18187
rect 48783 18164 48849 18187
rect 48463 18124 48472 18164
rect 48512 18124 48529 18164
rect 48615 18124 48636 18164
rect 48676 18124 48697 18164
rect 48783 18124 48800 18164
rect 48840 18124 48849 18164
rect 48463 18101 48529 18124
rect 48615 18101 48697 18124
rect 48783 18101 48849 18124
rect 48463 18082 48849 18101
rect 63583 18187 63969 18206
rect 63583 18164 63649 18187
rect 63735 18164 63817 18187
rect 63903 18164 63969 18187
rect 63583 18124 63592 18164
rect 63632 18124 63649 18164
rect 63735 18124 63756 18164
rect 63796 18124 63817 18164
rect 63903 18124 63920 18164
rect 63960 18124 63969 18164
rect 63583 18101 63649 18124
rect 63735 18101 63817 18124
rect 63903 18101 63969 18124
rect 63583 18082 63969 18101
rect 78703 18187 79089 18206
rect 78703 18164 78769 18187
rect 78855 18164 78937 18187
rect 79023 18164 79089 18187
rect 78703 18124 78712 18164
rect 78752 18124 78769 18164
rect 78855 18124 78876 18164
rect 78916 18124 78937 18164
rect 79023 18124 79040 18164
rect 79080 18124 79089 18164
rect 78703 18101 78769 18124
rect 78855 18101 78937 18124
rect 79023 18101 79089 18124
rect 78703 18082 79089 18101
rect 4343 17431 4729 17450
rect 4343 17408 4409 17431
rect 4495 17408 4577 17431
rect 4663 17408 4729 17431
rect 4343 17368 4352 17408
rect 4392 17368 4409 17408
rect 4495 17368 4516 17408
rect 4556 17368 4577 17408
rect 4663 17368 4680 17408
rect 4720 17368 4729 17408
rect 4343 17345 4409 17368
rect 4495 17345 4577 17368
rect 4663 17345 4729 17368
rect 4343 17326 4729 17345
rect 19463 17431 19849 17450
rect 19463 17408 19529 17431
rect 19615 17408 19697 17431
rect 19783 17408 19849 17431
rect 19463 17368 19472 17408
rect 19512 17368 19529 17408
rect 19615 17368 19636 17408
rect 19676 17368 19697 17408
rect 19783 17368 19800 17408
rect 19840 17368 19849 17408
rect 19463 17345 19529 17368
rect 19615 17345 19697 17368
rect 19783 17345 19849 17368
rect 19463 17326 19849 17345
rect 34583 17431 34969 17450
rect 34583 17408 34649 17431
rect 34735 17408 34817 17431
rect 34903 17408 34969 17431
rect 34583 17368 34592 17408
rect 34632 17368 34649 17408
rect 34735 17368 34756 17408
rect 34796 17368 34817 17408
rect 34903 17368 34920 17408
rect 34960 17368 34969 17408
rect 34583 17345 34649 17368
rect 34735 17345 34817 17368
rect 34903 17345 34969 17368
rect 34583 17326 34969 17345
rect 49703 17431 50089 17450
rect 49703 17408 49769 17431
rect 49855 17408 49937 17431
rect 50023 17408 50089 17431
rect 49703 17368 49712 17408
rect 49752 17368 49769 17408
rect 49855 17368 49876 17408
rect 49916 17368 49937 17408
rect 50023 17368 50040 17408
rect 50080 17368 50089 17408
rect 49703 17345 49769 17368
rect 49855 17345 49937 17368
rect 50023 17345 50089 17368
rect 49703 17326 50089 17345
rect 64823 17431 65209 17450
rect 64823 17408 64889 17431
rect 64975 17408 65057 17431
rect 65143 17408 65209 17431
rect 64823 17368 64832 17408
rect 64872 17368 64889 17408
rect 64975 17368 64996 17408
rect 65036 17368 65057 17408
rect 65143 17368 65160 17408
rect 65200 17368 65209 17408
rect 64823 17345 64889 17368
rect 64975 17345 65057 17368
rect 65143 17345 65209 17368
rect 64823 17326 65209 17345
rect 79943 17431 80329 17450
rect 79943 17408 80009 17431
rect 80095 17408 80177 17431
rect 80263 17408 80329 17431
rect 79943 17368 79952 17408
rect 79992 17368 80009 17408
rect 80095 17368 80116 17408
rect 80156 17368 80177 17408
rect 80263 17368 80280 17408
rect 80320 17368 80329 17408
rect 79943 17345 80009 17368
rect 80095 17345 80177 17368
rect 80263 17345 80329 17368
rect 79943 17326 80329 17345
rect 3103 16675 3489 16694
rect 3103 16652 3169 16675
rect 3255 16652 3337 16675
rect 3423 16652 3489 16675
rect 3103 16612 3112 16652
rect 3152 16612 3169 16652
rect 3255 16612 3276 16652
rect 3316 16612 3337 16652
rect 3423 16612 3440 16652
rect 3480 16612 3489 16652
rect 3103 16589 3169 16612
rect 3255 16589 3337 16612
rect 3423 16589 3489 16612
rect 3103 16570 3489 16589
rect 18223 16675 18609 16694
rect 18223 16652 18289 16675
rect 18375 16652 18457 16675
rect 18543 16652 18609 16675
rect 18223 16612 18232 16652
rect 18272 16612 18289 16652
rect 18375 16612 18396 16652
rect 18436 16612 18457 16652
rect 18543 16612 18560 16652
rect 18600 16612 18609 16652
rect 18223 16589 18289 16612
rect 18375 16589 18457 16612
rect 18543 16589 18609 16612
rect 18223 16570 18609 16589
rect 33343 16675 33729 16694
rect 33343 16652 33409 16675
rect 33495 16652 33577 16675
rect 33663 16652 33729 16675
rect 33343 16612 33352 16652
rect 33392 16612 33409 16652
rect 33495 16612 33516 16652
rect 33556 16612 33577 16652
rect 33663 16612 33680 16652
rect 33720 16612 33729 16652
rect 33343 16589 33409 16612
rect 33495 16589 33577 16612
rect 33663 16589 33729 16612
rect 33343 16570 33729 16589
rect 48463 16675 48849 16694
rect 48463 16652 48529 16675
rect 48615 16652 48697 16675
rect 48783 16652 48849 16675
rect 48463 16612 48472 16652
rect 48512 16612 48529 16652
rect 48615 16612 48636 16652
rect 48676 16612 48697 16652
rect 48783 16612 48800 16652
rect 48840 16612 48849 16652
rect 48463 16589 48529 16612
rect 48615 16589 48697 16612
rect 48783 16589 48849 16612
rect 48463 16570 48849 16589
rect 63583 16675 63969 16694
rect 63583 16652 63649 16675
rect 63735 16652 63817 16675
rect 63903 16652 63969 16675
rect 63583 16612 63592 16652
rect 63632 16612 63649 16652
rect 63735 16612 63756 16652
rect 63796 16612 63817 16652
rect 63903 16612 63920 16652
rect 63960 16612 63969 16652
rect 63583 16589 63649 16612
rect 63735 16589 63817 16612
rect 63903 16589 63969 16612
rect 63583 16570 63969 16589
rect 78703 16675 79089 16694
rect 78703 16652 78769 16675
rect 78855 16652 78937 16675
rect 79023 16652 79089 16675
rect 78703 16612 78712 16652
rect 78752 16612 78769 16652
rect 78855 16612 78876 16652
rect 78916 16612 78937 16652
rect 79023 16612 79040 16652
rect 79080 16612 79089 16652
rect 78703 16589 78769 16612
rect 78855 16589 78937 16612
rect 79023 16589 79089 16612
rect 78703 16570 79089 16589
rect 4343 15919 4729 15938
rect 4343 15896 4409 15919
rect 4495 15896 4577 15919
rect 4663 15896 4729 15919
rect 4343 15856 4352 15896
rect 4392 15856 4409 15896
rect 4495 15856 4516 15896
rect 4556 15856 4577 15896
rect 4663 15856 4680 15896
rect 4720 15856 4729 15896
rect 4343 15833 4409 15856
rect 4495 15833 4577 15856
rect 4663 15833 4729 15856
rect 4343 15814 4729 15833
rect 19463 15919 19849 15938
rect 19463 15896 19529 15919
rect 19615 15896 19697 15919
rect 19783 15896 19849 15919
rect 19463 15856 19472 15896
rect 19512 15856 19529 15896
rect 19615 15856 19636 15896
rect 19676 15856 19697 15896
rect 19783 15856 19800 15896
rect 19840 15856 19849 15896
rect 19463 15833 19529 15856
rect 19615 15833 19697 15856
rect 19783 15833 19849 15856
rect 19463 15814 19849 15833
rect 34583 15919 34969 15938
rect 34583 15896 34649 15919
rect 34735 15896 34817 15919
rect 34903 15896 34969 15919
rect 34583 15856 34592 15896
rect 34632 15856 34649 15896
rect 34735 15856 34756 15896
rect 34796 15856 34817 15896
rect 34903 15856 34920 15896
rect 34960 15856 34969 15896
rect 34583 15833 34649 15856
rect 34735 15833 34817 15856
rect 34903 15833 34969 15856
rect 34583 15814 34969 15833
rect 49703 15919 50089 15938
rect 49703 15896 49769 15919
rect 49855 15896 49937 15919
rect 50023 15896 50089 15919
rect 49703 15856 49712 15896
rect 49752 15856 49769 15896
rect 49855 15856 49876 15896
rect 49916 15856 49937 15896
rect 50023 15856 50040 15896
rect 50080 15856 50089 15896
rect 49703 15833 49769 15856
rect 49855 15833 49937 15856
rect 50023 15833 50089 15856
rect 49703 15814 50089 15833
rect 64823 15919 65209 15938
rect 64823 15896 64889 15919
rect 64975 15896 65057 15919
rect 65143 15896 65209 15919
rect 64823 15856 64832 15896
rect 64872 15856 64889 15896
rect 64975 15856 64996 15896
rect 65036 15856 65057 15896
rect 65143 15856 65160 15896
rect 65200 15856 65209 15896
rect 64823 15833 64889 15856
rect 64975 15833 65057 15856
rect 65143 15833 65209 15856
rect 64823 15814 65209 15833
rect 79943 15919 80329 15938
rect 79943 15896 80009 15919
rect 80095 15896 80177 15919
rect 80263 15896 80329 15919
rect 79943 15856 79952 15896
rect 79992 15856 80009 15896
rect 80095 15856 80116 15896
rect 80156 15856 80177 15896
rect 80263 15856 80280 15896
rect 80320 15856 80329 15896
rect 79943 15833 80009 15856
rect 80095 15833 80177 15856
rect 80263 15833 80329 15856
rect 79943 15814 80329 15833
rect 3103 15163 3489 15182
rect 3103 15140 3169 15163
rect 3255 15140 3337 15163
rect 3423 15140 3489 15163
rect 3103 15100 3112 15140
rect 3152 15100 3169 15140
rect 3255 15100 3276 15140
rect 3316 15100 3337 15140
rect 3423 15100 3440 15140
rect 3480 15100 3489 15140
rect 3103 15077 3169 15100
rect 3255 15077 3337 15100
rect 3423 15077 3489 15100
rect 3103 15058 3489 15077
rect 18223 15163 18609 15182
rect 18223 15140 18289 15163
rect 18375 15140 18457 15163
rect 18543 15140 18609 15163
rect 18223 15100 18232 15140
rect 18272 15100 18289 15140
rect 18375 15100 18396 15140
rect 18436 15100 18457 15140
rect 18543 15100 18560 15140
rect 18600 15100 18609 15140
rect 18223 15077 18289 15100
rect 18375 15077 18457 15100
rect 18543 15077 18609 15100
rect 18223 15058 18609 15077
rect 33343 15163 33729 15182
rect 33343 15140 33409 15163
rect 33495 15140 33577 15163
rect 33663 15140 33729 15163
rect 33343 15100 33352 15140
rect 33392 15100 33409 15140
rect 33495 15100 33516 15140
rect 33556 15100 33577 15140
rect 33663 15100 33680 15140
rect 33720 15100 33729 15140
rect 33343 15077 33409 15100
rect 33495 15077 33577 15100
rect 33663 15077 33729 15100
rect 33343 15058 33729 15077
rect 48463 15163 48849 15182
rect 48463 15140 48529 15163
rect 48615 15140 48697 15163
rect 48783 15140 48849 15163
rect 48463 15100 48472 15140
rect 48512 15100 48529 15140
rect 48615 15100 48636 15140
rect 48676 15100 48697 15140
rect 48783 15100 48800 15140
rect 48840 15100 48849 15140
rect 48463 15077 48529 15100
rect 48615 15077 48697 15100
rect 48783 15077 48849 15100
rect 48463 15058 48849 15077
rect 63583 15163 63969 15182
rect 63583 15140 63649 15163
rect 63735 15140 63817 15163
rect 63903 15140 63969 15163
rect 63583 15100 63592 15140
rect 63632 15100 63649 15140
rect 63735 15100 63756 15140
rect 63796 15100 63817 15140
rect 63903 15100 63920 15140
rect 63960 15100 63969 15140
rect 63583 15077 63649 15100
rect 63735 15077 63817 15100
rect 63903 15077 63969 15100
rect 63583 15058 63969 15077
rect 78703 15163 79089 15182
rect 78703 15140 78769 15163
rect 78855 15140 78937 15163
rect 79023 15140 79089 15163
rect 78703 15100 78712 15140
rect 78752 15100 78769 15140
rect 78855 15100 78876 15140
rect 78916 15100 78937 15140
rect 79023 15100 79040 15140
rect 79080 15100 79089 15140
rect 78703 15077 78769 15100
rect 78855 15077 78937 15100
rect 79023 15077 79089 15100
rect 78703 15058 79089 15077
rect 4343 14407 4729 14426
rect 4343 14384 4409 14407
rect 4495 14384 4577 14407
rect 4663 14384 4729 14407
rect 4343 14344 4352 14384
rect 4392 14344 4409 14384
rect 4495 14344 4516 14384
rect 4556 14344 4577 14384
rect 4663 14344 4680 14384
rect 4720 14344 4729 14384
rect 4343 14321 4409 14344
rect 4495 14321 4577 14344
rect 4663 14321 4729 14344
rect 4343 14302 4729 14321
rect 19463 14407 19849 14426
rect 19463 14384 19529 14407
rect 19615 14384 19697 14407
rect 19783 14384 19849 14407
rect 19463 14344 19472 14384
rect 19512 14344 19529 14384
rect 19615 14344 19636 14384
rect 19676 14344 19697 14384
rect 19783 14344 19800 14384
rect 19840 14344 19849 14384
rect 19463 14321 19529 14344
rect 19615 14321 19697 14344
rect 19783 14321 19849 14344
rect 19463 14302 19849 14321
rect 34583 14407 34969 14426
rect 34583 14384 34649 14407
rect 34735 14384 34817 14407
rect 34903 14384 34969 14407
rect 34583 14344 34592 14384
rect 34632 14344 34649 14384
rect 34735 14344 34756 14384
rect 34796 14344 34817 14384
rect 34903 14344 34920 14384
rect 34960 14344 34969 14384
rect 34583 14321 34649 14344
rect 34735 14321 34817 14344
rect 34903 14321 34969 14344
rect 34583 14302 34969 14321
rect 49703 14407 50089 14426
rect 49703 14384 49769 14407
rect 49855 14384 49937 14407
rect 50023 14384 50089 14407
rect 49703 14344 49712 14384
rect 49752 14344 49769 14384
rect 49855 14344 49876 14384
rect 49916 14344 49937 14384
rect 50023 14344 50040 14384
rect 50080 14344 50089 14384
rect 49703 14321 49769 14344
rect 49855 14321 49937 14344
rect 50023 14321 50089 14344
rect 49703 14302 50089 14321
rect 64823 14407 65209 14426
rect 64823 14384 64889 14407
rect 64975 14384 65057 14407
rect 65143 14384 65209 14407
rect 64823 14344 64832 14384
rect 64872 14344 64889 14384
rect 64975 14344 64996 14384
rect 65036 14344 65057 14384
rect 65143 14344 65160 14384
rect 65200 14344 65209 14384
rect 64823 14321 64889 14344
rect 64975 14321 65057 14344
rect 65143 14321 65209 14344
rect 64823 14302 65209 14321
rect 79943 14407 80329 14426
rect 79943 14384 80009 14407
rect 80095 14384 80177 14407
rect 80263 14384 80329 14407
rect 79943 14344 79952 14384
rect 79992 14344 80009 14384
rect 80095 14344 80116 14384
rect 80156 14344 80177 14384
rect 80263 14344 80280 14384
rect 80320 14344 80329 14384
rect 79943 14321 80009 14344
rect 80095 14321 80177 14344
rect 80263 14321 80329 14344
rect 79943 14302 80329 14321
rect 3103 13651 3489 13670
rect 3103 13628 3169 13651
rect 3255 13628 3337 13651
rect 3423 13628 3489 13651
rect 3103 13588 3112 13628
rect 3152 13588 3169 13628
rect 3255 13588 3276 13628
rect 3316 13588 3337 13628
rect 3423 13588 3440 13628
rect 3480 13588 3489 13628
rect 3103 13565 3169 13588
rect 3255 13565 3337 13588
rect 3423 13565 3489 13588
rect 3103 13546 3489 13565
rect 18223 13651 18609 13670
rect 18223 13628 18289 13651
rect 18375 13628 18457 13651
rect 18543 13628 18609 13651
rect 18223 13588 18232 13628
rect 18272 13588 18289 13628
rect 18375 13588 18396 13628
rect 18436 13588 18457 13628
rect 18543 13588 18560 13628
rect 18600 13588 18609 13628
rect 18223 13565 18289 13588
rect 18375 13565 18457 13588
rect 18543 13565 18609 13588
rect 18223 13546 18609 13565
rect 33343 13651 33729 13670
rect 33343 13628 33409 13651
rect 33495 13628 33577 13651
rect 33663 13628 33729 13651
rect 33343 13588 33352 13628
rect 33392 13588 33409 13628
rect 33495 13588 33516 13628
rect 33556 13588 33577 13628
rect 33663 13588 33680 13628
rect 33720 13588 33729 13628
rect 33343 13565 33409 13588
rect 33495 13565 33577 13588
rect 33663 13565 33729 13588
rect 33343 13546 33729 13565
rect 48463 13651 48849 13670
rect 48463 13628 48529 13651
rect 48615 13628 48697 13651
rect 48783 13628 48849 13651
rect 48463 13588 48472 13628
rect 48512 13588 48529 13628
rect 48615 13588 48636 13628
rect 48676 13588 48697 13628
rect 48783 13588 48800 13628
rect 48840 13588 48849 13628
rect 48463 13565 48529 13588
rect 48615 13565 48697 13588
rect 48783 13565 48849 13588
rect 48463 13546 48849 13565
rect 63583 13651 63969 13670
rect 63583 13628 63649 13651
rect 63735 13628 63817 13651
rect 63903 13628 63969 13651
rect 63583 13588 63592 13628
rect 63632 13588 63649 13628
rect 63735 13588 63756 13628
rect 63796 13588 63817 13628
rect 63903 13588 63920 13628
rect 63960 13588 63969 13628
rect 63583 13565 63649 13588
rect 63735 13565 63817 13588
rect 63903 13565 63969 13588
rect 63583 13546 63969 13565
rect 78703 13651 79089 13670
rect 78703 13628 78769 13651
rect 78855 13628 78937 13651
rect 79023 13628 79089 13651
rect 78703 13588 78712 13628
rect 78752 13588 78769 13628
rect 78855 13588 78876 13628
rect 78916 13588 78937 13628
rect 79023 13588 79040 13628
rect 79080 13588 79089 13628
rect 78703 13565 78769 13588
rect 78855 13565 78937 13588
rect 79023 13565 79089 13588
rect 78703 13546 79089 13565
rect 4343 12895 4729 12914
rect 4343 12872 4409 12895
rect 4495 12872 4577 12895
rect 4663 12872 4729 12895
rect 4343 12832 4352 12872
rect 4392 12832 4409 12872
rect 4495 12832 4516 12872
rect 4556 12832 4577 12872
rect 4663 12832 4680 12872
rect 4720 12832 4729 12872
rect 4343 12809 4409 12832
rect 4495 12809 4577 12832
rect 4663 12809 4729 12832
rect 4343 12790 4729 12809
rect 19463 12895 19849 12914
rect 19463 12872 19529 12895
rect 19615 12872 19697 12895
rect 19783 12872 19849 12895
rect 19463 12832 19472 12872
rect 19512 12832 19529 12872
rect 19615 12832 19636 12872
rect 19676 12832 19697 12872
rect 19783 12832 19800 12872
rect 19840 12832 19849 12872
rect 19463 12809 19529 12832
rect 19615 12809 19697 12832
rect 19783 12809 19849 12832
rect 19463 12790 19849 12809
rect 34583 12895 34969 12914
rect 34583 12872 34649 12895
rect 34735 12872 34817 12895
rect 34903 12872 34969 12895
rect 34583 12832 34592 12872
rect 34632 12832 34649 12872
rect 34735 12832 34756 12872
rect 34796 12832 34817 12872
rect 34903 12832 34920 12872
rect 34960 12832 34969 12872
rect 34583 12809 34649 12832
rect 34735 12809 34817 12832
rect 34903 12809 34969 12832
rect 34583 12790 34969 12809
rect 49703 12895 50089 12914
rect 49703 12872 49769 12895
rect 49855 12872 49937 12895
rect 50023 12872 50089 12895
rect 49703 12832 49712 12872
rect 49752 12832 49769 12872
rect 49855 12832 49876 12872
rect 49916 12832 49937 12872
rect 50023 12832 50040 12872
rect 50080 12832 50089 12872
rect 49703 12809 49769 12832
rect 49855 12809 49937 12832
rect 50023 12809 50089 12832
rect 49703 12790 50089 12809
rect 64823 12895 65209 12914
rect 64823 12872 64889 12895
rect 64975 12872 65057 12895
rect 65143 12872 65209 12895
rect 64823 12832 64832 12872
rect 64872 12832 64889 12872
rect 64975 12832 64996 12872
rect 65036 12832 65057 12872
rect 65143 12832 65160 12872
rect 65200 12832 65209 12872
rect 64823 12809 64889 12832
rect 64975 12809 65057 12832
rect 65143 12809 65209 12832
rect 64823 12790 65209 12809
rect 79943 12895 80329 12914
rect 79943 12872 80009 12895
rect 80095 12872 80177 12895
rect 80263 12872 80329 12895
rect 79943 12832 79952 12872
rect 79992 12832 80009 12872
rect 80095 12832 80116 12872
rect 80156 12832 80177 12872
rect 80263 12832 80280 12872
rect 80320 12832 80329 12872
rect 79943 12809 80009 12832
rect 80095 12809 80177 12832
rect 80263 12809 80329 12832
rect 79943 12790 80329 12809
rect 3103 12139 3489 12158
rect 3103 12116 3169 12139
rect 3255 12116 3337 12139
rect 3423 12116 3489 12139
rect 3103 12076 3112 12116
rect 3152 12076 3169 12116
rect 3255 12076 3276 12116
rect 3316 12076 3337 12116
rect 3423 12076 3440 12116
rect 3480 12076 3489 12116
rect 3103 12053 3169 12076
rect 3255 12053 3337 12076
rect 3423 12053 3489 12076
rect 3103 12034 3489 12053
rect 18223 12139 18609 12158
rect 18223 12116 18289 12139
rect 18375 12116 18457 12139
rect 18543 12116 18609 12139
rect 18223 12076 18232 12116
rect 18272 12076 18289 12116
rect 18375 12076 18396 12116
rect 18436 12076 18457 12116
rect 18543 12076 18560 12116
rect 18600 12076 18609 12116
rect 18223 12053 18289 12076
rect 18375 12053 18457 12076
rect 18543 12053 18609 12076
rect 18223 12034 18609 12053
rect 33343 12139 33729 12158
rect 33343 12116 33409 12139
rect 33495 12116 33577 12139
rect 33663 12116 33729 12139
rect 33343 12076 33352 12116
rect 33392 12076 33409 12116
rect 33495 12076 33516 12116
rect 33556 12076 33577 12116
rect 33663 12076 33680 12116
rect 33720 12076 33729 12116
rect 33343 12053 33409 12076
rect 33495 12053 33577 12076
rect 33663 12053 33729 12076
rect 33343 12034 33729 12053
rect 48463 12139 48849 12158
rect 48463 12116 48529 12139
rect 48615 12116 48697 12139
rect 48783 12116 48849 12139
rect 48463 12076 48472 12116
rect 48512 12076 48529 12116
rect 48615 12076 48636 12116
rect 48676 12076 48697 12116
rect 48783 12076 48800 12116
rect 48840 12076 48849 12116
rect 48463 12053 48529 12076
rect 48615 12053 48697 12076
rect 48783 12053 48849 12076
rect 48463 12034 48849 12053
rect 63583 12139 63969 12158
rect 63583 12116 63649 12139
rect 63735 12116 63817 12139
rect 63903 12116 63969 12139
rect 63583 12076 63592 12116
rect 63632 12076 63649 12116
rect 63735 12076 63756 12116
rect 63796 12076 63817 12116
rect 63903 12076 63920 12116
rect 63960 12076 63969 12116
rect 63583 12053 63649 12076
rect 63735 12053 63817 12076
rect 63903 12053 63969 12076
rect 63583 12034 63969 12053
rect 78703 12139 79089 12158
rect 78703 12116 78769 12139
rect 78855 12116 78937 12139
rect 79023 12116 79089 12139
rect 78703 12076 78712 12116
rect 78752 12076 78769 12116
rect 78855 12076 78876 12116
rect 78916 12076 78937 12116
rect 79023 12076 79040 12116
rect 79080 12076 79089 12116
rect 78703 12053 78769 12076
rect 78855 12053 78937 12076
rect 79023 12053 79089 12076
rect 78703 12034 79089 12053
rect 4343 11383 4729 11402
rect 4343 11360 4409 11383
rect 4495 11360 4577 11383
rect 4663 11360 4729 11383
rect 4343 11320 4352 11360
rect 4392 11320 4409 11360
rect 4495 11320 4516 11360
rect 4556 11320 4577 11360
rect 4663 11320 4680 11360
rect 4720 11320 4729 11360
rect 4343 11297 4409 11320
rect 4495 11297 4577 11320
rect 4663 11297 4729 11320
rect 4343 11278 4729 11297
rect 19463 11383 19849 11402
rect 19463 11360 19529 11383
rect 19615 11360 19697 11383
rect 19783 11360 19849 11383
rect 19463 11320 19472 11360
rect 19512 11320 19529 11360
rect 19615 11320 19636 11360
rect 19676 11320 19697 11360
rect 19783 11320 19800 11360
rect 19840 11320 19849 11360
rect 19463 11297 19529 11320
rect 19615 11297 19697 11320
rect 19783 11297 19849 11320
rect 19463 11278 19849 11297
rect 34583 11383 34969 11402
rect 34583 11360 34649 11383
rect 34735 11360 34817 11383
rect 34903 11360 34969 11383
rect 34583 11320 34592 11360
rect 34632 11320 34649 11360
rect 34735 11320 34756 11360
rect 34796 11320 34817 11360
rect 34903 11320 34920 11360
rect 34960 11320 34969 11360
rect 34583 11297 34649 11320
rect 34735 11297 34817 11320
rect 34903 11297 34969 11320
rect 34583 11278 34969 11297
rect 49703 11383 50089 11402
rect 49703 11360 49769 11383
rect 49855 11360 49937 11383
rect 50023 11360 50089 11383
rect 49703 11320 49712 11360
rect 49752 11320 49769 11360
rect 49855 11320 49876 11360
rect 49916 11320 49937 11360
rect 50023 11320 50040 11360
rect 50080 11320 50089 11360
rect 49703 11297 49769 11320
rect 49855 11297 49937 11320
rect 50023 11297 50089 11320
rect 49703 11278 50089 11297
rect 64823 11383 65209 11402
rect 64823 11360 64889 11383
rect 64975 11360 65057 11383
rect 65143 11360 65209 11383
rect 64823 11320 64832 11360
rect 64872 11320 64889 11360
rect 64975 11320 64996 11360
rect 65036 11320 65057 11360
rect 65143 11320 65160 11360
rect 65200 11320 65209 11360
rect 64823 11297 64889 11320
rect 64975 11297 65057 11320
rect 65143 11297 65209 11320
rect 64823 11278 65209 11297
rect 79943 11383 80329 11402
rect 79943 11360 80009 11383
rect 80095 11360 80177 11383
rect 80263 11360 80329 11383
rect 79943 11320 79952 11360
rect 79992 11320 80009 11360
rect 80095 11320 80116 11360
rect 80156 11320 80177 11360
rect 80263 11320 80280 11360
rect 80320 11320 80329 11360
rect 79943 11297 80009 11320
rect 80095 11297 80177 11320
rect 80263 11297 80329 11320
rect 79943 11278 80329 11297
rect 3103 10627 3489 10646
rect 3103 10604 3169 10627
rect 3255 10604 3337 10627
rect 3423 10604 3489 10627
rect 3103 10564 3112 10604
rect 3152 10564 3169 10604
rect 3255 10564 3276 10604
rect 3316 10564 3337 10604
rect 3423 10564 3440 10604
rect 3480 10564 3489 10604
rect 3103 10541 3169 10564
rect 3255 10541 3337 10564
rect 3423 10541 3489 10564
rect 3103 10522 3489 10541
rect 18223 10627 18609 10646
rect 18223 10604 18289 10627
rect 18375 10604 18457 10627
rect 18543 10604 18609 10627
rect 18223 10564 18232 10604
rect 18272 10564 18289 10604
rect 18375 10564 18396 10604
rect 18436 10564 18457 10604
rect 18543 10564 18560 10604
rect 18600 10564 18609 10604
rect 18223 10541 18289 10564
rect 18375 10541 18457 10564
rect 18543 10541 18609 10564
rect 18223 10522 18609 10541
rect 33343 10627 33729 10646
rect 33343 10604 33409 10627
rect 33495 10604 33577 10627
rect 33663 10604 33729 10627
rect 33343 10564 33352 10604
rect 33392 10564 33409 10604
rect 33495 10564 33516 10604
rect 33556 10564 33577 10604
rect 33663 10564 33680 10604
rect 33720 10564 33729 10604
rect 33343 10541 33409 10564
rect 33495 10541 33577 10564
rect 33663 10541 33729 10564
rect 33343 10522 33729 10541
rect 48463 10627 48849 10646
rect 48463 10604 48529 10627
rect 48615 10604 48697 10627
rect 48783 10604 48849 10627
rect 48463 10564 48472 10604
rect 48512 10564 48529 10604
rect 48615 10564 48636 10604
rect 48676 10564 48697 10604
rect 48783 10564 48800 10604
rect 48840 10564 48849 10604
rect 48463 10541 48529 10564
rect 48615 10541 48697 10564
rect 48783 10541 48849 10564
rect 48463 10522 48849 10541
rect 63583 10627 63969 10646
rect 63583 10604 63649 10627
rect 63735 10604 63817 10627
rect 63903 10604 63969 10627
rect 63583 10564 63592 10604
rect 63632 10564 63649 10604
rect 63735 10564 63756 10604
rect 63796 10564 63817 10604
rect 63903 10564 63920 10604
rect 63960 10564 63969 10604
rect 63583 10541 63649 10564
rect 63735 10541 63817 10564
rect 63903 10541 63969 10564
rect 63583 10522 63969 10541
rect 78703 10627 79089 10646
rect 78703 10604 78769 10627
rect 78855 10604 78937 10627
rect 79023 10604 79089 10627
rect 78703 10564 78712 10604
rect 78752 10564 78769 10604
rect 78855 10564 78876 10604
rect 78916 10564 78937 10604
rect 79023 10564 79040 10604
rect 79080 10564 79089 10604
rect 78703 10541 78769 10564
rect 78855 10541 78937 10564
rect 79023 10541 79089 10564
rect 78703 10522 79089 10541
rect 4343 9871 4729 9890
rect 4343 9848 4409 9871
rect 4495 9848 4577 9871
rect 4663 9848 4729 9871
rect 4343 9808 4352 9848
rect 4392 9808 4409 9848
rect 4495 9808 4516 9848
rect 4556 9808 4577 9848
rect 4663 9808 4680 9848
rect 4720 9808 4729 9848
rect 4343 9785 4409 9808
rect 4495 9785 4577 9808
rect 4663 9785 4729 9808
rect 4343 9766 4729 9785
rect 19463 9871 19849 9890
rect 19463 9848 19529 9871
rect 19615 9848 19697 9871
rect 19783 9848 19849 9871
rect 19463 9808 19472 9848
rect 19512 9808 19529 9848
rect 19615 9808 19636 9848
rect 19676 9808 19697 9848
rect 19783 9808 19800 9848
rect 19840 9808 19849 9848
rect 19463 9785 19529 9808
rect 19615 9785 19697 9808
rect 19783 9785 19849 9808
rect 19463 9766 19849 9785
rect 34583 9871 34969 9890
rect 34583 9848 34649 9871
rect 34735 9848 34817 9871
rect 34903 9848 34969 9871
rect 34583 9808 34592 9848
rect 34632 9808 34649 9848
rect 34735 9808 34756 9848
rect 34796 9808 34817 9848
rect 34903 9808 34920 9848
rect 34960 9808 34969 9848
rect 34583 9785 34649 9808
rect 34735 9785 34817 9808
rect 34903 9785 34969 9808
rect 34583 9766 34969 9785
rect 49703 9871 50089 9890
rect 49703 9848 49769 9871
rect 49855 9848 49937 9871
rect 50023 9848 50089 9871
rect 49703 9808 49712 9848
rect 49752 9808 49769 9848
rect 49855 9808 49876 9848
rect 49916 9808 49937 9848
rect 50023 9808 50040 9848
rect 50080 9808 50089 9848
rect 49703 9785 49769 9808
rect 49855 9785 49937 9808
rect 50023 9785 50089 9808
rect 49703 9766 50089 9785
rect 64823 9871 65209 9890
rect 64823 9848 64889 9871
rect 64975 9848 65057 9871
rect 65143 9848 65209 9871
rect 64823 9808 64832 9848
rect 64872 9808 64889 9848
rect 64975 9808 64996 9848
rect 65036 9808 65057 9848
rect 65143 9808 65160 9848
rect 65200 9808 65209 9848
rect 64823 9785 64889 9808
rect 64975 9785 65057 9808
rect 65143 9785 65209 9808
rect 64823 9766 65209 9785
rect 79943 9871 80329 9890
rect 79943 9848 80009 9871
rect 80095 9848 80177 9871
rect 80263 9848 80329 9871
rect 79943 9808 79952 9848
rect 79992 9808 80009 9848
rect 80095 9808 80116 9848
rect 80156 9808 80177 9848
rect 80263 9808 80280 9848
rect 80320 9808 80329 9848
rect 79943 9785 80009 9808
rect 80095 9785 80177 9808
rect 80263 9785 80329 9808
rect 79943 9766 80329 9785
rect 3103 9115 3489 9134
rect 3103 9092 3169 9115
rect 3255 9092 3337 9115
rect 3423 9092 3489 9115
rect 3103 9052 3112 9092
rect 3152 9052 3169 9092
rect 3255 9052 3276 9092
rect 3316 9052 3337 9092
rect 3423 9052 3440 9092
rect 3480 9052 3489 9092
rect 3103 9029 3169 9052
rect 3255 9029 3337 9052
rect 3423 9029 3489 9052
rect 3103 9010 3489 9029
rect 18223 9115 18609 9134
rect 18223 9092 18289 9115
rect 18375 9092 18457 9115
rect 18543 9092 18609 9115
rect 18223 9052 18232 9092
rect 18272 9052 18289 9092
rect 18375 9052 18396 9092
rect 18436 9052 18457 9092
rect 18543 9052 18560 9092
rect 18600 9052 18609 9092
rect 18223 9029 18289 9052
rect 18375 9029 18457 9052
rect 18543 9029 18609 9052
rect 18223 9010 18609 9029
rect 33343 9115 33729 9134
rect 33343 9092 33409 9115
rect 33495 9092 33577 9115
rect 33663 9092 33729 9115
rect 33343 9052 33352 9092
rect 33392 9052 33409 9092
rect 33495 9052 33516 9092
rect 33556 9052 33577 9092
rect 33663 9052 33680 9092
rect 33720 9052 33729 9092
rect 33343 9029 33409 9052
rect 33495 9029 33577 9052
rect 33663 9029 33729 9052
rect 33343 9010 33729 9029
rect 48463 9115 48849 9134
rect 48463 9092 48529 9115
rect 48615 9092 48697 9115
rect 48783 9092 48849 9115
rect 48463 9052 48472 9092
rect 48512 9052 48529 9092
rect 48615 9052 48636 9092
rect 48676 9052 48697 9092
rect 48783 9052 48800 9092
rect 48840 9052 48849 9092
rect 48463 9029 48529 9052
rect 48615 9029 48697 9052
rect 48783 9029 48849 9052
rect 48463 9010 48849 9029
rect 63583 9115 63969 9134
rect 63583 9092 63649 9115
rect 63735 9092 63817 9115
rect 63903 9092 63969 9115
rect 63583 9052 63592 9092
rect 63632 9052 63649 9092
rect 63735 9052 63756 9092
rect 63796 9052 63817 9092
rect 63903 9052 63920 9092
rect 63960 9052 63969 9092
rect 63583 9029 63649 9052
rect 63735 9029 63817 9052
rect 63903 9029 63969 9052
rect 63583 9010 63969 9029
rect 78703 9115 79089 9134
rect 78703 9092 78769 9115
rect 78855 9092 78937 9115
rect 79023 9092 79089 9115
rect 78703 9052 78712 9092
rect 78752 9052 78769 9092
rect 78855 9052 78876 9092
rect 78916 9052 78937 9092
rect 79023 9052 79040 9092
rect 79080 9052 79089 9092
rect 78703 9029 78769 9052
rect 78855 9029 78937 9052
rect 79023 9029 79089 9052
rect 78703 9010 79089 9029
rect 4343 8359 4729 8378
rect 4343 8336 4409 8359
rect 4495 8336 4577 8359
rect 4663 8336 4729 8359
rect 4343 8296 4352 8336
rect 4392 8296 4409 8336
rect 4495 8296 4516 8336
rect 4556 8296 4577 8336
rect 4663 8296 4680 8336
rect 4720 8296 4729 8336
rect 4343 8273 4409 8296
rect 4495 8273 4577 8296
rect 4663 8273 4729 8296
rect 4343 8254 4729 8273
rect 19463 8359 19849 8378
rect 19463 8336 19529 8359
rect 19615 8336 19697 8359
rect 19783 8336 19849 8359
rect 19463 8296 19472 8336
rect 19512 8296 19529 8336
rect 19615 8296 19636 8336
rect 19676 8296 19697 8336
rect 19783 8296 19800 8336
rect 19840 8296 19849 8336
rect 19463 8273 19529 8296
rect 19615 8273 19697 8296
rect 19783 8273 19849 8296
rect 19463 8254 19849 8273
rect 34583 8359 34969 8378
rect 34583 8336 34649 8359
rect 34735 8336 34817 8359
rect 34903 8336 34969 8359
rect 34583 8296 34592 8336
rect 34632 8296 34649 8336
rect 34735 8296 34756 8336
rect 34796 8296 34817 8336
rect 34903 8296 34920 8336
rect 34960 8296 34969 8336
rect 34583 8273 34649 8296
rect 34735 8273 34817 8296
rect 34903 8273 34969 8296
rect 34583 8254 34969 8273
rect 49703 8359 50089 8378
rect 49703 8336 49769 8359
rect 49855 8336 49937 8359
rect 50023 8336 50089 8359
rect 49703 8296 49712 8336
rect 49752 8296 49769 8336
rect 49855 8296 49876 8336
rect 49916 8296 49937 8336
rect 50023 8296 50040 8336
rect 50080 8296 50089 8336
rect 49703 8273 49769 8296
rect 49855 8273 49937 8296
rect 50023 8273 50089 8296
rect 49703 8254 50089 8273
rect 64823 8359 65209 8378
rect 64823 8336 64889 8359
rect 64975 8336 65057 8359
rect 65143 8336 65209 8359
rect 64823 8296 64832 8336
rect 64872 8296 64889 8336
rect 64975 8296 64996 8336
rect 65036 8296 65057 8336
rect 65143 8296 65160 8336
rect 65200 8296 65209 8336
rect 64823 8273 64889 8296
rect 64975 8273 65057 8296
rect 65143 8273 65209 8296
rect 64823 8254 65209 8273
rect 79943 8359 80329 8378
rect 79943 8336 80009 8359
rect 80095 8336 80177 8359
rect 80263 8336 80329 8359
rect 79943 8296 79952 8336
rect 79992 8296 80009 8336
rect 80095 8296 80116 8336
rect 80156 8296 80177 8336
rect 80263 8296 80280 8336
rect 80320 8296 80329 8336
rect 79943 8273 80009 8296
rect 80095 8273 80177 8296
rect 80263 8273 80329 8296
rect 79943 8254 80329 8273
rect 3103 7603 3489 7622
rect 3103 7580 3169 7603
rect 3255 7580 3337 7603
rect 3423 7580 3489 7603
rect 3103 7540 3112 7580
rect 3152 7540 3169 7580
rect 3255 7540 3276 7580
rect 3316 7540 3337 7580
rect 3423 7540 3440 7580
rect 3480 7540 3489 7580
rect 3103 7517 3169 7540
rect 3255 7517 3337 7540
rect 3423 7517 3489 7540
rect 3103 7498 3489 7517
rect 18223 7603 18609 7622
rect 18223 7580 18289 7603
rect 18375 7580 18457 7603
rect 18543 7580 18609 7603
rect 18223 7540 18232 7580
rect 18272 7540 18289 7580
rect 18375 7540 18396 7580
rect 18436 7540 18457 7580
rect 18543 7540 18560 7580
rect 18600 7540 18609 7580
rect 18223 7517 18289 7540
rect 18375 7517 18457 7540
rect 18543 7517 18609 7540
rect 18223 7498 18609 7517
rect 33343 7603 33729 7622
rect 33343 7580 33409 7603
rect 33495 7580 33577 7603
rect 33663 7580 33729 7603
rect 33343 7540 33352 7580
rect 33392 7540 33409 7580
rect 33495 7540 33516 7580
rect 33556 7540 33577 7580
rect 33663 7540 33680 7580
rect 33720 7540 33729 7580
rect 33343 7517 33409 7540
rect 33495 7517 33577 7540
rect 33663 7517 33729 7540
rect 33343 7498 33729 7517
rect 48463 7603 48849 7622
rect 48463 7580 48529 7603
rect 48615 7580 48697 7603
rect 48783 7580 48849 7603
rect 48463 7540 48472 7580
rect 48512 7540 48529 7580
rect 48615 7540 48636 7580
rect 48676 7540 48697 7580
rect 48783 7540 48800 7580
rect 48840 7540 48849 7580
rect 48463 7517 48529 7540
rect 48615 7517 48697 7540
rect 48783 7517 48849 7540
rect 48463 7498 48849 7517
rect 63583 7603 63969 7622
rect 63583 7580 63649 7603
rect 63735 7580 63817 7603
rect 63903 7580 63969 7603
rect 63583 7540 63592 7580
rect 63632 7540 63649 7580
rect 63735 7540 63756 7580
rect 63796 7540 63817 7580
rect 63903 7540 63920 7580
rect 63960 7540 63969 7580
rect 63583 7517 63649 7540
rect 63735 7517 63817 7540
rect 63903 7517 63969 7540
rect 63583 7498 63969 7517
rect 78703 7603 79089 7622
rect 78703 7580 78769 7603
rect 78855 7580 78937 7603
rect 79023 7580 79089 7603
rect 78703 7540 78712 7580
rect 78752 7540 78769 7580
rect 78855 7540 78876 7580
rect 78916 7540 78937 7580
rect 79023 7540 79040 7580
rect 79080 7540 79089 7580
rect 78703 7517 78769 7540
rect 78855 7517 78937 7540
rect 79023 7517 79089 7540
rect 78703 7498 79089 7517
rect 4343 6847 4729 6866
rect 4343 6824 4409 6847
rect 4495 6824 4577 6847
rect 4663 6824 4729 6847
rect 4343 6784 4352 6824
rect 4392 6784 4409 6824
rect 4495 6784 4516 6824
rect 4556 6784 4577 6824
rect 4663 6784 4680 6824
rect 4720 6784 4729 6824
rect 4343 6761 4409 6784
rect 4495 6761 4577 6784
rect 4663 6761 4729 6784
rect 4343 6742 4729 6761
rect 19463 6847 19849 6866
rect 19463 6824 19529 6847
rect 19615 6824 19697 6847
rect 19783 6824 19849 6847
rect 19463 6784 19472 6824
rect 19512 6784 19529 6824
rect 19615 6784 19636 6824
rect 19676 6784 19697 6824
rect 19783 6784 19800 6824
rect 19840 6784 19849 6824
rect 19463 6761 19529 6784
rect 19615 6761 19697 6784
rect 19783 6761 19849 6784
rect 19463 6742 19849 6761
rect 34583 6847 34969 6866
rect 34583 6824 34649 6847
rect 34735 6824 34817 6847
rect 34903 6824 34969 6847
rect 34583 6784 34592 6824
rect 34632 6784 34649 6824
rect 34735 6784 34756 6824
rect 34796 6784 34817 6824
rect 34903 6784 34920 6824
rect 34960 6784 34969 6824
rect 34583 6761 34649 6784
rect 34735 6761 34817 6784
rect 34903 6761 34969 6784
rect 34583 6742 34969 6761
rect 49703 6847 50089 6866
rect 49703 6824 49769 6847
rect 49855 6824 49937 6847
rect 50023 6824 50089 6847
rect 49703 6784 49712 6824
rect 49752 6784 49769 6824
rect 49855 6784 49876 6824
rect 49916 6784 49937 6824
rect 50023 6784 50040 6824
rect 50080 6784 50089 6824
rect 49703 6761 49769 6784
rect 49855 6761 49937 6784
rect 50023 6761 50089 6784
rect 49703 6742 50089 6761
rect 64823 6847 65209 6866
rect 64823 6824 64889 6847
rect 64975 6824 65057 6847
rect 65143 6824 65209 6847
rect 64823 6784 64832 6824
rect 64872 6784 64889 6824
rect 64975 6784 64996 6824
rect 65036 6784 65057 6824
rect 65143 6784 65160 6824
rect 65200 6784 65209 6824
rect 64823 6761 64889 6784
rect 64975 6761 65057 6784
rect 65143 6761 65209 6784
rect 64823 6742 65209 6761
rect 79943 6847 80329 6866
rect 79943 6824 80009 6847
rect 80095 6824 80177 6847
rect 80263 6824 80329 6847
rect 79943 6784 79952 6824
rect 79992 6784 80009 6824
rect 80095 6784 80116 6824
rect 80156 6784 80177 6824
rect 80263 6784 80280 6824
rect 80320 6784 80329 6824
rect 79943 6761 80009 6784
rect 80095 6761 80177 6784
rect 80263 6761 80329 6784
rect 79943 6742 80329 6761
rect 3103 6091 3489 6110
rect 3103 6068 3169 6091
rect 3255 6068 3337 6091
rect 3423 6068 3489 6091
rect 3103 6028 3112 6068
rect 3152 6028 3169 6068
rect 3255 6028 3276 6068
rect 3316 6028 3337 6068
rect 3423 6028 3440 6068
rect 3480 6028 3489 6068
rect 3103 6005 3169 6028
rect 3255 6005 3337 6028
rect 3423 6005 3489 6028
rect 3103 5986 3489 6005
rect 18223 6091 18609 6110
rect 18223 6068 18289 6091
rect 18375 6068 18457 6091
rect 18543 6068 18609 6091
rect 18223 6028 18232 6068
rect 18272 6028 18289 6068
rect 18375 6028 18396 6068
rect 18436 6028 18457 6068
rect 18543 6028 18560 6068
rect 18600 6028 18609 6068
rect 18223 6005 18289 6028
rect 18375 6005 18457 6028
rect 18543 6005 18609 6028
rect 18223 5986 18609 6005
rect 33343 6091 33729 6110
rect 33343 6068 33409 6091
rect 33495 6068 33577 6091
rect 33663 6068 33729 6091
rect 33343 6028 33352 6068
rect 33392 6028 33409 6068
rect 33495 6028 33516 6068
rect 33556 6028 33577 6068
rect 33663 6028 33680 6068
rect 33720 6028 33729 6068
rect 33343 6005 33409 6028
rect 33495 6005 33577 6028
rect 33663 6005 33729 6028
rect 33343 5986 33729 6005
rect 48463 6091 48849 6110
rect 48463 6068 48529 6091
rect 48615 6068 48697 6091
rect 48783 6068 48849 6091
rect 48463 6028 48472 6068
rect 48512 6028 48529 6068
rect 48615 6028 48636 6068
rect 48676 6028 48697 6068
rect 48783 6028 48800 6068
rect 48840 6028 48849 6068
rect 48463 6005 48529 6028
rect 48615 6005 48697 6028
rect 48783 6005 48849 6028
rect 48463 5986 48849 6005
rect 63583 6091 63969 6110
rect 63583 6068 63649 6091
rect 63735 6068 63817 6091
rect 63903 6068 63969 6091
rect 63583 6028 63592 6068
rect 63632 6028 63649 6068
rect 63735 6028 63756 6068
rect 63796 6028 63817 6068
rect 63903 6028 63920 6068
rect 63960 6028 63969 6068
rect 63583 6005 63649 6028
rect 63735 6005 63817 6028
rect 63903 6005 63969 6028
rect 63583 5986 63969 6005
rect 78703 6091 79089 6110
rect 78703 6068 78769 6091
rect 78855 6068 78937 6091
rect 79023 6068 79089 6091
rect 78703 6028 78712 6068
rect 78752 6028 78769 6068
rect 78855 6028 78876 6068
rect 78916 6028 78937 6068
rect 79023 6028 79040 6068
rect 79080 6028 79089 6068
rect 78703 6005 78769 6028
rect 78855 6005 78937 6028
rect 79023 6005 79089 6028
rect 78703 5986 79089 6005
rect 4343 5335 4729 5354
rect 4343 5312 4409 5335
rect 4495 5312 4577 5335
rect 4663 5312 4729 5335
rect 4343 5272 4352 5312
rect 4392 5272 4409 5312
rect 4495 5272 4516 5312
rect 4556 5272 4577 5312
rect 4663 5272 4680 5312
rect 4720 5272 4729 5312
rect 4343 5249 4409 5272
rect 4495 5249 4577 5272
rect 4663 5249 4729 5272
rect 4343 5230 4729 5249
rect 19463 5335 19849 5354
rect 19463 5312 19529 5335
rect 19615 5312 19697 5335
rect 19783 5312 19849 5335
rect 19463 5272 19472 5312
rect 19512 5272 19529 5312
rect 19615 5272 19636 5312
rect 19676 5272 19697 5312
rect 19783 5272 19800 5312
rect 19840 5272 19849 5312
rect 19463 5249 19529 5272
rect 19615 5249 19697 5272
rect 19783 5249 19849 5272
rect 19463 5230 19849 5249
rect 34583 5335 34969 5354
rect 34583 5312 34649 5335
rect 34735 5312 34817 5335
rect 34903 5312 34969 5335
rect 34583 5272 34592 5312
rect 34632 5272 34649 5312
rect 34735 5272 34756 5312
rect 34796 5272 34817 5312
rect 34903 5272 34920 5312
rect 34960 5272 34969 5312
rect 34583 5249 34649 5272
rect 34735 5249 34817 5272
rect 34903 5249 34969 5272
rect 34583 5230 34969 5249
rect 49703 5335 50089 5354
rect 49703 5312 49769 5335
rect 49855 5312 49937 5335
rect 50023 5312 50089 5335
rect 49703 5272 49712 5312
rect 49752 5272 49769 5312
rect 49855 5272 49876 5312
rect 49916 5272 49937 5312
rect 50023 5272 50040 5312
rect 50080 5272 50089 5312
rect 49703 5249 49769 5272
rect 49855 5249 49937 5272
rect 50023 5249 50089 5272
rect 49703 5230 50089 5249
rect 64823 5335 65209 5354
rect 64823 5312 64889 5335
rect 64975 5312 65057 5335
rect 65143 5312 65209 5335
rect 64823 5272 64832 5312
rect 64872 5272 64889 5312
rect 64975 5272 64996 5312
rect 65036 5272 65057 5312
rect 65143 5272 65160 5312
rect 65200 5272 65209 5312
rect 64823 5249 64889 5272
rect 64975 5249 65057 5272
rect 65143 5249 65209 5272
rect 64823 5230 65209 5249
rect 79943 5335 80329 5354
rect 79943 5312 80009 5335
rect 80095 5312 80177 5335
rect 80263 5312 80329 5335
rect 79943 5272 79952 5312
rect 79992 5272 80009 5312
rect 80095 5272 80116 5312
rect 80156 5272 80177 5312
rect 80263 5272 80280 5312
rect 80320 5272 80329 5312
rect 79943 5249 80009 5272
rect 80095 5249 80177 5272
rect 80263 5249 80329 5272
rect 79943 5230 80329 5249
rect 3103 4579 3489 4598
rect 3103 4556 3169 4579
rect 3255 4556 3337 4579
rect 3423 4556 3489 4579
rect 3103 4516 3112 4556
rect 3152 4516 3169 4556
rect 3255 4516 3276 4556
rect 3316 4516 3337 4556
rect 3423 4516 3440 4556
rect 3480 4516 3489 4556
rect 3103 4493 3169 4516
rect 3255 4493 3337 4516
rect 3423 4493 3489 4516
rect 3103 4474 3489 4493
rect 18223 4579 18609 4598
rect 18223 4556 18289 4579
rect 18375 4556 18457 4579
rect 18543 4556 18609 4579
rect 18223 4516 18232 4556
rect 18272 4516 18289 4556
rect 18375 4516 18396 4556
rect 18436 4516 18457 4556
rect 18543 4516 18560 4556
rect 18600 4516 18609 4556
rect 18223 4493 18289 4516
rect 18375 4493 18457 4516
rect 18543 4493 18609 4516
rect 18223 4474 18609 4493
rect 33343 4579 33729 4598
rect 33343 4556 33409 4579
rect 33495 4556 33577 4579
rect 33663 4556 33729 4579
rect 33343 4516 33352 4556
rect 33392 4516 33409 4556
rect 33495 4516 33516 4556
rect 33556 4516 33577 4556
rect 33663 4516 33680 4556
rect 33720 4516 33729 4556
rect 33343 4493 33409 4516
rect 33495 4493 33577 4516
rect 33663 4493 33729 4516
rect 33343 4474 33729 4493
rect 48463 4579 48849 4598
rect 48463 4556 48529 4579
rect 48615 4556 48697 4579
rect 48783 4556 48849 4579
rect 48463 4516 48472 4556
rect 48512 4516 48529 4556
rect 48615 4516 48636 4556
rect 48676 4516 48697 4556
rect 48783 4516 48800 4556
rect 48840 4516 48849 4556
rect 48463 4493 48529 4516
rect 48615 4493 48697 4516
rect 48783 4493 48849 4516
rect 48463 4474 48849 4493
rect 63583 4579 63969 4598
rect 63583 4556 63649 4579
rect 63735 4556 63817 4579
rect 63903 4556 63969 4579
rect 63583 4516 63592 4556
rect 63632 4516 63649 4556
rect 63735 4516 63756 4556
rect 63796 4516 63817 4556
rect 63903 4516 63920 4556
rect 63960 4516 63969 4556
rect 63583 4493 63649 4516
rect 63735 4493 63817 4516
rect 63903 4493 63969 4516
rect 63583 4474 63969 4493
rect 78703 4579 79089 4598
rect 78703 4556 78769 4579
rect 78855 4556 78937 4579
rect 79023 4556 79089 4579
rect 78703 4516 78712 4556
rect 78752 4516 78769 4556
rect 78855 4516 78876 4556
rect 78916 4516 78937 4556
rect 79023 4516 79040 4556
rect 79080 4516 79089 4556
rect 78703 4493 78769 4516
rect 78855 4493 78937 4516
rect 79023 4493 79089 4516
rect 78703 4474 79089 4493
rect 4343 3823 4729 3842
rect 4343 3800 4409 3823
rect 4495 3800 4577 3823
rect 4663 3800 4729 3823
rect 4343 3760 4352 3800
rect 4392 3760 4409 3800
rect 4495 3760 4516 3800
rect 4556 3760 4577 3800
rect 4663 3760 4680 3800
rect 4720 3760 4729 3800
rect 4343 3737 4409 3760
rect 4495 3737 4577 3760
rect 4663 3737 4729 3760
rect 4343 3718 4729 3737
rect 19463 3823 19849 3842
rect 19463 3800 19529 3823
rect 19615 3800 19697 3823
rect 19783 3800 19849 3823
rect 19463 3760 19472 3800
rect 19512 3760 19529 3800
rect 19615 3760 19636 3800
rect 19676 3760 19697 3800
rect 19783 3760 19800 3800
rect 19840 3760 19849 3800
rect 19463 3737 19529 3760
rect 19615 3737 19697 3760
rect 19783 3737 19849 3760
rect 19463 3718 19849 3737
rect 34583 3823 34969 3842
rect 34583 3800 34649 3823
rect 34735 3800 34817 3823
rect 34903 3800 34969 3823
rect 34583 3760 34592 3800
rect 34632 3760 34649 3800
rect 34735 3760 34756 3800
rect 34796 3760 34817 3800
rect 34903 3760 34920 3800
rect 34960 3760 34969 3800
rect 34583 3737 34649 3760
rect 34735 3737 34817 3760
rect 34903 3737 34969 3760
rect 34583 3718 34969 3737
rect 49703 3823 50089 3842
rect 49703 3800 49769 3823
rect 49855 3800 49937 3823
rect 50023 3800 50089 3823
rect 49703 3760 49712 3800
rect 49752 3760 49769 3800
rect 49855 3760 49876 3800
rect 49916 3760 49937 3800
rect 50023 3760 50040 3800
rect 50080 3760 50089 3800
rect 49703 3737 49769 3760
rect 49855 3737 49937 3760
rect 50023 3737 50089 3760
rect 49703 3718 50089 3737
rect 64823 3823 65209 3842
rect 64823 3800 64889 3823
rect 64975 3800 65057 3823
rect 65143 3800 65209 3823
rect 64823 3760 64832 3800
rect 64872 3760 64889 3800
rect 64975 3760 64996 3800
rect 65036 3760 65057 3800
rect 65143 3760 65160 3800
rect 65200 3760 65209 3800
rect 64823 3737 64889 3760
rect 64975 3737 65057 3760
rect 65143 3737 65209 3760
rect 64823 3718 65209 3737
rect 79943 3823 80329 3842
rect 79943 3800 80009 3823
rect 80095 3800 80177 3823
rect 80263 3800 80329 3823
rect 79943 3760 79952 3800
rect 79992 3760 80009 3800
rect 80095 3760 80116 3800
rect 80156 3760 80177 3800
rect 80263 3760 80280 3800
rect 80320 3760 80329 3800
rect 79943 3737 80009 3760
rect 80095 3737 80177 3760
rect 80263 3737 80329 3760
rect 79943 3718 80329 3737
rect 3103 3067 3489 3086
rect 3103 3044 3169 3067
rect 3255 3044 3337 3067
rect 3423 3044 3489 3067
rect 3103 3004 3112 3044
rect 3152 3004 3169 3044
rect 3255 3004 3276 3044
rect 3316 3004 3337 3044
rect 3423 3004 3440 3044
rect 3480 3004 3489 3044
rect 3103 2981 3169 3004
rect 3255 2981 3337 3004
rect 3423 2981 3489 3004
rect 3103 2962 3489 2981
rect 18223 3067 18609 3086
rect 18223 3044 18289 3067
rect 18375 3044 18457 3067
rect 18543 3044 18609 3067
rect 18223 3004 18232 3044
rect 18272 3004 18289 3044
rect 18375 3004 18396 3044
rect 18436 3004 18457 3044
rect 18543 3004 18560 3044
rect 18600 3004 18609 3044
rect 18223 2981 18289 3004
rect 18375 2981 18457 3004
rect 18543 2981 18609 3004
rect 18223 2962 18609 2981
rect 33343 3067 33729 3086
rect 33343 3044 33409 3067
rect 33495 3044 33577 3067
rect 33663 3044 33729 3067
rect 33343 3004 33352 3044
rect 33392 3004 33409 3044
rect 33495 3004 33516 3044
rect 33556 3004 33577 3044
rect 33663 3004 33680 3044
rect 33720 3004 33729 3044
rect 33343 2981 33409 3004
rect 33495 2981 33577 3004
rect 33663 2981 33729 3004
rect 33343 2962 33729 2981
rect 48463 3067 48849 3086
rect 48463 3044 48529 3067
rect 48615 3044 48697 3067
rect 48783 3044 48849 3067
rect 48463 3004 48472 3044
rect 48512 3004 48529 3044
rect 48615 3004 48636 3044
rect 48676 3004 48697 3044
rect 48783 3004 48800 3044
rect 48840 3004 48849 3044
rect 48463 2981 48529 3004
rect 48615 2981 48697 3004
rect 48783 2981 48849 3004
rect 48463 2962 48849 2981
rect 63583 3067 63969 3086
rect 63583 3044 63649 3067
rect 63735 3044 63817 3067
rect 63903 3044 63969 3067
rect 63583 3004 63592 3044
rect 63632 3004 63649 3044
rect 63735 3004 63756 3044
rect 63796 3004 63817 3044
rect 63903 3004 63920 3044
rect 63960 3004 63969 3044
rect 63583 2981 63649 3004
rect 63735 2981 63817 3004
rect 63903 2981 63969 3004
rect 63583 2962 63969 2981
rect 78703 3067 79089 3086
rect 78703 3044 78769 3067
rect 78855 3044 78937 3067
rect 79023 3044 79089 3067
rect 78703 3004 78712 3044
rect 78752 3004 78769 3044
rect 78855 3004 78876 3044
rect 78916 3004 78937 3044
rect 79023 3004 79040 3044
rect 79080 3004 79089 3044
rect 78703 2981 78769 3004
rect 78855 2981 78937 3004
rect 79023 2981 79089 3004
rect 78703 2962 79089 2981
rect 4343 2311 4729 2330
rect 4343 2288 4409 2311
rect 4495 2288 4577 2311
rect 4663 2288 4729 2311
rect 4343 2248 4352 2288
rect 4392 2248 4409 2288
rect 4495 2248 4516 2288
rect 4556 2248 4577 2288
rect 4663 2248 4680 2288
rect 4720 2248 4729 2288
rect 4343 2225 4409 2248
rect 4495 2225 4577 2248
rect 4663 2225 4729 2248
rect 4343 2206 4729 2225
rect 19463 2311 19849 2330
rect 19463 2288 19529 2311
rect 19615 2288 19697 2311
rect 19783 2288 19849 2311
rect 19463 2248 19472 2288
rect 19512 2248 19529 2288
rect 19615 2248 19636 2288
rect 19676 2248 19697 2288
rect 19783 2248 19800 2288
rect 19840 2248 19849 2288
rect 19463 2225 19529 2248
rect 19615 2225 19697 2248
rect 19783 2225 19849 2248
rect 19463 2206 19849 2225
rect 34583 2311 34969 2330
rect 34583 2288 34649 2311
rect 34735 2288 34817 2311
rect 34903 2288 34969 2311
rect 34583 2248 34592 2288
rect 34632 2248 34649 2288
rect 34735 2248 34756 2288
rect 34796 2248 34817 2288
rect 34903 2248 34920 2288
rect 34960 2248 34969 2288
rect 34583 2225 34649 2248
rect 34735 2225 34817 2248
rect 34903 2225 34969 2248
rect 34583 2206 34969 2225
rect 49703 2311 50089 2330
rect 49703 2288 49769 2311
rect 49855 2288 49937 2311
rect 50023 2288 50089 2311
rect 49703 2248 49712 2288
rect 49752 2248 49769 2288
rect 49855 2248 49876 2288
rect 49916 2248 49937 2288
rect 50023 2248 50040 2288
rect 50080 2248 50089 2288
rect 49703 2225 49769 2248
rect 49855 2225 49937 2248
rect 50023 2225 50089 2248
rect 49703 2206 50089 2225
rect 64823 2311 65209 2330
rect 64823 2288 64889 2311
rect 64975 2288 65057 2311
rect 65143 2288 65209 2311
rect 64823 2248 64832 2288
rect 64872 2248 64889 2288
rect 64975 2248 64996 2288
rect 65036 2248 65057 2288
rect 65143 2248 65160 2288
rect 65200 2248 65209 2288
rect 64823 2225 64889 2248
rect 64975 2225 65057 2248
rect 65143 2225 65209 2248
rect 64823 2206 65209 2225
rect 79943 2311 80329 2330
rect 79943 2288 80009 2311
rect 80095 2288 80177 2311
rect 80263 2288 80329 2311
rect 79943 2248 79952 2288
rect 79992 2248 80009 2288
rect 80095 2248 80116 2288
rect 80156 2248 80177 2288
rect 80263 2248 80280 2288
rect 80320 2248 80329 2288
rect 79943 2225 80009 2248
rect 80095 2225 80177 2248
rect 80263 2225 80329 2248
rect 79943 2206 80329 2225
rect 3103 1555 3489 1574
rect 3103 1532 3169 1555
rect 3255 1532 3337 1555
rect 3423 1532 3489 1555
rect 3103 1492 3112 1532
rect 3152 1492 3169 1532
rect 3255 1492 3276 1532
rect 3316 1492 3337 1532
rect 3423 1492 3440 1532
rect 3480 1492 3489 1532
rect 3103 1469 3169 1492
rect 3255 1469 3337 1492
rect 3423 1469 3489 1492
rect 3103 1450 3489 1469
rect 18223 1555 18609 1574
rect 18223 1532 18289 1555
rect 18375 1532 18457 1555
rect 18543 1532 18609 1555
rect 18223 1492 18232 1532
rect 18272 1492 18289 1532
rect 18375 1492 18396 1532
rect 18436 1492 18457 1532
rect 18543 1492 18560 1532
rect 18600 1492 18609 1532
rect 18223 1469 18289 1492
rect 18375 1469 18457 1492
rect 18543 1469 18609 1492
rect 18223 1450 18609 1469
rect 33343 1555 33729 1574
rect 33343 1532 33409 1555
rect 33495 1532 33577 1555
rect 33663 1532 33729 1555
rect 33343 1492 33352 1532
rect 33392 1492 33409 1532
rect 33495 1492 33516 1532
rect 33556 1492 33577 1532
rect 33663 1492 33680 1532
rect 33720 1492 33729 1532
rect 33343 1469 33409 1492
rect 33495 1469 33577 1492
rect 33663 1469 33729 1492
rect 33343 1450 33729 1469
rect 48463 1555 48849 1574
rect 48463 1532 48529 1555
rect 48615 1532 48697 1555
rect 48783 1532 48849 1555
rect 48463 1492 48472 1532
rect 48512 1492 48529 1532
rect 48615 1492 48636 1532
rect 48676 1492 48697 1532
rect 48783 1492 48800 1532
rect 48840 1492 48849 1532
rect 48463 1469 48529 1492
rect 48615 1469 48697 1492
rect 48783 1469 48849 1492
rect 48463 1450 48849 1469
rect 63583 1555 63969 1574
rect 63583 1532 63649 1555
rect 63735 1532 63817 1555
rect 63903 1532 63969 1555
rect 63583 1492 63592 1532
rect 63632 1492 63649 1532
rect 63735 1492 63756 1532
rect 63796 1492 63817 1532
rect 63903 1492 63920 1532
rect 63960 1492 63969 1532
rect 63583 1469 63649 1492
rect 63735 1469 63817 1492
rect 63903 1469 63969 1492
rect 63583 1450 63969 1469
rect 78703 1555 79089 1574
rect 78703 1532 78769 1555
rect 78855 1532 78937 1555
rect 79023 1532 79089 1555
rect 78703 1492 78712 1532
rect 78752 1492 78769 1532
rect 78855 1492 78876 1532
rect 78916 1492 78937 1532
rect 79023 1492 79040 1532
rect 79080 1492 79089 1532
rect 78703 1469 78769 1492
rect 78855 1469 78937 1492
rect 79023 1469 79089 1492
rect 78703 1450 79089 1469
rect 4343 799 4729 818
rect 4343 776 4409 799
rect 4495 776 4577 799
rect 4663 776 4729 799
rect 4343 736 4352 776
rect 4392 736 4409 776
rect 4495 736 4516 776
rect 4556 736 4577 776
rect 4663 736 4680 776
rect 4720 736 4729 776
rect 4343 713 4409 736
rect 4495 713 4577 736
rect 4663 713 4729 736
rect 4343 694 4729 713
rect 19463 799 19849 818
rect 19463 776 19529 799
rect 19615 776 19697 799
rect 19783 776 19849 799
rect 19463 736 19472 776
rect 19512 736 19529 776
rect 19615 736 19636 776
rect 19676 736 19697 776
rect 19783 736 19800 776
rect 19840 736 19849 776
rect 19463 713 19529 736
rect 19615 713 19697 736
rect 19783 713 19849 736
rect 19463 694 19849 713
rect 34583 799 34969 818
rect 34583 776 34649 799
rect 34735 776 34817 799
rect 34903 776 34969 799
rect 34583 736 34592 776
rect 34632 736 34649 776
rect 34735 736 34756 776
rect 34796 736 34817 776
rect 34903 736 34920 776
rect 34960 736 34969 776
rect 34583 713 34649 736
rect 34735 713 34817 736
rect 34903 713 34969 736
rect 34583 694 34969 713
rect 49703 799 50089 818
rect 49703 776 49769 799
rect 49855 776 49937 799
rect 50023 776 50089 799
rect 49703 736 49712 776
rect 49752 736 49769 776
rect 49855 736 49876 776
rect 49916 736 49937 776
rect 50023 736 50040 776
rect 50080 736 50089 776
rect 49703 713 49769 736
rect 49855 713 49937 736
rect 50023 713 50089 736
rect 49703 694 50089 713
rect 64823 799 65209 818
rect 64823 776 64889 799
rect 64975 776 65057 799
rect 65143 776 65209 799
rect 64823 736 64832 776
rect 64872 736 64889 776
rect 64975 736 64996 776
rect 65036 736 65057 776
rect 65143 736 65160 776
rect 65200 736 65209 776
rect 64823 713 64889 736
rect 64975 713 65057 736
rect 65143 713 65209 736
rect 64823 694 65209 713
rect 79943 799 80329 818
rect 79943 776 80009 799
rect 80095 776 80177 799
rect 80263 776 80329 799
rect 79943 736 79952 776
rect 79992 736 80009 776
rect 80095 736 80116 776
rect 80156 736 80177 776
rect 80263 736 80280 776
rect 80320 736 80329 776
rect 79943 713 80009 736
rect 80095 713 80177 736
rect 80263 713 80329 736
rect 79943 694 80329 713
<< via5 >>
rect 4409 38576 4495 38599
rect 4577 38576 4663 38599
rect 4409 38536 4434 38576
rect 4434 38536 4474 38576
rect 4474 38536 4495 38576
rect 4577 38536 4598 38576
rect 4598 38536 4638 38576
rect 4638 38536 4663 38576
rect 4409 38513 4495 38536
rect 4577 38513 4663 38536
rect 19529 38576 19615 38599
rect 19697 38576 19783 38599
rect 19529 38536 19554 38576
rect 19554 38536 19594 38576
rect 19594 38536 19615 38576
rect 19697 38536 19718 38576
rect 19718 38536 19758 38576
rect 19758 38536 19783 38576
rect 19529 38513 19615 38536
rect 19697 38513 19783 38536
rect 34649 38576 34735 38599
rect 34817 38576 34903 38599
rect 34649 38536 34674 38576
rect 34674 38536 34714 38576
rect 34714 38536 34735 38576
rect 34817 38536 34838 38576
rect 34838 38536 34878 38576
rect 34878 38536 34903 38576
rect 34649 38513 34735 38536
rect 34817 38513 34903 38536
rect 49769 38576 49855 38599
rect 49937 38576 50023 38599
rect 49769 38536 49794 38576
rect 49794 38536 49834 38576
rect 49834 38536 49855 38576
rect 49937 38536 49958 38576
rect 49958 38536 49998 38576
rect 49998 38536 50023 38576
rect 49769 38513 49855 38536
rect 49937 38513 50023 38536
rect 64889 38576 64975 38599
rect 65057 38576 65143 38599
rect 64889 38536 64914 38576
rect 64914 38536 64954 38576
rect 64954 38536 64975 38576
rect 65057 38536 65078 38576
rect 65078 38536 65118 38576
rect 65118 38536 65143 38576
rect 64889 38513 64975 38536
rect 65057 38513 65143 38536
rect 80009 38576 80095 38599
rect 80177 38576 80263 38599
rect 80009 38536 80034 38576
rect 80034 38536 80074 38576
rect 80074 38536 80095 38576
rect 80177 38536 80198 38576
rect 80198 38536 80238 38576
rect 80238 38536 80263 38576
rect 80009 38513 80095 38536
rect 80177 38513 80263 38536
rect 3169 37820 3255 37843
rect 3337 37820 3423 37843
rect 3169 37780 3194 37820
rect 3194 37780 3234 37820
rect 3234 37780 3255 37820
rect 3337 37780 3358 37820
rect 3358 37780 3398 37820
rect 3398 37780 3423 37820
rect 3169 37757 3255 37780
rect 3337 37757 3423 37780
rect 18289 37820 18375 37843
rect 18457 37820 18543 37843
rect 18289 37780 18314 37820
rect 18314 37780 18354 37820
rect 18354 37780 18375 37820
rect 18457 37780 18478 37820
rect 18478 37780 18518 37820
rect 18518 37780 18543 37820
rect 18289 37757 18375 37780
rect 18457 37757 18543 37780
rect 33409 37820 33495 37843
rect 33577 37820 33663 37843
rect 33409 37780 33434 37820
rect 33434 37780 33474 37820
rect 33474 37780 33495 37820
rect 33577 37780 33598 37820
rect 33598 37780 33638 37820
rect 33638 37780 33663 37820
rect 33409 37757 33495 37780
rect 33577 37757 33663 37780
rect 48529 37820 48615 37843
rect 48697 37820 48783 37843
rect 48529 37780 48554 37820
rect 48554 37780 48594 37820
rect 48594 37780 48615 37820
rect 48697 37780 48718 37820
rect 48718 37780 48758 37820
rect 48758 37780 48783 37820
rect 48529 37757 48615 37780
rect 48697 37757 48783 37780
rect 63649 37820 63735 37843
rect 63817 37820 63903 37843
rect 63649 37780 63674 37820
rect 63674 37780 63714 37820
rect 63714 37780 63735 37820
rect 63817 37780 63838 37820
rect 63838 37780 63878 37820
rect 63878 37780 63903 37820
rect 63649 37757 63735 37780
rect 63817 37757 63903 37780
rect 78769 37820 78855 37843
rect 78937 37820 79023 37843
rect 78769 37780 78794 37820
rect 78794 37780 78834 37820
rect 78834 37780 78855 37820
rect 78937 37780 78958 37820
rect 78958 37780 78998 37820
rect 78998 37780 79023 37820
rect 78769 37757 78855 37780
rect 78937 37757 79023 37780
rect 4409 37064 4495 37087
rect 4577 37064 4663 37087
rect 4409 37024 4434 37064
rect 4434 37024 4474 37064
rect 4474 37024 4495 37064
rect 4577 37024 4598 37064
rect 4598 37024 4638 37064
rect 4638 37024 4663 37064
rect 4409 37001 4495 37024
rect 4577 37001 4663 37024
rect 19529 37064 19615 37087
rect 19697 37064 19783 37087
rect 19529 37024 19554 37064
rect 19554 37024 19594 37064
rect 19594 37024 19615 37064
rect 19697 37024 19718 37064
rect 19718 37024 19758 37064
rect 19758 37024 19783 37064
rect 19529 37001 19615 37024
rect 19697 37001 19783 37024
rect 34649 37064 34735 37087
rect 34817 37064 34903 37087
rect 34649 37024 34674 37064
rect 34674 37024 34714 37064
rect 34714 37024 34735 37064
rect 34817 37024 34838 37064
rect 34838 37024 34878 37064
rect 34878 37024 34903 37064
rect 34649 37001 34735 37024
rect 34817 37001 34903 37024
rect 49769 37064 49855 37087
rect 49937 37064 50023 37087
rect 49769 37024 49794 37064
rect 49794 37024 49834 37064
rect 49834 37024 49855 37064
rect 49937 37024 49958 37064
rect 49958 37024 49998 37064
rect 49998 37024 50023 37064
rect 49769 37001 49855 37024
rect 49937 37001 50023 37024
rect 64889 37064 64975 37087
rect 65057 37064 65143 37087
rect 64889 37024 64914 37064
rect 64914 37024 64954 37064
rect 64954 37024 64975 37064
rect 65057 37024 65078 37064
rect 65078 37024 65118 37064
rect 65118 37024 65143 37064
rect 64889 37001 64975 37024
rect 65057 37001 65143 37024
rect 80009 37064 80095 37087
rect 80177 37064 80263 37087
rect 80009 37024 80034 37064
rect 80034 37024 80074 37064
rect 80074 37024 80095 37064
rect 80177 37024 80198 37064
rect 80198 37024 80238 37064
rect 80238 37024 80263 37064
rect 80009 37001 80095 37024
rect 80177 37001 80263 37024
rect 3169 36308 3255 36331
rect 3337 36308 3423 36331
rect 3169 36268 3194 36308
rect 3194 36268 3234 36308
rect 3234 36268 3255 36308
rect 3337 36268 3358 36308
rect 3358 36268 3398 36308
rect 3398 36268 3423 36308
rect 3169 36245 3255 36268
rect 3337 36245 3423 36268
rect 18289 36308 18375 36331
rect 18457 36308 18543 36331
rect 18289 36268 18314 36308
rect 18314 36268 18354 36308
rect 18354 36268 18375 36308
rect 18457 36268 18478 36308
rect 18478 36268 18518 36308
rect 18518 36268 18543 36308
rect 18289 36245 18375 36268
rect 18457 36245 18543 36268
rect 33409 36308 33495 36331
rect 33577 36308 33663 36331
rect 33409 36268 33434 36308
rect 33434 36268 33474 36308
rect 33474 36268 33495 36308
rect 33577 36268 33598 36308
rect 33598 36268 33638 36308
rect 33638 36268 33663 36308
rect 33409 36245 33495 36268
rect 33577 36245 33663 36268
rect 48529 36308 48615 36331
rect 48697 36308 48783 36331
rect 48529 36268 48554 36308
rect 48554 36268 48594 36308
rect 48594 36268 48615 36308
rect 48697 36268 48718 36308
rect 48718 36268 48758 36308
rect 48758 36268 48783 36308
rect 48529 36245 48615 36268
rect 48697 36245 48783 36268
rect 63649 36308 63735 36331
rect 63817 36308 63903 36331
rect 63649 36268 63674 36308
rect 63674 36268 63714 36308
rect 63714 36268 63735 36308
rect 63817 36268 63838 36308
rect 63838 36268 63878 36308
rect 63878 36268 63903 36308
rect 63649 36245 63735 36268
rect 63817 36245 63903 36268
rect 78769 36308 78855 36331
rect 78937 36308 79023 36331
rect 78769 36268 78794 36308
rect 78794 36268 78834 36308
rect 78834 36268 78855 36308
rect 78937 36268 78958 36308
rect 78958 36268 78998 36308
rect 78998 36268 79023 36308
rect 78769 36245 78855 36268
rect 78937 36245 79023 36268
rect 4409 35552 4495 35575
rect 4577 35552 4663 35575
rect 4409 35512 4434 35552
rect 4434 35512 4474 35552
rect 4474 35512 4495 35552
rect 4577 35512 4598 35552
rect 4598 35512 4638 35552
rect 4638 35512 4663 35552
rect 4409 35489 4495 35512
rect 4577 35489 4663 35512
rect 19529 35552 19615 35575
rect 19697 35552 19783 35575
rect 19529 35512 19554 35552
rect 19554 35512 19594 35552
rect 19594 35512 19615 35552
rect 19697 35512 19718 35552
rect 19718 35512 19758 35552
rect 19758 35512 19783 35552
rect 19529 35489 19615 35512
rect 19697 35489 19783 35512
rect 34649 35552 34735 35575
rect 34817 35552 34903 35575
rect 34649 35512 34674 35552
rect 34674 35512 34714 35552
rect 34714 35512 34735 35552
rect 34817 35512 34838 35552
rect 34838 35512 34878 35552
rect 34878 35512 34903 35552
rect 34649 35489 34735 35512
rect 34817 35489 34903 35512
rect 49769 35552 49855 35575
rect 49937 35552 50023 35575
rect 49769 35512 49794 35552
rect 49794 35512 49834 35552
rect 49834 35512 49855 35552
rect 49937 35512 49958 35552
rect 49958 35512 49998 35552
rect 49998 35512 50023 35552
rect 49769 35489 49855 35512
rect 49937 35489 50023 35512
rect 64889 35552 64975 35575
rect 65057 35552 65143 35575
rect 64889 35512 64914 35552
rect 64914 35512 64954 35552
rect 64954 35512 64975 35552
rect 65057 35512 65078 35552
rect 65078 35512 65118 35552
rect 65118 35512 65143 35552
rect 64889 35489 64975 35512
rect 65057 35489 65143 35512
rect 80009 35552 80095 35575
rect 80177 35552 80263 35575
rect 80009 35512 80034 35552
rect 80034 35512 80074 35552
rect 80074 35512 80095 35552
rect 80177 35512 80198 35552
rect 80198 35512 80238 35552
rect 80238 35512 80263 35552
rect 80009 35489 80095 35512
rect 80177 35489 80263 35512
rect 3169 34796 3255 34819
rect 3337 34796 3423 34819
rect 3169 34756 3194 34796
rect 3194 34756 3234 34796
rect 3234 34756 3255 34796
rect 3337 34756 3358 34796
rect 3358 34756 3398 34796
rect 3398 34756 3423 34796
rect 3169 34733 3255 34756
rect 3337 34733 3423 34756
rect 18289 34796 18375 34819
rect 18457 34796 18543 34819
rect 18289 34756 18314 34796
rect 18314 34756 18354 34796
rect 18354 34756 18375 34796
rect 18457 34756 18478 34796
rect 18478 34756 18518 34796
rect 18518 34756 18543 34796
rect 18289 34733 18375 34756
rect 18457 34733 18543 34756
rect 33409 34796 33495 34819
rect 33577 34796 33663 34819
rect 33409 34756 33434 34796
rect 33434 34756 33474 34796
rect 33474 34756 33495 34796
rect 33577 34756 33598 34796
rect 33598 34756 33638 34796
rect 33638 34756 33663 34796
rect 33409 34733 33495 34756
rect 33577 34733 33663 34756
rect 48529 34796 48615 34819
rect 48697 34796 48783 34819
rect 48529 34756 48554 34796
rect 48554 34756 48594 34796
rect 48594 34756 48615 34796
rect 48697 34756 48718 34796
rect 48718 34756 48758 34796
rect 48758 34756 48783 34796
rect 48529 34733 48615 34756
rect 48697 34733 48783 34756
rect 63649 34796 63735 34819
rect 63817 34796 63903 34819
rect 63649 34756 63674 34796
rect 63674 34756 63714 34796
rect 63714 34756 63735 34796
rect 63817 34756 63838 34796
rect 63838 34756 63878 34796
rect 63878 34756 63903 34796
rect 63649 34733 63735 34756
rect 63817 34733 63903 34756
rect 78769 34796 78855 34819
rect 78937 34796 79023 34819
rect 78769 34756 78794 34796
rect 78794 34756 78834 34796
rect 78834 34756 78855 34796
rect 78937 34756 78958 34796
rect 78958 34756 78998 34796
rect 78998 34756 79023 34796
rect 78769 34733 78855 34756
rect 78937 34733 79023 34756
rect 4409 34040 4495 34063
rect 4577 34040 4663 34063
rect 4409 34000 4434 34040
rect 4434 34000 4474 34040
rect 4474 34000 4495 34040
rect 4577 34000 4598 34040
rect 4598 34000 4638 34040
rect 4638 34000 4663 34040
rect 4409 33977 4495 34000
rect 4577 33977 4663 34000
rect 19529 34040 19615 34063
rect 19697 34040 19783 34063
rect 19529 34000 19554 34040
rect 19554 34000 19594 34040
rect 19594 34000 19615 34040
rect 19697 34000 19718 34040
rect 19718 34000 19758 34040
rect 19758 34000 19783 34040
rect 19529 33977 19615 34000
rect 19697 33977 19783 34000
rect 34649 34040 34735 34063
rect 34817 34040 34903 34063
rect 34649 34000 34674 34040
rect 34674 34000 34714 34040
rect 34714 34000 34735 34040
rect 34817 34000 34838 34040
rect 34838 34000 34878 34040
rect 34878 34000 34903 34040
rect 34649 33977 34735 34000
rect 34817 33977 34903 34000
rect 49769 34040 49855 34063
rect 49937 34040 50023 34063
rect 49769 34000 49794 34040
rect 49794 34000 49834 34040
rect 49834 34000 49855 34040
rect 49937 34000 49958 34040
rect 49958 34000 49998 34040
rect 49998 34000 50023 34040
rect 49769 33977 49855 34000
rect 49937 33977 50023 34000
rect 64889 34040 64975 34063
rect 65057 34040 65143 34063
rect 64889 34000 64914 34040
rect 64914 34000 64954 34040
rect 64954 34000 64975 34040
rect 65057 34000 65078 34040
rect 65078 34000 65118 34040
rect 65118 34000 65143 34040
rect 64889 33977 64975 34000
rect 65057 33977 65143 34000
rect 80009 34040 80095 34063
rect 80177 34040 80263 34063
rect 80009 34000 80034 34040
rect 80034 34000 80074 34040
rect 80074 34000 80095 34040
rect 80177 34000 80198 34040
rect 80198 34000 80238 34040
rect 80238 34000 80263 34040
rect 80009 33977 80095 34000
rect 80177 33977 80263 34000
rect 3169 33284 3255 33307
rect 3337 33284 3423 33307
rect 3169 33244 3194 33284
rect 3194 33244 3234 33284
rect 3234 33244 3255 33284
rect 3337 33244 3358 33284
rect 3358 33244 3398 33284
rect 3398 33244 3423 33284
rect 3169 33221 3255 33244
rect 3337 33221 3423 33244
rect 18289 33284 18375 33307
rect 18457 33284 18543 33307
rect 18289 33244 18314 33284
rect 18314 33244 18354 33284
rect 18354 33244 18375 33284
rect 18457 33244 18478 33284
rect 18478 33244 18518 33284
rect 18518 33244 18543 33284
rect 18289 33221 18375 33244
rect 18457 33221 18543 33244
rect 33409 33284 33495 33307
rect 33577 33284 33663 33307
rect 33409 33244 33434 33284
rect 33434 33244 33474 33284
rect 33474 33244 33495 33284
rect 33577 33244 33598 33284
rect 33598 33244 33638 33284
rect 33638 33244 33663 33284
rect 33409 33221 33495 33244
rect 33577 33221 33663 33244
rect 48529 33284 48615 33307
rect 48697 33284 48783 33307
rect 48529 33244 48554 33284
rect 48554 33244 48594 33284
rect 48594 33244 48615 33284
rect 48697 33244 48718 33284
rect 48718 33244 48758 33284
rect 48758 33244 48783 33284
rect 48529 33221 48615 33244
rect 48697 33221 48783 33244
rect 63649 33284 63735 33307
rect 63817 33284 63903 33307
rect 63649 33244 63674 33284
rect 63674 33244 63714 33284
rect 63714 33244 63735 33284
rect 63817 33244 63838 33284
rect 63838 33244 63878 33284
rect 63878 33244 63903 33284
rect 63649 33221 63735 33244
rect 63817 33221 63903 33244
rect 78769 33284 78855 33307
rect 78937 33284 79023 33307
rect 78769 33244 78794 33284
rect 78794 33244 78834 33284
rect 78834 33244 78855 33284
rect 78937 33244 78958 33284
rect 78958 33244 78998 33284
rect 78998 33244 79023 33284
rect 78769 33221 78855 33244
rect 78937 33221 79023 33244
rect 4409 32528 4495 32551
rect 4577 32528 4663 32551
rect 4409 32488 4434 32528
rect 4434 32488 4474 32528
rect 4474 32488 4495 32528
rect 4577 32488 4598 32528
rect 4598 32488 4638 32528
rect 4638 32488 4663 32528
rect 4409 32465 4495 32488
rect 4577 32465 4663 32488
rect 19529 32528 19615 32551
rect 19697 32528 19783 32551
rect 19529 32488 19554 32528
rect 19554 32488 19594 32528
rect 19594 32488 19615 32528
rect 19697 32488 19718 32528
rect 19718 32488 19758 32528
rect 19758 32488 19783 32528
rect 19529 32465 19615 32488
rect 19697 32465 19783 32488
rect 34649 32528 34735 32551
rect 34817 32528 34903 32551
rect 34649 32488 34674 32528
rect 34674 32488 34714 32528
rect 34714 32488 34735 32528
rect 34817 32488 34838 32528
rect 34838 32488 34878 32528
rect 34878 32488 34903 32528
rect 34649 32465 34735 32488
rect 34817 32465 34903 32488
rect 49769 32528 49855 32551
rect 49937 32528 50023 32551
rect 49769 32488 49794 32528
rect 49794 32488 49834 32528
rect 49834 32488 49855 32528
rect 49937 32488 49958 32528
rect 49958 32488 49998 32528
rect 49998 32488 50023 32528
rect 49769 32465 49855 32488
rect 49937 32465 50023 32488
rect 64889 32528 64975 32551
rect 65057 32528 65143 32551
rect 64889 32488 64914 32528
rect 64914 32488 64954 32528
rect 64954 32488 64975 32528
rect 65057 32488 65078 32528
rect 65078 32488 65118 32528
rect 65118 32488 65143 32528
rect 64889 32465 64975 32488
rect 65057 32465 65143 32488
rect 80009 32528 80095 32551
rect 80177 32528 80263 32551
rect 80009 32488 80034 32528
rect 80034 32488 80074 32528
rect 80074 32488 80095 32528
rect 80177 32488 80198 32528
rect 80198 32488 80238 32528
rect 80238 32488 80263 32528
rect 80009 32465 80095 32488
rect 80177 32465 80263 32488
rect 3169 31772 3255 31795
rect 3337 31772 3423 31795
rect 3169 31732 3194 31772
rect 3194 31732 3234 31772
rect 3234 31732 3255 31772
rect 3337 31732 3358 31772
rect 3358 31732 3398 31772
rect 3398 31732 3423 31772
rect 3169 31709 3255 31732
rect 3337 31709 3423 31732
rect 18289 31772 18375 31795
rect 18457 31772 18543 31795
rect 18289 31732 18314 31772
rect 18314 31732 18354 31772
rect 18354 31732 18375 31772
rect 18457 31732 18478 31772
rect 18478 31732 18518 31772
rect 18518 31732 18543 31772
rect 18289 31709 18375 31732
rect 18457 31709 18543 31732
rect 33409 31772 33495 31795
rect 33577 31772 33663 31795
rect 33409 31732 33434 31772
rect 33434 31732 33474 31772
rect 33474 31732 33495 31772
rect 33577 31732 33598 31772
rect 33598 31732 33638 31772
rect 33638 31732 33663 31772
rect 33409 31709 33495 31732
rect 33577 31709 33663 31732
rect 48529 31772 48615 31795
rect 48697 31772 48783 31795
rect 48529 31732 48554 31772
rect 48554 31732 48594 31772
rect 48594 31732 48615 31772
rect 48697 31732 48718 31772
rect 48718 31732 48758 31772
rect 48758 31732 48783 31772
rect 48529 31709 48615 31732
rect 48697 31709 48783 31732
rect 63649 31772 63735 31795
rect 63817 31772 63903 31795
rect 63649 31732 63674 31772
rect 63674 31732 63714 31772
rect 63714 31732 63735 31772
rect 63817 31732 63838 31772
rect 63838 31732 63878 31772
rect 63878 31732 63903 31772
rect 63649 31709 63735 31732
rect 63817 31709 63903 31732
rect 78769 31772 78855 31795
rect 78937 31772 79023 31795
rect 78769 31732 78794 31772
rect 78794 31732 78834 31772
rect 78834 31732 78855 31772
rect 78937 31732 78958 31772
rect 78958 31732 78998 31772
rect 78998 31732 79023 31772
rect 78769 31709 78855 31732
rect 78937 31709 79023 31732
rect 4409 31016 4495 31039
rect 4577 31016 4663 31039
rect 4409 30976 4434 31016
rect 4434 30976 4474 31016
rect 4474 30976 4495 31016
rect 4577 30976 4598 31016
rect 4598 30976 4638 31016
rect 4638 30976 4663 31016
rect 4409 30953 4495 30976
rect 4577 30953 4663 30976
rect 19529 31016 19615 31039
rect 19697 31016 19783 31039
rect 19529 30976 19554 31016
rect 19554 30976 19594 31016
rect 19594 30976 19615 31016
rect 19697 30976 19718 31016
rect 19718 30976 19758 31016
rect 19758 30976 19783 31016
rect 19529 30953 19615 30976
rect 19697 30953 19783 30976
rect 34649 31016 34735 31039
rect 34817 31016 34903 31039
rect 34649 30976 34674 31016
rect 34674 30976 34714 31016
rect 34714 30976 34735 31016
rect 34817 30976 34838 31016
rect 34838 30976 34878 31016
rect 34878 30976 34903 31016
rect 34649 30953 34735 30976
rect 34817 30953 34903 30976
rect 49769 31016 49855 31039
rect 49937 31016 50023 31039
rect 49769 30976 49794 31016
rect 49794 30976 49834 31016
rect 49834 30976 49855 31016
rect 49937 30976 49958 31016
rect 49958 30976 49998 31016
rect 49998 30976 50023 31016
rect 49769 30953 49855 30976
rect 49937 30953 50023 30976
rect 64889 31016 64975 31039
rect 65057 31016 65143 31039
rect 64889 30976 64914 31016
rect 64914 30976 64954 31016
rect 64954 30976 64975 31016
rect 65057 30976 65078 31016
rect 65078 30976 65118 31016
rect 65118 30976 65143 31016
rect 64889 30953 64975 30976
rect 65057 30953 65143 30976
rect 80009 31016 80095 31039
rect 80177 31016 80263 31039
rect 80009 30976 80034 31016
rect 80034 30976 80074 31016
rect 80074 30976 80095 31016
rect 80177 30976 80198 31016
rect 80198 30976 80238 31016
rect 80238 30976 80263 31016
rect 80009 30953 80095 30976
rect 80177 30953 80263 30976
rect 3169 30260 3255 30283
rect 3337 30260 3423 30283
rect 3169 30220 3194 30260
rect 3194 30220 3234 30260
rect 3234 30220 3255 30260
rect 3337 30220 3358 30260
rect 3358 30220 3398 30260
rect 3398 30220 3423 30260
rect 3169 30197 3255 30220
rect 3337 30197 3423 30220
rect 18289 30260 18375 30283
rect 18457 30260 18543 30283
rect 18289 30220 18314 30260
rect 18314 30220 18354 30260
rect 18354 30220 18375 30260
rect 18457 30220 18478 30260
rect 18478 30220 18518 30260
rect 18518 30220 18543 30260
rect 18289 30197 18375 30220
rect 18457 30197 18543 30220
rect 33409 30260 33495 30283
rect 33577 30260 33663 30283
rect 33409 30220 33434 30260
rect 33434 30220 33474 30260
rect 33474 30220 33495 30260
rect 33577 30220 33598 30260
rect 33598 30220 33638 30260
rect 33638 30220 33663 30260
rect 33409 30197 33495 30220
rect 33577 30197 33663 30220
rect 48529 30260 48615 30283
rect 48697 30260 48783 30283
rect 48529 30220 48554 30260
rect 48554 30220 48594 30260
rect 48594 30220 48615 30260
rect 48697 30220 48718 30260
rect 48718 30220 48758 30260
rect 48758 30220 48783 30260
rect 48529 30197 48615 30220
rect 48697 30197 48783 30220
rect 63649 30260 63735 30283
rect 63817 30260 63903 30283
rect 63649 30220 63674 30260
rect 63674 30220 63714 30260
rect 63714 30220 63735 30260
rect 63817 30220 63838 30260
rect 63838 30220 63878 30260
rect 63878 30220 63903 30260
rect 63649 30197 63735 30220
rect 63817 30197 63903 30220
rect 78769 30260 78855 30283
rect 78937 30260 79023 30283
rect 78769 30220 78794 30260
rect 78794 30220 78834 30260
rect 78834 30220 78855 30260
rect 78937 30220 78958 30260
rect 78958 30220 78998 30260
rect 78998 30220 79023 30260
rect 78769 30197 78855 30220
rect 78937 30197 79023 30220
rect 4409 29504 4495 29527
rect 4577 29504 4663 29527
rect 4409 29464 4434 29504
rect 4434 29464 4474 29504
rect 4474 29464 4495 29504
rect 4577 29464 4598 29504
rect 4598 29464 4638 29504
rect 4638 29464 4663 29504
rect 4409 29441 4495 29464
rect 4577 29441 4663 29464
rect 19529 29504 19615 29527
rect 19697 29504 19783 29527
rect 19529 29464 19554 29504
rect 19554 29464 19594 29504
rect 19594 29464 19615 29504
rect 19697 29464 19718 29504
rect 19718 29464 19758 29504
rect 19758 29464 19783 29504
rect 19529 29441 19615 29464
rect 19697 29441 19783 29464
rect 34649 29504 34735 29527
rect 34817 29504 34903 29527
rect 34649 29464 34674 29504
rect 34674 29464 34714 29504
rect 34714 29464 34735 29504
rect 34817 29464 34838 29504
rect 34838 29464 34878 29504
rect 34878 29464 34903 29504
rect 34649 29441 34735 29464
rect 34817 29441 34903 29464
rect 49769 29504 49855 29527
rect 49937 29504 50023 29527
rect 49769 29464 49794 29504
rect 49794 29464 49834 29504
rect 49834 29464 49855 29504
rect 49937 29464 49958 29504
rect 49958 29464 49998 29504
rect 49998 29464 50023 29504
rect 49769 29441 49855 29464
rect 49937 29441 50023 29464
rect 64889 29504 64975 29527
rect 65057 29504 65143 29527
rect 64889 29464 64914 29504
rect 64914 29464 64954 29504
rect 64954 29464 64975 29504
rect 65057 29464 65078 29504
rect 65078 29464 65118 29504
rect 65118 29464 65143 29504
rect 64889 29441 64975 29464
rect 65057 29441 65143 29464
rect 80009 29504 80095 29527
rect 80177 29504 80263 29527
rect 80009 29464 80034 29504
rect 80034 29464 80074 29504
rect 80074 29464 80095 29504
rect 80177 29464 80198 29504
rect 80198 29464 80238 29504
rect 80238 29464 80263 29504
rect 80009 29441 80095 29464
rect 80177 29441 80263 29464
rect 3169 28748 3255 28771
rect 3337 28748 3423 28771
rect 3169 28708 3194 28748
rect 3194 28708 3234 28748
rect 3234 28708 3255 28748
rect 3337 28708 3358 28748
rect 3358 28708 3398 28748
rect 3398 28708 3423 28748
rect 3169 28685 3255 28708
rect 3337 28685 3423 28708
rect 18289 28748 18375 28771
rect 18457 28748 18543 28771
rect 18289 28708 18314 28748
rect 18314 28708 18354 28748
rect 18354 28708 18375 28748
rect 18457 28708 18478 28748
rect 18478 28708 18518 28748
rect 18518 28708 18543 28748
rect 18289 28685 18375 28708
rect 18457 28685 18543 28708
rect 33409 28748 33495 28771
rect 33577 28748 33663 28771
rect 33409 28708 33434 28748
rect 33434 28708 33474 28748
rect 33474 28708 33495 28748
rect 33577 28708 33598 28748
rect 33598 28708 33638 28748
rect 33638 28708 33663 28748
rect 33409 28685 33495 28708
rect 33577 28685 33663 28708
rect 48529 28748 48615 28771
rect 48697 28748 48783 28771
rect 48529 28708 48554 28748
rect 48554 28708 48594 28748
rect 48594 28708 48615 28748
rect 48697 28708 48718 28748
rect 48718 28708 48758 28748
rect 48758 28708 48783 28748
rect 48529 28685 48615 28708
rect 48697 28685 48783 28708
rect 63649 28748 63735 28771
rect 63817 28748 63903 28771
rect 63649 28708 63674 28748
rect 63674 28708 63714 28748
rect 63714 28708 63735 28748
rect 63817 28708 63838 28748
rect 63838 28708 63878 28748
rect 63878 28708 63903 28748
rect 63649 28685 63735 28708
rect 63817 28685 63903 28708
rect 78769 28748 78855 28771
rect 78937 28748 79023 28771
rect 78769 28708 78794 28748
rect 78794 28708 78834 28748
rect 78834 28708 78855 28748
rect 78937 28708 78958 28748
rect 78958 28708 78998 28748
rect 78998 28708 79023 28748
rect 78769 28685 78855 28708
rect 78937 28685 79023 28708
rect 4409 27992 4495 28015
rect 4577 27992 4663 28015
rect 4409 27952 4434 27992
rect 4434 27952 4474 27992
rect 4474 27952 4495 27992
rect 4577 27952 4598 27992
rect 4598 27952 4638 27992
rect 4638 27952 4663 27992
rect 4409 27929 4495 27952
rect 4577 27929 4663 27952
rect 19529 27992 19615 28015
rect 19697 27992 19783 28015
rect 19529 27952 19554 27992
rect 19554 27952 19594 27992
rect 19594 27952 19615 27992
rect 19697 27952 19718 27992
rect 19718 27952 19758 27992
rect 19758 27952 19783 27992
rect 19529 27929 19615 27952
rect 19697 27929 19783 27952
rect 34649 27992 34735 28015
rect 34817 27992 34903 28015
rect 34649 27952 34674 27992
rect 34674 27952 34714 27992
rect 34714 27952 34735 27992
rect 34817 27952 34838 27992
rect 34838 27952 34878 27992
rect 34878 27952 34903 27992
rect 34649 27929 34735 27952
rect 34817 27929 34903 27952
rect 49769 27992 49855 28015
rect 49937 27992 50023 28015
rect 49769 27952 49794 27992
rect 49794 27952 49834 27992
rect 49834 27952 49855 27992
rect 49937 27952 49958 27992
rect 49958 27952 49998 27992
rect 49998 27952 50023 27992
rect 49769 27929 49855 27952
rect 49937 27929 50023 27952
rect 64889 27992 64975 28015
rect 65057 27992 65143 28015
rect 64889 27952 64914 27992
rect 64914 27952 64954 27992
rect 64954 27952 64975 27992
rect 65057 27952 65078 27992
rect 65078 27952 65118 27992
rect 65118 27952 65143 27992
rect 64889 27929 64975 27952
rect 65057 27929 65143 27952
rect 80009 27992 80095 28015
rect 80177 27992 80263 28015
rect 80009 27952 80034 27992
rect 80034 27952 80074 27992
rect 80074 27952 80095 27992
rect 80177 27952 80198 27992
rect 80198 27952 80238 27992
rect 80238 27952 80263 27992
rect 80009 27929 80095 27952
rect 80177 27929 80263 27952
rect 3169 27236 3255 27259
rect 3337 27236 3423 27259
rect 3169 27196 3194 27236
rect 3194 27196 3234 27236
rect 3234 27196 3255 27236
rect 3337 27196 3358 27236
rect 3358 27196 3398 27236
rect 3398 27196 3423 27236
rect 3169 27173 3255 27196
rect 3337 27173 3423 27196
rect 18289 27236 18375 27259
rect 18457 27236 18543 27259
rect 18289 27196 18314 27236
rect 18314 27196 18354 27236
rect 18354 27196 18375 27236
rect 18457 27196 18478 27236
rect 18478 27196 18518 27236
rect 18518 27196 18543 27236
rect 18289 27173 18375 27196
rect 18457 27173 18543 27196
rect 33409 27236 33495 27259
rect 33577 27236 33663 27259
rect 33409 27196 33434 27236
rect 33434 27196 33474 27236
rect 33474 27196 33495 27236
rect 33577 27196 33598 27236
rect 33598 27196 33638 27236
rect 33638 27196 33663 27236
rect 33409 27173 33495 27196
rect 33577 27173 33663 27196
rect 48529 27236 48615 27259
rect 48697 27236 48783 27259
rect 48529 27196 48554 27236
rect 48554 27196 48594 27236
rect 48594 27196 48615 27236
rect 48697 27196 48718 27236
rect 48718 27196 48758 27236
rect 48758 27196 48783 27236
rect 48529 27173 48615 27196
rect 48697 27173 48783 27196
rect 63649 27236 63735 27259
rect 63817 27236 63903 27259
rect 63649 27196 63674 27236
rect 63674 27196 63714 27236
rect 63714 27196 63735 27236
rect 63817 27196 63838 27236
rect 63838 27196 63878 27236
rect 63878 27196 63903 27236
rect 63649 27173 63735 27196
rect 63817 27173 63903 27196
rect 78769 27236 78855 27259
rect 78937 27236 79023 27259
rect 78769 27196 78794 27236
rect 78794 27196 78834 27236
rect 78834 27196 78855 27236
rect 78937 27196 78958 27236
rect 78958 27196 78998 27236
rect 78998 27196 79023 27236
rect 78769 27173 78855 27196
rect 78937 27173 79023 27196
rect 4409 26480 4495 26503
rect 4577 26480 4663 26503
rect 4409 26440 4434 26480
rect 4434 26440 4474 26480
rect 4474 26440 4495 26480
rect 4577 26440 4598 26480
rect 4598 26440 4638 26480
rect 4638 26440 4663 26480
rect 4409 26417 4495 26440
rect 4577 26417 4663 26440
rect 19529 26480 19615 26503
rect 19697 26480 19783 26503
rect 19529 26440 19554 26480
rect 19554 26440 19594 26480
rect 19594 26440 19615 26480
rect 19697 26440 19718 26480
rect 19718 26440 19758 26480
rect 19758 26440 19783 26480
rect 19529 26417 19615 26440
rect 19697 26417 19783 26440
rect 34649 26480 34735 26503
rect 34817 26480 34903 26503
rect 34649 26440 34674 26480
rect 34674 26440 34714 26480
rect 34714 26440 34735 26480
rect 34817 26440 34838 26480
rect 34838 26440 34878 26480
rect 34878 26440 34903 26480
rect 34649 26417 34735 26440
rect 34817 26417 34903 26440
rect 49769 26480 49855 26503
rect 49937 26480 50023 26503
rect 49769 26440 49794 26480
rect 49794 26440 49834 26480
rect 49834 26440 49855 26480
rect 49937 26440 49958 26480
rect 49958 26440 49998 26480
rect 49998 26440 50023 26480
rect 49769 26417 49855 26440
rect 49937 26417 50023 26440
rect 64889 26480 64975 26503
rect 65057 26480 65143 26503
rect 64889 26440 64914 26480
rect 64914 26440 64954 26480
rect 64954 26440 64975 26480
rect 65057 26440 65078 26480
rect 65078 26440 65118 26480
rect 65118 26440 65143 26480
rect 64889 26417 64975 26440
rect 65057 26417 65143 26440
rect 80009 26480 80095 26503
rect 80177 26480 80263 26503
rect 80009 26440 80034 26480
rect 80034 26440 80074 26480
rect 80074 26440 80095 26480
rect 80177 26440 80198 26480
rect 80198 26440 80238 26480
rect 80238 26440 80263 26480
rect 80009 26417 80095 26440
rect 80177 26417 80263 26440
rect 3169 25724 3255 25747
rect 3337 25724 3423 25747
rect 3169 25684 3194 25724
rect 3194 25684 3234 25724
rect 3234 25684 3255 25724
rect 3337 25684 3358 25724
rect 3358 25684 3398 25724
rect 3398 25684 3423 25724
rect 3169 25661 3255 25684
rect 3337 25661 3423 25684
rect 18289 25724 18375 25747
rect 18457 25724 18543 25747
rect 18289 25684 18314 25724
rect 18314 25684 18354 25724
rect 18354 25684 18375 25724
rect 18457 25684 18478 25724
rect 18478 25684 18518 25724
rect 18518 25684 18543 25724
rect 18289 25661 18375 25684
rect 18457 25661 18543 25684
rect 33409 25724 33495 25747
rect 33577 25724 33663 25747
rect 33409 25684 33434 25724
rect 33434 25684 33474 25724
rect 33474 25684 33495 25724
rect 33577 25684 33598 25724
rect 33598 25684 33638 25724
rect 33638 25684 33663 25724
rect 33409 25661 33495 25684
rect 33577 25661 33663 25684
rect 48529 25724 48615 25747
rect 48697 25724 48783 25747
rect 48529 25684 48554 25724
rect 48554 25684 48594 25724
rect 48594 25684 48615 25724
rect 48697 25684 48718 25724
rect 48718 25684 48758 25724
rect 48758 25684 48783 25724
rect 48529 25661 48615 25684
rect 48697 25661 48783 25684
rect 63649 25724 63735 25747
rect 63817 25724 63903 25747
rect 63649 25684 63674 25724
rect 63674 25684 63714 25724
rect 63714 25684 63735 25724
rect 63817 25684 63838 25724
rect 63838 25684 63878 25724
rect 63878 25684 63903 25724
rect 63649 25661 63735 25684
rect 63817 25661 63903 25684
rect 78769 25724 78855 25747
rect 78937 25724 79023 25747
rect 78769 25684 78794 25724
rect 78794 25684 78834 25724
rect 78834 25684 78855 25724
rect 78937 25684 78958 25724
rect 78958 25684 78998 25724
rect 78998 25684 79023 25724
rect 78769 25661 78855 25684
rect 78937 25661 79023 25684
rect 4409 24968 4495 24991
rect 4577 24968 4663 24991
rect 4409 24928 4434 24968
rect 4434 24928 4474 24968
rect 4474 24928 4495 24968
rect 4577 24928 4598 24968
rect 4598 24928 4638 24968
rect 4638 24928 4663 24968
rect 4409 24905 4495 24928
rect 4577 24905 4663 24928
rect 19529 24968 19615 24991
rect 19697 24968 19783 24991
rect 19529 24928 19554 24968
rect 19554 24928 19594 24968
rect 19594 24928 19615 24968
rect 19697 24928 19718 24968
rect 19718 24928 19758 24968
rect 19758 24928 19783 24968
rect 19529 24905 19615 24928
rect 19697 24905 19783 24928
rect 34649 24968 34735 24991
rect 34817 24968 34903 24991
rect 34649 24928 34674 24968
rect 34674 24928 34714 24968
rect 34714 24928 34735 24968
rect 34817 24928 34838 24968
rect 34838 24928 34878 24968
rect 34878 24928 34903 24968
rect 34649 24905 34735 24928
rect 34817 24905 34903 24928
rect 49769 24968 49855 24991
rect 49937 24968 50023 24991
rect 49769 24928 49794 24968
rect 49794 24928 49834 24968
rect 49834 24928 49855 24968
rect 49937 24928 49958 24968
rect 49958 24928 49998 24968
rect 49998 24928 50023 24968
rect 49769 24905 49855 24928
rect 49937 24905 50023 24928
rect 64889 24968 64975 24991
rect 65057 24968 65143 24991
rect 64889 24928 64914 24968
rect 64914 24928 64954 24968
rect 64954 24928 64975 24968
rect 65057 24928 65078 24968
rect 65078 24928 65118 24968
rect 65118 24928 65143 24968
rect 64889 24905 64975 24928
rect 65057 24905 65143 24928
rect 80009 24968 80095 24991
rect 80177 24968 80263 24991
rect 80009 24928 80034 24968
rect 80034 24928 80074 24968
rect 80074 24928 80095 24968
rect 80177 24928 80198 24968
rect 80198 24928 80238 24968
rect 80238 24928 80263 24968
rect 80009 24905 80095 24928
rect 80177 24905 80263 24928
rect 3169 24212 3255 24235
rect 3337 24212 3423 24235
rect 3169 24172 3194 24212
rect 3194 24172 3234 24212
rect 3234 24172 3255 24212
rect 3337 24172 3358 24212
rect 3358 24172 3398 24212
rect 3398 24172 3423 24212
rect 3169 24149 3255 24172
rect 3337 24149 3423 24172
rect 18289 24212 18375 24235
rect 18457 24212 18543 24235
rect 18289 24172 18314 24212
rect 18314 24172 18354 24212
rect 18354 24172 18375 24212
rect 18457 24172 18478 24212
rect 18478 24172 18518 24212
rect 18518 24172 18543 24212
rect 18289 24149 18375 24172
rect 18457 24149 18543 24172
rect 33409 24212 33495 24235
rect 33577 24212 33663 24235
rect 33409 24172 33434 24212
rect 33434 24172 33474 24212
rect 33474 24172 33495 24212
rect 33577 24172 33598 24212
rect 33598 24172 33638 24212
rect 33638 24172 33663 24212
rect 33409 24149 33495 24172
rect 33577 24149 33663 24172
rect 48529 24212 48615 24235
rect 48697 24212 48783 24235
rect 48529 24172 48554 24212
rect 48554 24172 48594 24212
rect 48594 24172 48615 24212
rect 48697 24172 48718 24212
rect 48718 24172 48758 24212
rect 48758 24172 48783 24212
rect 48529 24149 48615 24172
rect 48697 24149 48783 24172
rect 63649 24212 63735 24235
rect 63817 24212 63903 24235
rect 63649 24172 63674 24212
rect 63674 24172 63714 24212
rect 63714 24172 63735 24212
rect 63817 24172 63838 24212
rect 63838 24172 63878 24212
rect 63878 24172 63903 24212
rect 63649 24149 63735 24172
rect 63817 24149 63903 24172
rect 78769 24212 78855 24235
rect 78937 24212 79023 24235
rect 78769 24172 78794 24212
rect 78794 24172 78834 24212
rect 78834 24172 78855 24212
rect 78937 24172 78958 24212
rect 78958 24172 78998 24212
rect 78998 24172 79023 24212
rect 78769 24149 78855 24172
rect 78937 24149 79023 24172
rect 4409 23456 4495 23479
rect 4577 23456 4663 23479
rect 4409 23416 4434 23456
rect 4434 23416 4474 23456
rect 4474 23416 4495 23456
rect 4577 23416 4598 23456
rect 4598 23416 4638 23456
rect 4638 23416 4663 23456
rect 4409 23393 4495 23416
rect 4577 23393 4663 23416
rect 19529 23456 19615 23479
rect 19697 23456 19783 23479
rect 19529 23416 19554 23456
rect 19554 23416 19594 23456
rect 19594 23416 19615 23456
rect 19697 23416 19718 23456
rect 19718 23416 19758 23456
rect 19758 23416 19783 23456
rect 19529 23393 19615 23416
rect 19697 23393 19783 23416
rect 34649 23456 34735 23479
rect 34817 23456 34903 23479
rect 34649 23416 34674 23456
rect 34674 23416 34714 23456
rect 34714 23416 34735 23456
rect 34817 23416 34838 23456
rect 34838 23416 34878 23456
rect 34878 23416 34903 23456
rect 34649 23393 34735 23416
rect 34817 23393 34903 23416
rect 49769 23456 49855 23479
rect 49937 23456 50023 23479
rect 49769 23416 49794 23456
rect 49794 23416 49834 23456
rect 49834 23416 49855 23456
rect 49937 23416 49958 23456
rect 49958 23416 49998 23456
rect 49998 23416 50023 23456
rect 49769 23393 49855 23416
rect 49937 23393 50023 23416
rect 64889 23456 64975 23479
rect 65057 23456 65143 23479
rect 64889 23416 64914 23456
rect 64914 23416 64954 23456
rect 64954 23416 64975 23456
rect 65057 23416 65078 23456
rect 65078 23416 65118 23456
rect 65118 23416 65143 23456
rect 64889 23393 64975 23416
rect 65057 23393 65143 23416
rect 80009 23456 80095 23479
rect 80177 23456 80263 23479
rect 80009 23416 80034 23456
rect 80034 23416 80074 23456
rect 80074 23416 80095 23456
rect 80177 23416 80198 23456
rect 80198 23416 80238 23456
rect 80238 23416 80263 23456
rect 80009 23393 80095 23416
rect 80177 23393 80263 23416
rect 3169 22700 3255 22723
rect 3337 22700 3423 22723
rect 3169 22660 3194 22700
rect 3194 22660 3234 22700
rect 3234 22660 3255 22700
rect 3337 22660 3358 22700
rect 3358 22660 3398 22700
rect 3398 22660 3423 22700
rect 3169 22637 3255 22660
rect 3337 22637 3423 22660
rect 18289 22700 18375 22723
rect 18457 22700 18543 22723
rect 18289 22660 18314 22700
rect 18314 22660 18354 22700
rect 18354 22660 18375 22700
rect 18457 22660 18478 22700
rect 18478 22660 18518 22700
rect 18518 22660 18543 22700
rect 18289 22637 18375 22660
rect 18457 22637 18543 22660
rect 33409 22700 33495 22723
rect 33577 22700 33663 22723
rect 33409 22660 33434 22700
rect 33434 22660 33474 22700
rect 33474 22660 33495 22700
rect 33577 22660 33598 22700
rect 33598 22660 33638 22700
rect 33638 22660 33663 22700
rect 33409 22637 33495 22660
rect 33577 22637 33663 22660
rect 48529 22700 48615 22723
rect 48697 22700 48783 22723
rect 48529 22660 48554 22700
rect 48554 22660 48594 22700
rect 48594 22660 48615 22700
rect 48697 22660 48718 22700
rect 48718 22660 48758 22700
rect 48758 22660 48783 22700
rect 48529 22637 48615 22660
rect 48697 22637 48783 22660
rect 63649 22700 63735 22723
rect 63817 22700 63903 22723
rect 63649 22660 63674 22700
rect 63674 22660 63714 22700
rect 63714 22660 63735 22700
rect 63817 22660 63838 22700
rect 63838 22660 63878 22700
rect 63878 22660 63903 22700
rect 63649 22637 63735 22660
rect 63817 22637 63903 22660
rect 78769 22700 78855 22723
rect 78937 22700 79023 22723
rect 78769 22660 78794 22700
rect 78794 22660 78834 22700
rect 78834 22660 78855 22700
rect 78937 22660 78958 22700
rect 78958 22660 78998 22700
rect 78998 22660 79023 22700
rect 78769 22637 78855 22660
rect 78937 22637 79023 22660
rect 4409 21944 4495 21967
rect 4577 21944 4663 21967
rect 4409 21904 4434 21944
rect 4434 21904 4474 21944
rect 4474 21904 4495 21944
rect 4577 21904 4598 21944
rect 4598 21904 4638 21944
rect 4638 21904 4663 21944
rect 4409 21881 4495 21904
rect 4577 21881 4663 21904
rect 19529 21944 19615 21967
rect 19697 21944 19783 21967
rect 19529 21904 19554 21944
rect 19554 21904 19594 21944
rect 19594 21904 19615 21944
rect 19697 21904 19718 21944
rect 19718 21904 19758 21944
rect 19758 21904 19783 21944
rect 19529 21881 19615 21904
rect 19697 21881 19783 21904
rect 34649 21944 34735 21967
rect 34817 21944 34903 21967
rect 34649 21904 34674 21944
rect 34674 21904 34714 21944
rect 34714 21904 34735 21944
rect 34817 21904 34838 21944
rect 34838 21904 34878 21944
rect 34878 21904 34903 21944
rect 34649 21881 34735 21904
rect 34817 21881 34903 21904
rect 49769 21944 49855 21967
rect 49937 21944 50023 21967
rect 49769 21904 49794 21944
rect 49794 21904 49834 21944
rect 49834 21904 49855 21944
rect 49937 21904 49958 21944
rect 49958 21904 49998 21944
rect 49998 21904 50023 21944
rect 49769 21881 49855 21904
rect 49937 21881 50023 21904
rect 64889 21944 64975 21967
rect 65057 21944 65143 21967
rect 64889 21904 64914 21944
rect 64914 21904 64954 21944
rect 64954 21904 64975 21944
rect 65057 21904 65078 21944
rect 65078 21904 65118 21944
rect 65118 21904 65143 21944
rect 64889 21881 64975 21904
rect 65057 21881 65143 21904
rect 80009 21944 80095 21967
rect 80177 21944 80263 21967
rect 80009 21904 80034 21944
rect 80034 21904 80074 21944
rect 80074 21904 80095 21944
rect 80177 21904 80198 21944
rect 80198 21904 80238 21944
rect 80238 21904 80263 21944
rect 80009 21881 80095 21904
rect 80177 21881 80263 21904
rect 3169 21188 3255 21211
rect 3337 21188 3423 21211
rect 3169 21148 3194 21188
rect 3194 21148 3234 21188
rect 3234 21148 3255 21188
rect 3337 21148 3358 21188
rect 3358 21148 3398 21188
rect 3398 21148 3423 21188
rect 3169 21125 3255 21148
rect 3337 21125 3423 21148
rect 18289 21188 18375 21211
rect 18457 21188 18543 21211
rect 18289 21148 18314 21188
rect 18314 21148 18354 21188
rect 18354 21148 18375 21188
rect 18457 21148 18478 21188
rect 18478 21148 18518 21188
rect 18518 21148 18543 21188
rect 18289 21125 18375 21148
rect 18457 21125 18543 21148
rect 33409 21188 33495 21211
rect 33577 21188 33663 21211
rect 33409 21148 33434 21188
rect 33434 21148 33474 21188
rect 33474 21148 33495 21188
rect 33577 21148 33598 21188
rect 33598 21148 33638 21188
rect 33638 21148 33663 21188
rect 33409 21125 33495 21148
rect 33577 21125 33663 21148
rect 48529 21188 48615 21211
rect 48697 21188 48783 21211
rect 48529 21148 48554 21188
rect 48554 21148 48594 21188
rect 48594 21148 48615 21188
rect 48697 21148 48718 21188
rect 48718 21148 48758 21188
rect 48758 21148 48783 21188
rect 48529 21125 48615 21148
rect 48697 21125 48783 21148
rect 63649 21188 63735 21211
rect 63817 21188 63903 21211
rect 63649 21148 63674 21188
rect 63674 21148 63714 21188
rect 63714 21148 63735 21188
rect 63817 21148 63838 21188
rect 63838 21148 63878 21188
rect 63878 21148 63903 21188
rect 63649 21125 63735 21148
rect 63817 21125 63903 21148
rect 78769 21188 78855 21211
rect 78937 21188 79023 21211
rect 78769 21148 78794 21188
rect 78794 21148 78834 21188
rect 78834 21148 78855 21188
rect 78937 21148 78958 21188
rect 78958 21148 78998 21188
rect 78998 21148 79023 21188
rect 78769 21125 78855 21148
rect 78937 21125 79023 21148
rect 4409 20432 4495 20455
rect 4577 20432 4663 20455
rect 4409 20392 4434 20432
rect 4434 20392 4474 20432
rect 4474 20392 4495 20432
rect 4577 20392 4598 20432
rect 4598 20392 4638 20432
rect 4638 20392 4663 20432
rect 4409 20369 4495 20392
rect 4577 20369 4663 20392
rect 19529 20432 19615 20455
rect 19697 20432 19783 20455
rect 19529 20392 19554 20432
rect 19554 20392 19594 20432
rect 19594 20392 19615 20432
rect 19697 20392 19718 20432
rect 19718 20392 19758 20432
rect 19758 20392 19783 20432
rect 19529 20369 19615 20392
rect 19697 20369 19783 20392
rect 34649 20432 34735 20455
rect 34817 20432 34903 20455
rect 34649 20392 34674 20432
rect 34674 20392 34714 20432
rect 34714 20392 34735 20432
rect 34817 20392 34838 20432
rect 34838 20392 34878 20432
rect 34878 20392 34903 20432
rect 34649 20369 34735 20392
rect 34817 20369 34903 20392
rect 49769 20432 49855 20455
rect 49937 20432 50023 20455
rect 49769 20392 49794 20432
rect 49794 20392 49834 20432
rect 49834 20392 49855 20432
rect 49937 20392 49958 20432
rect 49958 20392 49998 20432
rect 49998 20392 50023 20432
rect 49769 20369 49855 20392
rect 49937 20369 50023 20392
rect 64889 20432 64975 20455
rect 65057 20432 65143 20455
rect 64889 20392 64914 20432
rect 64914 20392 64954 20432
rect 64954 20392 64975 20432
rect 65057 20392 65078 20432
rect 65078 20392 65118 20432
rect 65118 20392 65143 20432
rect 64889 20369 64975 20392
rect 65057 20369 65143 20392
rect 80009 20432 80095 20455
rect 80177 20432 80263 20455
rect 80009 20392 80034 20432
rect 80034 20392 80074 20432
rect 80074 20392 80095 20432
rect 80177 20392 80198 20432
rect 80198 20392 80238 20432
rect 80238 20392 80263 20432
rect 80009 20369 80095 20392
rect 80177 20369 80263 20392
rect 3169 19676 3255 19699
rect 3337 19676 3423 19699
rect 3169 19636 3194 19676
rect 3194 19636 3234 19676
rect 3234 19636 3255 19676
rect 3337 19636 3358 19676
rect 3358 19636 3398 19676
rect 3398 19636 3423 19676
rect 3169 19613 3255 19636
rect 3337 19613 3423 19636
rect 18289 19676 18375 19699
rect 18457 19676 18543 19699
rect 18289 19636 18314 19676
rect 18314 19636 18354 19676
rect 18354 19636 18375 19676
rect 18457 19636 18478 19676
rect 18478 19636 18518 19676
rect 18518 19636 18543 19676
rect 18289 19613 18375 19636
rect 18457 19613 18543 19636
rect 33409 19676 33495 19699
rect 33577 19676 33663 19699
rect 33409 19636 33434 19676
rect 33434 19636 33474 19676
rect 33474 19636 33495 19676
rect 33577 19636 33598 19676
rect 33598 19636 33638 19676
rect 33638 19636 33663 19676
rect 33409 19613 33495 19636
rect 33577 19613 33663 19636
rect 48529 19676 48615 19699
rect 48697 19676 48783 19699
rect 48529 19636 48554 19676
rect 48554 19636 48594 19676
rect 48594 19636 48615 19676
rect 48697 19636 48718 19676
rect 48718 19636 48758 19676
rect 48758 19636 48783 19676
rect 48529 19613 48615 19636
rect 48697 19613 48783 19636
rect 63649 19676 63735 19699
rect 63817 19676 63903 19699
rect 63649 19636 63674 19676
rect 63674 19636 63714 19676
rect 63714 19636 63735 19676
rect 63817 19636 63838 19676
rect 63838 19636 63878 19676
rect 63878 19636 63903 19676
rect 63649 19613 63735 19636
rect 63817 19613 63903 19636
rect 78769 19676 78855 19699
rect 78937 19676 79023 19699
rect 78769 19636 78794 19676
rect 78794 19636 78834 19676
rect 78834 19636 78855 19676
rect 78937 19636 78958 19676
rect 78958 19636 78998 19676
rect 78998 19636 79023 19676
rect 78769 19613 78855 19636
rect 78937 19613 79023 19636
rect 4409 18920 4495 18943
rect 4577 18920 4663 18943
rect 4409 18880 4434 18920
rect 4434 18880 4474 18920
rect 4474 18880 4495 18920
rect 4577 18880 4598 18920
rect 4598 18880 4638 18920
rect 4638 18880 4663 18920
rect 4409 18857 4495 18880
rect 4577 18857 4663 18880
rect 19529 18920 19615 18943
rect 19697 18920 19783 18943
rect 19529 18880 19554 18920
rect 19554 18880 19594 18920
rect 19594 18880 19615 18920
rect 19697 18880 19718 18920
rect 19718 18880 19758 18920
rect 19758 18880 19783 18920
rect 19529 18857 19615 18880
rect 19697 18857 19783 18880
rect 34649 18920 34735 18943
rect 34817 18920 34903 18943
rect 34649 18880 34674 18920
rect 34674 18880 34714 18920
rect 34714 18880 34735 18920
rect 34817 18880 34838 18920
rect 34838 18880 34878 18920
rect 34878 18880 34903 18920
rect 34649 18857 34735 18880
rect 34817 18857 34903 18880
rect 49769 18920 49855 18943
rect 49937 18920 50023 18943
rect 49769 18880 49794 18920
rect 49794 18880 49834 18920
rect 49834 18880 49855 18920
rect 49937 18880 49958 18920
rect 49958 18880 49998 18920
rect 49998 18880 50023 18920
rect 49769 18857 49855 18880
rect 49937 18857 50023 18880
rect 64889 18920 64975 18943
rect 65057 18920 65143 18943
rect 64889 18880 64914 18920
rect 64914 18880 64954 18920
rect 64954 18880 64975 18920
rect 65057 18880 65078 18920
rect 65078 18880 65118 18920
rect 65118 18880 65143 18920
rect 64889 18857 64975 18880
rect 65057 18857 65143 18880
rect 80009 18920 80095 18943
rect 80177 18920 80263 18943
rect 80009 18880 80034 18920
rect 80034 18880 80074 18920
rect 80074 18880 80095 18920
rect 80177 18880 80198 18920
rect 80198 18880 80238 18920
rect 80238 18880 80263 18920
rect 80009 18857 80095 18880
rect 80177 18857 80263 18880
rect 3169 18164 3255 18187
rect 3337 18164 3423 18187
rect 3169 18124 3194 18164
rect 3194 18124 3234 18164
rect 3234 18124 3255 18164
rect 3337 18124 3358 18164
rect 3358 18124 3398 18164
rect 3398 18124 3423 18164
rect 3169 18101 3255 18124
rect 3337 18101 3423 18124
rect 18289 18164 18375 18187
rect 18457 18164 18543 18187
rect 18289 18124 18314 18164
rect 18314 18124 18354 18164
rect 18354 18124 18375 18164
rect 18457 18124 18478 18164
rect 18478 18124 18518 18164
rect 18518 18124 18543 18164
rect 18289 18101 18375 18124
rect 18457 18101 18543 18124
rect 33409 18164 33495 18187
rect 33577 18164 33663 18187
rect 33409 18124 33434 18164
rect 33434 18124 33474 18164
rect 33474 18124 33495 18164
rect 33577 18124 33598 18164
rect 33598 18124 33638 18164
rect 33638 18124 33663 18164
rect 33409 18101 33495 18124
rect 33577 18101 33663 18124
rect 48529 18164 48615 18187
rect 48697 18164 48783 18187
rect 48529 18124 48554 18164
rect 48554 18124 48594 18164
rect 48594 18124 48615 18164
rect 48697 18124 48718 18164
rect 48718 18124 48758 18164
rect 48758 18124 48783 18164
rect 48529 18101 48615 18124
rect 48697 18101 48783 18124
rect 63649 18164 63735 18187
rect 63817 18164 63903 18187
rect 63649 18124 63674 18164
rect 63674 18124 63714 18164
rect 63714 18124 63735 18164
rect 63817 18124 63838 18164
rect 63838 18124 63878 18164
rect 63878 18124 63903 18164
rect 63649 18101 63735 18124
rect 63817 18101 63903 18124
rect 78769 18164 78855 18187
rect 78937 18164 79023 18187
rect 78769 18124 78794 18164
rect 78794 18124 78834 18164
rect 78834 18124 78855 18164
rect 78937 18124 78958 18164
rect 78958 18124 78998 18164
rect 78998 18124 79023 18164
rect 78769 18101 78855 18124
rect 78937 18101 79023 18124
rect 4409 17408 4495 17431
rect 4577 17408 4663 17431
rect 4409 17368 4434 17408
rect 4434 17368 4474 17408
rect 4474 17368 4495 17408
rect 4577 17368 4598 17408
rect 4598 17368 4638 17408
rect 4638 17368 4663 17408
rect 4409 17345 4495 17368
rect 4577 17345 4663 17368
rect 19529 17408 19615 17431
rect 19697 17408 19783 17431
rect 19529 17368 19554 17408
rect 19554 17368 19594 17408
rect 19594 17368 19615 17408
rect 19697 17368 19718 17408
rect 19718 17368 19758 17408
rect 19758 17368 19783 17408
rect 19529 17345 19615 17368
rect 19697 17345 19783 17368
rect 34649 17408 34735 17431
rect 34817 17408 34903 17431
rect 34649 17368 34674 17408
rect 34674 17368 34714 17408
rect 34714 17368 34735 17408
rect 34817 17368 34838 17408
rect 34838 17368 34878 17408
rect 34878 17368 34903 17408
rect 34649 17345 34735 17368
rect 34817 17345 34903 17368
rect 49769 17408 49855 17431
rect 49937 17408 50023 17431
rect 49769 17368 49794 17408
rect 49794 17368 49834 17408
rect 49834 17368 49855 17408
rect 49937 17368 49958 17408
rect 49958 17368 49998 17408
rect 49998 17368 50023 17408
rect 49769 17345 49855 17368
rect 49937 17345 50023 17368
rect 64889 17408 64975 17431
rect 65057 17408 65143 17431
rect 64889 17368 64914 17408
rect 64914 17368 64954 17408
rect 64954 17368 64975 17408
rect 65057 17368 65078 17408
rect 65078 17368 65118 17408
rect 65118 17368 65143 17408
rect 64889 17345 64975 17368
rect 65057 17345 65143 17368
rect 80009 17408 80095 17431
rect 80177 17408 80263 17431
rect 80009 17368 80034 17408
rect 80034 17368 80074 17408
rect 80074 17368 80095 17408
rect 80177 17368 80198 17408
rect 80198 17368 80238 17408
rect 80238 17368 80263 17408
rect 80009 17345 80095 17368
rect 80177 17345 80263 17368
rect 3169 16652 3255 16675
rect 3337 16652 3423 16675
rect 3169 16612 3194 16652
rect 3194 16612 3234 16652
rect 3234 16612 3255 16652
rect 3337 16612 3358 16652
rect 3358 16612 3398 16652
rect 3398 16612 3423 16652
rect 3169 16589 3255 16612
rect 3337 16589 3423 16612
rect 18289 16652 18375 16675
rect 18457 16652 18543 16675
rect 18289 16612 18314 16652
rect 18314 16612 18354 16652
rect 18354 16612 18375 16652
rect 18457 16612 18478 16652
rect 18478 16612 18518 16652
rect 18518 16612 18543 16652
rect 18289 16589 18375 16612
rect 18457 16589 18543 16612
rect 33409 16652 33495 16675
rect 33577 16652 33663 16675
rect 33409 16612 33434 16652
rect 33434 16612 33474 16652
rect 33474 16612 33495 16652
rect 33577 16612 33598 16652
rect 33598 16612 33638 16652
rect 33638 16612 33663 16652
rect 33409 16589 33495 16612
rect 33577 16589 33663 16612
rect 48529 16652 48615 16675
rect 48697 16652 48783 16675
rect 48529 16612 48554 16652
rect 48554 16612 48594 16652
rect 48594 16612 48615 16652
rect 48697 16612 48718 16652
rect 48718 16612 48758 16652
rect 48758 16612 48783 16652
rect 48529 16589 48615 16612
rect 48697 16589 48783 16612
rect 63649 16652 63735 16675
rect 63817 16652 63903 16675
rect 63649 16612 63674 16652
rect 63674 16612 63714 16652
rect 63714 16612 63735 16652
rect 63817 16612 63838 16652
rect 63838 16612 63878 16652
rect 63878 16612 63903 16652
rect 63649 16589 63735 16612
rect 63817 16589 63903 16612
rect 78769 16652 78855 16675
rect 78937 16652 79023 16675
rect 78769 16612 78794 16652
rect 78794 16612 78834 16652
rect 78834 16612 78855 16652
rect 78937 16612 78958 16652
rect 78958 16612 78998 16652
rect 78998 16612 79023 16652
rect 78769 16589 78855 16612
rect 78937 16589 79023 16612
rect 4409 15896 4495 15919
rect 4577 15896 4663 15919
rect 4409 15856 4434 15896
rect 4434 15856 4474 15896
rect 4474 15856 4495 15896
rect 4577 15856 4598 15896
rect 4598 15856 4638 15896
rect 4638 15856 4663 15896
rect 4409 15833 4495 15856
rect 4577 15833 4663 15856
rect 19529 15896 19615 15919
rect 19697 15896 19783 15919
rect 19529 15856 19554 15896
rect 19554 15856 19594 15896
rect 19594 15856 19615 15896
rect 19697 15856 19718 15896
rect 19718 15856 19758 15896
rect 19758 15856 19783 15896
rect 19529 15833 19615 15856
rect 19697 15833 19783 15856
rect 34649 15896 34735 15919
rect 34817 15896 34903 15919
rect 34649 15856 34674 15896
rect 34674 15856 34714 15896
rect 34714 15856 34735 15896
rect 34817 15856 34838 15896
rect 34838 15856 34878 15896
rect 34878 15856 34903 15896
rect 34649 15833 34735 15856
rect 34817 15833 34903 15856
rect 49769 15896 49855 15919
rect 49937 15896 50023 15919
rect 49769 15856 49794 15896
rect 49794 15856 49834 15896
rect 49834 15856 49855 15896
rect 49937 15856 49958 15896
rect 49958 15856 49998 15896
rect 49998 15856 50023 15896
rect 49769 15833 49855 15856
rect 49937 15833 50023 15856
rect 64889 15896 64975 15919
rect 65057 15896 65143 15919
rect 64889 15856 64914 15896
rect 64914 15856 64954 15896
rect 64954 15856 64975 15896
rect 65057 15856 65078 15896
rect 65078 15856 65118 15896
rect 65118 15856 65143 15896
rect 64889 15833 64975 15856
rect 65057 15833 65143 15856
rect 80009 15896 80095 15919
rect 80177 15896 80263 15919
rect 80009 15856 80034 15896
rect 80034 15856 80074 15896
rect 80074 15856 80095 15896
rect 80177 15856 80198 15896
rect 80198 15856 80238 15896
rect 80238 15856 80263 15896
rect 80009 15833 80095 15856
rect 80177 15833 80263 15856
rect 3169 15140 3255 15163
rect 3337 15140 3423 15163
rect 3169 15100 3194 15140
rect 3194 15100 3234 15140
rect 3234 15100 3255 15140
rect 3337 15100 3358 15140
rect 3358 15100 3398 15140
rect 3398 15100 3423 15140
rect 3169 15077 3255 15100
rect 3337 15077 3423 15100
rect 18289 15140 18375 15163
rect 18457 15140 18543 15163
rect 18289 15100 18314 15140
rect 18314 15100 18354 15140
rect 18354 15100 18375 15140
rect 18457 15100 18478 15140
rect 18478 15100 18518 15140
rect 18518 15100 18543 15140
rect 18289 15077 18375 15100
rect 18457 15077 18543 15100
rect 33409 15140 33495 15163
rect 33577 15140 33663 15163
rect 33409 15100 33434 15140
rect 33434 15100 33474 15140
rect 33474 15100 33495 15140
rect 33577 15100 33598 15140
rect 33598 15100 33638 15140
rect 33638 15100 33663 15140
rect 33409 15077 33495 15100
rect 33577 15077 33663 15100
rect 48529 15140 48615 15163
rect 48697 15140 48783 15163
rect 48529 15100 48554 15140
rect 48554 15100 48594 15140
rect 48594 15100 48615 15140
rect 48697 15100 48718 15140
rect 48718 15100 48758 15140
rect 48758 15100 48783 15140
rect 48529 15077 48615 15100
rect 48697 15077 48783 15100
rect 63649 15140 63735 15163
rect 63817 15140 63903 15163
rect 63649 15100 63674 15140
rect 63674 15100 63714 15140
rect 63714 15100 63735 15140
rect 63817 15100 63838 15140
rect 63838 15100 63878 15140
rect 63878 15100 63903 15140
rect 63649 15077 63735 15100
rect 63817 15077 63903 15100
rect 78769 15140 78855 15163
rect 78937 15140 79023 15163
rect 78769 15100 78794 15140
rect 78794 15100 78834 15140
rect 78834 15100 78855 15140
rect 78937 15100 78958 15140
rect 78958 15100 78998 15140
rect 78998 15100 79023 15140
rect 78769 15077 78855 15100
rect 78937 15077 79023 15100
rect 4409 14384 4495 14407
rect 4577 14384 4663 14407
rect 4409 14344 4434 14384
rect 4434 14344 4474 14384
rect 4474 14344 4495 14384
rect 4577 14344 4598 14384
rect 4598 14344 4638 14384
rect 4638 14344 4663 14384
rect 4409 14321 4495 14344
rect 4577 14321 4663 14344
rect 19529 14384 19615 14407
rect 19697 14384 19783 14407
rect 19529 14344 19554 14384
rect 19554 14344 19594 14384
rect 19594 14344 19615 14384
rect 19697 14344 19718 14384
rect 19718 14344 19758 14384
rect 19758 14344 19783 14384
rect 19529 14321 19615 14344
rect 19697 14321 19783 14344
rect 34649 14384 34735 14407
rect 34817 14384 34903 14407
rect 34649 14344 34674 14384
rect 34674 14344 34714 14384
rect 34714 14344 34735 14384
rect 34817 14344 34838 14384
rect 34838 14344 34878 14384
rect 34878 14344 34903 14384
rect 34649 14321 34735 14344
rect 34817 14321 34903 14344
rect 49769 14384 49855 14407
rect 49937 14384 50023 14407
rect 49769 14344 49794 14384
rect 49794 14344 49834 14384
rect 49834 14344 49855 14384
rect 49937 14344 49958 14384
rect 49958 14344 49998 14384
rect 49998 14344 50023 14384
rect 49769 14321 49855 14344
rect 49937 14321 50023 14344
rect 64889 14384 64975 14407
rect 65057 14384 65143 14407
rect 64889 14344 64914 14384
rect 64914 14344 64954 14384
rect 64954 14344 64975 14384
rect 65057 14344 65078 14384
rect 65078 14344 65118 14384
rect 65118 14344 65143 14384
rect 64889 14321 64975 14344
rect 65057 14321 65143 14344
rect 80009 14384 80095 14407
rect 80177 14384 80263 14407
rect 80009 14344 80034 14384
rect 80034 14344 80074 14384
rect 80074 14344 80095 14384
rect 80177 14344 80198 14384
rect 80198 14344 80238 14384
rect 80238 14344 80263 14384
rect 80009 14321 80095 14344
rect 80177 14321 80263 14344
rect 3169 13628 3255 13651
rect 3337 13628 3423 13651
rect 3169 13588 3194 13628
rect 3194 13588 3234 13628
rect 3234 13588 3255 13628
rect 3337 13588 3358 13628
rect 3358 13588 3398 13628
rect 3398 13588 3423 13628
rect 3169 13565 3255 13588
rect 3337 13565 3423 13588
rect 18289 13628 18375 13651
rect 18457 13628 18543 13651
rect 18289 13588 18314 13628
rect 18314 13588 18354 13628
rect 18354 13588 18375 13628
rect 18457 13588 18478 13628
rect 18478 13588 18518 13628
rect 18518 13588 18543 13628
rect 18289 13565 18375 13588
rect 18457 13565 18543 13588
rect 33409 13628 33495 13651
rect 33577 13628 33663 13651
rect 33409 13588 33434 13628
rect 33434 13588 33474 13628
rect 33474 13588 33495 13628
rect 33577 13588 33598 13628
rect 33598 13588 33638 13628
rect 33638 13588 33663 13628
rect 33409 13565 33495 13588
rect 33577 13565 33663 13588
rect 48529 13628 48615 13651
rect 48697 13628 48783 13651
rect 48529 13588 48554 13628
rect 48554 13588 48594 13628
rect 48594 13588 48615 13628
rect 48697 13588 48718 13628
rect 48718 13588 48758 13628
rect 48758 13588 48783 13628
rect 48529 13565 48615 13588
rect 48697 13565 48783 13588
rect 63649 13628 63735 13651
rect 63817 13628 63903 13651
rect 63649 13588 63674 13628
rect 63674 13588 63714 13628
rect 63714 13588 63735 13628
rect 63817 13588 63838 13628
rect 63838 13588 63878 13628
rect 63878 13588 63903 13628
rect 63649 13565 63735 13588
rect 63817 13565 63903 13588
rect 78769 13628 78855 13651
rect 78937 13628 79023 13651
rect 78769 13588 78794 13628
rect 78794 13588 78834 13628
rect 78834 13588 78855 13628
rect 78937 13588 78958 13628
rect 78958 13588 78998 13628
rect 78998 13588 79023 13628
rect 78769 13565 78855 13588
rect 78937 13565 79023 13588
rect 4409 12872 4495 12895
rect 4577 12872 4663 12895
rect 4409 12832 4434 12872
rect 4434 12832 4474 12872
rect 4474 12832 4495 12872
rect 4577 12832 4598 12872
rect 4598 12832 4638 12872
rect 4638 12832 4663 12872
rect 4409 12809 4495 12832
rect 4577 12809 4663 12832
rect 19529 12872 19615 12895
rect 19697 12872 19783 12895
rect 19529 12832 19554 12872
rect 19554 12832 19594 12872
rect 19594 12832 19615 12872
rect 19697 12832 19718 12872
rect 19718 12832 19758 12872
rect 19758 12832 19783 12872
rect 19529 12809 19615 12832
rect 19697 12809 19783 12832
rect 34649 12872 34735 12895
rect 34817 12872 34903 12895
rect 34649 12832 34674 12872
rect 34674 12832 34714 12872
rect 34714 12832 34735 12872
rect 34817 12832 34838 12872
rect 34838 12832 34878 12872
rect 34878 12832 34903 12872
rect 34649 12809 34735 12832
rect 34817 12809 34903 12832
rect 49769 12872 49855 12895
rect 49937 12872 50023 12895
rect 49769 12832 49794 12872
rect 49794 12832 49834 12872
rect 49834 12832 49855 12872
rect 49937 12832 49958 12872
rect 49958 12832 49998 12872
rect 49998 12832 50023 12872
rect 49769 12809 49855 12832
rect 49937 12809 50023 12832
rect 64889 12872 64975 12895
rect 65057 12872 65143 12895
rect 64889 12832 64914 12872
rect 64914 12832 64954 12872
rect 64954 12832 64975 12872
rect 65057 12832 65078 12872
rect 65078 12832 65118 12872
rect 65118 12832 65143 12872
rect 64889 12809 64975 12832
rect 65057 12809 65143 12832
rect 80009 12872 80095 12895
rect 80177 12872 80263 12895
rect 80009 12832 80034 12872
rect 80034 12832 80074 12872
rect 80074 12832 80095 12872
rect 80177 12832 80198 12872
rect 80198 12832 80238 12872
rect 80238 12832 80263 12872
rect 80009 12809 80095 12832
rect 80177 12809 80263 12832
rect 3169 12116 3255 12139
rect 3337 12116 3423 12139
rect 3169 12076 3194 12116
rect 3194 12076 3234 12116
rect 3234 12076 3255 12116
rect 3337 12076 3358 12116
rect 3358 12076 3398 12116
rect 3398 12076 3423 12116
rect 3169 12053 3255 12076
rect 3337 12053 3423 12076
rect 18289 12116 18375 12139
rect 18457 12116 18543 12139
rect 18289 12076 18314 12116
rect 18314 12076 18354 12116
rect 18354 12076 18375 12116
rect 18457 12076 18478 12116
rect 18478 12076 18518 12116
rect 18518 12076 18543 12116
rect 18289 12053 18375 12076
rect 18457 12053 18543 12076
rect 33409 12116 33495 12139
rect 33577 12116 33663 12139
rect 33409 12076 33434 12116
rect 33434 12076 33474 12116
rect 33474 12076 33495 12116
rect 33577 12076 33598 12116
rect 33598 12076 33638 12116
rect 33638 12076 33663 12116
rect 33409 12053 33495 12076
rect 33577 12053 33663 12076
rect 48529 12116 48615 12139
rect 48697 12116 48783 12139
rect 48529 12076 48554 12116
rect 48554 12076 48594 12116
rect 48594 12076 48615 12116
rect 48697 12076 48718 12116
rect 48718 12076 48758 12116
rect 48758 12076 48783 12116
rect 48529 12053 48615 12076
rect 48697 12053 48783 12076
rect 63649 12116 63735 12139
rect 63817 12116 63903 12139
rect 63649 12076 63674 12116
rect 63674 12076 63714 12116
rect 63714 12076 63735 12116
rect 63817 12076 63838 12116
rect 63838 12076 63878 12116
rect 63878 12076 63903 12116
rect 63649 12053 63735 12076
rect 63817 12053 63903 12076
rect 78769 12116 78855 12139
rect 78937 12116 79023 12139
rect 78769 12076 78794 12116
rect 78794 12076 78834 12116
rect 78834 12076 78855 12116
rect 78937 12076 78958 12116
rect 78958 12076 78998 12116
rect 78998 12076 79023 12116
rect 78769 12053 78855 12076
rect 78937 12053 79023 12076
rect 4409 11360 4495 11383
rect 4577 11360 4663 11383
rect 4409 11320 4434 11360
rect 4434 11320 4474 11360
rect 4474 11320 4495 11360
rect 4577 11320 4598 11360
rect 4598 11320 4638 11360
rect 4638 11320 4663 11360
rect 4409 11297 4495 11320
rect 4577 11297 4663 11320
rect 19529 11360 19615 11383
rect 19697 11360 19783 11383
rect 19529 11320 19554 11360
rect 19554 11320 19594 11360
rect 19594 11320 19615 11360
rect 19697 11320 19718 11360
rect 19718 11320 19758 11360
rect 19758 11320 19783 11360
rect 19529 11297 19615 11320
rect 19697 11297 19783 11320
rect 34649 11360 34735 11383
rect 34817 11360 34903 11383
rect 34649 11320 34674 11360
rect 34674 11320 34714 11360
rect 34714 11320 34735 11360
rect 34817 11320 34838 11360
rect 34838 11320 34878 11360
rect 34878 11320 34903 11360
rect 34649 11297 34735 11320
rect 34817 11297 34903 11320
rect 49769 11360 49855 11383
rect 49937 11360 50023 11383
rect 49769 11320 49794 11360
rect 49794 11320 49834 11360
rect 49834 11320 49855 11360
rect 49937 11320 49958 11360
rect 49958 11320 49998 11360
rect 49998 11320 50023 11360
rect 49769 11297 49855 11320
rect 49937 11297 50023 11320
rect 64889 11360 64975 11383
rect 65057 11360 65143 11383
rect 64889 11320 64914 11360
rect 64914 11320 64954 11360
rect 64954 11320 64975 11360
rect 65057 11320 65078 11360
rect 65078 11320 65118 11360
rect 65118 11320 65143 11360
rect 64889 11297 64975 11320
rect 65057 11297 65143 11320
rect 80009 11360 80095 11383
rect 80177 11360 80263 11383
rect 80009 11320 80034 11360
rect 80034 11320 80074 11360
rect 80074 11320 80095 11360
rect 80177 11320 80198 11360
rect 80198 11320 80238 11360
rect 80238 11320 80263 11360
rect 80009 11297 80095 11320
rect 80177 11297 80263 11320
rect 3169 10604 3255 10627
rect 3337 10604 3423 10627
rect 3169 10564 3194 10604
rect 3194 10564 3234 10604
rect 3234 10564 3255 10604
rect 3337 10564 3358 10604
rect 3358 10564 3398 10604
rect 3398 10564 3423 10604
rect 3169 10541 3255 10564
rect 3337 10541 3423 10564
rect 18289 10604 18375 10627
rect 18457 10604 18543 10627
rect 18289 10564 18314 10604
rect 18314 10564 18354 10604
rect 18354 10564 18375 10604
rect 18457 10564 18478 10604
rect 18478 10564 18518 10604
rect 18518 10564 18543 10604
rect 18289 10541 18375 10564
rect 18457 10541 18543 10564
rect 33409 10604 33495 10627
rect 33577 10604 33663 10627
rect 33409 10564 33434 10604
rect 33434 10564 33474 10604
rect 33474 10564 33495 10604
rect 33577 10564 33598 10604
rect 33598 10564 33638 10604
rect 33638 10564 33663 10604
rect 33409 10541 33495 10564
rect 33577 10541 33663 10564
rect 48529 10604 48615 10627
rect 48697 10604 48783 10627
rect 48529 10564 48554 10604
rect 48554 10564 48594 10604
rect 48594 10564 48615 10604
rect 48697 10564 48718 10604
rect 48718 10564 48758 10604
rect 48758 10564 48783 10604
rect 48529 10541 48615 10564
rect 48697 10541 48783 10564
rect 63649 10604 63735 10627
rect 63817 10604 63903 10627
rect 63649 10564 63674 10604
rect 63674 10564 63714 10604
rect 63714 10564 63735 10604
rect 63817 10564 63838 10604
rect 63838 10564 63878 10604
rect 63878 10564 63903 10604
rect 63649 10541 63735 10564
rect 63817 10541 63903 10564
rect 78769 10604 78855 10627
rect 78937 10604 79023 10627
rect 78769 10564 78794 10604
rect 78794 10564 78834 10604
rect 78834 10564 78855 10604
rect 78937 10564 78958 10604
rect 78958 10564 78998 10604
rect 78998 10564 79023 10604
rect 78769 10541 78855 10564
rect 78937 10541 79023 10564
rect 4409 9848 4495 9871
rect 4577 9848 4663 9871
rect 4409 9808 4434 9848
rect 4434 9808 4474 9848
rect 4474 9808 4495 9848
rect 4577 9808 4598 9848
rect 4598 9808 4638 9848
rect 4638 9808 4663 9848
rect 4409 9785 4495 9808
rect 4577 9785 4663 9808
rect 19529 9848 19615 9871
rect 19697 9848 19783 9871
rect 19529 9808 19554 9848
rect 19554 9808 19594 9848
rect 19594 9808 19615 9848
rect 19697 9808 19718 9848
rect 19718 9808 19758 9848
rect 19758 9808 19783 9848
rect 19529 9785 19615 9808
rect 19697 9785 19783 9808
rect 34649 9848 34735 9871
rect 34817 9848 34903 9871
rect 34649 9808 34674 9848
rect 34674 9808 34714 9848
rect 34714 9808 34735 9848
rect 34817 9808 34838 9848
rect 34838 9808 34878 9848
rect 34878 9808 34903 9848
rect 34649 9785 34735 9808
rect 34817 9785 34903 9808
rect 49769 9848 49855 9871
rect 49937 9848 50023 9871
rect 49769 9808 49794 9848
rect 49794 9808 49834 9848
rect 49834 9808 49855 9848
rect 49937 9808 49958 9848
rect 49958 9808 49998 9848
rect 49998 9808 50023 9848
rect 49769 9785 49855 9808
rect 49937 9785 50023 9808
rect 64889 9848 64975 9871
rect 65057 9848 65143 9871
rect 64889 9808 64914 9848
rect 64914 9808 64954 9848
rect 64954 9808 64975 9848
rect 65057 9808 65078 9848
rect 65078 9808 65118 9848
rect 65118 9808 65143 9848
rect 64889 9785 64975 9808
rect 65057 9785 65143 9808
rect 80009 9848 80095 9871
rect 80177 9848 80263 9871
rect 80009 9808 80034 9848
rect 80034 9808 80074 9848
rect 80074 9808 80095 9848
rect 80177 9808 80198 9848
rect 80198 9808 80238 9848
rect 80238 9808 80263 9848
rect 80009 9785 80095 9808
rect 80177 9785 80263 9808
rect 3169 9092 3255 9115
rect 3337 9092 3423 9115
rect 3169 9052 3194 9092
rect 3194 9052 3234 9092
rect 3234 9052 3255 9092
rect 3337 9052 3358 9092
rect 3358 9052 3398 9092
rect 3398 9052 3423 9092
rect 3169 9029 3255 9052
rect 3337 9029 3423 9052
rect 18289 9092 18375 9115
rect 18457 9092 18543 9115
rect 18289 9052 18314 9092
rect 18314 9052 18354 9092
rect 18354 9052 18375 9092
rect 18457 9052 18478 9092
rect 18478 9052 18518 9092
rect 18518 9052 18543 9092
rect 18289 9029 18375 9052
rect 18457 9029 18543 9052
rect 33409 9092 33495 9115
rect 33577 9092 33663 9115
rect 33409 9052 33434 9092
rect 33434 9052 33474 9092
rect 33474 9052 33495 9092
rect 33577 9052 33598 9092
rect 33598 9052 33638 9092
rect 33638 9052 33663 9092
rect 33409 9029 33495 9052
rect 33577 9029 33663 9052
rect 48529 9092 48615 9115
rect 48697 9092 48783 9115
rect 48529 9052 48554 9092
rect 48554 9052 48594 9092
rect 48594 9052 48615 9092
rect 48697 9052 48718 9092
rect 48718 9052 48758 9092
rect 48758 9052 48783 9092
rect 48529 9029 48615 9052
rect 48697 9029 48783 9052
rect 63649 9092 63735 9115
rect 63817 9092 63903 9115
rect 63649 9052 63674 9092
rect 63674 9052 63714 9092
rect 63714 9052 63735 9092
rect 63817 9052 63838 9092
rect 63838 9052 63878 9092
rect 63878 9052 63903 9092
rect 63649 9029 63735 9052
rect 63817 9029 63903 9052
rect 78769 9092 78855 9115
rect 78937 9092 79023 9115
rect 78769 9052 78794 9092
rect 78794 9052 78834 9092
rect 78834 9052 78855 9092
rect 78937 9052 78958 9092
rect 78958 9052 78998 9092
rect 78998 9052 79023 9092
rect 78769 9029 78855 9052
rect 78937 9029 79023 9052
rect 4409 8336 4495 8359
rect 4577 8336 4663 8359
rect 4409 8296 4434 8336
rect 4434 8296 4474 8336
rect 4474 8296 4495 8336
rect 4577 8296 4598 8336
rect 4598 8296 4638 8336
rect 4638 8296 4663 8336
rect 4409 8273 4495 8296
rect 4577 8273 4663 8296
rect 19529 8336 19615 8359
rect 19697 8336 19783 8359
rect 19529 8296 19554 8336
rect 19554 8296 19594 8336
rect 19594 8296 19615 8336
rect 19697 8296 19718 8336
rect 19718 8296 19758 8336
rect 19758 8296 19783 8336
rect 19529 8273 19615 8296
rect 19697 8273 19783 8296
rect 34649 8336 34735 8359
rect 34817 8336 34903 8359
rect 34649 8296 34674 8336
rect 34674 8296 34714 8336
rect 34714 8296 34735 8336
rect 34817 8296 34838 8336
rect 34838 8296 34878 8336
rect 34878 8296 34903 8336
rect 34649 8273 34735 8296
rect 34817 8273 34903 8296
rect 49769 8336 49855 8359
rect 49937 8336 50023 8359
rect 49769 8296 49794 8336
rect 49794 8296 49834 8336
rect 49834 8296 49855 8336
rect 49937 8296 49958 8336
rect 49958 8296 49998 8336
rect 49998 8296 50023 8336
rect 49769 8273 49855 8296
rect 49937 8273 50023 8296
rect 64889 8336 64975 8359
rect 65057 8336 65143 8359
rect 64889 8296 64914 8336
rect 64914 8296 64954 8336
rect 64954 8296 64975 8336
rect 65057 8296 65078 8336
rect 65078 8296 65118 8336
rect 65118 8296 65143 8336
rect 64889 8273 64975 8296
rect 65057 8273 65143 8296
rect 80009 8336 80095 8359
rect 80177 8336 80263 8359
rect 80009 8296 80034 8336
rect 80034 8296 80074 8336
rect 80074 8296 80095 8336
rect 80177 8296 80198 8336
rect 80198 8296 80238 8336
rect 80238 8296 80263 8336
rect 80009 8273 80095 8296
rect 80177 8273 80263 8296
rect 3169 7580 3255 7603
rect 3337 7580 3423 7603
rect 3169 7540 3194 7580
rect 3194 7540 3234 7580
rect 3234 7540 3255 7580
rect 3337 7540 3358 7580
rect 3358 7540 3398 7580
rect 3398 7540 3423 7580
rect 3169 7517 3255 7540
rect 3337 7517 3423 7540
rect 18289 7580 18375 7603
rect 18457 7580 18543 7603
rect 18289 7540 18314 7580
rect 18314 7540 18354 7580
rect 18354 7540 18375 7580
rect 18457 7540 18478 7580
rect 18478 7540 18518 7580
rect 18518 7540 18543 7580
rect 18289 7517 18375 7540
rect 18457 7517 18543 7540
rect 33409 7580 33495 7603
rect 33577 7580 33663 7603
rect 33409 7540 33434 7580
rect 33434 7540 33474 7580
rect 33474 7540 33495 7580
rect 33577 7540 33598 7580
rect 33598 7540 33638 7580
rect 33638 7540 33663 7580
rect 33409 7517 33495 7540
rect 33577 7517 33663 7540
rect 48529 7580 48615 7603
rect 48697 7580 48783 7603
rect 48529 7540 48554 7580
rect 48554 7540 48594 7580
rect 48594 7540 48615 7580
rect 48697 7540 48718 7580
rect 48718 7540 48758 7580
rect 48758 7540 48783 7580
rect 48529 7517 48615 7540
rect 48697 7517 48783 7540
rect 63649 7580 63735 7603
rect 63817 7580 63903 7603
rect 63649 7540 63674 7580
rect 63674 7540 63714 7580
rect 63714 7540 63735 7580
rect 63817 7540 63838 7580
rect 63838 7540 63878 7580
rect 63878 7540 63903 7580
rect 63649 7517 63735 7540
rect 63817 7517 63903 7540
rect 78769 7580 78855 7603
rect 78937 7580 79023 7603
rect 78769 7540 78794 7580
rect 78794 7540 78834 7580
rect 78834 7540 78855 7580
rect 78937 7540 78958 7580
rect 78958 7540 78998 7580
rect 78998 7540 79023 7580
rect 78769 7517 78855 7540
rect 78937 7517 79023 7540
rect 4409 6824 4495 6847
rect 4577 6824 4663 6847
rect 4409 6784 4434 6824
rect 4434 6784 4474 6824
rect 4474 6784 4495 6824
rect 4577 6784 4598 6824
rect 4598 6784 4638 6824
rect 4638 6784 4663 6824
rect 4409 6761 4495 6784
rect 4577 6761 4663 6784
rect 19529 6824 19615 6847
rect 19697 6824 19783 6847
rect 19529 6784 19554 6824
rect 19554 6784 19594 6824
rect 19594 6784 19615 6824
rect 19697 6784 19718 6824
rect 19718 6784 19758 6824
rect 19758 6784 19783 6824
rect 19529 6761 19615 6784
rect 19697 6761 19783 6784
rect 34649 6824 34735 6847
rect 34817 6824 34903 6847
rect 34649 6784 34674 6824
rect 34674 6784 34714 6824
rect 34714 6784 34735 6824
rect 34817 6784 34838 6824
rect 34838 6784 34878 6824
rect 34878 6784 34903 6824
rect 34649 6761 34735 6784
rect 34817 6761 34903 6784
rect 49769 6824 49855 6847
rect 49937 6824 50023 6847
rect 49769 6784 49794 6824
rect 49794 6784 49834 6824
rect 49834 6784 49855 6824
rect 49937 6784 49958 6824
rect 49958 6784 49998 6824
rect 49998 6784 50023 6824
rect 49769 6761 49855 6784
rect 49937 6761 50023 6784
rect 64889 6824 64975 6847
rect 65057 6824 65143 6847
rect 64889 6784 64914 6824
rect 64914 6784 64954 6824
rect 64954 6784 64975 6824
rect 65057 6784 65078 6824
rect 65078 6784 65118 6824
rect 65118 6784 65143 6824
rect 64889 6761 64975 6784
rect 65057 6761 65143 6784
rect 80009 6824 80095 6847
rect 80177 6824 80263 6847
rect 80009 6784 80034 6824
rect 80034 6784 80074 6824
rect 80074 6784 80095 6824
rect 80177 6784 80198 6824
rect 80198 6784 80238 6824
rect 80238 6784 80263 6824
rect 80009 6761 80095 6784
rect 80177 6761 80263 6784
rect 3169 6068 3255 6091
rect 3337 6068 3423 6091
rect 3169 6028 3194 6068
rect 3194 6028 3234 6068
rect 3234 6028 3255 6068
rect 3337 6028 3358 6068
rect 3358 6028 3398 6068
rect 3398 6028 3423 6068
rect 3169 6005 3255 6028
rect 3337 6005 3423 6028
rect 18289 6068 18375 6091
rect 18457 6068 18543 6091
rect 18289 6028 18314 6068
rect 18314 6028 18354 6068
rect 18354 6028 18375 6068
rect 18457 6028 18478 6068
rect 18478 6028 18518 6068
rect 18518 6028 18543 6068
rect 18289 6005 18375 6028
rect 18457 6005 18543 6028
rect 33409 6068 33495 6091
rect 33577 6068 33663 6091
rect 33409 6028 33434 6068
rect 33434 6028 33474 6068
rect 33474 6028 33495 6068
rect 33577 6028 33598 6068
rect 33598 6028 33638 6068
rect 33638 6028 33663 6068
rect 33409 6005 33495 6028
rect 33577 6005 33663 6028
rect 48529 6068 48615 6091
rect 48697 6068 48783 6091
rect 48529 6028 48554 6068
rect 48554 6028 48594 6068
rect 48594 6028 48615 6068
rect 48697 6028 48718 6068
rect 48718 6028 48758 6068
rect 48758 6028 48783 6068
rect 48529 6005 48615 6028
rect 48697 6005 48783 6028
rect 63649 6068 63735 6091
rect 63817 6068 63903 6091
rect 63649 6028 63674 6068
rect 63674 6028 63714 6068
rect 63714 6028 63735 6068
rect 63817 6028 63838 6068
rect 63838 6028 63878 6068
rect 63878 6028 63903 6068
rect 63649 6005 63735 6028
rect 63817 6005 63903 6028
rect 78769 6068 78855 6091
rect 78937 6068 79023 6091
rect 78769 6028 78794 6068
rect 78794 6028 78834 6068
rect 78834 6028 78855 6068
rect 78937 6028 78958 6068
rect 78958 6028 78998 6068
rect 78998 6028 79023 6068
rect 78769 6005 78855 6028
rect 78937 6005 79023 6028
rect 4409 5312 4495 5335
rect 4577 5312 4663 5335
rect 4409 5272 4434 5312
rect 4434 5272 4474 5312
rect 4474 5272 4495 5312
rect 4577 5272 4598 5312
rect 4598 5272 4638 5312
rect 4638 5272 4663 5312
rect 4409 5249 4495 5272
rect 4577 5249 4663 5272
rect 19529 5312 19615 5335
rect 19697 5312 19783 5335
rect 19529 5272 19554 5312
rect 19554 5272 19594 5312
rect 19594 5272 19615 5312
rect 19697 5272 19718 5312
rect 19718 5272 19758 5312
rect 19758 5272 19783 5312
rect 19529 5249 19615 5272
rect 19697 5249 19783 5272
rect 34649 5312 34735 5335
rect 34817 5312 34903 5335
rect 34649 5272 34674 5312
rect 34674 5272 34714 5312
rect 34714 5272 34735 5312
rect 34817 5272 34838 5312
rect 34838 5272 34878 5312
rect 34878 5272 34903 5312
rect 34649 5249 34735 5272
rect 34817 5249 34903 5272
rect 49769 5312 49855 5335
rect 49937 5312 50023 5335
rect 49769 5272 49794 5312
rect 49794 5272 49834 5312
rect 49834 5272 49855 5312
rect 49937 5272 49958 5312
rect 49958 5272 49998 5312
rect 49998 5272 50023 5312
rect 49769 5249 49855 5272
rect 49937 5249 50023 5272
rect 64889 5312 64975 5335
rect 65057 5312 65143 5335
rect 64889 5272 64914 5312
rect 64914 5272 64954 5312
rect 64954 5272 64975 5312
rect 65057 5272 65078 5312
rect 65078 5272 65118 5312
rect 65118 5272 65143 5312
rect 64889 5249 64975 5272
rect 65057 5249 65143 5272
rect 80009 5312 80095 5335
rect 80177 5312 80263 5335
rect 80009 5272 80034 5312
rect 80034 5272 80074 5312
rect 80074 5272 80095 5312
rect 80177 5272 80198 5312
rect 80198 5272 80238 5312
rect 80238 5272 80263 5312
rect 80009 5249 80095 5272
rect 80177 5249 80263 5272
rect 3169 4556 3255 4579
rect 3337 4556 3423 4579
rect 3169 4516 3194 4556
rect 3194 4516 3234 4556
rect 3234 4516 3255 4556
rect 3337 4516 3358 4556
rect 3358 4516 3398 4556
rect 3398 4516 3423 4556
rect 3169 4493 3255 4516
rect 3337 4493 3423 4516
rect 18289 4556 18375 4579
rect 18457 4556 18543 4579
rect 18289 4516 18314 4556
rect 18314 4516 18354 4556
rect 18354 4516 18375 4556
rect 18457 4516 18478 4556
rect 18478 4516 18518 4556
rect 18518 4516 18543 4556
rect 18289 4493 18375 4516
rect 18457 4493 18543 4516
rect 33409 4556 33495 4579
rect 33577 4556 33663 4579
rect 33409 4516 33434 4556
rect 33434 4516 33474 4556
rect 33474 4516 33495 4556
rect 33577 4516 33598 4556
rect 33598 4516 33638 4556
rect 33638 4516 33663 4556
rect 33409 4493 33495 4516
rect 33577 4493 33663 4516
rect 48529 4556 48615 4579
rect 48697 4556 48783 4579
rect 48529 4516 48554 4556
rect 48554 4516 48594 4556
rect 48594 4516 48615 4556
rect 48697 4516 48718 4556
rect 48718 4516 48758 4556
rect 48758 4516 48783 4556
rect 48529 4493 48615 4516
rect 48697 4493 48783 4516
rect 63649 4556 63735 4579
rect 63817 4556 63903 4579
rect 63649 4516 63674 4556
rect 63674 4516 63714 4556
rect 63714 4516 63735 4556
rect 63817 4516 63838 4556
rect 63838 4516 63878 4556
rect 63878 4516 63903 4556
rect 63649 4493 63735 4516
rect 63817 4493 63903 4516
rect 78769 4556 78855 4579
rect 78937 4556 79023 4579
rect 78769 4516 78794 4556
rect 78794 4516 78834 4556
rect 78834 4516 78855 4556
rect 78937 4516 78958 4556
rect 78958 4516 78998 4556
rect 78998 4516 79023 4556
rect 78769 4493 78855 4516
rect 78937 4493 79023 4516
rect 4409 3800 4495 3823
rect 4577 3800 4663 3823
rect 4409 3760 4434 3800
rect 4434 3760 4474 3800
rect 4474 3760 4495 3800
rect 4577 3760 4598 3800
rect 4598 3760 4638 3800
rect 4638 3760 4663 3800
rect 4409 3737 4495 3760
rect 4577 3737 4663 3760
rect 19529 3800 19615 3823
rect 19697 3800 19783 3823
rect 19529 3760 19554 3800
rect 19554 3760 19594 3800
rect 19594 3760 19615 3800
rect 19697 3760 19718 3800
rect 19718 3760 19758 3800
rect 19758 3760 19783 3800
rect 19529 3737 19615 3760
rect 19697 3737 19783 3760
rect 34649 3800 34735 3823
rect 34817 3800 34903 3823
rect 34649 3760 34674 3800
rect 34674 3760 34714 3800
rect 34714 3760 34735 3800
rect 34817 3760 34838 3800
rect 34838 3760 34878 3800
rect 34878 3760 34903 3800
rect 34649 3737 34735 3760
rect 34817 3737 34903 3760
rect 49769 3800 49855 3823
rect 49937 3800 50023 3823
rect 49769 3760 49794 3800
rect 49794 3760 49834 3800
rect 49834 3760 49855 3800
rect 49937 3760 49958 3800
rect 49958 3760 49998 3800
rect 49998 3760 50023 3800
rect 49769 3737 49855 3760
rect 49937 3737 50023 3760
rect 64889 3800 64975 3823
rect 65057 3800 65143 3823
rect 64889 3760 64914 3800
rect 64914 3760 64954 3800
rect 64954 3760 64975 3800
rect 65057 3760 65078 3800
rect 65078 3760 65118 3800
rect 65118 3760 65143 3800
rect 64889 3737 64975 3760
rect 65057 3737 65143 3760
rect 80009 3800 80095 3823
rect 80177 3800 80263 3823
rect 80009 3760 80034 3800
rect 80034 3760 80074 3800
rect 80074 3760 80095 3800
rect 80177 3760 80198 3800
rect 80198 3760 80238 3800
rect 80238 3760 80263 3800
rect 80009 3737 80095 3760
rect 80177 3737 80263 3760
rect 3169 3044 3255 3067
rect 3337 3044 3423 3067
rect 3169 3004 3194 3044
rect 3194 3004 3234 3044
rect 3234 3004 3255 3044
rect 3337 3004 3358 3044
rect 3358 3004 3398 3044
rect 3398 3004 3423 3044
rect 3169 2981 3255 3004
rect 3337 2981 3423 3004
rect 18289 3044 18375 3067
rect 18457 3044 18543 3067
rect 18289 3004 18314 3044
rect 18314 3004 18354 3044
rect 18354 3004 18375 3044
rect 18457 3004 18478 3044
rect 18478 3004 18518 3044
rect 18518 3004 18543 3044
rect 18289 2981 18375 3004
rect 18457 2981 18543 3004
rect 33409 3044 33495 3067
rect 33577 3044 33663 3067
rect 33409 3004 33434 3044
rect 33434 3004 33474 3044
rect 33474 3004 33495 3044
rect 33577 3004 33598 3044
rect 33598 3004 33638 3044
rect 33638 3004 33663 3044
rect 33409 2981 33495 3004
rect 33577 2981 33663 3004
rect 48529 3044 48615 3067
rect 48697 3044 48783 3067
rect 48529 3004 48554 3044
rect 48554 3004 48594 3044
rect 48594 3004 48615 3044
rect 48697 3004 48718 3044
rect 48718 3004 48758 3044
rect 48758 3004 48783 3044
rect 48529 2981 48615 3004
rect 48697 2981 48783 3004
rect 63649 3044 63735 3067
rect 63817 3044 63903 3067
rect 63649 3004 63674 3044
rect 63674 3004 63714 3044
rect 63714 3004 63735 3044
rect 63817 3004 63838 3044
rect 63838 3004 63878 3044
rect 63878 3004 63903 3044
rect 63649 2981 63735 3004
rect 63817 2981 63903 3004
rect 78769 3044 78855 3067
rect 78937 3044 79023 3067
rect 78769 3004 78794 3044
rect 78794 3004 78834 3044
rect 78834 3004 78855 3044
rect 78937 3004 78958 3044
rect 78958 3004 78998 3044
rect 78998 3004 79023 3044
rect 78769 2981 78855 3004
rect 78937 2981 79023 3004
rect 4409 2288 4495 2311
rect 4577 2288 4663 2311
rect 4409 2248 4434 2288
rect 4434 2248 4474 2288
rect 4474 2248 4495 2288
rect 4577 2248 4598 2288
rect 4598 2248 4638 2288
rect 4638 2248 4663 2288
rect 4409 2225 4495 2248
rect 4577 2225 4663 2248
rect 19529 2288 19615 2311
rect 19697 2288 19783 2311
rect 19529 2248 19554 2288
rect 19554 2248 19594 2288
rect 19594 2248 19615 2288
rect 19697 2248 19718 2288
rect 19718 2248 19758 2288
rect 19758 2248 19783 2288
rect 19529 2225 19615 2248
rect 19697 2225 19783 2248
rect 34649 2288 34735 2311
rect 34817 2288 34903 2311
rect 34649 2248 34674 2288
rect 34674 2248 34714 2288
rect 34714 2248 34735 2288
rect 34817 2248 34838 2288
rect 34838 2248 34878 2288
rect 34878 2248 34903 2288
rect 34649 2225 34735 2248
rect 34817 2225 34903 2248
rect 49769 2288 49855 2311
rect 49937 2288 50023 2311
rect 49769 2248 49794 2288
rect 49794 2248 49834 2288
rect 49834 2248 49855 2288
rect 49937 2248 49958 2288
rect 49958 2248 49998 2288
rect 49998 2248 50023 2288
rect 49769 2225 49855 2248
rect 49937 2225 50023 2248
rect 64889 2288 64975 2311
rect 65057 2288 65143 2311
rect 64889 2248 64914 2288
rect 64914 2248 64954 2288
rect 64954 2248 64975 2288
rect 65057 2248 65078 2288
rect 65078 2248 65118 2288
rect 65118 2248 65143 2288
rect 64889 2225 64975 2248
rect 65057 2225 65143 2248
rect 80009 2288 80095 2311
rect 80177 2288 80263 2311
rect 80009 2248 80034 2288
rect 80034 2248 80074 2288
rect 80074 2248 80095 2288
rect 80177 2248 80198 2288
rect 80198 2248 80238 2288
rect 80238 2248 80263 2288
rect 80009 2225 80095 2248
rect 80177 2225 80263 2248
rect 3169 1532 3255 1555
rect 3337 1532 3423 1555
rect 3169 1492 3194 1532
rect 3194 1492 3234 1532
rect 3234 1492 3255 1532
rect 3337 1492 3358 1532
rect 3358 1492 3398 1532
rect 3398 1492 3423 1532
rect 3169 1469 3255 1492
rect 3337 1469 3423 1492
rect 18289 1532 18375 1555
rect 18457 1532 18543 1555
rect 18289 1492 18314 1532
rect 18314 1492 18354 1532
rect 18354 1492 18375 1532
rect 18457 1492 18478 1532
rect 18478 1492 18518 1532
rect 18518 1492 18543 1532
rect 18289 1469 18375 1492
rect 18457 1469 18543 1492
rect 33409 1532 33495 1555
rect 33577 1532 33663 1555
rect 33409 1492 33434 1532
rect 33434 1492 33474 1532
rect 33474 1492 33495 1532
rect 33577 1492 33598 1532
rect 33598 1492 33638 1532
rect 33638 1492 33663 1532
rect 33409 1469 33495 1492
rect 33577 1469 33663 1492
rect 48529 1532 48615 1555
rect 48697 1532 48783 1555
rect 48529 1492 48554 1532
rect 48554 1492 48594 1532
rect 48594 1492 48615 1532
rect 48697 1492 48718 1532
rect 48718 1492 48758 1532
rect 48758 1492 48783 1532
rect 48529 1469 48615 1492
rect 48697 1469 48783 1492
rect 63649 1532 63735 1555
rect 63817 1532 63903 1555
rect 63649 1492 63674 1532
rect 63674 1492 63714 1532
rect 63714 1492 63735 1532
rect 63817 1492 63838 1532
rect 63838 1492 63878 1532
rect 63878 1492 63903 1532
rect 63649 1469 63735 1492
rect 63817 1469 63903 1492
rect 78769 1532 78855 1555
rect 78937 1532 79023 1555
rect 78769 1492 78794 1532
rect 78794 1492 78834 1532
rect 78834 1492 78855 1532
rect 78937 1492 78958 1532
rect 78958 1492 78998 1532
rect 78998 1492 79023 1532
rect 78769 1469 78855 1492
rect 78937 1469 79023 1492
rect 4409 776 4495 799
rect 4577 776 4663 799
rect 4409 736 4434 776
rect 4434 736 4474 776
rect 4474 736 4495 776
rect 4577 736 4598 776
rect 4598 736 4638 776
rect 4638 736 4663 776
rect 4409 713 4495 736
rect 4577 713 4663 736
rect 19529 776 19615 799
rect 19697 776 19783 799
rect 19529 736 19554 776
rect 19554 736 19594 776
rect 19594 736 19615 776
rect 19697 736 19718 776
rect 19718 736 19758 776
rect 19758 736 19783 776
rect 19529 713 19615 736
rect 19697 713 19783 736
rect 34649 776 34735 799
rect 34817 776 34903 799
rect 34649 736 34674 776
rect 34674 736 34714 776
rect 34714 736 34735 776
rect 34817 736 34838 776
rect 34838 736 34878 776
rect 34878 736 34903 776
rect 34649 713 34735 736
rect 34817 713 34903 736
rect 49769 776 49855 799
rect 49937 776 50023 799
rect 49769 736 49794 776
rect 49794 736 49834 776
rect 49834 736 49855 776
rect 49937 736 49958 776
rect 49958 736 49998 776
rect 49998 736 50023 776
rect 49769 713 49855 736
rect 49937 713 50023 736
rect 64889 776 64975 799
rect 65057 776 65143 799
rect 64889 736 64914 776
rect 64914 736 64954 776
rect 64954 736 64975 776
rect 65057 736 65078 776
rect 65078 736 65118 776
rect 65118 736 65143 776
rect 64889 713 64975 736
rect 65057 713 65143 736
rect 80009 776 80095 799
rect 80177 776 80263 799
rect 80009 736 80034 776
rect 80034 736 80074 776
rect 80074 736 80095 776
rect 80177 736 80198 776
rect 80198 736 80238 776
rect 80238 736 80263 776
rect 80009 713 80095 736
rect 80177 713 80263 736
<< metal6 >>
rect 3076 37843 3516 38600
rect 3076 37757 3169 37843
rect 3255 37757 3337 37843
rect 3423 37757 3516 37843
rect 3076 36331 3516 37757
rect 3076 36245 3169 36331
rect 3255 36245 3337 36331
rect 3423 36245 3516 36331
rect 3076 34819 3516 36245
rect 3076 34733 3169 34819
rect 3255 34733 3337 34819
rect 3423 34733 3516 34819
rect 3076 33307 3516 34733
rect 3076 33221 3169 33307
rect 3255 33221 3337 33307
rect 3423 33221 3516 33307
rect 3076 31795 3516 33221
rect 3076 31709 3169 31795
rect 3255 31709 3337 31795
rect 3423 31709 3516 31795
rect 3076 30283 3516 31709
rect 3076 30197 3169 30283
rect 3255 30197 3337 30283
rect 3423 30197 3516 30283
rect 3076 28771 3516 30197
rect 3076 28685 3169 28771
rect 3255 28685 3337 28771
rect 3423 28685 3516 28771
rect 3076 27259 3516 28685
rect 3076 27173 3169 27259
rect 3255 27173 3337 27259
rect 3423 27173 3516 27259
rect 3076 25747 3516 27173
rect 3076 25661 3169 25747
rect 3255 25661 3337 25747
rect 3423 25661 3516 25747
rect 3076 24235 3516 25661
rect 3076 24149 3169 24235
rect 3255 24149 3337 24235
rect 3423 24149 3516 24235
rect 3076 22723 3516 24149
rect 3076 22637 3169 22723
rect 3255 22637 3337 22723
rect 3423 22637 3516 22723
rect 3076 21211 3516 22637
rect 3076 21125 3169 21211
rect 3255 21125 3337 21211
rect 3423 21125 3516 21211
rect 3076 19699 3516 21125
rect 3076 19613 3169 19699
rect 3255 19613 3337 19699
rect 3423 19613 3516 19699
rect 3076 18187 3516 19613
rect 3076 18101 3169 18187
rect 3255 18101 3337 18187
rect 3423 18101 3516 18187
rect 3076 16675 3516 18101
rect 3076 16589 3169 16675
rect 3255 16589 3337 16675
rect 3423 16589 3516 16675
rect 3076 15163 3516 16589
rect 3076 15077 3169 15163
rect 3255 15077 3337 15163
rect 3423 15077 3516 15163
rect 3076 13651 3516 15077
rect 3076 13565 3169 13651
rect 3255 13565 3337 13651
rect 3423 13565 3516 13651
rect 3076 12139 3516 13565
rect 3076 12053 3169 12139
rect 3255 12053 3337 12139
rect 3423 12053 3516 12139
rect 3076 10627 3516 12053
rect 3076 10541 3169 10627
rect 3255 10541 3337 10627
rect 3423 10541 3516 10627
rect 3076 9115 3516 10541
rect 3076 9029 3169 9115
rect 3255 9029 3337 9115
rect 3423 9029 3516 9115
rect 3076 7603 3516 9029
rect 3076 7517 3169 7603
rect 3255 7517 3337 7603
rect 3423 7517 3516 7603
rect 3076 6091 3516 7517
rect 3076 6005 3169 6091
rect 3255 6005 3337 6091
rect 3423 6005 3516 6091
rect 3076 4579 3516 6005
rect 3076 4493 3169 4579
rect 3255 4493 3337 4579
rect 3423 4493 3516 4579
rect 3076 3067 3516 4493
rect 3076 2981 3169 3067
rect 3255 2981 3337 3067
rect 3423 2981 3516 3067
rect 3076 1555 3516 2981
rect 3076 1469 3169 1555
rect 3255 1469 3337 1555
rect 3423 1469 3516 1555
rect 3076 712 3516 1469
rect 4316 38599 4756 38682
rect 4316 38513 4409 38599
rect 4495 38513 4577 38599
rect 4663 38513 4756 38599
rect 4316 37087 4756 38513
rect 4316 37001 4409 37087
rect 4495 37001 4577 37087
rect 4663 37001 4756 37087
rect 4316 35575 4756 37001
rect 4316 35489 4409 35575
rect 4495 35489 4577 35575
rect 4663 35489 4756 35575
rect 4316 34063 4756 35489
rect 4316 33977 4409 34063
rect 4495 33977 4577 34063
rect 4663 33977 4756 34063
rect 4316 32551 4756 33977
rect 4316 32465 4409 32551
rect 4495 32465 4577 32551
rect 4663 32465 4756 32551
rect 4316 31039 4756 32465
rect 4316 30953 4409 31039
rect 4495 30953 4577 31039
rect 4663 30953 4756 31039
rect 4316 29527 4756 30953
rect 4316 29441 4409 29527
rect 4495 29441 4577 29527
rect 4663 29441 4756 29527
rect 4316 28015 4756 29441
rect 4316 27929 4409 28015
rect 4495 27929 4577 28015
rect 4663 27929 4756 28015
rect 4316 26503 4756 27929
rect 4316 26417 4409 26503
rect 4495 26417 4577 26503
rect 4663 26417 4756 26503
rect 4316 24991 4756 26417
rect 4316 24905 4409 24991
rect 4495 24905 4577 24991
rect 4663 24905 4756 24991
rect 4316 23479 4756 24905
rect 4316 23393 4409 23479
rect 4495 23393 4577 23479
rect 4663 23393 4756 23479
rect 4316 21967 4756 23393
rect 4316 21881 4409 21967
rect 4495 21881 4577 21967
rect 4663 21881 4756 21967
rect 4316 20455 4756 21881
rect 4316 20369 4409 20455
rect 4495 20369 4577 20455
rect 4663 20369 4756 20455
rect 4316 18943 4756 20369
rect 4316 18857 4409 18943
rect 4495 18857 4577 18943
rect 4663 18857 4756 18943
rect 4316 17431 4756 18857
rect 4316 17345 4409 17431
rect 4495 17345 4577 17431
rect 4663 17345 4756 17431
rect 4316 15919 4756 17345
rect 4316 15833 4409 15919
rect 4495 15833 4577 15919
rect 4663 15833 4756 15919
rect 4316 14407 4756 15833
rect 4316 14321 4409 14407
rect 4495 14321 4577 14407
rect 4663 14321 4756 14407
rect 4316 12895 4756 14321
rect 4316 12809 4409 12895
rect 4495 12809 4577 12895
rect 4663 12809 4756 12895
rect 4316 11383 4756 12809
rect 4316 11297 4409 11383
rect 4495 11297 4577 11383
rect 4663 11297 4756 11383
rect 4316 9871 4756 11297
rect 4316 9785 4409 9871
rect 4495 9785 4577 9871
rect 4663 9785 4756 9871
rect 4316 8359 4756 9785
rect 4316 8273 4409 8359
rect 4495 8273 4577 8359
rect 4663 8273 4756 8359
rect 4316 6847 4756 8273
rect 4316 6761 4409 6847
rect 4495 6761 4577 6847
rect 4663 6761 4756 6847
rect 4316 5335 4756 6761
rect 4316 5249 4409 5335
rect 4495 5249 4577 5335
rect 4663 5249 4756 5335
rect 4316 3823 4756 5249
rect 4316 3737 4409 3823
rect 4495 3737 4577 3823
rect 4663 3737 4756 3823
rect 4316 2311 4756 3737
rect 4316 2225 4409 2311
rect 4495 2225 4577 2311
rect 4663 2225 4756 2311
rect 4316 799 4756 2225
rect 4316 713 4409 799
rect 4495 713 4577 799
rect 4663 713 4756 799
rect 4316 630 4756 713
rect 18196 37843 18636 38600
rect 18196 37757 18289 37843
rect 18375 37757 18457 37843
rect 18543 37757 18636 37843
rect 18196 36331 18636 37757
rect 18196 36245 18289 36331
rect 18375 36245 18457 36331
rect 18543 36245 18636 36331
rect 18196 34819 18636 36245
rect 18196 34733 18289 34819
rect 18375 34733 18457 34819
rect 18543 34733 18636 34819
rect 18196 33307 18636 34733
rect 18196 33221 18289 33307
rect 18375 33221 18457 33307
rect 18543 33221 18636 33307
rect 18196 31795 18636 33221
rect 18196 31709 18289 31795
rect 18375 31709 18457 31795
rect 18543 31709 18636 31795
rect 18196 30283 18636 31709
rect 18196 30197 18289 30283
rect 18375 30197 18457 30283
rect 18543 30197 18636 30283
rect 18196 28771 18636 30197
rect 18196 28685 18289 28771
rect 18375 28685 18457 28771
rect 18543 28685 18636 28771
rect 18196 27259 18636 28685
rect 18196 27173 18289 27259
rect 18375 27173 18457 27259
rect 18543 27173 18636 27259
rect 18196 25747 18636 27173
rect 18196 25661 18289 25747
rect 18375 25661 18457 25747
rect 18543 25661 18636 25747
rect 18196 24235 18636 25661
rect 18196 24149 18289 24235
rect 18375 24149 18457 24235
rect 18543 24149 18636 24235
rect 18196 22723 18636 24149
rect 18196 22637 18289 22723
rect 18375 22637 18457 22723
rect 18543 22637 18636 22723
rect 18196 21211 18636 22637
rect 18196 21125 18289 21211
rect 18375 21125 18457 21211
rect 18543 21125 18636 21211
rect 18196 19699 18636 21125
rect 18196 19613 18289 19699
rect 18375 19613 18457 19699
rect 18543 19613 18636 19699
rect 18196 18187 18636 19613
rect 18196 18101 18289 18187
rect 18375 18101 18457 18187
rect 18543 18101 18636 18187
rect 18196 16675 18636 18101
rect 18196 16589 18289 16675
rect 18375 16589 18457 16675
rect 18543 16589 18636 16675
rect 18196 15163 18636 16589
rect 18196 15077 18289 15163
rect 18375 15077 18457 15163
rect 18543 15077 18636 15163
rect 18196 13651 18636 15077
rect 18196 13565 18289 13651
rect 18375 13565 18457 13651
rect 18543 13565 18636 13651
rect 18196 12139 18636 13565
rect 18196 12053 18289 12139
rect 18375 12053 18457 12139
rect 18543 12053 18636 12139
rect 18196 10627 18636 12053
rect 18196 10541 18289 10627
rect 18375 10541 18457 10627
rect 18543 10541 18636 10627
rect 18196 9115 18636 10541
rect 18196 9029 18289 9115
rect 18375 9029 18457 9115
rect 18543 9029 18636 9115
rect 18196 7603 18636 9029
rect 18196 7517 18289 7603
rect 18375 7517 18457 7603
rect 18543 7517 18636 7603
rect 18196 6091 18636 7517
rect 18196 6005 18289 6091
rect 18375 6005 18457 6091
rect 18543 6005 18636 6091
rect 18196 4579 18636 6005
rect 18196 4493 18289 4579
rect 18375 4493 18457 4579
rect 18543 4493 18636 4579
rect 18196 3067 18636 4493
rect 18196 2981 18289 3067
rect 18375 2981 18457 3067
rect 18543 2981 18636 3067
rect 18196 1555 18636 2981
rect 18196 1469 18289 1555
rect 18375 1469 18457 1555
rect 18543 1469 18636 1555
rect 18196 712 18636 1469
rect 19436 38599 19876 38682
rect 19436 38513 19529 38599
rect 19615 38513 19697 38599
rect 19783 38513 19876 38599
rect 19436 37087 19876 38513
rect 19436 37001 19529 37087
rect 19615 37001 19697 37087
rect 19783 37001 19876 37087
rect 19436 35575 19876 37001
rect 19436 35489 19529 35575
rect 19615 35489 19697 35575
rect 19783 35489 19876 35575
rect 19436 34063 19876 35489
rect 19436 33977 19529 34063
rect 19615 33977 19697 34063
rect 19783 33977 19876 34063
rect 19436 32551 19876 33977
rect 19436 32465 19529 32551
rect 19615 32465 19697 32551
rect 19783 32465 19876 32551
rect 19436 31039 19876 32465
rect 19436 30953 19529 31039
rect 19615 30953 19697 31039
rect 19783 30953 19876 31039
rect 19436 29527 19876 30953
rect 19436 29441 19529 29527
rect 19615 29441 19697 29527
rect 19783 29441 19876 29527
rect 19436 28015 19876 29441
rect 19436 27929 19529 28015
rect 19615 27929 19697 28015
rect 19783 27929 19876 28015
rect 19436 26503 19876 27929
rect 19436 26417 19529 26503
rect 19615 26417 19697 26503
rect 19783 26417 19876 26503
rect 19436 24991 19876 26417
rect 19436 24905 19529 24991
rect 19615 24905 19697 24991
rect 19783 24905 19876 24991
rect 19436 23479 19876 24905
rect 19436 23393 19529 23479
rect 19615 23393 19697 23479
rect 19783 23393 19876 23479
rect 19436 21967 19876 23393
rect 19436 21881 19529 21967
rect 19615 21881 19697 21967
rect 19783 21881 19876 21967
rect 19436 20455 19876 21881
rect 19436 20369 19529 20455
rect 19615 20369 19697 20455
rect 19783 20369 19876 20455
rect 19436 18943 19876 20369
rect 19436 18857 19529 18943
rect 19615 18857 19697 18943
rect 19783 18857 19876 18943
rect 19436 17431 19876 18857
rect 19436 17345 19529 17431
rect 19615 17345 19697 17431
rect 19783 17345 19876 17431
rect 19436 15919 19876 17345
rect 19436 15833 19529 15919
rect 19615 15833 19697 15919
rect 19783 15833 19876 15919
rect 19436 14407 19876 15833
rect 19436 14321 19529 14407
rect 19615 14321 19697 14407
rect 19783 14321 19876 14407
rect 19436 12895 19876 14321
rect 19436 12809 19529 12895
rect 19615 12809 19697 12895
rect 19783 12809 19876 12895
rect 19436 11383 19876 12809
rect 19436 11297 19529 11383
rect 19615 11297 19697 11383
rect 19783 11297 19876 11383
rect 19436 9871 19876 11297
rect 19436 9785 19529 9871
rect 19615 9785 19697 9871
rect 19783 9785 19876 9871
rect 19436 8359 19876 9785
rect 19436 8273 19529 8359
rect 19615 8273 19697 8359
rect 19783 8273 19876 8359
rect 19436 6847 19876 8273
rect 19436 6761 19529 6847
rect 19615 6761 19697 6847
rect 19783 6761 19876 6847
rect 19436 5335 19876 6761
rect 19436 5249 19529 5335
rect 19615 5249 19697 5335
rect 19783 5249 19876 5335
rect 19436 3823 19876 5249
rect 19436 3737 19529 3823
rect 19615 3737 19697 3823
rect 19783 3737 19876 3823
rect 19436 2311 19876 3737
rect 19436 2225 19529 2311
rect 19615 2225 19697 2311
rect 19783 2225 19876 2311
rect 19436 799 19876 2225
rect 19436 713 19529 799
rect 19615 713 19697 799
rect 19783 713 19876 799
rect 19436 630 19876 713
rect 33316 37843 33756 38600
rect 33316 37757 33409 37843
rect 33495 37757 33577 37843
rect 33663 37757 33756 37843
rect 33316 36331 33756 37757
rect 33316 36245 33409 36331
rect 33495 36245 33577 36331
rect 33663 36245 33756 36331
rect 33316 34819 33756 36245
rect 33316 34733 33409 34819
rect 33495 34733 33577 34819
rect 33663 34733 33756 34819
rect 33316 33307 33756 34733
rect 33316 33221 33409 33307
rect 33495 33221 33577 33307
rect 33663 33221 33756 33307
rect 33316 31795 33756 33221
rect 33316 31709 33409 31795
rect 33495 31709 33577 31795
rect 33663 31709 33756 31795
rect 33316 30283 33756 31709
rect 33316 30197 33409 30283
rect 33495 30197 33577 30283
rect 33663 30197 33756 30283
rect 33316 28771 33756 30197
rect 33316 28685 33409 28771
rect 33495 28685 33577 28771
rect 33663 28685 33756 28771
rect 33316 27259 33756 28685
rect 33316 27173 33409 27259
rect 33495 27173 33577 27259
rect 33663 27173 33756 27259
rect 33316 25747 33756 27173
rect 33316 25661 33409 25747
rect 33495 25661 33577 25747
rect 33663 25661 33756 25747
rect 33316 24235 33756 25661
rect 33316 24149 33409 24235
rect 33495 24149 33577 24235
rect 33663 24149 33756 24235
rect 33316 22723 33756 24149
rect 33316 22637 33409 22723
rect 33495 22637 33577 22723
rect 33663 22637 33756 22723
rect 33316 21211 33756 22637
rect 33316 21125 33409 21211
rect 33495 21125 33577 21211
rect 33663 21125 33756 21211
rect 33316 19699 33756 21125
rect 33316 19613 33409 19699
rect 33495 19613 33577 19699
rect 33663 19613 33756 19699
rect 33316 18187 33756 19613
rect 33316 18101 33409 18187
rect 33495 18101 33577 18187
rect 33663 18101 33756 18187
rect 33316 16675 33756 18101
rect 33316 16589 33409 16675
rect 33495 16589 33577 16675
rect 33663 16589 33756 16675
rect 33316 15163 33756 16589
rect 33316 15077 33409 15163
rect 33495 15077 33577 15163
rect 33663 15077 33756 15163
rect 33316 13651 33756 15077
rect 33316 13565 33409 13651
rect 33495 13565 33577 13651
rect 33663 13565 33756 13651
rect 33316 12139 33756 13565
rect 33316 12053 33409 12139
rect 33495 12053 33577 12139
rect 33663 12053 33756 12139
rect 33316 10627 33756 12053
rect 33316 10541 33409 10627
rect 33495 10541 33577 10627
rect 33663 10541 33756 10627
rect 33316 9115 33756 10541
rect 33316 9029 33409 9115
rect 33495 9029 33577 9115
rect 33663 9029 33756 9115
rect 33316 7603 33756 9029
rect 33316 7517 33409 7603
rect 33495 7517 33577 7603
rect 33663 7517 33756 7603
rect 33316 6091 33756 7517
rect 33316 6005 33409 6091
rect 33495 6005 33577 6091
rect 33663 6005 33756 6091
rect 33316 4579 33756 6005
rect 33316 4493 33409 4579
rect 33495 4493 33577 4579
rect 33663 4493 33756 4579
rect 33316 3067 33756 4493
rect 33316 2981 33409 3067
rect 33495 2981 33577 3067
rect 33663 2981 33756 3067
rect 33316 1555 33756 2981
rect 33316 1469 33409 1555
rect 33495 1469 33577 1555
rect 33663 1469 33756 1555
rect 33316 712 33756 1469
rect 34556 38599 34996 38682
rect 34556 38513 34649 38599
rect 34735 38513 34817 38599
rect 34903 38513 34996 38599
rect 34556 37087 34996 38513
rect 34556 37001 34649 37087
rect 34735 37001 34817 37087
rect 34903 37001 34996 37087
rect 34556 35575 34996 37001
rect 34556 35489 34649 35575
rect 34735 35489 34817 35575
rect 34903 35489 34996 35575
rect 34556 34063 34996 35489
rect 34556 33977 34649 34063
rect 34735 33977 34817 34063
rect 34903 33977 34996 34063
rect 34556 32551 34996 33977
rect 34556 32465 34649 32551
rect 34735 32465 34817 32551
rect 34903 32465 34996 32551
rect 34556 31039 34996 32465
rect 34556 30953 34649 31039
rect 34735 30953 34817 31039
rect 34903 30953 34996 31039
rect 34556 29527 34996 30953
rect 34556 29441 34649 29527
rect 34735 29441 34817 29527
rect 34903 29441 34996 29527
rect 34556 28015 34996 29441
rect 34556 27929 34649 28015
rect 34735 27929 34817 28015
rect 34903 27929 34996 28015
rect 34556 26503 34996 27929
rect 34556 26417 34649 26503
rect 34735 26417 34817 26503
rect 34903 26417 34996 26503
rect 34556 24991 34996 26417
rect 34556 24905 34649 24991
rect 34735 24905 34817 24991
rect 34903 24905 34996 24991
rect 34556 23479 34996 24905
rect 34556 23393 34649 23479
rect 34735 23393 34817 23479
rect 34903 23393 34996 23479
rect 34556 21967 34996 23393
rect 34556 21881 34649 21967
rect 34735 21881 34817 21967
rect 34903 21881 34996 21967
rect 34556 20455 34996 21881
rect 34556 20369 34649 20455
rect 34735 20369 34817 20455
rect 34903 20369 34996 20455
rect 34556 18943 34996 20369
rect 34556 18857 34649 18943
rect 34735 18857 34817 18943
rect 34903 18857 34996 18943
rect 34556 17431 34996 18857
rect 34556 17345 34649 17431
rect 34735 17345 34817 17431
rect 34903 17345 34996 17431
rect 34556 15919 34996 17345
rect 34556 15833 34649 15919
rect 34735 15833 34817 15919
rect 34903 15833 34996 15919
rect 34556 14407 34996 15833
rect 34556 14321 34649 14407
rect 34735 14321 34817 14407
rect 34903 14321 34996 14407
rect 34556 12895 34996 14321
rect 34556 12809 34649 12895
rect 34735 12809 34817 12895
rect 34903 12809 34996 12895
rect 34556 11383 34996 12809
rect 34556 11297 34649 11383
rect 34735 11297 34817 11383
rect 34903 11297 34996 11383
rect 34556 9871 34996 11297
rect 34556 9785 34649 9871
rect 34735 9785 34817 9871
rect 34903 9785 34996 9871
rect 34556 8359 34996 9785
rect 34556 8273 34649 8359
rect 34735 8273 34817 8359
rect 34903 8273 34996 8359
rect 34556 6847 34996 8273
rect 34556 6761 34649 6847
rect 34735 6761 34817 6847
rect 34903 6761 34996 6847
rect 34556 5335 34996 6761
rect 34556 5249 34649 5335
rect 34735 5249 34817 5335
rect 34903 5249 34996 5335
rect 34556 3823 34996 5249
rect 34556 3737 34649 3823
rect 34735 3737 34817 3823
rect 34903 3737 34996 3823
rect 34556 2311 34996 3737
rect 34556 2225 34649 2311
rect 34735 2225 34817 2311
rect 34903 2225 34996 2311
rect 34556 799 34996 2225
rect 34556 713 34649 799
rect 34735 713 34817 799
rect 34903 713 34996 799
rect 34556 630 34996 713
rect 48436 37843 48876 38600
rect 48436 37757 48529 37843
rect 48615 37757 48697 37843
rect 48783 37757 48876 37843
rect 48436 36331 48876 37757
rect 48436 36245 48529 36331
rect 48615 36245 48697 36331
rect 48783 36245 48876 36331
rect 48436 34819 48876 36245
rect 48436 34733 48529 34819
rect 48615 34733 48697 34819
rect 48783 34733 48876 34819
rect 48436 33307 48876 34733
rect 48436 33221 48529 33307
rect 48615 33221 48697 33307
rect 48783 33221 48876 33307
rect 48436 31795 48876 33221
rect 48436 31709 48529 31795
rect 48615 31709 48697 31795
rect 48783 31709 48876 31795
rect 48436 30283 48876 31709
rect 48436 30197 48529 30283
rect 48615 30197 48697 30283
rect 48783 30197 48876 30283
rect 48436 28771 48876 30197
rect 48436 28685 48529 28771
rect 48615 28685 48697 28771
rect 48783 28685 48876 28771
rect 48436 27259 48876 28685
rect 48436 27173 48529 27259
rect 48615 27173 48697 27259
rect 48783 27173 48876 27259
rect 48436 25747 48876 27173
rect 48436 25661 48529 25747
rect 48615 25661 48697 25747
rect 48783 25661 48876 25747
rect 48436 24235 48876 25661
rect 48436 24149 48529 24235
rect 48615 24149 48697 24235
rect 48783 24149 48876 24235
rect 48436 22723 48876 24149
rect 48436 22637 48529 22723
rect 48615 22637 48697 22723
rect 48783 22637 48876 22723
rect 48436 21211 48876 22637
rect 48436 21125 48529 21211
rect 48615 21125 48697 21211
rect 48783 21125 48876 21211
rect 48436 19699 48876 21125
rect 48436 19613 48529 19699
rect 48615 19613 48697 19699
rect 48783 19613 48876 19699
rect 48436 18187 48876 19613
rect 48436 18101 48529 18187
rect 48615 18101 48697 18187
rect 48783 18101 48876 18187
rect 48436 16675 48876 18101
rect 48436 16589 48529 16675
rect 48615 16589 48697 16675
rect 48783 16589 48876 16675
rect 48436 15163 48876 16589
rect 48436 15077 48529 15163
rect 48615 15077 48697 15163
rect 48783 15077 48876 15163
rect 48436 13651 48876 15077
rect 48436 13565 48529 13651
rect 48615 13565 48697 13651
rect 48783 13565 48876 13651
rect 48436 12139 48876 13565
rect 48436 12053 48529 12139
rect 48615 12053 48697 12139
rect 48783 12053 48876 12139
rect 48436 10627 48876 12053
rect 48436 10541 48529 10627
rect 48615 10541 48697 10627
rect 48783 10541 48876 10627
rect 48436 9115 48876 10541
rect 48436 9029 48529 9115
rect 48615 9029 48697 9115
rect 48783 9029 48876 9115
rect 48436 7603 48876 9029
rect 48436 7517 48529 7603
rect 48615 7517 48697 7603
rect 48783 7517 48876 7603
rect 48436 6091 48876 7517
rect 48436 6005 48529 6091
rect 48615 6005 48697 6091
rect 48783 6005 48876 6091
rect 48436 4579 48876 6005
rect 48436 4493 48529 4579
rect 48615 4493 48697 4579
rect 48783 4493 48876 4579
rect 48436 3067 48876 4493
rect 48436 2981 48529 3067
rect 48615 2981 48697 3067
rect 48783 2981 48876 3067
rect 48436 1555 48876 2981
rect 48436 1469 48529 1555
rect 48615 1469 48697 1555
rect 48783 1469 48876 1555
rect 48436 712 48876 1469
rect 49676 38599 50116 38682
rect 49676 38513 49769 38599
rect 49855 38513 49937 38599
rect 50023 38513 50116 38599
rect 49676 37087 50116 38513
rect 49676 37001 49769 37087
rect 49855 37001 49937 37087
rect 50023 37001 50116 37087
rect 49676 35575 50116 37001
rect 49676 35489 49769 35575
rect 49855 35489 49937 35575
rect 50023 35489 50116 35575
rect 49676 34063 50116 35489
rect 49676 33977 49769 34063
rect 49855 33977 49937 34063
rect 50023 33977 50116 34063
rect 49676 32551 50116 33977
rect 49676 32465 49769 32551
rect 49855 32465 49937 32551
rect 50023 32465 50116 32551
rect 49676 31039 50116 32465
rect 49676 30953 49769 31039
rect 49855 30953 49937 31039
rect 50023 30953 50116 31039
rect 49676 29527 50116 30953
rect 49676 29441 49769 29527
rect 49855 29441 49937 29527
rect 50023 29441 50116 29527
rect 49676 28015 50116 29441
rect 49676 27929 49769 28015
rect 49855 27929 49937 28015
rect 50023 27929 50116 28015
rect 49676 26503 50116 27929
rect 49676 26417 49769 26503
rect 49855 26417 49937 26503
rect 50023 26417 50116 26503
rect 49676 24991 50116 26417
rect 49676 24905 49769 24991
rect 49855 24905 49937 24991
rect 50023 24905 50116 24991
rect 49676 23479 50116 24905
rect 49676 23393 49769 23479
rect 49855 23393 49937 23479
rect 50023 23393 50116 23479
rect 49676 21967 50116 23393
rect 49676 21881 49769 21967
rect 49855 21881 49937 21967
rect 50023 21881 50116 21967
rect 49676 20455 50116 21881
rect 49676 20369 49769 20455
rect 49855 20369 49937 20455
rect 50023 20369 50116 20455
rect 49676 18943 50116 20369
rect 49676 18857 49769 18943
rect 49855 18857 49937 18943
rect 50023 18857 50116 18943
rect 49676 17431 50116 18857
rect 49676 17345 49769 17431
rect 49855 17345 49937 17431
rect 50023 17345 50116 17431
rect 49676 15919 50116 17345
rect 49676 15833 49769 15919
rect 49855 15833 49937 15919
rect 50023 15833 50116 15919
rect 49676 14407 50116 15833
rect 49676 14321 49769 14407
rect 49855 14321 49937 14407
rect 50023 14321 50116 14407
rect 49676 12895 50116 14321
rect 49676 12809 49769 12895
rect 49855 12809 49937 12895
rect 50023 12809 50116 12895
rect 49676 11383 50116 12809
rect 49676 11297 49769 11383
rect 49855 11297 49937 11383
rect 50023 11297 50116 11383
rect 49676 9871 50116 11297
rect 49676 9785 49769 9871
rect 49855 9785 49937 9871
rect 50023 9785 50116 9871
rect 49676 8359 50116 9785
rect 49676 8273 49769 8359
rect 49855 8273 49937 8359
rect 50023 8273 50116 8359
rect 49676 6847 50116 8273
rect 49676 6761 49769 6847
rect 49855 6761 49937 6847
rect 50023 6761 50116 6847
rect 49676 5335 50116 6761
rect 49676 5249 49769 5335
rect 49855 5249 49937 5335
rect 50023 5249 50116 5335
rect 49676 3823 50116 5249
rect 49676 3737 49769 3823
rect 49855 3737 49937 3823
rect 50023 3737 50116 3823
rect 49676 2311 50116 3737
rect 49676 2225 49769 2311
rect 49855 2225 49937 2311
rect 50023 2225 50116 2311
rect 49676 799 50116 2225
rect 49676 713 49769 799
rect 49855 713 49937 799
rect 50023 713 50116 799
rect 49676 630 50116 713
rect 63556 37843 63996 38600
rect 63556 37757 63649 37843
rect 63735 37757 63817 37843
rect 63903 37757 63996 37843
rect 63556 36331 63996 37757
rect 63556 36245 63649 36331
rect 63735 36245 63817 36331
rect 63903 36245 63996 36331
rect 63556 34819 63996 36245
rect 63556 34733 63649 34819
rect 63735 34733 63817 34819
rect 63903 34733 63996 34819
rect 63556 33307 63996 34733
rect 63556 33221 63649 33307
rect 63735 33221 63817 33307
rect 63903 33221 63996 33307
rect 63556 31795 63996 33221
rect 63556 31709 63649 31795
rect 63735 31709 63817 31795
rect 63903 31709 63996 31795
rect 63556 30283 63996 31709
rect 63556 30197 63649 30283
rect 63735 30197 63817 30283
rect 63903 30197 63996 30283
rect 63556 28771 63996 30197
rect 63556 28685 63649 28771
rect 63735 28685 63817 28771
rect 63903 28685 63996 28771
rect 63556 27259 63996 28685
rect 63556 27173 63649 27259
rect 63735 27173 63817 27259
rect 63903 27173 63996 27259
rect 63556 25747 63996 27173
rect 63556 25661 63649 25747
rect 63735 25661 63817 25747
rect 63903 25661 63996 25747
rect 63556 24235 63996 25661
rect 63556 24149 63649 24235
rect 63735 24149 63817 24235
rect 63903 24149 63996 24235
rect 63556 22723 63996 24149
rect 63556 22637 63649 22723
rect 63735 22637 63817 22723
rect 63903 22637 63996 22723
rect 63556 21211 63996 22637
rect 63556 21125 63649 21211
rect 63735 21125 63817 21211
rect 63903 21125 63996 21211
rect 63556 19699 63996 21125
rect 63556 19613 63649 19699
rect 63735 19613 63817 19699
rect 63903 19613 63996 19699
rect 63556 18187 63996 19613
rect 63556 18101 63649 18187
rect 63735 18101 63817 18187
rect 63903 18101 63996 18187
rect 63556 16675 63996 18101
rect 63556 16589 63649 16675
rect 63735 16589 63817 16675
rect 63903 16589 63996 16675
rect 63556 15163 63996 16589
rect 63556 15077 63649 15163
rect 63735 15077 63817 15163
rect 63903 15077 63996 15163
rect 63556 13651 63996 15077
rect 63556 13565 63649 13651
rect 63735 13565 63817 13651
rect 63903 13565 63996 13651
rect 63556 12139 63996 13565
rect 63556 12053 63649 12139
rect 63735 12053 63817 12139
rect 63903 12053 63996 12139
rect 63556 10627 63996 12053
rect 63556 10541 63649 10627
rect 63735 10541 63817 10627
rect 63903 10541 63996 10627
rect 63556 9115 63996 10541
rect 63556 9029 63649 9115
rect 63735 9029 63817 9115
rect 63903 9029 63996 9115
rect 63556 7603 63996 9029
rect 63556 7517 63649 7603
rect 63735 7517 63817 7603
rect 63903 7517 63996 7603
rect 63556 6091 63996 7517
rect 63556 6005 63649 6091
rect 63735 6005 63817 6091
rect 63903 6005 63996 6091
rect 63556 4579 63996 6005
rect 63556 4493 63649 4579
rect 63735 4493 63817 4579
rect 63903 4493 63996 4579
rect 63556 3067 63996 4493
rect 63556 2981 63649 3067
rect 63735 2981 63817 3067
rect 63903 2981 63996 3067
rect 63556 1555 63996 2981
rect 63556 1469 63649 1555
rect 63735 1469 63817 1555
rect 63903 1469 63996 1555
rect 63556 712 63996 1469
rect 64796 38599 65236 38682
rect 64796 38513 64889 38599
rect 64975 38513 65057 38599
rect 65143 38513 65236 38599
rect 64796 37087 65236 38513
rect 64796 37001 64889 37087
rect 64975 37001 65057 37087
rect 65143 37001 65236 37087
rect 64796 35575 65236 37001
rect 64796 35489 64889 35575
rect 64975 35489 65057 35575
rect 65143 35489 65236 35575
rect 64796 34063 65236 35489
rect 64796 33977 64889 34063
rect 64975 33977 65057 34063
rect 65143 33977 65236 34063
rect 64796 32551 65236 33977
rect 64796 32465 64889 32551
rect 64975 32465 65057 32551
rect 65143 32465 65236 32551
rect 64796 31039 65236 32465
rect 64796 30953 64889 31039
rect 64975 30953 65057 31039
rect 65143 30953 65236 31039
rect 64796 29527 65236 30953
rect 64796 29441 64889 29527
rect 64975 29441 65057 29527
rect 65143 29441 65236 29527
rect 64796 28015 65236 29441
rect 64796 27929 64889 28015
rect 64975 27929 65057 28015
rect 65143 27929 65236 28015
rect 64796 26503 65236 27929
rect 64796 26417 64889 26503
rect 64975 26417 65057 26503
rect 65143 26417 65236 26503
rect 64796 24991 65236 26417
rect 64796 24905 64889 24991
rect 64975 24905 65057 24991
rect 65143 24905 65236 24991
rect 64796 23479 65236 24905
rect 64796 23393 64889 23479
rect 64975 23393 65057 23479
rect 65143 23393 65236 23479
rect 64796 21967 65236 23393
rect 64796 21881 64889 21967
rect 64975 21881 65057 21967
rect 65143 21881 65236 21967
rect 64796 20455 65236 21881
rect 64796 20369 64889 20455
rect 64975 20369 65057 20455
rect 65143 20369 65236 20455
rect 64796 18943 65236 20369
rect 64796 18857 64889 18943
rect 64975 18857 65057 18943
rect 65143 18857 65236 18943
rect 64796 17431 65236 18857
rect 64796 17345 64889 17431
rect 64975 17345 65057 17431
rect 65143 17345 65236 17431
rect 64796 15919 65236 17345
rect 64796 15833 64889 15919
rect 64975 15833 65057 15919
rect 65143 15833 65236 15919
rect 64796 14407 65236 15833
rect 64796 14321 64889 14407
rect 64975 14321 65057 14407
rect 65143 14321 65236 14407
rect 64796 12895 65236 14321
rect 64796 12809 64889 12895
rect 64975 12809 65057 12895
rect 65143 12809 65236 12895
rect 64796 11383 65236 12809
rect 64796 11297 64889 11383
rect 64975 11297 65057 11383
rect 65143 11297 65236 11383
rect 64796 9871 65236 11297
rect 64796 9785 64889 9871
rect 64975 9785 65057 9871
rect 65143 9785 65236 9871
rect 64796 8359 65236 9785
rect 64796 8273 64889 8359
rect 64975 8273 65057 8359
rect 65143 8273 65236 8359
rect 64796 6847 65236 8273
rect 64796 6761 64889 6847
rect 64975 6761 65057 6847
rect 65143 6761 65236 6847
rect 64796 5335 65236 6761
rect 64796 5249 64889 5335
rect 64975 5249 65057 5335
rect 65143 5249 65236 5335
rect 64796 3823 65236 5249
rect 64796 3737 64889 3823
rect 64975 3737 65057 3823
rect 65143 3737 65236 3823
rect 64796 2311 65236 3737
rect 64796 2225 64889 2311
rect 64975 2225 65057 2311
rect 65143 2225 65236 2311
rect 64796 799 65236 2225
rect 64796 713 64889 799
rect 64975 713 65057 799
rect 65143 713 65236 799
rect 64796 630 65236 713
rect 78676 37843 79116 38600
rect 78676 37757 78769 37843
rect 78855 37757 78937 37843
rect 79023 37757 79116 37843
rect 78676 36331 79116 37757
rect 78676 36245 78769 36331
rect 78855 36245 78937 36331
rect 79023 36245 79116 36331
rect 78676 34819 79116 36245
rect 78676 34733 78769 34819
rect 78855 34733 78937 34819
rect 79023 34733 79116 34819
rect 78676 33307 79116 34733
rect 78676 33221 78769 33307
rect 78855 33221 78937 33307
rect 79023 33221 79116 33307
rect 78676 31795 79116 33221
rect 78676 31709 78769 31795
rect 78855 31709 78937 31795
rect 79023 31709 79116 31795
rect 78676 30283 79116 31709
rect 78676 30197 78769 30283
rect 78855 30197 78937 30283
rect 79023 30197 79116 30283
rect 78676 28771 79116 30197
rect 78676 28685 78769 28771
rect 78855 28685 78937 28771
rect 79023 28685 79116 28771
rect 78676 27259 79116 28685
rect 78676 27173 78769 27259
rect 78855 27173 78937 27259
rect 79023 27173 79116 27259
rect 78676 25747 79116 27173
rect 78676 25661 78769 25747
rect 78855 25661 78937 25747
rect 79023 25661 79116 25747
rect 78676 24235 79116 25661
rect 78676 24149 78769 24235
rect 78855 24149 78937 24235
rect 79023 24149 79116 24235
rect 78676 22723 79116 24149
rect 78676 22637 78769 22723
rect 78855 22637 78937 22723
rect 79023 22637 79116 22723
rect 78676 21211 79116 22637
rect 78676 21125 78769 21211
rect 78855 21125 78937 21211
rect 79023 21125 79116 21211
rect 78676 19699 79116 21125
rect 78676 19613 78769 19699
rect 78855 19613 78937 19699
rect 79023 19613 79116 19699
rect 78676 18187 79116 19613
rect 78676 18101 78769 18187
rect 78855 18101 78937 18187
rect 79023 18101 79116 18187
rect 78676 16675 79116 18101
rect 78676 16589 78769 16675
rect 78855 16589 78937 16675
rect 79023 16589 79116 16675
rect 78676 15163 79116 16589
rect 78676 15077 78769 15163
rect 78855 15077 78937 15163
rect 79023 15077 79116 15163
rect 78676 13651 79116 15077
rect 78676 13565 78769 13651
rect 78855 13565 78937 13651
rect 79023 13565 79116 13651
rect 78676 12139 79116 13565
rect 78676 12053 78769 12139
rect 78855 12053 78937 12139
rect 79023 12053 79116 12139
rect 78676 10627 79116 12053
rect 78676 10541 78769 10627
rect 78855 10541 78937 10627
rect 79023 10541 79116 10627
rect 78676 9115 79116 10541
rect 78676 9029 78769 9115
rect 78855 9029 78937 9115
rect 79023 9029 79116 9115
rect 78676 7603 79116 9029
rect 78676 7517 78769 7603
rect 78855 7517 78937 7603
rect 79023 7517 79116 7603
rect 78676 6091 79116 7517
rect 78676 6005 78769 6091
rect 78855 6005 78937 6091
rect 79023 6005 79116 6091
rect 78676 4579 79116 6005
rect 78676 4493 78769 4579
rect 78855 4493 78937 4579
rect 79023 4493 79116 4579
rect 78676 3067 79116 4493
rect 78676 2981 78769 3067
rect 78855 2981 78937 3067
rect 79023 2981 79116 3067
rect 78676 1555 79116 2981
rect 78676 1469 78769 1555
rect 78855 1469 78937 1555
rect 79023 1469 79116 1555
rect 78676 712 79116 1469
rect 79916 38599 80356 38682
rect 79916 38513 80009 38599
rect 80095 38513 80177 38599
rect 80263 38513 80356 38599
rect 79916 37087 80356 38513
rect 79916 37001 80009 37087
rect 80095 37001 80177 37087
rect 80263 37001 80356 37087
rect 79916 35575 80356 37001
rect 79916 35489 80009 35575
rect 80095 35489 80177 35575
rect 80263 35489 80356 35575
rect 79916 34063 80356 35489
rect 79916 33977 80009 34063
rect 80095 33977 80177 34063
rect 80263 33977 80356 34063
rect 79916 32551 80356 33977
rect 79916 32465 80009 32551
rect 80095 32465 80177 32551
rect 80263 32465 80356 32551
rect 79916 31039 80356 32465
rect 79916 30953 80009 31039
rect 80095 30953 80177 31039
rect 80263 30953 80356 31039
rect 79916 29527 80356 30953
rect 79916 29441 80009 29527
rect 80095 29441 80177 29527
rect 80263 29441 80356 29527
rect 79916 28015 80356 29441
rect 79916 27929 80009 28015
rect 80095 27929 80177 28015
rect 80263 27929 80356 28015
rect 79916 26503 80356 27929
rect 79916 26417 80009 26503
rect 80095 26417 80177 26503
rect 80263 26417 80356 26503
rect 79916 24991 80356 26417
rect 79916 24905 80009 24991
rect 80095 24905 80177 24991
rect 80263 24905 80356 24991
rect 79916 23479 80356 24905
rect 79916 23393 80009 23479
rect 80095 23393 80177 23479
rect 80263 23393 80356 23479
rect 79916 21967 80356 23393
rect 79916 21881 80009 21967
rect 80095 21881 80177 21967
rect 80263 21881 80356 21967
rect 79916 20455 80356 21881
rect 79916 20369 80009 20455
rect 80095 20369 80177 20455
rect 80263 20369 80356 20455
rect 79916 18943 80356 20369
rect 79916 18857 80009 18943
rect 80095 18857 80177 18943
rect 80263 18857 80356 18943
rect 79916 17431 80356 18857
rect 79916 17345 80009 17431
rect 80095 17345 80177 17431
rect 80263 17345 80356 17431
rect 79916 15919 80356 17345
rect 79916 15833 80009 15919
rect 80095 15833 80177 15919
rect 80263 15833 80356 15919
rect 79916 14407 80356 15833
rect 79916 14321 80009 14407
rect 80095 14321 80177 14407
rect 80263 14321 80356 14407
rect 79916 12895 80356 14321
rect 79916 12809 80009 12895
rect 80095 12809 80177 12895
rect 80263 12809 80356 12895
rect 79916 11383 80356 12809
rect 79916 11297 80009 11383
rect 80095 11297 80177 11383
rect 80263 11297 80356 11383
rect 79916 9871 80356 11297
rect 79916 9785 80009 9871
rect 80095 9785 80177 9871
rect 80263 9785 80356 9871
rect 79916 8359 80356 9785
rect 79916 8273 80009 8359
rect 80095 8273 80177 8359
rect 80263 8273 80356 8359
rect 79916 6847 80356 8273
rect 79916 6761 80009 6847
rect 80095 6761 80177 6847
rect 80263 6761 80356 6847
rect 79916 5335 80356 6761
rect 79916 5249 80009 5335
rect 80095 5249 80177 5335
rect 80263 5249 80356 5335
rect 79916 3823 80356 5249
rect 79916 3737 80009 3823
rect 80095 3737 80177 3823
rect 80263 3737 80356 3823
rect 79916 2311 80356 3737
rect 79916 2225 80009 2311
rect 80095 2225 80177 2311
rect 80263 2225 80356 2311
rect 79916 799 80356 2225
rect 79916 713 80009 799
rect 80095 713 80177 799
rect 80263 713 80356 799
rect 79916 630 80356 713
use sg13g2_and2_1  _29_
timestamp 1676901763
transform 1 0 3936 0 1 20412
box -48 -56 528 834
use sg13g2_and2_1  _30_
timestamp 1676901763
transform 1 0 7968 0 1 18900
box -48 -56 528 834
use sg13g2_xor2_1  _31_
timestamp 1677577977
transform -1 0 9216 0 -1 20412
box -48 -56 816 834
use sg13g2_xor2_1  _32_
timestamp 1677577977
transform -1 0 8448 0 -1 20412
box -48 -56 816 834
use sg13g2_a21oi_2  _33_
timestamp 1685174172
transform 1 0 8256 0 1 20412
box -48 -56 816 834
use sg13g2_and2_1  _34_
timestamp 1676901763
transform -1 0 12480 0 -1 23436
box -48 -56 528 834
use sg13g2_xnor2_1  _35_
timestamp 1677516600
transform -1 0 12576 0 1 21924
box -48 -56 816 834
use sg13g2_nor2_1  _36_
timestamp 1676627187
transform 1 0 11136 0 1 23436
box -48 -56 432 834
use sg13g2_xor2_1  _37_
timestamp 1677577977
transform -1 0 11712 0 1 21924
box -48 -56 816 834
use sg13g2_or2_1  _38_
timestamp 1684236171
transform 1 0 10656 0 1 26460
box -48 -56 528 834
use sg13g2_and2_1  _39_
timestamp 1676901763
transform -1 0 11520 0 -1 27972
box -48 -56 528 834
use sg13g2_xor2_1  _40_
timestamp 1677577977
transform 1 0 11136 0 1 26460
box -48 -56 816 834
use sg13g2_nor2_1  _41_
timestamp 1676627187
transform 1 0 11904 0 -1 24948
box -48 -56 432 834
use sg13g2_xnor2_1  _42_
timestamp 1677516600
transform -1 0 13056 0 1 24948
box -48 -56 816 834
use sg13g2_nand2b_1  _43_
timestamp 1676567195
transform -1 0 11232 0 -1 24948
box -48 -56 528 834
use sg13g2_a21oi_1  _44_
timestamp 1683973020
transform 1 0 11040 0 -1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  _45_
timestamp 1685175443
transform -1 0 10176 0 -1 24948
box -48 -56 538 834
use sg13g2_nand2_1  _46_
timestamp 1676557249
transform 1 0 1728 0 1 23436
box -48 -56 432 834
use sg13g2_xor2_1  _47_
timestamp 1677577977
transform 1 0 2112 0 1 23436
box -48 -56 816 834
use sg13g2_inv_1  _48_
timestamp 1676382929
transform 1 0 4608 0 -1 24948
box -48 -56 336 834
use sg13g2_nand2_1  _49_
timestamp 1676557249
transform -1 0 4416 0 1 23436
box -48 -56 432 834
use sg13g2_xnor2_1  _50_
timestamp 1677516600
transform -1 0 7008 0 -1 24948
box -48 -56 816 834
use sg13g2_nor2_1  _51_
timestamp 1676627187
transform 1 0 3360 0 1 26460
box -48 -56 432 834
use sg13g2_xnor2_1  _52_
timestamp 1677516600
transform 1 0 4512 0 1 26460
box -48 -56 816 834
use sg13g2_nand2_1  _53_
timestamp 1676557249
transform 1 0 4032 0 -1 24948
box -48 -56 432 834
use sg13g2_xnor2_1  _54_
timestamp 1677516600
transform -1 0 5952 0 -1 24948
box -48 -56 816 834
use sg13g2_nor2_1  _55_
timestamp 1676627187
transform -1 0 5472 0 -1 26460
box -48 -56 432 834
use sg13g2_nor2_1  _56_
timestamp 1676627187
transform 1 0 3360 0 -1 26460
box -48 -56 432 834
use sg13g2_a221oi_1  _57_
timestamp 1685197497
transform 1 0 3744 0 1 26460
box -48 -56 816 834
use sg13g2_nand2_1  _58_
timestamp 1676557249
transform 1 0 2976 0 -1 30996
box -48 -56 432 834
use sg13g2_nor2_1  _59_
timestamp 1676627187
transform 1 0 2592 0 -1 30996
box -48 -56 432 834
use sg13g2_xor2_1  _60_
timestamp 1677577977
transform 1 0 2208 0 1 29484
box -48 -56 816 834
use sg13g2_xnor2_1  _61_
timestamp 1677516600
transform -1 0 3744 0 1 29484
box -48 -56 816 834
use sg13g2_o21ai_1  _62_
timestamp 1685175443
transform 1 0 3456 0 -1 30996
box -48 -56 538 834
use sg13g2_xnor2_1  _63_
timestamp 1677516600
transform 1 0 3936 0 1 32508
box -48 -56 816 834
use sg13g2_xnor2_1  _64_
timestamp 1677516600
transform -1 0 4800 0 -1 32508
box -48 -56 816 834
use sg13g2_xor2_1  _65_
timestamp 1677577977
transform -1 0 3936 0 1 20412
box -48 -56 816 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1679581782
transform 1 0 576 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1679581782
transform 1 0 1248 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1679581782
transform 1 0 1920 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_21
timestamp 1679581782
transform 1 0 2592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_28
timestamp 1679581782
transform 1 0 3264 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_35
timestamp 1679581782
transform 1 0 3936 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_42
timestamp 1679581782
transform 1 0 4608 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_49
timestamp 1679581782
transform 1 0 5280 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_56
timestamp 1679581782
transform 1 0 5952 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_63
timestamp 1679581782
transform 1 0 6624 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_70
timestamp 1679581782
transform 1 0 7296 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_77
timestamp 1679581782
transform 1 0 7968 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_84
timestamp 1679581782
transform 1 0 8640 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_91
timestamp 1679581782
transform 1 0 9312 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_98
timestamp 1679581782
transform 1 0 9984 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_105
timestamp 1679581782
transform 1 0 10656 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_112
timestamp 1679581782
transform 1 0 11328 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_119
timestamp 1679581782
transform 1 0 12000 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_126
timestamp 1679581782
transform 1 0 12672 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_133
timestamp 1679581782
transform 1 0 13344 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_140
timestamp 1679581782
transform 1 0 14016 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_147
timestamp 1679581782
transform 1 0 14688 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_154
timestamp 1679581782
transform 1 0 15360 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_161
timestamp 1679581782
transform 1 0 16032 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_168
timestamp 1679581782
transform 1 0 16704 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_175
timestamp 1679581782
transform 1 0 17376 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_182
timestamp 1679581782
transform 1 0 18048 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_189
timestamp 1679581782
transform 1 0 18720 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_196
timestamp 1679581782
transform 1 0 19392 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_203
timestamp 1679581782
transform 1 0 20064 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_210
timestamp 1679581782
transform 1 0 20736 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_217
timestamp 1679581782
transform 1 0 21408 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_224
timestamp 1679581782
transform 1 0 22080 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_231
timestamp 1679581782
transform 1 0 22752 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_238
timestamp 1679581782
transform 1 0 23424 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_245
timestamp 1679581782
transform 1 0 24096 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_252
timestamp 1679581782
transform 1 0 24768 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_259
timestamp 1679581782
transform 1 0 25440 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_266
timestamp 1679581782
transform 1 0 26112 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_273
timestamp 1679581782
transform 1 0 26784 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_280
timestamp 1679581782
transform 1 0 27456 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_287
timestamp 1679581782
transform 1 0 28128 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_294
timestamp 1679581782
transform 1 0 28800 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_301
timestamp 1679581782
transform 1 0 29472 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_308
timestamp 1679581782
transform 1 0 30144 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_315
timestamp 1679581782
transform 1 0 30816 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_322
timestamp 1679581782
transform 1 0 31488 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_329
timestamp 1679581782
transform 1 0 32160 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_336
timestamp 1679581782
transform 1 0 32832 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_343
timestamp 1679581782
transform 1 0 33504 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_350
timestamp 1679581782
transform 1 0 34176 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_357
timestamp 1679581782
transform 1 0 34848 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_364
timestamp 1679581782
transform 1 0 35520 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_371
timestamp 1679581782
transform 1 0 36192 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_378
timestamp 1679581782
transform 1 0 36864 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_385
timestamp 1679581782
transform 1 0 37536 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_392
timestamp 1679581782
transform 1 0 38208 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_399
timestamp 1679581782
transform 1 0 38880 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_406
timestamp 1679581782
transform 1 0 39552 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_413
timestamp 1679581782
transform 1 0 40224 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_420
timestamp 1679581782
transform 1 0 40896 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_427
timestamp 1679581782
transform 1 0 41568 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_434
timestamp 1679581782
transform 1 0 42240 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_441
timestamp 1679581782
transform 1 0 42912 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_448
timestamp 1679581782
transform 1 0 43584 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_455
timestamp 1679581782
transform 1 0 44256 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_462
timestamp 1679581782
transform 1 0 44928 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_469
timestamp 1679581782
transform 1 0 45600 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_476
timestamp 1679581782
transform 1 0 46272 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_483
timestamp 1679581782
transform 1 0 46944 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_490
timestamp 1679581782
transform 1 0 47616 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_497
timestamp 1679581782
transform 1 0 48288 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_504
timestamp 1679581782
transform 1 0 48960 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_511
timestamp 1679581782
transform 1 0 49632 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_518
timestamp 1679581782
transform 1 0 50304 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_525
timestamp 1679581782
transform 1 0 50976 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_532
timestamp 1679581782
transform 1 0 51648 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_539
timestamp 1679581782
transform 1 0 52320 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_546
timestamp 1679581782
transform 1 0 52992 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_553
timestamp 1679581782
transform 1 0 53664 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_560
timestamp 1679581782
transform 1 0 54336 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_567
timestamp 1679581782
transform 1 0 55008 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_574
timestamp 1679581782
transform 1 0 55680 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_581
timestamp 1679581782
transform 1 0 56352 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_588
timestamp 1679581782
transform 1 0 57024 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_595
timestamp 1679581782
transform 1 0 57696 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_602
timestamp 1679581782
transform 1 0 58368 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_609
timestamp 1679581782
transform 1 0 59040 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_616
timestamp 1679581782
transform 1 0 59712 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_623
timestamp 1679581782
transform 1 0 60384 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_630
timestamp 1679581782
transform 1 0 61056 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_637
timestamp 1679581782
transform 1 0 61728 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_644
timestamp 1679581782
transform 1 0 62400 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_651
timestamp 1679581782
transform 1 0 63072 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_658
timestamp 1679581782
transform 1 0 63744 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_665
timestamp 1679581782
transform 1 0 64416 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_672
timestamp 1679581782
transform 1 0 65088 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_679
timestamp 1679581782
transform 1 0 65760 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_686
timestamp 1679581782
transform 1 0 66432 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_693
timestamp 1679581782
transform 1 0 67104 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_700
timestamp 1679581782
transform 1 0 67776 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_707
timestamp 1679581782
transform 1 0 68448 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_714
timestamp 1679581782
transform 1 0 69120 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_721
timestamp 1679581782
transform 1 0 69792 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_728
timestamp 1679581782
transform 1 0 70464 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_735
timestamp 1679581782
transform 1 0 71136 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_742
timestamp 1679581782
transform 1 0 71808 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_749
timestamp 1679581782
transform 1 0 72480 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_756
timestamp 1679581782
transform 1 0 73152 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_763
timestamp 1679581782
transform 1 0 73824 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_770
timestamp 1679581782
transform 1 0 74496 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_777
timestamp 1679581782
transform 1 0 75168 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_784
timestamp 1679581782
transform 1 0 75840 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_791
timestamp 1679581782
transform 1 0 76512 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_798
timestamp 1679581782
transform 1 0 77184 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_805
timestamp 1679581782
transform 1 0 77856 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_812
timestamp 1679581782
transform 1 0 78528 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_819
timestamp 1679581782
transform 1 0 79200 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_826
timestamp 1679581782
transform 1 0 79872 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_833
timestamp 1679581782
transform 1 0 80544 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_840
timestamp 1679581782
transform 1 0 81216 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_847
timestamp 1679581782
transform 1 0 81888 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_854
timestamp 1679581782
transform 1 0 82560 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_861
timestamp 1679581782
transform 1 0 83232 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_868
timestamp 1679581782
transform 1 0 83904 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_875
timestamp 1679581782
transform 1 0 84576 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_882
timestamp 1679581782
transform 1 0 85248 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_889
timestamp 1679581782
transform 1 0 85920 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_896
timestamp 1679581782
transform 1 0 86592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_903
timestamp 1679581782
transform 1 0 87264 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_910
timestamp 1679581782
transform 1 0 87936 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_917
timestamp 1679581782
transform 1 0 88608 0 1 756
box -48 -56 720 834
use sg13g2_fill_1  FILLER_0_924
timestamp 1677579658
transform 1 0 89280 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679581782
transform 1 0 576 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_7
timestamp 1679581782
transform 1 0 1248 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_14
timestamp 1679581782
transform 1 0 1920 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_21
timestamp 1679581782
transform 1 0 2592 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_28
timestamp 1679581782
transform 1 0 3264 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_35
timestamp 1679581782
transform 1 0 3936 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_42
timestamp 1679581782
transform 1 0 4608 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_49
timestamp 1679581782
transform 1 0 5280 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_56
timestamp 1679581782
transform 1 0 5952 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_63
timestamp 1679581782
transform 1 0 6624 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_70
timestamp 1679581782
transform 1 0 7296 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_77
timestamp 1679581782
transform 1 0 7968 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_84
timestamp 1679581782
transform 1 0 8640 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_91
timestamp 1679581782
transform 1 0 9312 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_98
timestamp 1679581782
transform 1 0 9984 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_105
timestamp 1679581782
transform 1 0 10656 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_112
timestamp 1679581782
transform 1 0 11328 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_119
timestamp 1679581782
transform 1 0 12000 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_126
timestamp 1679581782
transform 1 0 12672 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_133
timestamp 1679581782
transform 1 0 13344 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_140
timestamp 1679581782
transform 1 0 14016 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_147
timestamp 1679581782
transform 1 0 14688 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_154
timestamp 1679581782
transform 1 0 15360 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_161
timestamp 1679581782
transform 1 0 16032 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_168
timestamp 1679581782
transform 1 0 16704 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_175
timestamp 1679581782
transform 1 0 17376 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_182
timestamp 1679581782
transform 1 0 18048 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_189
timestamp 1679581782
transform 1 0 18720 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_196
timestamp 1679581782
transform 1 0 19392 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_203
timestamp 1679581782
transform 1 0 20064 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_210
timestamp 1679581782
transform 1 0 20736 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_217
timestamp 1679581782
transform 1 0 21408 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_224
timestamp 1679581782
transform 1 0 22080 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_231
timestamp 1679581782
transform 1 0 22752 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_238
timestamp 1679581782
transform 1 0 23424 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_245
timestamp 1679581782
transform 1 0 24096 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_252
timestamp 1679581782
transform 1 0 24768 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_259
timestamp 1679581782
transform 1 0 25440 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_266
timestamp 1679581782
transform 1 0 26112 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_273
timestamp 1679581782
transform 1 0 26784 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_280
timestamp 1679581782
transform 1 0 27456 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_287
timestamp 1679581782
transform 1 0 28128 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_294
timestamp 1679581782
transform 1 0 28800 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_301
timestamp 1679581782
transform 1 0 29472 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_308
timestamp 1679581782
transform 1 0 30144 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_315
timestamp 1679581782
transform 1 0 30816 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_322
timestamp 1679581782
transform 1 0 31488 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_329
timestamp 1679581782
transform 1 0 32160 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_336
timestamp 1679581782
transform 1 0 32832 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_343
timestamp 1679581782
transform 1 0 33504 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_350
timestamp 1679581782
transform 1 0 34176 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_357
timestamp 1679581782
transform 1 0 34848 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_364
timestamp 1679581782
transform 1 0 35520 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_371
timestamp 1679581782
transform 1 0 36192 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_378
timestamp 1679581782
transform 1 0 36864 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_385
timestamp 1679581782
transform 1 0 37536 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_392
timestamp 1679581782
transform 1 0 38208 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_399
timestamp 1679581782
transform 1 0 38880 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_406
timestamp 1679581782
transform 1 0 39552 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_413
timestamp 1679581782
transform 1 0 40224 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_420
timestamp 1679581782
transform 1 0 40896 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_427
timestamp 1679581782
transform 1 0 41568 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_434
timestamp 1679581782
transform 1 0 42240 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_441
timestamp 1679581782
transform 1 0 42912 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_448
timestamp 1679581782
transform 1 0 43584 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_455
timestamp 1679581782
transform 1 0 44256 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_462
timestamp 1679581782
transform 1 0 44928 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_469
timestamp 1679581782
transform 1 0 45600 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_476
timestamp 1679581782
transform 1 0 46272 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_483
timestamp 1679581782
transform 1 0 46944 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_490
timestamp 1679581782
transform 1 0 47616 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_497
timestamp 1679581782
transform 1 0 48288 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_504
timestamp 1679581782
transform 1 0 48960 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_511
timestamp 1679581782
transform 1 0 49632 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_518
timestamp 1679581782
transform 1 0 50304 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_525
timestamp 1679581782
transform 1 0 50976 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_532
timestamp 1679581782
transform 1 0 51648 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_539
timestamp 1679581782
transform 1 0 52320 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_546
timestamp 1679581782
transform 1 0 52992 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_553
timestamp 1679581782
transform 1 0 53664 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_560
timestamp 1679581782
transform 1 0 54336 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_567
timestamp 1679581782
transform 1 0 55008 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_574
timestamp 1679581782
transform 1 0 55680 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_581
timestamp 1679581782
transform 1 0 56352 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_588
timestamp 1679581782
transform 1 0 57024 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_595
timestamp 1679581782
transform 1 0 57696 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_602
timestamp 1679581782
transform 1 0 58368 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_609
timestamp 1679581782
transform 1 0 59040 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_616
timestamp 1679581782
transform 1 0 59712 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_623
timestamp 1679581782
transform 1 0 60384 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_630
timestamp 1679581782
transform 1 0 61056 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_637
timestamp 1679581782
transform 1 0 61728 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_644
timestamp 1679581782
transform 1 0 62400 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_651
timestamp 1679581782
transform 1 0 63072 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_658
timestamp 1679581782
transform 1 0 63744 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_665
timestamp 1679581782
transform 1 0 64416 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_672
timestamp 1679581782
transform 1 0 65088 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_679
timestamp 1679581782
transform 1 0 65760 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_686
timestamp 1679581782
transform 1 0 66432 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_693
timestamp 1679581782
transform 1 0 67104 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_700
timestamp 1679581782
transform 1 0 67776 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_707
timestamp 1679581782
transform 1 0 68448 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_714
timestamp 1679581782
transform 1 0 69120 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_721
timestamp 1679581782
transform 1 0 69792 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_728
timestamp 1679581782
transform 1 0 70464 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_735
timestamp 1679581782
transform 1 0 71136 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_742
timestamp 1679581782
transform 1 0 71808 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_749
timestamp 1679581782
transform 1 0 72480 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_756
timestamp 1679581782
transform 1 0 73152 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_763
timestamp 1679581782
transform 1 0 73824 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_770
timestamp 1679581782
transform 1 0 74496 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_777
timestamp 1679581782
transform 1 0 75168 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_784
timestamp 1679581782
transform 1 0 75840 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_791
timestamp 1679581782
transform 1 0 76512 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_798
timestamp 1679581782
transform 1 0 77184 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_805
timestamp 1679581782
transform 1 0 77856 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_812
timestamp 1679581782
transform 1 0 78528 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_819
timestamp 1679581782
transform 1 0 79200 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_826
timestamp 1679581782
transform 1 0 79872 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_833
timestamp 1679581782
transform 1 0 80544 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_840
timestamp 1679581782
transform 1 0 81216 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_847
timestamp 1679581782
transform 1 0 81888 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_854
timestamp 1679581782
transform 1 0 82560 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_861
timestamp 1679581782
transform 1 0 83232 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_868
timestamp 1679581782
transform 1 0 83904 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_875
timestamp 1679581782
transform 1 0 84576 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_882
timestamp 1679581782
transform 1 0 85248 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_889
timestamp 1679581782
transform 1 0 85920 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_896
timestamp 1679581782
transform 1 0 86592 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_903
timestamp 1679581782
transform 1 0 87264 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_910
timestamp 1679581782
transform 1 0 87936 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_917
timestamp 1679581782
transform 1 0 88608 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_1_924
timestamp 1677579658
transform 1 0 89280 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_4
timestamp 1679581782
transform 1 0 960 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_11
timestamp 1679581782
transform 1 0 1632 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_18
timestamp 1679581782
transform 1 0 2304 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_25
timestamp 1679581782
transform 1 0 2976 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_32
timestamp 1679581782
transform 1 0 3648 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_39
timestamp 1679581782
transform 1 0 4320 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_46
timestamp 1679581782
transform 1 0 4992 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_53
timestamp 1679581782
transform 1 0 5664 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_60
timestamp 1679581782
transform 1 0 6336 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_67
timestamp 1679581782
transform 1 0 7008 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_74
timestamp 1679581782
transform 1 0 7680 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_81
timestamp 1679581782
transform 1 0 8352 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_88
timestamp 1679581782
transform 1 0 9024 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_95
timestamp 1679581782
transform 1 0 9696 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_102
timestamp 1679581782
transform 1 0 10368 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_109
timestamp 1679581782
transform 1 0 11040 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_116
timestamp 1679581782
transform 1 0 11712 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_123
timestamp 1679581782
transform 1 0 12384 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_130
timestamp 1679581782
transform 1 0 13056 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_137
timestamp 1679581782
transform 1 0 13728 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_144
timestamp 1679581782
transform 1 0 14400 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_151
timestamp 1679581782
transform 1 0 15072 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_158
timestamp 1679581782
transform 1 0 15744 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_165
timestamp 1679581782
transform 1 0 16416 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_172
timestamp 1679581782
transform 1 0 17088 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_179
timestamp 1679581782
transform 1 0 17760 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_186
timestamp 1679581782
transform 1 0 18432 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_193
timestamp 1679581782
transform 1 0 19104 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_200
timestamp 1679581782
transform 1 0 19776 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_207
timestamp 1679581782
transform 1 0 20448 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_214
timestamp 1679581782
transform 1 0 21120 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_221
timestamp 1679581782
transform 1 0 21792 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_228
timestamp 1679581782
transform 1 0 22464 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_235
timestamp 1679581782
transform 1 0 23136 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_242
timestamp 1679581782
transform 1 0 23808 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_249
timestamp 1679581782
transform 1 0 24480 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_256
timestamp 1679581782
transform 1 0 25152 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_263
timestamp 1679581782
transform 1 0 25824 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_270
timestamp 1679581782
transform 1 0 26496 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_277
timestamp 1679581782
transform 1 0 27168 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_284
timestamp 1679581782
transform 1 0 27840 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_291
timestamp 1679581782
transform 1 0 28512 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_298
timestamp 1679581782
transform 1 0 29184 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_305
timestamp 1679581782
transform 1 0 29856 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_312
timestamp 1679581782
transform 1 0 30528 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_319
timestamp 1679581782
transform 1 0 31200 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_326
timestamp 1679581782
transform 1 0 31872 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_333
timestamp 1679581782
transform 1 0 32544 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_340
timestamp 1679581782
transform 1 0 33216 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_347
timestamp 1679581782
transform 1 0 33888 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_354
timestamp 1679581782
transform 1 0 34560 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_361
timestamp 1679581782
transform 1 0 35232 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_368
timestamp 1679581782
transform 1 0 35904 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_375
timestamp 1679581782
transform 1 0 36576 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_382
timestamp 1679581782
transform 1 0 37248 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_389
timestamp 1679581782
transform 1 0 37920 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_396
timestamp 1679581782
transform 1 0 38592 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_403
timestamp 1679581782
transform 1 0 39264 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_410
timestamp 1679581782
transform 1 0 39936 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_417
timestamp 1679581782
transform 1 0 40608 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_424
timestamp 1679581782
transform 1 0 41280 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_431
timestamp 1679581782
transform 1 0 41952 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_438
timestamp 1679581782
transform 1 0 42624 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_445
timestamp 1679581782
transform 1 0 43296 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_452
timestamp 1679581782
transform 1 0 43968 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_459
timestamp 1679581782
transform 1 0 44640 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_466
timestamp 1679581782
transform 1 0 45312 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_473
timestamp 1679581782
transform 1 0 45984 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_480
timestamp 1679581782
transform 1 0 46656 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_487
timestamp 1679581782
transform 1 0 47328 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_494
timestamp 1679581782
transform 1 0 48000 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_501
timestamp 1679581782
transform 1 0 48672 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_508
timestamp 1679581782
transform 1 0 49344 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_515
timestamp 1679581782
transform 1 0 50016 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_522
timestamp 1679581782
transform 1 0 50688 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_529
timestamp 1679581782
transform 1 0 51360 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_536
timestamp 1679581782
transform 1 0 52032 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_543
timestamp 1679581782
transform 1 0 52704 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_550
timestamp 1679581782
transform 1 0 53376 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_557
timestamp 1679581782
transform 1 0 54048 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_564
timestamp 1679581782
transform 1 0 54720 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_571
timestamp 1679581782
transform 1 0 55392 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_578
timestamp 1679581782
transform 1 0 56064 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_585
timestamp 1679581782
transform 1 0 56736 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_592
timestamp 1679581782
transform 1 0 57408 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_599
timestamp 1679581782
transform 1 0 58080 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_606
timestamp 1679581782
transform 1 0 58752 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_613
timestamp 1679581782
transform 1 0 59424 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_620
timestamp 1679581782
transform 1 0 60096 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_627
timestamp 1679581782
transform 1 0 60768 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_634
timestamp 1679581782
transform 1 0 61440 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_641
timestamp 1679581782
transform 1 0 62112 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_648
timestamp 1679581782
transform 1 0 62784 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_655
timestamp 1679581782
transform 1 0 63456 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_662
timestamp 1679581782
transform 1 0 64128 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_669
timestamp 1679581782
transform 1 0 64800 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_676
timestamp 1679581782
transform 1 0 65472 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_683
timestamp 1679581782
transform 1 0 66144 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_690
timestamp 1679581782
transform 1 0 66816 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_697
timestamp 1679581782
transform 1 0 67488 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_704
timestamp 1679581782
transform 1 0 68160 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_711
timestamp 1679581782
transform 1 0 68832 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_718
timestamp 1679581782
transform 1 0 69504 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_725
timestamp 1679581782
transform 1 0 70176 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_732
timestamp 1679581782
transform 1 0 70848 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_739
timestamp 1679581782
transform 1 0 71520 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_746
timestamp 1679581782
transform 1 0 72192 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_753
timestamp 1679581782
transform 1 0 72864 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_760
timestamp 1679581782
transform 1 0 73536 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_767
timestamp 1679581782
transform 1 0 74208 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_774
timestamp 1679581782
transform 1 0 74880 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_781
timestamp 1679581782
transform 1 0 75552 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_788
timestamp 1679581782
transform 1 0 76224 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_795
timestamp 1679581782
transform 1 0 76896 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_802
timestamp 1679581782
transform 1 0 77568 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_809
timestamp 1679581782
transform 1 0 78240 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_816
timestamp 1679581782
transform 1 0 78912 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_823
timestamp 1679581782
transform 1 0 79584 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_830
timestamp 1679581782
transform 1 0 80256 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_837
timestamp 1679581782
transform 1 0 80928 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_844
timestamp 1679581782
transform 1 0 81600 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_851
timestamp 1679581782
transform 1 0 82272 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_858
timestamp 1679581782
transform 1 0 82944 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_865
timestamp 1679581782
transform 1 0 83616 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_872
timestamp 1679581782
transform 1 0 84288 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_879
timestamp 1679581782
transform 1 0 84960 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_886
timestamp 1679581782
transform 1 0 85632 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_893
timestamp 1679581782
transform 1 0 86304 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_900
timestamp 1679581782
transform 1 0 86976 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_907
timestamp 1679581782
transform 1 0 87648 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_914
timestamp 1679581782
transform 1 0 88320 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_921
timestamp 1679577901
transform 1 0 88992 0 1 2268
box -48 -56 432 834
use sg13g2_decap_8  FILLER_3_4
timestamp 1679581782
transform 1 0 960 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_11
timestamp 1679581782
transform 1 0 1632 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_18
timestamp 1679581782
transform 1 0 2304 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_25
timestamp 1679581782
transform 1 0 2976 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_32
timestamp 1679581782
transform 1 0 3648 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_39
timestamp 1679581782
transform 1 0 4320 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_46
timestamp 1679581782
transform 1 0 4992 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_53
timestamp 1679581782
transform 1 0 5664 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_60
timestamp 1679581782
transform 1 0 6336 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_67
timestamp 1679581782
transform 1 0 7008 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_74
timestamp 1679581782
transform 1 0 7680 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_81
timestamp 1679581782
transform 1 0 8352 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_88
timestamp 1679581782
transform 1 0 9024 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_95
timestamp 1679581782
transform 1 0 9696 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_102
timestamp 1679581782
transform 1 0 10368 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_109
timestamp 1679581782
transform 1 0 11040 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_116
timestamp 1679581782
transform 1 0 11712 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_123
timestamp 1679581782
transform 1 0 12384 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_130
timestamp 1679581782
transform 1 0 13056 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_137
timestamp 1679581782
transform 1 0 13728 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_144
timestamp 1679581782
transform 1 0 14400 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_151
timestamp 1679581782
transform 1 0 15072 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_158
timestamp 1679581782
transform 1 0 15744 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_165
timestamp 1679581782
transform 1 0 16416 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_172
timestamp 1679581782
transform 1 0 17088 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_179
timestamp 1679581782
transform 1 0 17760 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_186
timestamp 1679581782
transform 1 0 18432 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_193
timestamp 1679581782
transform 1 0 19104 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_200
timestamp 1679581782
transform 1 0 19776 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_207
timestamp 1679581782
transform 1 0 20448 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_214
timestamp 1679581782
transform 1 0 21120 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_221
timestamp 1679581782
transform 1 0 21792 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_228
timestamp 1679581782
transform 1 0 22464 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_235
timestamp 1679581782
transform 1 0 23136 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_242
timestamp 1679581782
transform 1 0 23808 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_249
timestamp 1679581782
transform 1 0 24480 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_256
timestamp 1679581782
transform 1 0 25152 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_263
timestamp 1679581782
transform 1 0 25824 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_270
timestamp 1679581782
transform 1 0 26496 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_277
timestamp 1679581782
transform 1 0 27168 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_284
timestamp 1679581782
transform 1 0 27840 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_291
timestamp 1679581782
transform 1 0 28512 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_298
timestamp 1679581782
transform 1 0 29184 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_305
timestamp 1679581782
transform 1 0 29856 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_312
timestamp 1679581782
transform 1 0 30528 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_319
timestamp 1679581782
transform 1 0 31200 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_326
timestamp 1679581782
transform 1 0 31872 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_333
timestamp 1679581782
transform 1 0 32544 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_340
timestamp 1679581782
transform 1 0 33216 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_347
timestamp 1679581782
transform 1 0 33888 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_354
timestamp 1679581782
transform 1 0 34560 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_361
timestamp 1679581782
transform 1 0 35232 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_368
timestamp 1679581782
transform 1 0 35904 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_375
timestamp 1679581782
transform 1 0 36576 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_382
timestamp 1679581782
transform 1 0 37248 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_389
timestamp 1679581782
transform 1 0 37920 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_396
timestamp 1679581782
transform 1 0 38592 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_403
timestamp 1679581782
transform 1 0 39264 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_410
timestamp 1679581782
transform 1 0 39936 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_417
timestamp 1679581782
transform 1 0 40608 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_424
timestamp 1679581782
transform 1 0 41280 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_431
timestamp 1679581782
transform 1 0 41952 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_438
timestamp 1679581782
transform 1 0 42624 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_445
timestamp 1679581782
transform 1 0 43296 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_452
timestamp 1679581782
transform 1 0 43968 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_459
timestamp 1679581782
transform 1 0 44640 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_466
timestamp 1679581782
transform 1 0 45312 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_473
timestamp 1679581782
transform 1 0 45984 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_480
timestamp 1679581782
transform 1 0 46656 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_487
timestamp 1679581782
transform 1 0 47328 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_494
timestamp 1679581782
transform 1 0 48000 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_501
timestamp 1679581782
transform 1 0 48672 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_508
timestamp 1679581782
transform 1 0 49344 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_515
timestamp 1679581782
transform 1 0 50016 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_522
timestamp 1679581782
transform 1 0 50688 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_529
timestamp 1679581782
transform 1 0 51360 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_536
timestamp 1679581782
transform 1 0 52032 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_543
timestamp 1679581782
transform 1 0 52704 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_550
timestamp 1679581782
transform 1 0 53376 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_557
timestamp 1679581782
transform 1 0 54048 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_564
timestamp 1679581782
transform 1 0 54720 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_571
timestamp 1679581782
transform 1 0 55392 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_578
timestamp 1679581782
transform 1 0 56064 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_585
timestamp 1679581782
transform 1 0 56736 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_592
timestamp 1679581782
transform 1 0 57408 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_599
timestamp 1679581782
transform 1 0 58080 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_606
timestamp 1679581782
transform 1 0 58752 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_613
timestamp 1679581782
transform 1 0 59424 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_620
timestamp 1679581782
transform 1 0 60096 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_627
timestamp 1679581782
transform 1 0 60768 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_634
timestamp 1679581782
transform 1 0 61440 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_641
timestamp 1679581782
transform 1 0 62112 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_648
timestamp 1679581782
transform 1 0 62784 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_655
timestamp 1679581782
transform 1 0 63456 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_662
timestamp 1679581782
transform 1 0 64128 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_669
timestamp 1679581782
transform 1 0 64800 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_676
timestamp 1679581782
transform 1 0 65472 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_683
timestamp 1679581782
transform 1 0 66144 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_690
timestamp 1679581782
transform 1 0 66816 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_697
timestamp 1679581782
transform 1 0 67488 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_704
timestamp 1679581782
transform 1 0 68160 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_711
timestamp 1679581782
transform 1 0 68832 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_718
timestamp 1679581782
transform 1 0 69504 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_725
timestamp 1679581782
transform 1 0 70176 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_732
timestamp 1679581782
transform 1 0 70848 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_739
timestamp 1679581782
transform 1 0 71520 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_746
timestamp 1679581782
transform 1 0 72192 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_753
timestamp 1679581782
transform 1 0 72864 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_760
timestamp 1679581782
transform 1 0 73536 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_767
timestamp 1679581782
transform 1 0 74208 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_774
timestamp 1679581782
transform 1 0 74880 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_781
timestamp 1679581782
transform 1 0 75552 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_788
timestamp 1679581782
transform 1 0 76224 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_795
timestamp 1679581782
transform 1 0 76896 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_802
timestamp 1679581782
transform 1 0 77568 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_809
timestamp 1679581782
transform 1 0 78240 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_816
timestamp 1679581782
transform 1 0 78912 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_823
timestamp 1679581782
transform 1 0 79584 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_830
timestamp 1679581782
transform 1 0 80256 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_837
timestamp 1679581782
transform 1 0 80928 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_844
timestamp 1679581782
transform 1 0 81600 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_851
timestamp 1679581782
transform 1 0 82272 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_858
timestamp 1679581782
transform 1 0 82944 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_865
timestamp 1679581782
transform 1 0 83616 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_872
timestamp 1679581782
transform 1 0 84288 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_879
timestamp 1679581782
transform 1 0 84960 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_886
timestamp 1679581782
transform 1 0 85632 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_893
timestamp 1679581782
transform 1 0 86304 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_900
timestamp 1679581782
transform 1 0 86976 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_907
timestamp 1679581782
transform 1 0 87648 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_914
timestamp 1679581782
transform 1 0 88320 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_921
timestamp 1679577901
transform 1 0 88992 0 -1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_4_4
timestamp 1679581782
transform 1 0 960 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_11
timestamp 1679581782
transform 1 0 1632 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_18
timestamp 1679581782
transform 1 0 2304 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_25
timestamp 1679581782
transform 1 0 2976 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_32
timestamp 1679581782
transform 1 0 3648 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_39
timestamp 1679581782
transform 1 0 4320 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_46
timestamp 1679581782
transform 1 0 4992 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_53
timestamp 1679581782
transform 1 0 5664 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_60
timestamp 1679581782
transform 1 0 6336 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_67
timestamp 1679581782
transform 1 0 7008 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_74
timestamp 1679581782
transform 1 0 7680 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_81
timestamp 1679581782
transform 1 0 8352 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_88
timestamp 1679581782
transform 1 0 9024 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_95
timestamp 1679581782
transform 1 0 9696 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_102
timestamp 1679581782
transform 1 0 10368 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_109
timestamp 1679581782
transform 1 0 11040 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_116
timestamp 1679581782
transform 1 0 11712 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_123
timestamp 1679581782
transform 1 0 12384 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_130
timestamp 1679581782
transform 1 0 13056 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_137
timestamp 1679581782
transform 1 0 13728 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_144
timestamp 1679581782
transform 1 0 14400 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_151
timestamp 1679581782
transform 1 0 15072 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_158
timestamp 1679581782
transform 1 0 15744 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_165
timestamp 1679581782
transform 1 0 16416 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_172
timestamp 1679581782
transform 1 0 17088 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_179
timestamp 1679581782
transform 1 0 17760 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_186
timestamp 1679581782
transform 1 0 18432 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_193
timestamp 1679581782
transform 1 0 19104 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_200
timestamp 1679581782
transform 1 0 19776 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_207
timestamp 1679581782
transform 1 0 20448 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_214
timestamp 1679581782
transform 1 0 21120 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_221
timestamp 1679581782
transform 1 0 21792 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_228
timestamp 1679581782
transform 1 0 22464 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_235
timestamp 1679581782
transform 1 0 23136 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_242
timestamp 1679581782
transform 1 0 23808 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_249
timestamp 1679581782
transform 1 0 24480 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_256
timestamp 1679581782
transform 1 0 25152 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_263
timestamp 1679581782
transform 1 0 25824 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_270
timestamp 1679581782
transform 1 0 26496 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_277
timestamp 1679581782
transform 1 0 27168 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_284
timestamp 1679581782
transform 1 0 27840 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_291
timestamp 1679581782
transform 1 0 28512 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_298
timestamp 1679581782
transform 1 0 29184 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_305
timestamp 1679581782
transform 1 0 29856 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_312
timestamp 1679581782
transform 1 0 30528 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_319
timestamp 1679581782
transform 1 0 31200 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_326
timestamp 1679581782
transform 1 0 31872 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_333
timestamp 1679581782
transform 1 0 32544 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_340
timestamp 1679581782
transform 1 0 33216 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_347
timestamp 1679581782
transform 1 0 33888 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_354
timestamp 1679581782
transform 1 0 34560 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_361
timestamp 1679581782
transform 1 0 35232 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_368
timestamp 1679581782
transform 1 0 35904 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_375
timestamp 1679581782
transform 1 0 36576 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_382
timestamp 1679581782
transform 1 0 37248 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_389
timestamp 1679581782
transform 1 0 37920 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_396
timestamp 1679581782
transform 1 0 38592 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_403
timestamp 1679581782
transform 1 0 39264 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_410
timestamp 1679581782
transform 1 0 39936 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_417
timestamp 1679581782
transform 1 0 40608 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_424
timestamp 1679581782
transform 1 0 41280 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_431
timestamp 1679581782
transform 1 0 41952 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_438
timestamp 1679581782
transform 1 0 42624 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_445
timestamp 1679581782
transform 1 0 43296 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_452
timestamp 1679581782
transform 1 0 43968 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_459
timestamp 1679581782
transform 1 0 44640 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_466
timestamp 1679581782
transform 1 0 45312 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_473
timestamp 1679581782
transform 1 0 45984 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_480
timestamp 1679581782
transform 1 0 46656 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_487
timestamp 1679581782
transform 1 0 47328 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_494
timestamp 1679581782
transform 1 0 48000 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_501
timestamp 1679581782
transform 1 0 48672 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_508
timestamp 1679581782
transform 1 0 49344 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_515
timestamp 1679581782
transform 1 0 50016 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_522
timestamp 1679581782
transform 1 0 50688 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_529
timestamp 1679581782
transform 1 0 51360 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_536
timestamp 1679581782
transform 1 0 52032 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_543
timestamp 1679581782
transform 1 0 52704 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_550
timestamp 1679581782
transform 1 0 53376 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_557
timestamp 1679581782
transform 1 0 54048 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_564
timestamp 1679581782
transform 1 0 54720 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_571
timestamp 1679581782
transform 1 0 55392 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_578
timestamp 1679581782
transform 1 0 56064 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_585
timestamp 1679581782
transform 1 0 56736 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_592
timestamp 1679581782
transform 1 0 57408 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_599
timestamp 1679581782
transform 1 0 58080 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_606
timestamp 1679581782
transform 1 0 58752 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_613
timestamp 1679581782
transform 1 0 59424 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_620
timestamp 1679581782
transform 1 0 60096 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_627
timestamp 1679581782
transform 1 0 60768 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_634
timestamp 1679581782
transform 1 0 61440 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_641
timestamp 1679581782
transform 1 0 62112 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_648
timestamp 1679581782
transform 1 0 62784 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_655
timestamp 1679581782
transform 1 0 63456 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_662
timestamp 1679581782
transform 1 0 64128 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_669
timestamp 1679581782
transform 1 0 64800 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_676
timestamp 1679581782
transform 1 0 65472 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_683
timestamp 1679581782
transform 1 0 66144 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_690
timestamp 1679581782
transform 1 0 66816 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_697
timestamp 1679581782
transform 1 0 67488 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_704
timestamp 1679581782
transform 1 0 68160 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_711
timestamp 1679581782
transform 1 0 68832 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_718
timestamp 1679581782
transform 1 0 69504 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_725
timestamp 1679581782
transform 1 0 70176 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_732
timestamp 1679581782
transform 1 0 70848 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_739
timestamp 1679581782
transform 1 0 71520 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_746
timestamp 1679581782
transform 1 0 72192 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_753
timestamp 1679581782
transform 1 0 72864 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_760
timestamp 1679581782
transform 1 0 73536 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_767
timestamp 1679581782
transform 1 0 74208 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_774
timestamp 1679581782
transform 1 0 74880 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_781
timestamp 1679581782
transform 1 0 75552 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_788
timestamp 1679581782
transform 1 0 76224 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_795
timestamp 1679581782
transform 1 0 76896 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_802
timestamp 1679581782
transform 1 0 77568 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_809
timestamp 1679581782
transform 1 0 78240 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_816
timestamp 1679581782
transform 1 0 78912 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_823
timestamp 1679581782
transform 1 0 79584 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_830
timestamp 1679581782
transform 1 0 80256 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_837
timestamp 1679581782
transform 1 0 80928 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_844
timestamp 1679581782
transform 1 0 81600 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_851
timestamp 1679581782
transform 1 0 82272 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_858
timestamp 1679581782
transform 1 0 82944 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_865
timestamp 1679581782
transform 1 0 83616 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_872
timestamp 1679581782
transform 1 0 84288 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_879
timestamp 1679581782
transform 1 0 84960 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_886
timestamp 1679581782
transform 1 0 85632 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_893
timestamp 1679581782
transform 1 0 86304 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_900
timestamp 1679581782
transform 1 0 86976 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_907
timestamp 1679581782
transform 1 0 87648 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_914
timestamp 1679581782
transform 1 0 88320 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_921
timestamp 1679577901
transform 1 0 88992 0 1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_5_4
timestamp 1679581782
transform 1 0 960 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_11
timestamp 1679581782
transform 1 0 1632 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_18
timestamp 1679581782
transform 1 0 2304 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_25
timestamp 1679581782
transform 1 0 2976 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_32
timestamp 1679581782
transform 1 0 3648 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_39
timestamp 1679581782
transform 1 0 4320 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_46
timestamp 1679581782
transform 1 0 4992 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_53
timestamp 1679581782
transform 1 0 5664 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_60
timestamp 1679581782
transform 1 0 6336 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_67
timestamp 1679581782
transform 1 0 7008 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_74
timestamp 1679581782
transform 1 0 7680 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_81
timestamp 1679581782
transform 1 0 8352 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_88
timestamp 1679581782
transform 1 0 9024 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_95
timestamp 1679581782
transform 1 0 9696 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_102
timestamp 1679581782
transform 1 0 10368 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_109
timestamp 1679581782
transform 1 0 11040 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_116
timestamp 1679581782
transform 1 0 11712 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_123
timestamp 1679581782
transform 1 0 12384 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_130
timestamp 1679581782
transform 1 0 13056 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_137
timestamp 1679581782
transform 1 0 13728 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_144
timestamp 1679581782
transform 1 0 14400 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_151
timestamp 1679581782
transform 1 0 15072 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_158
timestamp 1679581782
transform 1 0 15744 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_165
timestamp 1679581782
transform 1 0 16416 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_172
timestamp 1679581782
transform 1 0 17088 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_179
timestamp 1679581782
transform 1 0 17760 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_186
timestamp 1679581782
transform 1 0 18432 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_193
timestamp 1679581782
transform 1 0 19104 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_200
timestamp 1679581782
transform 1 0 19776 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_207
timestamp 1679581782
transform 1 0 20448 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_214
timestamp 1679581782
transform 1 0 21120 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_221
timestamp 1679581782
transform 1 0 21792 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_228
timestamp 1679581782
transform 1 0 22464 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_235
timestamp 1679581782
transform 1 0 23136 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_242
timestamp 1679581782
transform 1 0 23808 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_249
timestamp 1679581782
transform 1 0 24480 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_256
timestamp 1679581782
transform 1 0 25152 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_263
timestamp 1679581782
transform 1 0 25824 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_270
timestamp 1679581782
transform 1 0 26496 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_277
timestamp 1679581782
transform 1 0 27168 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_284
timestamp 1679581782
transform 1 0 27840 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_291
timestamp 1679581782
transform 1 0 28512 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_298
timestamp 1679581782
transform 1 0 29184 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_305
timestamp 1679581782
transform 1 0 29856 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_312
timestamp 1679581782
transform 1 0 30528 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_319
timestamp 1679581782
transform 1 0 31200 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_326
timestamp 1679581782
transform 1 0 31872 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_333
timestamp 1679581782
transform 1 0 32544 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_340
timestamp 1679581782
transform 1 0 33216 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_347
timestamp 1679581782
transform 1 0 33888 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_354
timestamp 1679581782
transform 1 0 34560 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_361
timestamp 1679581782
transform 1 0 35232 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_368
timestamp 1679581782
transform 1 0 35904 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_375
timestamp 1679581782
transform 1 0 36576 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_382
timestamp 1679581782
transform 1 0 37248 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_389
timestamp 1679581782
transform 1 0 37920 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_396
timestamp 1679581782
transform 1 0 38592 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_403
timestamp 1679581782
transform 1 0 39264 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_410
timestamp 1679581782
transform 1 0 39936 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_417
timestamp 1679581782
transform 1 0 40608 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_424
timestamp 1679581782
transform 1 0 41280 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_431
timestamp 1679581782
transform 1 0 41952 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_438
timestamp 1679581782
transform 1 0 42624 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_445
timestamp 1679581782
transform 1 0 43296 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_452
timestamp 1679581782
transform 1 0 43968 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_459
timestamp 1679581782
transform 1 0 44640 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_466
timestamp 1679581782
transform 1 0 45312 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_473
timestamp 1679581782
transform 1 0 45984 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_480
timestamp 1679581782
transform 1 0 46656 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_487
timestamp 1679581782
transform 1 0 47328 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_494
timestamp 1679581782
transform 1 0 48000 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_501
timestamp 1679581782
transform 1 0 48672 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_508
timestamp 1679581782
transform 1 0 49344 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_515
timestamp 1679581782
transform 1 0 50016 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_522
timestamp 1679581782
transform 1 0 50688 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_529
timestamp 1679581782
transform 1 0 51360 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_536
timestamp 1679581782
transform 1 0 52032 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_543
timestamp 1679581782
transform 1 0 52704 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_550
timestamp 1679581782
transform 1 0 53376 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_557
timestamp 1679581782
transform 1 0 54048 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_564
timestamp 1679581782
transform 1 0 54720 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_571
timestamp 1679581782
transform 1 0 55392 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_578
timestamp 1679581782
transform 1 0 56064 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_585
timestamp 1679581782
transform 1 0 56736 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_592
timestamp 1679581782
transform 1 0 57408 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_599
timestamp 1679581782
transform 1 0 58080 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_606
timestamp 1679581782
transform 1 0 58752 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_613
timestamp 1679581782
transform 1 0 59424 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_620
timestamp 1679581782
transform 1 0 60096 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_627
timestamp 1679581782
transform 1 0 60768 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_634
timestamp 1679581782
transform 1 0 61440 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_641
timestamp 1679581782
transform 1 0 62112 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_648
timestamp 1679581782
transform 1 0 62784 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_655
timestamp 1679581782
transform 1 0 63456 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_662
timestamp 1679581782
transform 1 0 64128 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_669
timestamp 1679581782
transform 1 0 64800 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_676
timestamp 1679581782
transform 1 0 65472 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_683
timestamp 1679581782
transform 1 0 66144 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_690
timestamp 1679581782
transform 1 0 66816 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_697
timestamp 1679581782
transform 1 0 67488 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_704
timestamp 1679581782
transform 1 0 68160 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_711
timestamp 1679581782
transform 1 0 68832 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_718
timestamp 1679581782
transform 1 0 69504 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_725
timestamp 1679581782
transform 1 0 70176 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_732
timestamp 1679581782
transform 1 0 70848 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_739
timestamp 1679581782
transform 1 0 71520 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_746
timestamp 1679581782
transform 1 0 72192 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_753
timestamp 1679581782
transform 1 0 72864 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_760
timestamp 1679581782
transform 1 0 73536 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_767
timestamp 1679581782
transform 1 0 74208 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_774
timestamp 1679581782
transform 1 0 74880 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_781
timestamp 1679581782
transform 1 0 75552 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_788
timestamp 1679581782
transform 1 0 76224 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_795
timestamp 1679581782
transform 1 0 76896 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_802
timestamp 1679581782
transform 1 0 77568 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_809
timestamp 1679581782
transform 1 0 78240 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_816
timestamp 1679581782
transform 1 0 78912 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_823
timestamp 1679581782
transform 1 0 79584 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_830
timestamp 1679581782
transform 1 0 80256 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_837
timestamp 1679581782
transform 1 0 80928 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_844
timestamp 1679581782
transform 1 0 81600 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_851
timestamp 1679581782
transform 1 0 82272 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_858
timestamp 1679581782
transform 1 0 82944 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_865
timestamp 1679581782
transform 1 0 83616 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_872
timestamp 1679581782
transform 1 0 84288 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_879
timestamp 1679581782
transform 1 0 84960 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_886
timestamp 1679581782
transform 1 0 85632 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_893
timestamp 1679581782
transform 1 0 86304 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_900
timestamp 1679581782
transform 1 0 86976 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_907
timestamp 1679581782
transform 1 0 87648 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_914
timestamp 1679581782
transform 1 0 88320 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_921
timestamp 1679577901
transform 1 0 88992 0 -1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_6_4
timestamp 1679581782
transform 1 0 960 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_11
timestamp 1679581782
transform 1 0 1632 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_18
timestamp 1679581782
transform 1 0 2304 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_25
timestamp 1679581782
transform 1 0 2976 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_32
timestamp 1679581782
transform 1 0 3648 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_39
timestamp 1679581782
transform 1 0 4320 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_46
timestamp 1679581782
transform 1 0 4992 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_53
timestamp 1679581782
transform 1 0 5664 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_60
timestamp 1679581782
transform 1 0 6336 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_67
timestamp 1679581782
transform 1 0 7008 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_74
timestamp 1679581782
transform 1 0 7680 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_81
timestamp 1679581782
transform 1 0 8352 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_88
timestamp 1679581782
transform 1 0 9024 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_95
timestamp 1679581782
transform 1 0 9696 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_102
timestamp 1679581782
transform 1 0 10368 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_109
timestamp 1679581782
transform 1 0 11040 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_116
timestamp 1679581782
transform 1 0 11712 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_123
timestamp 1679581782
transform 1 0 12384 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_130
timestamp 1679581782
transform 1 0 13056 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_137
timestamp 1679581782
transform 1 0 13728 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_144
timestamp 1679581782
transform 1 0 14400 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_151
timestamp 1679581782
transform 1 0 15072 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_158
timestamp 1679581782
transform 1 0 15744 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_165
timestamp 1679581782
transform 1 0 16416 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_172
timestamp 1679581782
transform 1 0 17088 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_179
timestamp 1679581782
transform 1 0 17760 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_186
timestamp 1679581782
transform 1 0 18432 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_193
timestamp 1679581782
transform 1 0 19104 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_200
timestamp 1679581782
transform 1 0 19776 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_207
timestamp 1679581782
transform 1 0 20448 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_214
timestamp 1679581782
transform 1 0 21120 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_221
timestamp 1679581782
transform 1 0 21792 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_228
timestamp 1679581782
transform 1 0 22464 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_235
timestamp 1679581782
transform 1 0 23136 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_242
timestamp 1679581782
transform 1 0 23808 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_249
timestamp 1679581782
transform 1 0 24480 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_256
timestamp 1679581782
transform 1 0 25152 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_263
timestamp 1679581782
transform 1 0 25824 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_270
timestamp 1679581782
transform 1 0 26496 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_277
timestamp 1679581782
transform 1 0 27168 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_284
timestamp 1679581782
transform 1 0 27840 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_291
timestamp 1679581782
transform 1 0 28512 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_298
timestamp 1679581782
transform 1 0 29184 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_305
timestamp 1679581782
transform 1 0 29856 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_312
timestamp 1679581782
transform 1 0 30528 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_319
timestamp 1679581782
transform 1 0 31200 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_326
timestamp 1679581782
transform 1 0 31872 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_333
timestamp 1679581782
transform 1 0 32544 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_340
timestamp 1679581782
transform 1 0 33216 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_347
timestamp 1679581782
transform 1 0 33888 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_354
timestamp 1679581782
transform 1 0 34560 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_361
timestamp 1679581782
transform 1 0 35232 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_368
timestamp 1679581782
transform 1 0 35904 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_375
timestamp 1679581782
transform 1 0 36576 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_382
timestamp 1679581782
transform 1 0 37248 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_389
timestamp 1679581782
transform 1 0 37920 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_396
timestamp 1679581782
transform 1 0 38592 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_403
timestamp 1679581782
transform 1 0 39264 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_410
timestamp 1679581782
transform 1 0 39936 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_417
timestamp 1679581782
transform 1 0 40608 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_424
timestamp 1679581782
transform 1 0 41280 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_431
timestamp 1679581782
transform 1 0 41952 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_438
timestamp 1679581782
transform 1 0 42624 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_445
timestamp 1679581782
transform 1 0 43296 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_452
timestamp 1679581782
transform 1 0 43968 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_459
timestamp 1679581782
transform 1 0 44640 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_466
timestamp 1679581782
transform 1 0 45312 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_473
timestamp 1679581782
transform 1 0 45984 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_480
timestamp 1679581782
transform 1 0 46656 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_487
timestamp 1679581782
transform 1 0 47328 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_494
timestamp 1679581782
transform 1 0 48000 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_501
timestamp 1679581782
transform 1 0 48672 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_508
timestamp 1679581782
transform 1 0 49344 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_515
timestamp 1679581782
transform 1 0 50016 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_522
timestamp 1679581782
transform 1 0 50688 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_529
timestamp 1679581782
transform 1 0 51360 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_536
timestamp 1679581782
transform 1 0 52032 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_543
timestamp 1679581782
transform 1 0 52704 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_550
timestamp 1679581782
transform 1 0 53376 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_557
timestamp 1679581782
transform 1 0 54048 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_564
timestamp 1679581782
transform 1 0 54720 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_571
timestamp 1679581782
transform 1 0 55392 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_578
timestamp 1679581782
transform 1 0 56064 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_585
timestamp 1679581782
transform 1 0 56736 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_592
timestamp 1679581782
transform 1 0 57408 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_599
timestamp 1679581782
transform 1 0 58080 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_606
timestamp 1679581782
transform 1 0 58752 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_613
timestamp 1679581782
transform 1 0 59424 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_620
timestamp 1679581782
transform 1 0 60096 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_627
timestamp 1679581782
transform 1 0 60768 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_634
timestamp 1679581782
transform 1 0 61440 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_641
timestamp 1679581782
transform 1 0 62112 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_648
timestamp 1679581782
transform 1 0 62784 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_655
timestamp 1679581782
transform 1 0 63456 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_662
timestamp 1679581782
transform 1 0 64128 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_669
timestamp 1679581782
transform 1 0 64800 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_676
timestamp 1679581782
transform 1 0 65472 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_683
timestamp 1679581782
transform 1 0 66144 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_690
timestamp 1679581782
transform 1 0 66816 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_697
timestamp 1679581782
transform 1 0 67488 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_704
timestamp 1679581782
transform 1 0 68160 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_711
timestamp 1679581782
transform 1 0 68832 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_718
timestamp 1679581782
transform 1 0 69504 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_725
timestamp 1679581782
transform 1 0 70176 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_732
timestamp 1679581782
transform 1 0 70848 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_739
timestamp 1679581782
transform 1 0 71520 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_746
timestamp 1679581782
transform 1 0 72192 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_753
timestamp 1679581782
transform 1 0 72864 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_760
timestamp 1679581782
transform 1 0 73536 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_767
timestamp 1679581782
transform 1 0 74208 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_774
timestamp 1679581782
transform 1 0 74880 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_781
timestamp 1679581782
transform 1 0 75552 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_788
timestamp 1679581782
transform 1 0 76224 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_795
timestamp 1679581782
transform 1 0 76896 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_802
timestamp 1679581782
transform 1 0 77568 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_809
timestamp 1679581782
transform 1 0 78240 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_816
timestamp 1679581782
transform 1 0 78912 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_823
timestamp 1679581782
transform 1 0 79584 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_830
timestamp 1679581782
transform 1 0 80256 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_837
timestamp 1679581782
transform 1 0 80928 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_844
timestamp 1679581782
transform 1 0 81600 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_851
timestamp 1679581782
transform 1 0 82272 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_858
timestamp 1679581782
transform 1 0 82944 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_865
timestamp 1679581782
transform 1 0 83616 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_872
timestamp 1679581782
transform 1 0 84288 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_879
timestamp 1679581782
transform 1 0 84960 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_886
timestamp 1679581782
transform 1 0 85632 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_893
timestamp 1679581782
transform 1 0 86304 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_900
timestamp 1679581782
transform 1 0 86976 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_907
timestamp 1679581782
transform 1 0 87648 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_914
timestamp 1679581782
transform 1 0 88320 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_921
timestamp 1679577901
transform 1 0 88992 0 1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_7_0
timestamp 1679581782
transform 1 0 576 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_7
timestamp 1679581782
transform 1 0 1248 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_14
timestamp 1679581782
transform 1 0 1920 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_21
timestamp 1679581782
transform 1 0 2592 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_28
timestamp 1679581782
transform 1 0 3264 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_35
timestamp 1679581782
transform 1 0 3936 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_42
timestamp 1679581782
transform 1 0 4608 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_49
timestamp 1679581782
transform 1 0 5280 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_56
timestamp 1679581782
transform 1 0 5952 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_63
timestamp 1679581782
transform 1 0 6624 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_70
timestamp 1679581782
transform 1 0 7296 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_77
timestamp 1679581782
transform 1 0 7968 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_84
timestamp 1679581782
transform 1 0 8640 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_91
timestamp 1679581782
transform 1 0 9312 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_98
timestamp 1679581782
transform 1 0 9984 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_105
timestamp 1679581782
transform 1 0 10656 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_112
timestamp 1679581782
transform 1 0 11328 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_119
timestamp 1679581782
transform 1 0 12000 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_126
timestamp 1679581782
transform 1 0 12672 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_133
timestamp 1679581782
transform 1 0 13344 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_140
timestamp 1679581782
transform 1 0 14016 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_147
timestamp 1679581782
transform 1 0 14688 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_154
timestamp 1679581782
transform 1 0 15360 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_161
timestamp 1679581782
transform 1 0 16032 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_168
timestamp 1679581782
transform 1 0 16704 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_175
timestamp 1679581782
transform 1 0 17376 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_182
timestamp 1679581782
transform 1 0 18048 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_189
timestamp 1679581782
transform 1 0 18720 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_196
timestamp 1679581782
transform 1 0 19392 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_203
timestamp 1679581782
transform 1 0 20064 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_210
timestamp 1679581782
transform 1 0 20736 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_217
timestamp 1679581782
transform 1 0 21408 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_224
timestamp 1679581782
transform 1 0 22080 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_231
timestamp 1679581782
transform 1 0 22752 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_238
timestamp 1679581782
transform 1 0 23424 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_245
timestamp 1679581782
transform 1 0 24096 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_252
timestamp 1679581782
transform 1 0 24768 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_259
timestamp 1679581782
transform 1 0 25440 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_266
timestamp 1679581782
transform 1 0 26112 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_273
timestamp 1679581782
transform 1 0 26784 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_280
timestamp 1679581782
transform 1 0 27456 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_287
timestamp 1679581782
transform 1 0 28128 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_294
timestamp 1679581782
transform 1 0 28800 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_301
timestamp 1679581782
transform 1 0 29472 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_308
timestamp 1679581782
transform 1 0 30144 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_315
timestamp 1679581782
transform 1 0 30816 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_322
timestamp 1679581782
transform 1 0 31488 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_329
timestamp 1679581782
transform 1 0 32160 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_336
timestamp 1679581782
transform 1 0 32832 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_343
timestamp 1679581782
transform 1 0 33504 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_350
timestamp 1679581782
transform 1 0 34176 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_357
timestamp 1679581782
transform 1 0 34848 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_364
timestamp 1679581782
transform 1 0 35520 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_371
timestamp 1679581782
transform 1 0 36192 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_378
timestamp 1679581782
transform 1 0 36864 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_385
timestamp 1679581782
transform 1 0 37536 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_392
timestamp 1679581782
transform 1 0 38208 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_399
timestamp 1679581782
transform 1 0 38880 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_406
timestamp 1679581782
transform 1 0 39552 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_413
timestamp 1679581782
transform 1 0 40224 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_420
timestamp 1679581782
transform 1 0 40896 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_427
timestamp 1679581782
transform 1 0 41568 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_434
timestamp 1679581782
transform 1 0 42240 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_441
timestamp 1679581782
transform 1 0 42912 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_448
timestamp 1679581782
transform 1 0 43584 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_455
timestamp 1679581782
transform 1 0 44256 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_462
timestamp 1679581782
transform 1 0 44928 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_469
timestamp 1679581782
transform 1 0 45600 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_476
timestamp 1679581782
transform 1 0 46272 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_483
timestamp 1679581782
transform 1 0 46944 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_490
timestamp 1679581782
transform 1 0 47616 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_497
timestamp 1679581782
transform 1 0 48288 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_504
timestamp 1679581782
transform 1 0 48960 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_511
timestamp 1679581782
transform 1 0 49632 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_518
timestamp 1679581782
transform 1 0 50304 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_525
timestamp 1679581782
transform 1 0 50976 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_532
timestamp 1679581782
transform 1 0 51648 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_539
timestamp 1679581782
transform 1 0 52320 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_546
timestamp 1679581782
transform 1 0 52992 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_553
timestamp 1679581782
transform 1 0 53664 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_560
timestamp 1679581782
transform 1 0 54336 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_567
timestamp 1679581782
transform 1 0 55008 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_574
timestamp 1679581782
transform 1 0 55680 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_581
timestamp 1679581782
transform 1 0 56352 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_588
timestamp 1679581782
transform 1 0 57024 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_595
timestamp 1679581782
transform 1 0 57696 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_602
timestamp 1679581782
transform 1 0 58368 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_609
timestamp 1679581782
transform 1 0 59040 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_616
timestamp 1679581782
transform 1 0 59712 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_623
timestamp 1679581782
transform 1 0 60384 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_630
timestamp 1679581782
transform 1 0 61056 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_637
timestamp 1679581782
transform 1 0 61728 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_644
timestamp 1679581782
transform 1 0 62400 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_651
timestamp 1679581782
transform 1 0 63072 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_658
timestamp 1679581782
transform 1 0 63744 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_665
timestamp 1679581782
transform 1 0 64416 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_672
timestamp 1679581782
transform 1 0 65088 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_679
timestamp 1679581782
transform 1 0 65760 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_686
timestamp 1679581782
transform 1 0 66432 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_693
timestamp 1679581782
transform 1 0 67104 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_700
timestamp 1679581782
transform 1 0 67776 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_707
timestamp 1679581782
transform 1 0 68448 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_714
timestamp 1679581782
transform 1 0 69120 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_721
timestamp 1679581782
transform 1 0 69792 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_728
timestamp 1679581782
transform 1 0 70464 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_735
timestamp 1679581782
transform 1 0 71136 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_742
timestamp 1679581782
transform 1 0 71808 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_749
timestamp 1679581782
transform 1 0 72480 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_756
timestamp 1679581782
transform 1 0 73152 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_763
timestamp 1679581782
transform 1 0 73824 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_770
timestamp 1679581782
transform 1 0 74496 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_777
timestamp 1679581782
transform 1 0 75168 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_784
timestamp 1679581782
transform 1 0 75840 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_791
timestamp 1679581782
transform 1 0 76512 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_798
timestamp 1679581782
transform 1 0 77184 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_805
timestamp 1679581782
transform 1 0 77856 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_812
timestamp 1679581782
transform 1 0 78528 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_819
timestamp 1679581782
transform 1 0 79200 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_826
timestamp 1679581782
transform 1 0 79872 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_833
timestamp 1679581782
transform 1 0 80544 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_840
timestamp 1679581782
transform 1 0 81216 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_847
timestamp 1679581782
transform 1 0 81888 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_854
timestamp 1679581782
transform 1 0 82560 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_861
timestamp 1679581782
transform 1 0 83232 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_868
timestamp 1679581782
transform 1 0 83904 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_875
timestamp 1679581782
transform 1 0 84576 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_882
timestamp 1679581782
transform 1 0 85248 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_889
timestamp 1679581782
transform 1 0 85920 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_896
timestamp 1679581782
transform 1 0 86592 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_903
timestamp 1679581782
transform 1 0 87264 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_910
timestamp 1679581782
transform 1 0 87936 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_917
timestamp 1679581782
transform 1 0 88608 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_924
timestamp 1677579658
transform 1 0 89280 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_4
timestamp 1679581782
transform 1 0 960 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_11
timestamp 1679581782
transform 1 0 1632 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_18
timestamp 1679581782
transform 1 0 2304 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_25
timestamp 1679581782
transform 1 0 2976 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_32
timestamp 1679581782
transform 1 0 3648 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_39
timestamp 1679581782
transform 1 0 4320 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_46
timestamp 1679581782
transform 1 0 4992 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_53
timestamp 1679581782
transform 1 0 5664 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_60
timestamp 1679581782
transform 1 0 6336 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_67
timestamp 1679581782
transform 1 0 7008 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_74
timestamp 1679581782
transform 1 0 7680 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_81
timestamp 1679581782
transform 1 0 8352 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_88
timestamp 1679581782
transform 1 0 9024 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_95
timestamp 1679581782
transform 1 0 9696 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_102
timestamp 1679581782
transform 1 0 10368 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_109
timestamp 1679581782
transform 1 0 11040 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_116
timestamp 1679581782
transform 1 0 11712 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_123
timestamp 1679581782
transform 1 0 12384 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_130
timestamp 1679581782
transform 1 0 13056 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_137
timestamp 1679581782
transform 1 0 13728 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_144
timestamp 1679581782
transform 1 0 14400 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_151
timestamp 1679581782
transform 1 0 15072 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_158
timestamp 1679581782
transform 1 0 15744 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_165
timestamp 1679581782
transform 1 0 16416 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_172
timestamp 1679581782
transform 1 0 17088 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_179
timestamp 1679581782
transform 1 0 17760 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_186
timestamp 1679581782
transform 1 0 18432 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_193
timestamp 1679581782
transform 1 0 19104 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_200
timestamp 1679581782
transform 1 0 19776 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_207
timestamp 1679581782
transform 1 0 20448 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_214
timestamp 1679581782
transform 1 0 21120 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_221
timestamp 1679581782
transform 1 0 21792 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_228
timestamp 1679581782
transform 1 0 22464 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_235
timestamp 1679581782
transform 1 0 23136 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_242
timestamp 1679581782
transform 1 0 23808 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_249
timestamp 1679581782
transform 1 0 24480 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_256
timestamp 1679581782
transform 1 0 25152 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_263
timestamp 1679581782
transform 1 0 25824 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_270
timestamp 1679581782
transform 1 0 26496 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_277
timestamp 1679581782
transform 1 0 27168 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_284
timestamp 1679581782
transform 1 0 27840 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_291
timestamp 1679581782
transform 1 0 28512 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_298
timestamp 1679581782
transform 1 0 29184 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_305
timestamp 1679581782
transform 1 0 29856 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_312
timestamp 1679581782
transform 1 0 30528 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_319
timestamp 1679581782
transform 1 0 31200 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_326
timestamp 1679581782
transform 1 0 31872 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_333
timestamp 1679581782
transform 1 0 32544 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_340
timestamp 1679581782
transform 1 0 33216 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_347
timestamp 1679581782
transform 1 0 33888 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_354
timestamp 1679581782
transform 1 0 34560 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_361
timestamp 1679581782
transform 1 0 35232 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_368
timestamp 1679581782
transform 1 0 35904 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_375
timestamp 1679581782
transform 1 0 36576 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_382
timestamp 1679581782
transform 1 0 37248 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_389
timestamp 1679581782
transform 1 0 37920 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_396
timestamp 1679581782
transform 1 0 38592 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_403
timestamp 1679581782
transform 1 0 39264 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_410
timestamp 1679581782
transform 1 0 39936 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_417
timestamp 1679581782
transform 1 0 40608 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_424
timestamp 1679581782
transform 1 0 41280 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_431
timestamp 1679581782
transform 1 0 41952 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_438
timestamp 1679581782
transform 1 0 42624 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_445
timestamp 1679581782
transform 1 0 43296 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_452
timestamp 1679581782
transform 1 0 43968 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_459
timestamp 1679581782
transform 1 0 44640 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_466
timestamp 1679581782
transform 1 0 45312 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_473
timestamp 1679581782
transform 1 0 45984 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_480
timestamp 1679581782
transform 1 0 46656 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_487
timestamp 1679581782
transform 1 0 47328 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_494
timestamp 1679581782
transform 1 0 48000 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_501
timestamp 1679581782
transform 1 0 48672 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_508
timestamp 1679581782
transform 1 0 49344 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_515
timestamp 1679581782
transform 1 0 50016 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_522
timestamp 1679581782
transform 1 0 50688 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_529
timestamp 1679581782
transform 1 0 51360 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_536
timestamp 1679581782
transform 1 0 52032 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_543
timestamp 1679581782
transform 1 0 52704 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_550
timestamp 1679581782
transform 1 0 53376 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_557
timestamp 1679581782
transform 1 0 54048 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_564
timestamp 1679581782
transform 1 0 54720 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_571
timestamp 1679581782
transform 1 0 55392 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_578
timestamp 1679581782
transform 1 0 56064 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_585
timestamp 1679581782
transform 1 0 56736 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_592
timestamp 1679581782
transform 1 0 57408 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_599
timestamp 1679581782
transform 1 0 58080 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_606
timestamp 1679581782
transform 1 0 58752 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_613
timestamp 1679581782
transform 1 0 59424 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_620
timestamp 1679581782
transform 1 0 60096 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_627
timestamp 1679581782
transform 1 0 60768 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_634
timestamp 1679581782
transform 1 0 61440 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_641
timestamp 1679581782
transform 1 0 62112 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_648
timestamp 1679581782
transform 1 0 62784 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_655
timestamp 1679581782
transform 1 0 63456 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_662
timestamp 1679581782
transform 1 0 64128 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_669
timestamp 1679581782
transform 1 0 64800 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_676
timestamp 1679581782
transform 1 0 65472 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_683
timestamp 1679581782
transform 1 0 66144 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_690
timestamp 1679581782
transform 1 0 66816 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_697
timestamp 1679581782
transform 1 0 67488 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_704
timestamp 1679581782
transform 1 0 68160 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_711
timestamp 1679581782
transform 1 0 68832 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_718
timestamp 1679581782
transform 1 0 69504 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_725
timestamp 1679581782
transform 1 0 70176 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_732
timestamp 1679581782
transform 1 0 70848 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_739
timestamp 1679581782
transform 1 0 71520 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_746
timestamp 1679581782
transform 1 0 72192 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_753
timestamp 1679581782
transform 1 0 72864 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_760
timestamp 1679581782
transform 1 0 73536 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_767
timestamp 1679581782
transform 1 0 74208 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_774
timestamp 1679581782
transform 1 0 74880 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_781
timestamp 1679581782
transform 1 0 75552 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_788
timestamp 1679581782
transform 1 0 76224 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_795
timestamp 1679581782
transform 1 0 76896 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_802
timestamp 1679581782
transform 1 0 77568 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_809
timestamp 1679581782
transform 1 0 78240 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_816
timestamp 1679581782
transform 1 0 78912 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_823
timestamp 1679581782
transform 1 0 79584 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_830
timestamp 1679581782
transform 1 0 80256 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_837
timestamp 1679581782
transform 1 0 80928 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_844
timestamp 1679581782
transform 1 0 81600 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_851
timestamp 1679581782
transform 1 0 82272 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_858
timestamp 1679581782
transform 1 0 82944 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_865
timestamp 1679581782
transform 1 0 83616 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_872
timestamp 1679581782
transform 1 0 84288 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_879
timestamp 1679581782
transform 1 0 84960 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_886
timestamp 1679581782
transform 1 0 85632 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_893
timestamp 1679581782
transform 1 0 86304 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_900
timestamp 1679581782
transform 1 0 86976 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_907
timestamp 1679581782
transform 1 0 87648 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_914
timestamp 1679581782
transform 1 0 88320 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_921
timestamp 1679577901
transform 1 0 88992 0 1 6804
box -48 -56 432 834
use sg13g2_decap_8  FILLER_9_4
timestamp 1679581782
transform 1 0 960 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_11
timestamp 1679581782
transform 1 0 1632 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_18
timestamp 1679581782
transform 1 0 2304 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_25
timestamp 1679581782
transform 1 0 2976 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_32
timestamp 1679581782
transform 1 0 3648 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_39
timestamp 1679581782
transform 1 0 4320 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_46
timestamp 1679581782
transform 1 0 4992 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_53
timestamp 1679581782
transform 1 0 5664 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_60
timestamp 1679581782
transform 1 0 6336 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_67
timestamp 1679581782
transform 1 0 7008 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_74
timestamp 1679581782
transform 1 0 7680 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_81
timestamp 1679581782
transform 1 0 8352 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_88
timestamp 1679581782
transform 1 0 9024 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_95
timestamp 1679581782
transform 1 0 9696 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_102
timestamp 1679581782
transform 1 0 10368 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_109
timestamp 1679581782
transform 1 0 11040 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_116
timestamp 1679581782
transform 1 0 11712 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_123
timestamp 1679581782
transform 1 0 12384 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_130
timestamp 1679581782
transform 1 0 13056 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_137
timestamp 1679581782
transform 1 0 13728 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_144
timestamp 1679581782
transform 1 0 14400 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_151
timestamp 1679581782
transform 1 0 15072 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_158
timestamp 1679581782
transform 1 0 15744 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_165
timestamp 1679581782
transform 1 0 16416 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_172
timestamp 1679581782
transform 1 0 17088 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_179
timestamp 1679581782
transform 1 0 17760 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_186
timestamp 1679581782
transform 1 0 18432 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_193
timestamp 1679581782
transform 1 0 19104 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_200
timestamp 1679581782
transform 1 0 19776 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_207
timestamp 1679581782
transform 1 0 20448 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_214
timestamp 1679581782
transform 1 0 21120 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_221
timestamp 1679581782
transform 1 0 21792 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_228
timestamp 1679581782
transform 1 0 22464 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_235
timestamp 1679581782
transform 1 0 23136 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_242
timestamp 1679581782
transform 1 0 23808 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_249
timestamp 1679581782
transform 1 0 24480 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_256
timestamp 1679581782
transform 1 0 25152 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_263
timestamp 1679581782
transform 1 0 25824 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_270
timestamp 1679581782
transform 1 0 26496 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_277
timestamp 1679581782
transform 1 0 27168 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_284
timestamp 1679581782
transform 1 0 27840 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_291
timestamp 1679581782
transform 1 0 28512 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_298
timestamp 1679581782
transform 1 0 29184 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_305
timestamp 1679581782
transform 1 0 29856 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_312
timestamp 1679581782
transform 1 0 30528 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_319
timestamp 1679581782
transform 1 0 31200 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_326
timestamp 1679581782
transform 1 0 31872 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_333
timestamp 1679581782
transform 1 0 32544 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_340
timestamp 1679581782
transform 1 0 33216 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_347
timestamp 1679581782
transform 1 0 33888 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_354
timestamp 1679581782
transform 1 0 34560 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_361
timestamp 1679581782
transform 1 0 35232 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_368
timestamp 1679581782
transform 1 0 35904 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_375
timestamp 1679581782
transform 1 0 36576 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_382
timestamp 1679581782
transform 1 0 37248 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_389
timestamp 1679581782
transform 1 0 37920 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_396
timestamp 1679581782
transform 1 0 38592 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_403
timestamp 1679581782
transform 1 0 39264 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_410
timestamp 1679581782
transform 1 0 39936 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_417
timestamp 1679581782
transform 1 0 40608 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_424
timestamp 1679581782
transform 1 0 41280 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_431
timestamp 1679581782
transform 1 0 41952 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_438
timestamp 1679581782
transform 1 0 42624 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_445
timestamp 1679581782
transform 1 0 43296 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_452
timestamp 1679581782
transform 1 0 43968 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_459
timestamp 1679581782
transform 1 0 44640 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_466
timestamp 1679581782
transform 1 0 45312 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_473
timestamp 1679581782
transform 1 0 45984 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_480
timestamp 1679581782
transform 1 0 46656 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_487
timestamp 1679581782
transform 1 0 47328 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_494
timestamp 1679581782
transform 1 0 48000 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_501
timestamp 1679581782
transform 1 0 48672 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_508
timestamp 1679581782
transform 1 0 49344 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_515
timestamp 1679581782
transform 1 0 50016 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_522
timestamp 1679581782
transform 1 0 50688 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_529
timestamp 1679581782
transform 1 0 51360 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_536
timestamp 1679581782
transform 1 0 52032 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_543
timestamp 1679581782
transform 1 0 52704 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_550
timestamp 1679581782
transform 1 0 53376 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_557
timestamp 1679581782
transform 1 0 54048 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_564
timestamp 1679581782
transform 1 0 54720 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_571
timestamp 1679581782
transform 1 0 55392 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_578
timestamp 1679581782
transform 1 0 56064 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_585
timestamp 1679581782
transform 1 0 56736 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_592
timestamp 1679581782
transform 1 0 57408 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_599
timestamp 1679581782
transform 1 0 58080 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_606
timestamp 1679581782
transform 1 0 58752 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_613
timestamp 1679581782
transform 1 0 59424 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_620
timestamp 1679581782
transform 1 0 60096 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_627
timestamp 1679581782
transform 1 0 60768 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_634
timestamp 1679581782
transform 1 0 61440 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_641
timestamp 1679581782
transform 1 0 62112 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_648
timestamp 1679581782
transform 1 0 62784 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_655
timestamp 1679581782
transform 1 0 63456 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_662
timestamp 1679581782
transform 1 0 64128 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_669
timestamp 1679581782
transform 1 0 64800 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_676
timestamp 1679581782
transform 1 0 65472 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_683
timestamp 1679581782
transform 1 0 66144 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_690
timestamp 1679581782
transform 1 0 66816 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_697
timestamp 1679581782
transform 1 0 67488 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_704
timestamp 1679581782
transform 1 0 68160 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_711
timestamp 1679581782
transform 1 0 68832 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_718
timestamp 1679581782
transform 1 0 69504 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_725
timestamp 1679581782
transform 1 0 70176 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_732
timestamp 1679581782
transform 1 0 70848 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_739
timestamp 1679581782
transform 1 0 71520 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_746
timestamp 1679581782
transform 1 0 72192 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_753
timestamp 1679581782
transform 1 0 72864 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_760
timestamp 1679581782
transform 1 0 73536 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_767
timestamp 1679581782
transform 1 0 74208 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_774
timestamp 1679581782
transform 1 0 74880 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_781
timestamp 1679581782
transform 1 0 75552 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_788
timestamp 1679581782
transform 1 0 76224 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_795
timestamp 1679581782
transform 1 0 76896 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_802
timestamp 1679581782
transform 1 0 77568 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_809
timestamp 1679581782
transform 1 0 78240 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_816
timestamp 1679581782
transform 1 0 78912 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_823
timestamp 1679581782
transform 1 0 79584 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_830
timestamp 1679581782
transform 1 0 80256 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_837
timestamp 1679581782
transform 1 0 80928 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_844
timestamp 1679581782
transform 1 0 81600 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_851
timestamp 1679581782
transform 1 0 82272 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_858
timestamp 1679581782
transform 1 0 82944 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_865
timestamp 1679581782
transform 1 0 83616 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_872
timestamp 1679581782
transform 1 0 84288 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_879
timestamp 1679581782
transform 1 0 84960 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_886
timestamp 1679581782
transform 1 0 85632 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_893
timestamp 1679581782
transform 1 0 86304 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_900
timestamp 1679581782
transform 1 0 86976 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_907
timestamp 1679581782
transform 1 0 87648 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_914
timestamp 1679581782
transform 1 0 88320 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_921
timestamp 1679577901
transform 1 0 88992 0 -1 8316
box -48 -56 432 834
use sg13g2_decap_8  FILLER_10_4
timestamp 1679581782
transform 1 0 960 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_11
timestamp 1679581782
transform 1 0 1632 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_18
timestamp 1679581782
transform 1 0 2304 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_25
timestamp 1679581782
transform 1 0 2976 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_32
timestamp 1679581782
transform 1 0 3648 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_39
timestamp 1679581782
transform 1 0 4320 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_46
timestamp 1679581782
transform 1 0 4992 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_53
timestamp 1679581782
transform 1 0 5664 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_60
timestamp 1679581782
transform 1 0 6336 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_67
timestamp 1679581782
transform 1 0 7008 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_74
timestamp 1679581782
transform 1 0 7680 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_81
timestamp 1679581782
transform 1 0 8352 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_88
timestamp 1679581782
transform 1 0 9024 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_95
timestamp 1679581782
transform 1 0 9696 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_102
timestamp 1679581782
transform 1 0 10368 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_109
timestamp 1679581782
transform 1 0 11040 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_116
timestamp 1679581782
transform 1 0 11712 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_123
timestamp 1679581782
transform 1 0 12384 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_130
timestamp 1679581782
transform 1 0 13056 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_137
timestamp 1679581782
transform 1 0 13728 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_144
timestamp 1679581782
transform 1 0 14400 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_151
timestamp 1679581782
transform 1 0 15072 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_158
timestamp 1679581782
transform 1 0 15744 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_165
timestamp 1679581782
transform 1 0 16416 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_172
timestamp 1679581782
transform 1 0 17088 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_179
timestamp 1679581782
transform 1 0 17760 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_186
timestamp 1679581782
transform 1 0 18432 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_193
timestamp 1679581782
transform 1 0 19104 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_200
timestamp 1679581782
transform 1 0 19776 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_207
timestamp 1679581782
transform 1 0 20448 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_214
timestamp 1679581782
transform 1 0 21120 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_221
timestamp 1679581782
transform 1 0 21792 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_228
timestamp 1679581782
transform 1 0 22464 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_235
timestamp 1679581782
transform 1 0 23136 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_242
timestamp 1679581782
transform 1 0 23808 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_249
timestamp 1679581782
transform 1 0 24480 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_256
timestamp 1679581782
transform 1 0 25152 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_263
timestamp 1679581782
transform 1 0 25824 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_270
timestamp 1679581782
transform 1 0 26496 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_277
timestamp 1679581782
transform 1 0 27168 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_284
timestamp 1679581782
transform 1 0 27840 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_291
timestamp 1679581782
transform 1 0 28512 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_298
timestamp 1679581782
transform 1 0 29184 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_305
timestamp 1679581782
transform 1 0 29856 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_312
timestamp 1679581782
transform 1 0 30528 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_319
timestamp 1679581782
transform 1 0 31200 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_326
timestamp 1679581782
transform 1 0 31872 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_333
timestamp 1679581782
transform 1 0 32544 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_340
timestamp 1679581782
transform 1 0 33216 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_347
timestamp 1679581782
transform 1 0 33888 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_354
timestamp 1679581782
transform 1 0 34560 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_361
timestamp 1679581782
transform 1 0 35232 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_368
timestamp 1679581782
transform 1 0 35904 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_375
timestamp 1679581782
transform 1 0 36576 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_382
timestamp 1679581782
transform 1 0 37248 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_389
timestamp 1679581782
transform 1 0 37920 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_396
timestamp 1679581782
transform 1 0 38592 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_403
timestamp 1679581782
transform 1 0 39264 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_410
timestamp 1679581782
transform 1 0 39936 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_417
timestamp 1679581782
transform 1 0 40608 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_424
timestamp 1679581782
transform 1 0 41280 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_431
timestamp 1679581782
transform 1 0 41952 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_438
timestamp 1679581782
transform 1 0 42624 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_445
timestamp 1679581782
transform 1 0 43296 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_452
timestamp 1679581782
transform 1 0 43968 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_459
timestamp 1679581782
transform 1 0 44640 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_466
timestamp 1679581782
transform 1 0 45312 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_473
timestamp 1679581782
transform 1 0 45984 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_480
timestamp 1679581782
transform 1 0 46656 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_487
timestamp 1679581782
transform 1 0 47328 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_494
timestamp 1679581782
transform 1 0 48000 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_501
timestamp 1679581782
transform 1 0 48672 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_508
timestamp 1679581782
transform 1 0 49344 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_515
timestamp 1679581782
transform 1 0 50016 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_522
timestamp 1679581782
transform 1 0 50688 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_529
timestamp 1679581782
transform 1 0 51360 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_536
timestamp 1679581782
transform 1 0 52032 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_543
timestamp 1679581782
transform 1 0 52704 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_550
timestamp 1679581782
transform 1 0 53376 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_557
timestamp 1679581782
transform 1 0 54048 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_564
timestamp 1679581782
transform 1 0 54720 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_571
timestamp 1679581782
transform 1 0 55392 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_578
timestamp 1679581782
transform 1 0 56064 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_585
timestamp 1679581782
transform 1 0 56736 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_592
timestamp 1679581782
transform 1 0 57408 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_599
timestamp 1679581782
transform 1 0 58080 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_606
timestamp 1679581782
transform 1 0 58752 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_613
timestamp 1679581782
transform 1 0 59424 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_620
timestamp 1679581782
transform 1 0 60096 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_627
timestamp 1679581782
transform 1 0 60768 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_634
timestamp 1679581782
transform 1 0 61440 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_641
timestamp 1679581782
transform 1 0 62112 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_648
timestamp 1679581782
transform 1 0 62784 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_655
timestamp 1679581782
transform 1 0 63456 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_662
timestamp 1679581782
transform 1 0 64128 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_669
timestamp 1679581782
transform 1 0 64800 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_676
timestamp 1679581782
transform 1 0 65472 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_683
timestamp 1679581782
transform 1 0 66144 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_690
timestamp 1679581782
transform 1 0 66816 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_697
timestamp 1679581782
transform 1 0 67488 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_704
timestamp 1679581782
transform 1 0 68160 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_711
timestamp 1679581782
transform 1 0 68832 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_718
timestamp 1679581782
transform 1 0 69504 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_725
timestamp 1679581782
transform 1 0 70176 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_732
timestamp 1679581782
transform 1 0 70848 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_739
timestamp 1679581782
transform 1 0 71520 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_746
timestamp 1679581782
transform 1 0 72192 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_753
timestamp 1679581782
transform 1 0 72864 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_760
timestamp 1679581782
transform 1 0 73536 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_767
timestamp 1679581782
transform 1 0 74208 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_774
timestamp 1679581782
transform 1 0 74880 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_781
timestamp 1679581782
transform 1 0 75552 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_788
timestamp 1679581782
transform 1 0 76224 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_795
timestamp 1679581782
transform 1 0 76896 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_802
timestamp 1679581782
transform 1 0 77568 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_809
timestamp 1679581782
transform 1 0 78240 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_816
timestamp 1679581782
transform 1 0 78912 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_823
timestamp 1679581782
transform 1 0 79584 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_830
timestamp 1679581782
transform 1 0 80256 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_837
timestamp 1679581782
transform 1 0 80928 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_844
timestamp 1679581782
transform 1 0 81600 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_851
timestamp 1679581782
transform 1 0 82272 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_858
timestamp 1679581782
transform 1 0 82944 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_865
timestamp 1679581782
transform 1 0 83616 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_872
timestamp 1679581782
transform 1 0 84288 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_879
timestamp 1679581782
transform 1 0 84960 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_886
timestamp 1679581782
transform 1 0 85632 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_893
timestamp 1679581782
transform 1 0 86304 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_900
timestamp 1679581782
transform 1 0 86976 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_907
timestamp 1679581782
transform 1 0 87648 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_914
timestamp 1679581782
transform 1 0 88320 0 1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_921
timestamp 1679577901
transform 1 0 88992 0 1 8316
box -48 -56 432 834
use sg13g2_decap_8  FILLER_11_4
timestamp 1679581782
transform 1 0 960 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_11
timestamp 1679581782
transform 1 0 1632 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_18
timestamp 1679581782
transform 1 0 2304 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_25
timestamp 1679581782
transform 1 0 2976 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_32
timestamp 1679581782
transform 1 0 3648 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_39
timestamp 1679581782
transform 1 0 4320 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_46
timestamp 1679581782
transform 1 0 4992 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_53
timestamp 1679581782
transform 1 0 5664 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_60
timestamp 1679581782
transform 1 0 6336 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_67
timestamp 1679581782
transform 1 0 7008 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_74
timestamp 1679581782
transform 1 0 7680 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_81
timestamp 1679581782
transform 1 0 8352 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_88
timestamp 1679581782
transform 1 0 9024 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_95
timestamp 1679581782
transform 1 0 9696 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_102
timestamp 1679581782
transform 1 0 10368 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_109
timestamp 1679581782
transform 1 0 11040 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_116
timestamp 1679581782
transform 1 0 11712 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_123
timestamp 1679581782
transform 1 0 12384 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_130
timestamp 1679581782
transform 1 0 13056 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_137
timestamp 1679581782
transform 1 0 13728 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_144
timestamp 1679581782
transform 1 0 14400 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_151
timestamp 1679581782
transform 1 0 15072 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_158
timestamp 1679581782
transform 1 0 15744 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_165
timestamp 1679581782
transform 1 0 16416 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_172
timestamp 1679581782
transform 1 0 17088 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_179
timestamp 1679581782
transform 1 0 17760 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_186
timestamp 1679581782
transform 1 0 18432 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_193
timestamp 1679581782
transform 1 0 19104 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_200
timestamp 1679581782
transform 1 0 19776 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_207
timestamp 1679581782
transform 1 0 20448 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_214
timestamp 1679581782
transform 1 0 21120 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_221
timestamp 1679581782
transform 1 0 21792 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_228
timestamp 1679581782
transform 1 0 22464 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_235
timestamp 1679581782
transform 1 0 23136 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_242
timestamp 1679581782
transform 1 0 23808 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_249
timestamp 1679581782
transform 1 0 24480 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_256
timestamp 1679581782
transform 1 0 25152 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_263
timestamp 1679581782
transform 1 0 25824 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_270
timestamp 1679581782
transform 1 0 26496 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_277
timestamp 1679581782
transform 1 0 27168 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_284
timestamp 1679581782
transform 1 0 27840 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_291
timestamp 1679581782
transform 1 0 28512 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_298
timestamp 1679581782
transform 1 0 29184 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_305
timestamp 1679581782
transform 1 0 29856 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_312
timestamp 1679581782
transform 1 0 30528 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_319
timestamp 1679581782
transform 1 0 31200 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_326
timestamp 1679581782
transform 1 0 31872 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_333
timestamp 1679581782
transform 1 0 32544 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_340
timestamp 1679581782
transform 1 0 33216 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_347
timestamp 1679581782
transform 1 0 33888 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_354
timestamp 1679581782
transform 1 0 34560 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_361
timestamp 1679581782
transform 1 0 35232 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_368
timestamp 1679581782
transform 1 0 35904 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_375
timestamp 1679581782
transform 1 0 36576 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_382
timestamp 1679581782
transform 1 0 37248 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_389
timestamp 1679581782
transform 1 0 37920 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_396
timestamp 1679581782
transform 1 0 38592 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_403
timestamp 1679581782
transform 1 0 39264 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_410
timestamp 1679581782
transform 1 0 39936 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_417
timestamp 1679581782
transform 1 0 40608 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_424
timestamp 1679581782
transform 1 0 41280 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_431
timestamp 1679581782
transform 1 0 41952 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_438
timestamp 1679581782
transform 1 0 42624 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_445
timestamp 1679581782
transform 1 0 43296 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_452
timestamp 1679581782
transform 1 0 43968 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_459
timestamp 1679581782
transform 1 0 44640 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_466
timestamp 1679581782
transform 1 0 45312 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_473
timestamp 1679581782
transform 1 0 45984 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_480
timestamp 1679581782
transform 1 0 46656 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_487
timestamp 1679581782
transform 1 0 47328 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_494
timestamp 1679581782
transform 1 0 48000 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_501
timestamp 1679581782
transform 1 0 48672 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_508
timestamp 1679581782
transform 1 0 49344 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_515
timestamp 1679581782
transform 1 0 50016 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_522
timestamp 1679581782
transform 1 0 50688 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_529
timestamp 1679581782
transform 1 0 51360 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_536
timestamp 1679581782
transform 1 0 52032 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_543
timestamp 1679581782
transform 1 0 52704 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_550
timestamp 1679581782
transform 1 0 53376 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_557
timestamp 1679581782
transform 1 0 54048 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_564
timestamp 1679581782
transform 1 0 54720 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_571
timestamp 1679581782
transform 1 0 55392 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_578
timestamp 1679581782
transform 1 0 56064 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_585
timestamp 1679581782
transform 1 0 56736 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_592
timestamp 1679581782
transform 1 0 57408 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_599
timestamp 1679581782
transform 1 0 58080 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_606
timestamp 1679581782
transform 1 0 58752 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_613
timestamp 1679581782
transform 1 0 59424 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_620
timestamp 1679581782
transform 1 0 60096 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_627
timestamp 1679581782
transform 1 0 60768 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_634
timestamp 1679581782
transform 1 0 61440 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_641
timestamp 1679581782
transform 1 0 62112 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_648
timestamp 1679581782
transform 1 0 62784 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_655
timestamp 1679581782
transform 1 0 63456 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_662
timestamp 1679581782
transform 1 0 64128 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_669
timestamp 1679581782
transform 1 0 64800 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_676
timestamp 1679581782
transform 1 0 65472 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_683
timestamp 1679581782
transform 1 0 66144 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_690
timestamp 1679581782
transform 1 0 66816 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_697
timestamp 1679581782
transform 1 0 67488 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_704
timestamp 1679581782
transform 1 0 68160 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_711
timestamp 1679581782
transform 1 0 68832 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_718
timestamp 1679581782
transform 1 0 69504 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_725
timestamp 1679581782
transform 1 0 70176 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_732
timestamp 1679581782
transform 1 0 70848 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_739
timestamp 1679581782
transform 1 0 71520 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_746
timestamp 1679581782
transform 1 0 72192 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_753
timestamp 1679581782
transform 1 0 72864 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_760
timestamp 1679581782
transform 1 0 73536 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_767
timestamp 1679581782
transform 1 0 74208 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_774
timestamp 1679581782
transform 1 0 74880 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_781
timestamp 1679581782
transform 1 0 75552 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_788
timestamp 1679581782
transform 1 0 76224 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_795
timestamp 1679581782
transform 1 0 76896 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_802
timestamp 1679581782
transform 1 0 77568 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_809
timestamp 1679581782
transform 1 0 78240 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_816
timestamp 1679581782
transform 1 0 78912 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_823
timestamp 1679581782
transform 1 0 79584 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_830
timestamp 1679581782
transform 1 0 80256 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_837
timestamp 1679581782
transform 1 0 80928 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_844
timestamp 1679581782
transform 1 0 81600 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_851
timestamp 1679581782
transform 1 0 82272 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_858
timestamp 1679581782
transform 1 0 82944 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_865
timestamp 1679581782
transform 1 0 83616 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_872
timestamp 1679581782
transform 1 0 84288 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_879
timestamp 1679581782
transform 1 0 84960 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_886
timestamp 1679581782
transform 1 0 85632 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_893
timestamp 1679581782
transform 1 0 86304 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_900
timestamp 1679581782
transform 1 0 86976 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_907
timestamp 1679581782
transform 1 0 87648 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_914
timestamp 1679581782
transform 1 0 88320 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_921
timestamp 1679577901
transform 1 0 88992 0 -1 9828
box -48 -56 432 834
use sg13g2_decap_8  FILLER_12_4
timestamp 1679581782
transform 1 0 960 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_11
timestamp 1679581782
transform 1 0 1632 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_18
timestamp 1679581782
transform 1 0 2304 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_25
timestamp 1679581782
transform 1 0 2976 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_32
timestamp 1679581782
transform 1 0 3648 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_39
timestamp 1679581782
transform 1 0 4320 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_46
timestamp 1679581782
transform 1 0 4992 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_53
timestamp 1679581782
transform 1 0 5664 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_60
timestamp 1679581782
transform 1 0 6336 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_67
timestamp 1679581782
transform 1 0 7008 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_74
timestamp 1679581782
transform 1 0 7680 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_81
timestamp 1679581782
transform 1 0 8352 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_88
timestamp 1679581782
transform 1 0 9024 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_95
timestamp 1679581782
transform 1 0 9696 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_102
timestamp 1679581782
transform 1 0 10368 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_109
timestamp 1679581782
transform 1 0 11040 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_116
timestamp 1679581782
transform 1 0 11712 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_123
timestamp 1679581782
transform 1 0 12384 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_130
timestamp 1679581782
transform 1 0 13056 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_137
timestamp 1679581782
transform 1 0 13728 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_144
timestamp 1679581782
transform 1 0 14400 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_151
timestamp 1679581782
transform 1 0 15072 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_158
timestamp 1679581782
transform 1 0 15744 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_165
timestamp 1679581782
transform 1 0 16416 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_172
timestamp 1679581782
transform 1 0 17088 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_179
timestamp 1679581782
transform 1 0 17760 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_186
timestamp 1679581782
transform 1 0 18432 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_193
timestamp 1679581782
transform 1 0 19104 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_200
timestamp 1679581782
transform 1 0 19776 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_207
timestamp 1679581782
transform 1 0 20448 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_214
timestamp 1679581782
transform 1 0 21120 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_221
timestamp 1679581782
transform 1 0 21792 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_228
timestamp 1679581782
transform 1 0 22464 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_235
timestamp 1679581782
transform 1 0 23136 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_242
timestamp 1679581782
transform 1 0 23808 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_249
timestamp 1679581782
transform 1 0 24480 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_256
timestamp 1679581782
transform 1 0 25152 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_263
timestamp 1679581782
transform 1 0 25824 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_270
timestamp 1679581782
transform 1 0 26496 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_277
timestamp 1679581782
transform 1 0 27168 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_284
timestamp 1679581782
transform 1 0 27840 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_291
timestamp 1679581782
transform 1 0 28512 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_298
timestamp 1679581782
transform 1 0 29184 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_305
timestamp 1679581782
transform 1 0 29856 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_312
timestamp 1679581782
transform 1 0 30528 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_319
timestamp 1679581782
transform 1 0 31200 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_326
timestamp 1679581782
transform 1 0 31872 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_333
timestamp 1679581782
transform 1 0 32544 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_340
timestamp 1679581782
transform 1 0 33216 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_347
timestamp 1679581782
transform 1 0 33888 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_354
timestamp 1679581782
transform 1 0 34560 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_361
timestamp 1679581782
transform 1 0 35232 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_368
timestamp 1679581782
transform 1 0 35904 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_375
timestamp 1679581782
transform 1 0 36576 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_382
timestamp 1679581782
transform 1 0 37248 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_389
timestamp 1679581782
transform 1 0 37920 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_396
timestamp 1679581782
transform 1 0 38592 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_403
timestamp 1679581782
transform 1 0 39264 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_410
timestamp 1679581782
transform 1 0 39936 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_417
timestamp 1679581782
transform 1 0 40608 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_424
timestamp 1679581782
transform 1 0 41280 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_431
timestamp 1679581782
transform 1 0 41952 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_438
timestamp 1679581782
transform 1 0 42624 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_445
timestamp 1679581782
transform 1 0 43296 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_452
timestamp 1679581782
transform 1 0 43968 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_459
timestamp 1679581782
transform 1 0 44640 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_466
timestamp 1679581782
transform 1 0 45312 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_473
timestamp 1679581782
transform 1 0 45984 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_480
timestamp 1679581782
transform 1 0 46656 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_487
timestamp 1679581782
transform 1 0 47328 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_494
timestamp 1679581782
transform 1 0 48000 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_501
timestamp 1679581782
transform 1 0 48672 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_508
timestamp 1679581782
transform 1 0 49344 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_515
timestamp 1679581782
transform 1 0 50016 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_522
timestamp 1679581782
transform 1 0 50688 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_529
timestamp 1679581782
transform 1 0 51360 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_536
timestamp 1679581782
transform 1 0 52032 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_543
timestamp 1679581782
transform 1 0 52704 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_550
timestamp 1679581782
transform 1 0 53376 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_557
timestamp 1679581782
transform 1 0 54048 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_564
timestamp 1679581782
transform 1 0 54720 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_571
timestamp 1679581782
transform 1 0 55392 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_578
timestamp 1679581782
transform 1 0 56064 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_585
timestamp 1679581782
transform 1 0 56736 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_592
timestamp 1679581782
transform 1 0 57408 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_599
timestamp 1679581782
transform 1 0 58080 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_606
timestamp 1679581782
transform 1 0 58752 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_613
timestamp 1679581782
transform 1 0 59424 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_620
timestamp 1679581782
transform 1 0 60096 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_627
timestamp 1679581782
transform 1 0 60768 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_634
timestamp 1679581782
transform 1 0 61440 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_641
timestamp 1679581782
transform 1 0 62112 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_648
timestamp 1679581782
transform 1 0 62784 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_655
timestamp 1679581782
transform 1 0 63456 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_662
timestamp 1679581782
transform 1 0 64128 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_669
timestamp 1679581782
transform 1 0 64800 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_676
timestamp 1679581782
transform 1 0 65472 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_683
timestamp 1679581782
transform 1 0 66144 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_690
timestamp 1679581782
transform 1 0 66816 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_697
timestamp 1679581782
transform 1 0 67488 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_704
timestamp 1679581782
transform 1 0 68160 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_711
timestamp 1679581782
transform 1 0 68832 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_718
timestamp 1679581782
transform 1 0 69504 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_725
timestamp 1679581782
transform 1 0 70176 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_732
timestamp 1679581782
transform 1 0 70848 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_739
timestamp 1679581782
transform 1 0 71520 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_746
timestamp 1679581782
transform 1 0 72192 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_753
timestamp 1679581782
transform 1 0 72864 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_760
timestamp 1679581782
transform 1 0 73536 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_767
timestamp 1679581782
transform 1 0 74208 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_774
timestamp 1679581782
transform 1 0 74880 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_781
timestamp 1679581782
transform 1 0 75552 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_788
timestamp 1679581782
transform 1 0 76224 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_795
timestamp 1679581782
transform 1 0 76896 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_802
timestamp 1679581782
transform 1 0 77568 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_809
timestamp 1679581782
transform 1 0 78240 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_816
timestamp 1679581782
transform 1 0 78912 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_823
timestamp 1679581782
transform 1 0 79584 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_830
timestamp 1679581782
transform 1 0 80256 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_837
timestamp 1679581782
transform 1 0 80928 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_844
timestamp 1679581782
transform 1 0 81600 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_851
timestamp 1679581782
transform 1 0 82272 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_858
timestamp 1679581782
transform 1 0 82944 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_865
timestamp 1679581782
transform 1 0 83616 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_872
timestamp 1679581782
transform 1 0 84288 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_879
timestamp 1679581782
transform 1 0 84960 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_886
timestamp 1679581782
transform 1 0 85632 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_893
timestamp 1679581782
transform 1 0 86304 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_900
timestamp 1679581782
transform 1 0 86976 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_907
timestamp 1679581782
transform 1 0 87648 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_914
timestamp 1679581782
transform 1 0 88320 0 1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_12_921
timestamp 1679577901
transform 1 0 88992 0 1 9828
box -48 -56 432 834
use sg13g2_decap_8  FILLER_13_4
timestamp 1679581782
transform 1 0 960 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_11
timestamp 1679581782
transform 1 0 1632 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_18
timestamp 1679581782
transform 1 0 2304 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_25
timestamp 1679581782
transform 1 0 2976 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_32
timestamp 1679581782
transform 1 0 3648 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_39
timestamp 1679581782
transform 1 0 4320 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_46
timestamp 1679581782
transform 1 0 4992 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_53
timestamp 1679581782
transform 1 0 5664 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_60
timestamp 1679581782
transform 1 0 6336 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_67
timestamp 1679581782
transform 1 0 7008 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_74
timestamp 1679581782
transform 1 0 7680 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_81
timestamp 1679581782
transform 1 0 8352 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_88
timestamp 1679581782
transform 1 0 9024 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_95
timestamp 1679581782
transform 1 0 9696 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_102
timestamp 1679581782
transform 1 0 10368 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_109
timestamp 1679581782
transform 1 0 11040 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_116
timestamp 1679581782
transform 1 0 11712 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_123
timestamp 1679581782
transform 1 0 12384 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_130
timestamp 1679581782
transform 1 0 13056 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_137
timestamp 1679581782
transform 1 0 13728 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_144
timestamp 1679581782
transform 1 0 14400 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_151
timestamp 1679581782
transform 1 0 15072 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_158
timestamp 1679581782
transform 1 0 15744 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_165
timestamp 1679581782
transform 1 0 16416 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_172
timestamp 1679581782
transform 1 0 17088 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_179
timestamp 1679581782
transform 1 0 17760 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_186
timestamp 1679581782
transform 1 0 18432 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_193
timestamp 1679581782
transform 1 0 19104 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_200
timestamp 1679581782
transform 1 0 19776 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_207
timestamp 1679581782
transform 1 0 20448 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_214
timestamp 1679581782
transform 1 0 21120 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_221
timestamp 1679581782
transform 1 0 21792 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_228
timestamp 1679581782
transform 1 0 22464 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_235
timestamp 1679581782
transform 1 0 23136 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_242
timestamp 1679581782
transform 1 0 23808 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_249
timestamp 1679581782
transform 1 0 24480 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_256
timestamp 1679581782
transform 1 0 25152 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_263
timestamp 1679581782
transform 1 0 25824 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_270
timestamp 1679581782
transform 1 0 26496 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_277
timestamp 1679581782
transform 1 0 27168 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_284
timestamp 1679581782
transform 1 0 27840 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_291
timestamp 1679581782
transform 1 0 28512 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_298
timestamp 1679581782
transform 1 0 29184 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_305
timestamp 1679581782
transform 1 0 29856 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_312
timestamp 1679581782
transform 1 0 30528 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_319
timestamp 1679581782
transform 1 0 31200 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_326
timestamp 1679581782
transform 1 0 31872 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_333
timestamp 1679581782
transform 1 0 32544 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_340
timestamp 1679581782
transform 1 0 33216 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_347
timestamp 1679581782
transform 1 0 33888 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_354
timestamp 1679581782
transform 1 0 34560 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_361
timestamp 1679581782
transform 1 0 35232 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_368
timestamp 1679581782
transform 1 0 35904 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_375
timestamp 1679581782
transform 1 0 36576 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_382
timestamp 1679581782
transform 1 0 37248 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_389
timestamp 1679581782
transform 1 0 37920 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_396
timestamp 1679581782
transform 1 0 38592 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_403
timestamp 1679581782
transform 1 0 39264 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_410
timestamp 1679581782
transform 1 0 39936 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_417
timestamp 1679581782
transform 1 0 40608 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_424
timestamp 1679581782
transform 1 0 41280 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_431
timestamp 1679581782
transform 1 0 41952 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_438
timestamp 1679581782
transform 1 0 42624 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_445
timestamp 1679581782
transform 1 0 43296 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_452
timestamp 1679581782
transform 1 0 43968 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_459
timestamp 1679581782
transform 1 0 44640 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_466
timestamp 1679581782
transform 1 0 45312 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_473
timestamp 1679581782
transform 1 0 45984 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_480
timestamp 1679581782
transform 1 0 46656 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_487
timestamp 1679581782
transform 1 0 47328 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_494
timestamp 1679581782
transform 1 0 48000 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_501
timestamp 1679581782
transform 1 0 48672 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_508
timestamp 1679581782
transform 1 0 49344 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_515
timestamp 1679581782
transform 1 0 50016 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_522
timestamp 1679581782
transform 1 0 50688 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_529
timestamp 1679581782
transform 1 0 51360 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_536
timestamp 1679581782
transform 1 0 52032 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_543
timestamp 1679581782
transform 1 0 52704 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_550
timestamp 1679581782
transform 1 0 53376 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_557
timestamp 1679581782
transform 1 0 54048 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_564
timestamp 1679581782
transform 1 0 54720 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_571
timestamp 1679581782
transform 1 0 55392 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_578
timestamp 1679581782
transform 1 0 56064 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_585
timestamp 1679581782
transform 1 0 56736 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_592
timestamp 1679581782
transform 1 0 57408 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_599
timestamp 1679581782
transform 1 0 58080 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_606
timestamp 1679581782
transform 1 0 58752 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_613
timestamp 1679581782
transform 1 0 59424 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_620
timestamp 1679581782
transform 1 0 60096 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_627
timestamp 1679581782
transform 1 0 60768 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_634
timestamp 1679581782
transform 1 0 61440 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_641
timestamp 1679581782
transform 1 0 62112 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_648
timestamp 1679581782
transform 1 0 62784 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_655
timestamp 1679581782
transform 1 0 63456 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_662
timestamp 1679581782
transform 1 0 64128 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_669
timestamp 1679581782
transform 1 0 64800 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_676
timestamp 1679581782
transform 1 0 65472 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_683
timestamp 1679581782
transform 1 0 66144 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_690
timestamp 1679581782
transform 1 0 66816 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_697
timestamp 1679581782
transform 1 0 67488 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_704
timestamp 1679581782
transform 1 0 68160 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_711
timestamp 1679581782
transform 1 0 68832 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_718
timestamp 1679581782
transform 1 0 69504 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_725
timestamp 1679581782
transform 1 0 70176 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_732
timestamp 1679581782
transform 1 0 70848 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_739
timestamp 1679581782
transform 1 0 71520 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_746
timestamp 1679581782
transform 1 0 72192 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_753
timestamp 1679581782
transform 1 0 72864 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_760
timestamp 1679581782
transform 1 0 73536 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_767
timestamp 1679581782
transform 1 0 74208 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_774
timestamp 1679581782
transform 1 0 74880 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_781
timestamp 1679581782
transform 1 0 75552 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_788
timestamp 1679581782
transform 1 0 76224 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_795
timestamp 1679581782
transform 1 0 76896 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_802
timestamp 1679581782
transform 1 0 77568 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_809
timestamp 1679581782
transform 1 0 78240 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_816
timestamp 1679581782
transform 1 0 78912 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_823
timestamp 1679581782
transform 1 0 79584 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_830
timestamp 1679581782
transform 1 0 80256 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_837
timestamp 1679581782
transform 1 0 80928 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_844
timestamp 1679581782
transform 1 0 81600 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_851
timestamp 1679581782
transform 1 0 82272 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_858
timestamp 1679581782
transform 1 0 82944 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_865
timestamp 1679581782
transform 1 0 83616 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_872
timestamp 1679581782
transform 1 0 84288 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_879
timestamp 1679581782
transform 1 0 84960 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_886
timestamp 1679581782
transform 1 0 85632 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_893
timestamp 1679581782
transform 1 0 86304 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_900
timestamp 1679581782
transform 1 0 86976 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_907
timestamp 1679581782
transform 1 0 87648 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_914
timestamp 1679581782
transform 1 0 88320 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_921
timestamp 1679577901
transform 1 0 88992 0 -1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_14_4
timestamp 1679581782
transform 1 0 960 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_11
timestamp 1679581782
transform 1 0 1632 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_18
timestamp 1679581782
transform 1 0 2304 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_25
timestamp 1679581782
transform 1 0 2976 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_32
timestamp 1679581782
transform 1 0 3648 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_39
timestamp 1679581782
transform 1 0 4320 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_46
timestamp 1679581782
transform 1 0 4992 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_53
timestamp 1679581782
transform 1 0 5664 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_60
timestamp 1679581782
transform 1 0 6336 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_67
timestamp 1679581782
transform 1 0 7008 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_74
timestamp 1679581782
transform 1 0 7680 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_81
timestamp 1679581782
transform 1 0 8352 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_88
timestamp 1679581782
transform 1 0 9024 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_95
timestamp 1679581782
transform 1 0 9696 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_102
timestamp 1679581782
transform 1 0 10368 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_109
timestamp 1679581782
transform 1 0 11040 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_116
timestamp 1679581782
transform 1 0 11712 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_123
timestamp 1679581782
transform 1 0 12384 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_130
timestamp 1679581782
transform 1 0 13056 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_137
timestamp 1679581782
transform 1 0 13728 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_144
timestamp 1679581782
transform 1 0 14400 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_151
timestamp 1679581782
transform 1 0 15072 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_158
timestamp 1679581782
transform 1 0 15744 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_165
timestamp 1679581782
transform 1 0 16416 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_172
timestamp 1679581782
transform 1 0 17088 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_179
timestamp 1679581782
transform 1 0 17760 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_186
timestamp 1679581782
transform 1 0 18432 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_193
timestamp 1679581782
transform 1 0 19104 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_200
timestamp 1679581782
transform 1 0 19776 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_207
timestamp 1679581782
transform 1 0 20448 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_214
timestamp 1679581782
transform 1 0 21120 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_221
timestamp 1679581782
transform 1 0 21792 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_228
timestamp 1679581782
transform 1 0 22464 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_235
timestamp 1679581782
transform 1 0 23136 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_242
timestamp 1679581782
transform 1 0 23808 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_249
timestamp 1679581782
transform 1 0 24480 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_256
timestamp 1679581782
transform 1 0 25152 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_263
timestamp 1679581782
transform 1 0 25824 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_270
timestamp 1679581782
transform 1 0 26496 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_277
timestamp 1679581782
transform 1 0 27168 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_284
timestamp 1679581782
transform 1 0 27840 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_291
timestamp 1679581782
transform 1 0 28512 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_298
timestamp 1679581782
transform 1 0 29184 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_305
timestamp 1679581782
transform 1 0 29856 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_312
timestamp 1679581782
transform 1 0 30528 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_319
timestamp 1679581782
transform 1 0 31200 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_326
timestamp 1679581782
transform 1 0 31872 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_333
timestamp 1679581782
transform 1 0 32544 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_340
timestamp 1679581782
transform 1 0 33216 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_347
timestamp 1679581782
transform 1 0 33888 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_354
timestamp 1679581782
transform 1 0 34560 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_361
timestamp 1679581782
transform 1 0 35232 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_368
timestamp 1679581782
transform 1 0 35904 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_375
timestamp 1679581782
transform 1 0 36576 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_382
timestamp 1679581782
transform 1 0 37248 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_389
timestamp 1679581782
transform 1 0 37920 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_396
timestamp 1679581782
transform 1 0 38592 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_403
timestamp 1679581782
transform 1 0 39264 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_410
timestamp 1679581782
transform 1 0 39936 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_417
timestamp 1679581782
transform 1 0 40608 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_424
timestamp 1679581782
transform 1 0 41280 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_431
timestamp 1679581782
transform 1 0 41952 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_438
timestamp 1679581782
transform 1 0 42624 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_445
timestamp 1679581782
transform 1 0 43296 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_452
timestamp 1679581782
transform 1 0 43968 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_459
timestamp 1679581782
transform 1 0 44640 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_466
timestamp 1679581782
transform 1 0 45312 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_473
timestamp 1679581782
transform 1 0 45984 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_480
timestamp 1679581782
transform 1 0 46656 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_487
timestamp 1679581782
transform 1 0 47328 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_494
timestamp 1679581782
transform 1 0 48000 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_501
timestamp 1679581782
transform 1 0 48672 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_508
timestamp 1679581782
transform 1 0 49344 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_515
timestamp 1679581782
transform 1 0 50016 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_522
timestamp 1679581782
transform 1 0 50688 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_529
timestamp 1679581782
transform 1 0 51360 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_536
timestamp 1679581782
transform 1 0 52032 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_543
timestamp 1679581782
transform 1 0 52704 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_550
timestamp 1679581782
transform 1 0 53376 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_557
timestamp 1679581782
transform 1 0 54048 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_564
timestamp 1679581782
transform 1 0 54720 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_571
timestamp 1679581782
transform 1 0 55392 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_578
timestamp 1679581782
transform 1 0 56064 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_585
timestamp 1679581782
transform 1 0 56736 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_592
timestamp 1679581782
transform 1 0 57408 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_599
timestamp 1679581782
transform 1 0 58080 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_606
timestamp 1679581782
transform 1 0 58752 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_613
timestamp 1679581782
transform 1 0 59424 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_620
timestamp 1679581782
transform 1 0 60096 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_627
timestamp 1679581782
transform 1 0 60768 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_634
timestamp 1679581782
transform 1 0 61440 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_641
timestamp 1679581782
transform 1 0 62112 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_648
timestamp 1679581782
transform 1 0 62784 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_655
timestamp 1679581782
transform 1 0 63456 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_662
timestamp 1679581782
transform 1 0 64128 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_669
timestamp 1679581782
transform 1 0 64800 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_676
timestamp 1679581782
transform 1 0 65472 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_683
timestamp 1679581782
transform 1 0 66144 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_690
timestamp 1679581782
transform 1 0 66816 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_697
timestamp 1679581782
transform 1 0 67488 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_704
timestamp 1679581782
transform 1 0 68160 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_711
timestamp 1679581782
transform 1 0 68832 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_718
timestamp 1679581782
transform 1 0 69504 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_725
timestamp 1679581782
transform 1 0 70176 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_732
timestamp 1679581782
transform 1 0 70848 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_739
timestamp 1679581782
transform 1 0 71520 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_746
timestamp 1679581782
transform 1 0 72192 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_753
timestamp 1679581782
transform 1 0 72864 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_760
timestamp 1679581782
transform 1 0 73536 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_767
timestamp 1679581782
transform 1 0 74208 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_774
timestamp 1679581782
transform 1 0 74880 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_781
timestamp 1679581782
transform 1 0 75552 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_788
timestamp 1679581782
transform 1 0 76224 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_795
timestamp 1679581782
transform 1 0 76896 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_802
timestamp 1679581782
transform 1 0 77568 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_809
timestamp 1679581782
transform 1 0 78240 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_816
timestamp 1679581782
transform 1 0 78912 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_823
timestamp 1679581782
transform 1 0 79584 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_830
timestamp 1679581782
transform 1 0 80256 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_837
timestamp 1679581782
transform 1 0 80928 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_844
timestamp 1679581782
transform 1 0 81600 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_851
timestamp 1679581782
transform 1 0 82272 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_858
timestamp 1679581782
transform 1 0 82944 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_865
timestamp 1679581782
transform 1 0 83616 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_872
timestamp 1679581782
transform 1 0 84288 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_879
timestamp 1679581782
transform 1 0 84960 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_886
timestamp 1679581782
transform 1 0 85632 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_893
timestamp 1679581782
transform 1 0 86304 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_900
timestamp 1679581782
transform 1 0 86976 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_907
timestamp 1679581782
transform 1 0 87648 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_914
timestamp 1679581782
transform 1 0 88320 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_921
timestamp 1679577901
transform 1 0 88992 0 1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_15_4
timestamp 1679581782
transform 1 0 960 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_11
timestamp 1679581782
transform 1 0 1632 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_18
timestamp 1679581782
transform 1 0 2304 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_25
timestamp 1679581782
transform 1 0 2976 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_32
timestamp 1679581782
transform 1 0 3648 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_39
timestamp 1679581782
transform 1 0 4320 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_46
timestamp 1679581782
transform 1 0 4992 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_53
timestamp 1679581782
transform 1 0 5664 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_60
timestamp 1679581782
transform 1 0 6336 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_67
timestamp 1679581782
transform 1 0 7008 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_74
timestamp 1679581782
transform 1 0 7680 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_81
timestamp 1679581782
transform 1 0 8352 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_88
timestamp 1679581782
transform 1 0 9024 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_95
timestamp 1679581782
transform 1 0 9696 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_102
timestamp 1679581782
transform 1 0 10368 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_109
timestamp 1679581782
transform 1 0 11040 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_116
timestamp 1679581782
transform 1 0 11712 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_123
timestamp 1679581782
transform 1 0 12384 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_130
timestamp 1679581782
transform 1 0 13056 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_137
timestamp 1679581782
transform 1 0 13728 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_144
timestamp 1679581782
transform 1 0 14400 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_151
timestamp 1679581782
transform 1 0 15072 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_158
timestamp 1679581782
transform 1 0 15744 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_165
timestamp 1679581782
transform 1 0 16416 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_172
timestamp 1679581782
transform 1 0 17088 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_179
timestamp 1679581782
transform 1 0 17760 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_186
timestamp 1679581782
transform 1 0 18432 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_193
timestamp 1679581782
transform 1 0 19104 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_200
timestamp 1679581782
transform 1 0 19776 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_207
timestamp 1679581782
transform 1 0 20448 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_214
timestamp 1679581782
transform 1 0 21120 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_221
timestamp 1679581782
transform 1 0 21792 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_228
timestamp 1679581782
transform 1 0 22464 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_235
timestamp 1679581782
transform 1 0 23136 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_242
timestamp 1679581782
transform 1 0 23808 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_249
timestamp 1679581782
transform 1 0 24480 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_256
timestamp 1679581782
transform 1 0 25152 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_263
timestamp 1679581782
transform 1 0 25824 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_270
timestamp 1679581782
transform 1 0 26496 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_277
timestamp 1679581782
transform 1 0 27168 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_284
timestamp 1679581782
transform 1 0 27840 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_291
timestamp 1679581782
transform 1 0 28512 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_298
timestamp 1679581782
transform 1 0 29184 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_305
timestamp 1679581782
transform 1 0 29856 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_312
timestamp 1679581782
transform 1 0 30528 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_319
timestamp 1679581782
transform 1 0 31200 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_326
timestamp 1679581782
transform 1 0 31872 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_333
timestamp 1679581782
transform 1 0 32544 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_340
timestamp 1679581782
transform 1 0 33216 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_347
timestamp 1679581782
transform 1 0 33888 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_354
timestamp 1679581782
transform 1 0 34560 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_361
timestamp 1679581782
transform 1 0 35232 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_368
timestamp 1679581782
transform 1 0 35904 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_375
timestamp 1679581782
transform 1 0 36576 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_382
timestamp 1679581782
transform 1 0 37248 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_389
timestamp 1679581782
transform 1 0 37920 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_396
timestamp 1679581782
transform 1 0 38592 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_403
timestamp 1679581782
transform 1 0 39264 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_410
timestamp 1679581782
transform 1 0 39936 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_417
timestamp 1679581782
transform 1 0 40608 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_424
timestamp 1679581782
transform 1 0 41280 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_431
timestamp 1679581782
transform 1 0 41952 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_438
timestamp 1679581782
transform 1 0 42624 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_445
timestamp 1679581782
transform 1 0 43296 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_452
timestamp 1679581782
transform 1 0 43968 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_459
timestamp 1679581782
transform 1 0 44640 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_466
timestamp 1679581782
transform 1 0 45312 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_473
timestamp 1679581782
transform 1 0 45984 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_480
timestamp 1679581782
transform 1 0 46656 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_487
timestamp 1679581782
transform 1 0 47328 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_494
timestamp 1679581782
transform 1 0 48000 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_501
timestamp 1679581782
transform 1 0 48672 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_508
timestamp 1679581782
transform 1 0 49344 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_515
timestamp 1679581782
transform 1 0 50016 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_522
timestamp 1679581782
transform 1 0 50688 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_529
timestamp 1679581782
transform 1 0 51360 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_536
timestamp 1679581782
transform 1 0 52032 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_543
timestamp 1679581782
transform 1 0 52704 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_550
timestamp 1679581782
transform 1 0 53376 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_557
timestamp 1679581782
transform 1 0 54048 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_564
timestamp 1679581782
transform 1 0 54720 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_571
timestamp 1679581782
transform 1 0 55392 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_578
timestamp 1679581782
transform 1 0 56064 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_585
timestamp 1679581782
transform 1 0 56736 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_592
timestamp 1679581782
transform 1 0 57408 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_599
timestamp 1679581782
transform 1 0 58080 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_606
timestamp 1679581782
transform 1 0 58752 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_613
timestamp 1679581782
transform 1 0 59424 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_620
timestamp 1679581782
transform 1 0 60096 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_627
timestamp 1679581782
transform 1 0 60768 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_634
timestamp 1679581782
transform 1 0 61440 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_641
timestamp 1679581782
transform 1 0 62112 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_648
timestamp 1679581782
transform 1 0 62784 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_655
timestamp 1679581782
transform 1 0 63456 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_662
timestamp 1679581782
transform 1 0 64128 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_669
timestamp 1679581782
transform 1 0 64800 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_676
timestamp 1679581782
transform 1 0 65472 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_683
timestamp 1679581782
transform 1 0 66144 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_690
timestamp 1679581782
transform 1 0 66816 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_697
timestamp 1679581782
transform 1 0 67488 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_704
timestamp 1679581782
transform 1 0 68160 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_711
timestamp 1679581782
transform 1 0 68832 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_718
timestamp 1679581782
transform 1 0 69504 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_725
timestamp 1679581782
transform 1 0 70176 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_732
timestamp 1679581782
transform 1 0 70848 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_739
timestamp 1679581782
transform 1 0 71520 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_746
timestamp 1679581782
transform 1 0 72192 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_753
timestamp 1679581782
transform 1 0 72864 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_760
timestamp 1679581782
transform 1 0 73536 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_767
timestamp 1679581782
transform 1 0 74208 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_774
timestamp 1679581782
transform 1 0 74880 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_781
timestamp 1679581782
transform 1 0 75552 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_788
timestamp 1679581782
transform 1 0 76224 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_795
timestamp 1679581782
transform 1 0 76896 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_802
timestamp 1679581782
transform 1 0 77568 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_809
timestamp 1679581782
transform 1 0 78240 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_816
timestamp 1679581782
transform 1 0 78912 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_823
timestamp 1679581782
transform 1 0 79584 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_830
timestamp 1679581782
transform 1 0 80256 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_837
timestamp 1679581782
transform 1 0 80928 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_844
timestamp 1679581782
transform 1 0 81600 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_851
timestamp 1679581782
transform 1 0 82272 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_858
timestamp 1679581782
transform 1 0 82944 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_865
timestamp 1679581782
transform 1 0 83616 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_872
timestamp 1679581782
transform 1 0 84288 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_879
timestamp 1679581782
transform 1 0 84960 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_886
timestamp 1679581782
transform 1 0 85632 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_893
timestamp 1679581782
transform 1 0 86304 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_900
timestamp 1679581782
transform 1 0 86976 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_907
timestamp 1679581782
transform 1 0 87648 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_914
timestamp 1679581782
transform 1 0 88320 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_15_921
timestamp 1679577901
transform 1 0 88992 0 -1 12852
box -48 -56 432 834
use sg13g2_decap_8  FILLER_16_4
timestamp 1679581782
transform 1 0 960 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_11
timestamp 1679581782
transform 1 0 1632 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_18
timestamp 1679581782
transform 1 0 2304 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_25
timestamp 1679581782
transform 1 0 2976 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_32
timestamp 1679581782
transform 1 0 3648 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_39
timestamp 1679581782
transform 1 0 4320 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_46
timestamp 1679581782
transform 1 0 4992 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_53
timestamp 1679581782
transform 1 0 5664 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_60
timestamp 1679581782
transform 1 0 6336 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_67
timestamp 1679581782
transform 1 0 7008 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_74
timestamp 1679581782
transform 1 0 7680 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_81
timestamp 1679581782
transform 1 0 8352 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_88
timestamp 1679581782
transform 1 0 9024 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_95
timestamp 1679581782
transform 1 0 9696 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_102
timestamp 1679581782
transform 1 0 10368 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_109
timestamp 1679581782
transform 1 0 11040 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_116
timestamp 1679581782
transform 1 0 11712 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_123
timestamp 1679581782
transform 1 0 12384 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_130
timestamp 1679581782
transform 1 0 13056 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_137
timestamp 1679581782
transform 1 0 13728 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_144
timestamp 1679581782
transform 1 0 14400 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_151
timestamp 1679581782
transform 1 0 15072 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_158
timestamp 1679581782
transform 1 0 15744 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_165
timestamp 1679581782
transform 1 0 16416 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_172
timestamp 1679581782
transform 1 0 17088 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_179
timestamp 1679581782
transform 1 0 17760 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_186
timestamp 1679581782
transform 1 0 18432 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_193
timestamp 1679581782
transform 1 0 19104 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_200
timestamp 1679581782
transform 1 0 19776 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_207
timestamp 1679581782
transform 1 0 20448 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_214
timestamp 1679581782
transform 1 0 21120 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_221
timestamp 1679581782
transform 1 0 21792 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_228
timestamp 1679581782
transform 1 0 22464 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_235
timestamp 1679581782
transform 1 0 23136 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_242
timestamp 1679581782
transform 1 0 23808 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_249
timestamp 1679581782
transform 1 0 24480 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_256
timestamp 1679581782
transform 1 0 25152 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_263
timestamp 1679581782
transform 1 0 25824 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_270
timestamp 1679581782
transform 1 0 26496 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_277
timestamp 1679581782
transform 1 0 27168 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_284
timestamp 1679581782
transform 1 0 27840 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_291
timestamp 1679581782
transform 1 0 28512 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_298
timestamp 1679581782
transform 1 0 29184 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_305
timestamp 1679581782
transform 1 0 29856 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_312
timestamp 1679581782
transform 1 0 30528 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_319
timestamp 1679581782
transform 1 0 31200 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_326
timestamp 1679581782
transform 1 0 31872 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_333
timestamp 1679581782
transform 1 0 32544 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_340
timestamp 1679581782
transform 1 0 33216 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_347
timestamp 1679581782
transform 1 0 33888 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_354
timestamp 1679581782
transform 1 0 34560 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_361
timestamp 1679581782
transform 1 0 35232 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_368
timestamp 1679581782
transform 1 0 35904 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_375
timestamp 1679581782
transform 1 0 36576 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_382
timestamp 1679581782
transform 1 0 37248 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_389
timestamp 1679581782
transform 1 0 37920 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_396
timestamp 1679581782
transform 1 0 38592 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_403
timestamp 1679581782
transform 1 0 39264 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_410
timestamp 1679581782
transform 1 0 39936 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_417
timestamp 1679581782
transform 1 0 40608 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_424
timestamp 1679581782
transform 1 0 41280 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_431
timestamp 1679581782
transform 1 0 41952 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_438
timestamp 1679581782
transform 1 0 42624 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_445
timestamp 1679581782
transform 1 0 43296 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_452
timestamp 1679581782
transform 1 0 43968 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_459
timestamp 1679581782
transform 1 0 44640 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_466
timestamp 1679581782
transform 1 0 45312 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_473
timestamp 1679581782
transform 1 0 45984 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_480
timestamp 1679581782
transform 1 0 46656 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_487
timestamp 1679581782
transform 1 0 47328 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_494
timestamp 1679581782
transform 1 0 48000 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_501
timestamp 1679581782
transform 1 0 48672 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_508
timestamp 1679581782
transform 1 0 49344 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_515
timestamp 1679581782
transform 1 0 50016 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_522
timestamp 1679581782
transform 1 0 50688 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_529
timestamp 1679581782
transform 1 0 51360 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_536
timestamp 1679581782
transform 1 0 52032 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_543
timestamp 1679581782
transform 1 0 52704 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_550
timestamp 1679581782
transform 1 0 53376 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_557
timestamp 1679581782
transform 1 0 54048 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_564
timestamp 1679581782
transform 1 0 54720 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_571
timestamp 1679581782
transform 1 0 55392 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_578
timestamp 1679581782
transform 1 0 56064 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_585
timestamp 1679581782
transform 1 0 56736 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_592
timestamp 1679581782
transform 1 0 57408 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_599
timestamp 1679581782
transform 1 0 58080 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_606
timestamp 1679581782
transform 1 0 58752 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_613
timestamp 1679581782
transform 1 0 59424 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_620
timestamp 1679581782
transform 1 0 60096 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_627
timestamp 1679581782
transform 1 0 60768 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_634
timestamp 1679581782
transform 1 0 61440 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_641
timestamp 1679581782
transform 1 0 62112 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_648
timestamp 1679581782
transform 1 0 62784 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_655
timestamp 1679581782
transform 1 0 63456 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_662
timestamp 1679581782
transform 1 0 64128 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_669
timestamp 1679581782
transform 1 0 64800 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_676
timestamp 1679581782
transform 1 0 65472 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_683
timestamp 1679581782
transform 1 0 66144 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_690
timestamp 1679581782
transform 1 0 66816 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_697
timestamp 1679581782
transform 1 0 67488 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_704
timestamp 1679581782
transform 1 0 68160 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_711
timestamp 1679581782
transform 1 0 68832 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_718
timestamp 1679581782
transform 1 0 69504 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_725
timestamp 1679581782
transform 1 0 70176 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_732
timestamp 1679581782
transform 1 0 70848 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_739
timestamp 1679581782
transform 1 0 71520 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_746
timestamp 1679581782
transform 1 0 72192 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_753
timestamp 1679581782
transform 1 0 72864 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_760
timestamp 1679581782
transform 1 0 73536 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_767
timestamp 1679581782
transform 1 0 74208 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_774
timestamp 1679581782
transform 1 0 74880 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_781
timestamp 1679581782
transform 1 0 75552 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_788
timestamp 1679581782
transform 1 0 76224 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_795
timestamp 1679581782
transform 1 0 76896 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_802
timestamp 1679581782
transform 1 0 77568 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_809
timestamp 1679581782
transform 1 0 78240 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_816
timestamp 1679581782
transform 1 0 78912 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_823
timestamp 1679581782
transform 1 0 79584 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_830
timestamp 1679581782
transform 1 0 80256 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_837
timestamp 1679581782
transform 1 0 80928 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_844
timestamp 1679581782
transform 1 0 81600 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_851
timestamp 1679581782
transform 1 0 82272 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_858
timestamp 1679581782
transform 1 0 82944 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_865
timestamp 1679581782
transform 1 0 83616 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_872
timestamp 1679581782
transform 1 0 84288 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_879
timestamp 1679581782
transform 1 0 84960 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_886
timestamp 1679581782
transform 1 0 85632 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_893
timestamp 1679581782
transform 1 0 86304 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_900
timestamp 1679581782
transform 1 0 86976 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_907
timestamp 1679581782
transform 1 0 87648 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_914
timestamp 1679581782
transform 1 0 88320 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_921
timestamp 1679577901
transform 1 0 88992 0 1 12852
box -48 -56 432 834
use sg13g2_decap_8  FILLER_17_0
timestamp 1679581782
transform 1 0 576 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_7
timestamp 1679581782
transform 1 0 1248 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_14
timestamp 1679581782
transform 1 0 1920 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_21
timestamp 1679581782
transform 1 0 2592 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_28
timestamp 1679581782
transform 1 0 3264 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_35
timestamp 1679581782
transform 1 0 3936 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_42
timestamp 1679581782
transform 1 0 4608 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_49
timestamp 1679581782
transform 1 0 5280 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_56
timestamp 1679581782
transform 1 0 5952 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_63
timestamp 1679581782
transform 1 0 6624 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_70
timestamp 1679581782
transform 1 0 7296 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_77
timestamp 1679581782
transform 1 0 7968 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_84
timestamp 1679581782
transform 1 0 8640 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_91
timestamp 1679581782
transform 1 0 9312 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_98
timestamp 1679581782
transform 1 0 9984 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_105
timestamp 1679581782
transform 1 0 10656 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_112
timestamp 1679581782
transform 1 0 11328 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_119
timestamp 1679581782
transform 1 0 12000 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_126
timestamp 1679581782
transform 1 0 12672 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_133
timestamp 1679581782
transform 1 0 13344 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_140
timestamp 1679581782
transform 1 0 14016 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_147
timestamp 1679581782
transform 1 0 14688 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_154
timestamp 1679581782
transform 1 0 15360 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_161
timestamp 1679581782
transform 1 0 16032 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_168
timestamp 1679581782
transform 1 0 16704 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_175
timestamp 1679581782
transform 1 0 17376 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_182
timestamp 1679581782
transform 1 0 18048 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_189
timestamp 1679581782
transform 1 0 18720 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_196
timestamp 1679581782
transform 1 0 19392 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_203
timestamp 1679581782
transform 1 0 20064 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_210
timestamp 1679581782
transform 1 0 20736 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_217
timestamp 1679581782
transform 1 0 21408 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_224
timestamp 1679581782
transform 1 0 22080 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_231
timestamp 1679581782
transform 1 0 22752 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_238
timestamp 1679581782
transform 1 0 23424 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_245
timestamp 1679581782
transform 1 0 24096 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_252
timestamp 1679581782
transform 1 0 24768 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_259
timestamp 1679581782
transform 1 0 25440 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_266
timestamp 1679581782
transform 1 0 26112 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_273
timestamp 1679581782
transform 1 0 26784 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_280
timestamp 1679581782
transform 1 0 27456 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_287
timestamp 1679581782
transform 1 0 28128 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_294
timestamp 1679581782
transform 1 0 28800 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_301
timestamp 1679581782
transform 1 0 29472 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_308
timestamp 1679581782
transform 1 0 30144 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_315
timestamp 1679581782
transform 1 0 30816 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_322
timestamp 1679581782
transform 1 0 31488 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_329
timestamp 1679581782
transform 1 0 32160 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_336
timestamp 1679581782
transform 1 0 32832 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_343
timestamp 1679581782
transform 1 0 33504 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_350
timestamp 1679581782
transform 1 0 34176 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_357
timestamp 1679581782
transform 1 0 34848 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_364
timestamp 1679581782
transform 1 0 35520 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_371
timestamp 1679581782
transform 1 0 36192 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_378
timestamp 1679581782
transform 1 0 36864 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_385
timestamp 1679581782
transform 1 0 37536 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_392
timestamp 1679581782
transform 1 0 38208 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_399
timestamp 1679581782
transform 1 0 38880 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_406
timestamp 1679581782
transform 1 0 39552 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_413
timestamp 1679581782
transform 1 0 40224 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_420
timestamp 1679581782
transform 1 0 40896 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_427
timestamp 1679581782
transform 1 0 41568 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_434
timestamp 1679581782
transform 1 0 42240 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_441
timestamp 1679581782
transform 1 0 42912 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_448
timestamp 1679581782
transform 1 0 43584 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_455
timestamp 1679581782
transform 1 0 44256 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_462
timestamp 1679581782
transform 1 0 44928 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_469
timestamp 1679581782
transform 1 0 45600 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_476
timestamp 1679581782
transform 1 0 46272 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_483
timestamp 1679581782
transform 1 0 46944 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_490
timestamp 1679581782
transform 1 0 47616 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_497
timestamp 1679581782
transform 1 0 48288 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_504
timestamp 1679581782
transform 1 0 48960 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_511
timestamp 1679581782
transform 1 0 49632 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_518
timestamp 1679581782
transform 1 0 50304 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_525
timestamp 1679581782
transform 1 0 50976 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_532
timestamp 1679581782
transform 1 0 51648 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_539
timestamp 1679581782
transform 1 0 52320 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_546
timestamp 1679581782
transform 1 0 52992 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_553
timestamp 1679581782
transform 1 0 53664 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_560
timestamp 1679581782
transform 1 0 54336 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_567
timestamp 1679581782
transform 1 0 55008 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_574
timestamp 1679581782
transform 1 0 55680 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_581
timestamp 1679581782
transform 1 0 56352 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_588
timestamp 1679581782
transform 1 0 57024 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_595
timestamp 1679581782
transform 1 0 57696 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_602
timestamp 1679581782
transform 1 0 58368 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_609
timestamp 1679581782
transform 1 0 59040 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_616
timestamp 1679581782
transform 1 0 59712 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_623
timestamp 1679581782
transform 1 0 60384 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_630
timestamp 1679581782
transform 1 0 61056 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_637
timestamp 1679581782
transform 1 0 61728 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_644
timestamp 1679581782
transform 1 0 62400 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_651
timestamp 1679581782
transform 1 0 63072 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_658
timestamp 1679581782
transform 1 0 63744 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_665
timestamp 1679581782
transform 1 0 64416 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_672
timestamp 1679581782
transform 1 0 65088 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_679
timestamp 1679581782
transform 1 0 65760 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_686
timestamp 1679581782
transform 1 0 66432 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_693
timestamp 1679581782
transform 1 0 67104 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_700
timestamp 1679581782
transform 1 0 67776 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_707
timestamp 1679581782
transform 1 0 68448 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_714
timestamp 1679581782
transform 1 0 69120 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_721
timestamp 1679581782
transform 1 0 69792 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_728
timestamp 1679581782
transform 1 0 70464 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_735
timestamp 1679581782
transform 1 0 71136 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_742
timestamp 1679581782
transform 1 0 71808 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_749
timestamp 1679581782
transform 1 0 72480 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_756
timestamp 1679581782
transform 1 0 73152 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_763
timestamp 1679581782
transform 1 0 73824 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_770
timestamp 1679581782
transform 1 0 74496 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_777
timestamp 1679581782
transform 1 0 75168 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_784
timestamp 1679581782
transform 1 0 75840 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_791
timestamp 1679581782
transform 1 0 76512 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_798
timestamp 1679581782
transform 1 0 77184 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_805
timestamp 1679581782
transform 1 0 77856 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_812
timestamp 1679581782
transform 1 0 78528 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_819
timestamp 1679581782
transform 1 0 79200 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_826
timestamp 1679581782
transform 1 0 79872 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_833
timestamp 1679581782
transform 1 0 80544 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_840
timestamp 1679581782
transform 1 0 81216 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_847
timestamp 1679581782
transform 1 0 81888 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_854
timestamp 1679581782
transform 1 0 82560 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_861
timestamp 1679581782
transform 1 0 83232 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_868
timestamp 1679581782
transform 1 0 83904 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_875
timestamp 1679581782
transform 1 0 84576 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_882
timestamp 1679581782
transform 1 0 85248 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_889
timestamp 1679581782
transform 1 0 85920 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_896
timestamp 1679581782
transform 1 0 86592 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_903
timestamp 1679581782
transform 1 0 87264 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_910
timestamp 1679581782
transform 1 0 87936 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_917
timestamp 1679581782
transform 1 0 88608 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_17_924
timestamp 1677579658
transform 1 0 89280 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_4
timestamp 1679581782
transform 1 0 960 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_11
timestamp 1679581782
transform 1 0 1632 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_18
timestamp 1679581782
transform 1 0 2304 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_25
timestamp 1679581782
transform 1 0 2976 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_32
timestamp 1679581782
transform 1 0 3648 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_39
timestamp 1679581782
transform 1 0 4320 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_46
timestamp 1679581782
transform 1 0 4992 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_53
timestamp 1679581782
transform 1 0 5664 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_60
timestamp 1679581782
transform 1 0 6336 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_67
timestamp 1679581782
transform 1 0 7008 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_74
timestamp 1679581782
transform 1 0 7680 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_81
timestamp 1679581782
transform 1 0 8352 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_88
timestamp 1679581782
transform 1 0 9024 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_95
timestamp 1679581782
transform 1 0 9696 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_102
timestamp 1679581782
transform 1 0 10368 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_109
timestamp 1679581782
transform 1 0 11040 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_116
timestamp 1679581782
transform 1 0 11712 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_123
timestamp 1679581782
transform 1 0 12384 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_130
timestamp 1679581782
transform 1 0 13056 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_137
timestamp 1679581782
transform 1 0 13728 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_144
timestamp 1679581782
transform 1 0 14400 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_151
timestamp 1679581782
transform 1 0 15072 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_158
timestamp 1679581782
transform 1 0 15744 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_165
timestamp 1679581782
transform 1 0 16416 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_172
timestamp 1679581782
transform 1 0 17088 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_179
timestamp 1679581782
transform 1 0 17760 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_186
timestamp 1679581782
transform 1 0 18432 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_193
timestamp 1679581782
transform 1 0 19104 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_200
timestamp 1679581782
transform 1 0 19776 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_207
timestamp 1679581782
transform 1 0 20448 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_214
timestamp 1679581782
transform 1 0 21120 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_221
timestamp 1679581782
transform 1 0 21792 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_228
timestamp 1679581782
transform 1 0 22464 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_235
timestamp 1679581782
transform 1 0 23136 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_242
timestamp 1679581782
transform 1 0 23808 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_249
timestamp 1679581782
transform 1 0 24480 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_256
timestamp 1679581782
transform 1 0 25152 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_263
timestamp 1679581782
transform 1 0 25824 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_270
timestamp 1679581782
transform 1 0 26496 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_277
timestamp 1679581782
transform 1 0 27168 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_284
timestamp 1679581782
transform 1 0 27840 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_291
timestamp 1679581782
transform 1 0 28512 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_298
timestamp 1679581782
transform 1 0 29184 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_305
timestamp 1679581782
transform 1 0 29856 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_312
timestamp 1679581782
transform 1 0 30528 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_319
timestamp 1679581782
transform 1 0 31200 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_326
timestamp 1679581782
transform 1 0 31872 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_333
timestamp 1679581782
transform 1 0 32544 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_340
timestamp 1679581782
transform 1 0 33216 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_347
timestamp 1679581782
transform 1 0 33888 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_354
timestamp 1679581782
transform 1 0 34560 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_361
timestamp 1679581782
transform 1 0 35232 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_368
timestamp 1679581782
transform 1 0 35904 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_375
timestamp 1679581782
transform 1 0 36576 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_382
timestamp 1679581782
transform 1 0 37248 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_389
timestamp 1679581782
transform 1 0 37920 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_396
timestamp 1679581782
transform 1 0 38592 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_403
timestamp 1679581782
transform 1 0 39264 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_410
timestamp 1679581782
transform 1 0 39936 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_417
timestamp 1679581782
transform 1 0 40608 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_424
timestamp 1679581782
transform 1 0 41280 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_431
timestamp 1679581782
transform 1 0 41952 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_438
timestamp 1679581782
transform 1 0 42624 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_445
timestamp 1679581782
transform 1 0 43296 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_452
timestamp 1679581782
transform 1 0 43968 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_459
timestamp 1679581782
transform 1 0 44640 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_466
timestamp 1679581782
transform 1 0 45312 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_473
timestamp 1679581782
transform 1 0 45984 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_480
timestamp 1679581782
transform 1 0 46656 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_487
timestamp 1679581782
transform 1 0 47328 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_494
timestamp 1679581782
transform 1 0 48000 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_501
timestamp 1679581782
transform 1 0 48672 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_508
timestamp 1679581782
transform 1 0 49344 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_515
timestamp 1679581782
transform 1 0 50016 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_522
timestamp 1679581782
transform 1 0 50688 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_529
timestamp 1679581782
transform 1 0 51360 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_536
timestamp 1679581782
transform 1 0 52032 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_543
timestamp 1679581782
transform 1 0 52704 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_550
timestamp 1679581782
transform 1 0 53376 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_557
timestamp 1679581782
transform 1 0 54048 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_564
timestamp 1679581782
transform 1 0 54720 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_571
timestamp 1679581782
transform 1 0 55392 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_578
timestamp 1679581782
transform 1 0 56064 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_585
timestamp 1679581782
transform 1 0 56736 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_592
timestamp 1679581782
transform 1 0 57408 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_599
timestamp 1679581782
transform 1 0 58080 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_606
timestamp 1679581782
transform 1 0 58752 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_613
timestamp 1679581782
transform 1 0 59424 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_620
timestamp 1679581782
transform 1 0 60096 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_627
timestamp 1679581782
transform 1 0 60768 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_634
timestamp 1679581782
transform 1 0 61440 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_641
timestamp 1679581782
transform 1 0 62112 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_648
timestamp 1679581782
transform 1 0 62784 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_655
timestamp 1679581782
transform 1 0 63456 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_662
timestamp 1679581782
transform 1 0 64128 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_669
timestamp 1679581782
transform 1 0 64800 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_676
timestamp 1679581782
transform 1 0 65472 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_683
timestamp 1679581782
transform 1 0 66144 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_690
timestamp 1679581782
transform 1 0 66816 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_697
timestamp 1679581782
transform 1 0 67488 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_704
timestamp 1679581782
transform 1 0 68160 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_711
timestamp 1679581782
transform 1 0 68832 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_718
timestamp 1679581782
transform 1 0 69504 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_725
timestamp 1679581782
transform 1 0 70176 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_732
timestamp 1679581782
transform 1 0 70848 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_739
timestamp 1679581782
transform 1 0 71520 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_746
timestamp 1679581782
transform 1 0 72192 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_753
timestamp 1679581782
transform 1 0 72864 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_760
timestamp 1679581782
transform 1 0 73536 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_767
timestamp 1679581782
transform 1 0 74208 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_774
timestamp 1679581782
transform 1 0 74880 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_781
timestamp 1679581782
transform 1 0 75552 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_788
timestamp 1679581782
transform 1 0 76224 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_795
timestamp 1679581782
transform 1 0 76896 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_802
timestamp 1679581782
transform 1 0 77568 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_809
timestamp 1679581782
transform 1 0 78240 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_816
timestamp 1679581782
transform 1 0 78912 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_823
timestamp 1679581782
transform 1 0 79584 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_830
timestamp 1679581782
transform 1 0 80256 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_837
timestamp 1679581782
transform 1 0 80928 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_844
timestamp 1679581782
transform 1 0 81600 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_851
timestamp 1679581782
transform 1 0 82272 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_858
timestamp 1679581782
transform 1 0 82944 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_865
timestamp 1679581782
transform 1 0 83616 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_872
timestamp 1679581782
transform 1 0 84288 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_879
timestamp 1679581782
transform 1 0 84960 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_886
timestamp 1679581782
transform 1 0 85632 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_893
timestamp 1679581782
transform 1 0 86304 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_900
timestamp 1679581782
transform 1 0 86976 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_907
timestamp 1679581782
transform 1 0 87648 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_914
timestamp 1679581782
transform 1 0 88320 0 1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_18_921
timestamp 1679577901
transform 1 0 88992 0 1 14364
box -48 -56 432 834
use sg13g2_decap_8  FILLER_19_4
timestamp 1679581782
transform 1 0 960 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_11
timestamp 1679581782
transform 1 0 1632 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_18
timestamp 1679581782
transform 1 0 2304 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_25
timestamp 1679581782
transform 1 0 2976 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_32
timestamp 1679581782
transform 1 0 3648 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_39
timestamp 1679581782
transform 1 0 4320 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_46
timestamp 1679581782
transform 1 0 4992 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_53
timestamp 1679581782
transform 1 0 5664 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_60
timestamp 1679581782
transform 1 0 6336 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_67
timestamp 1679581782
transform 1 0 7008 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_74
timestamp 1679581782
transform 1 0 7680 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_81
timestamp 1679581782
transform 1 0 8352 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_88
timestamp 1679581782
transform 1 0 9024 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_95
timestamp 1679581782
transform 1 0 9696 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_102
timestamp 1679581782
transform 1 0 10368 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_109
timestamp 1679581782
transform 1 0 11040 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_116
timestamp 1679581782
transform 1 0 11712 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_123
timestamp 1679581782
transform 1 0 12384 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_130
timestamp 1679581782
transform 1 0 13056 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_137
timestamp 1679581782
transform 1 0 13728 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_144
timestamp 1679581782
transform 1 0 14400 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_151
timestamp 1679581782
transform 1 0 15072 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_158
timestamp 1679581782
transform 1 0 15744 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_165
timestamp 1679581782
transform 1 0 16416 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_172
timestamp 1679581782
transform 1 0 17088 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_179
timestamp 1679581782
transform 1 0 17760 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_186
timestamp 1679581782
transform 1 0 18432 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_193
timestamp 1679581782
transform 1 0 19104 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_200
timestamp 1679581782
transform 1 0 19776 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_207
timestamp 1679581782
transform 1 0 20448 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_214
timestamp 1679581782
transform 1 0 21120 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_221
timestamp 1679581782
transform 1 0 21792 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_228
timestamp 1679581782
transform 1 0 22464 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_235
timestamp 1679581782
transform 1 0 23136 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_242
timestamp 1679581782
transform 1 0 23808 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_249
timestamp 1679581782
transform 1 0 24480 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_256
timestamp 1679581782
transform 1 0 25152 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_263
timestamp 1679581782
transform 1 0 25824 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_270
timestamp 1679581782
transform 1 0 26496 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_277
timestamp 1679581782
transform 1 0 27168 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_284
timestamp 1679581782
transform 1 0 27840 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_291
timestamp 1679581782
transform 1 0 28512 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_298
timestamp 1679581782
transform 1 0 29184 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_305
timestamp 1679581782
transform 1 0 29856 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_312
timestamp 1679581782
transform 1 0 30528 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_319
timestamp 1679581782
transform 1 0 31200 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_326
timestamp 1679581782
transform 1 0 31872 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_333
timestamp 1679581782
transform 1 0 32544 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_340
timestamp 1679581782
transform 1 0 33216 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_347
timestamp 1679581782
transform 1 0 33888 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_354
timestamp 1679581782
transform 1 0 34560 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_361
timestamp 1679581782
transform 1 0 35232 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_368
timestamp 1679581782
transform 1 0 35904 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_375
timestamp 1679581782
transform 1 0 36576 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_382
timestamp 1679581782
transform 1 0 37248 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_389
timestamp 1679581782
transform 1 0 37920 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_396
timestamp 1679581782
transform 1 0 38592 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_403
timestamp 1679581782
transform 1 0 39264 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_410
timestamp 1679581782
transform 1 0 39936 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_417
timestamp 1679581782
transform 1 0 40608 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_424
timestamp 1679581782
transform 1 0 41280 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_431
timestamp 1679581782
transform 1 0 41952 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_438
timestamp 1679581782
transform 1 0 42624 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_445
timestamp 1679581782
transform 1 0 43296 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_452
timestamp 1679581782
transform 1 0 43968 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_459
timestamp 1679581782
transform 1 0 44640 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_466
timestamp 1679581782
transform 1 0 45312 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_473
timestamp 1679581782
transform 1 0 45984 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_480
timestamp 1679581782
transform 1 0 46656 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_487
timestamp 1679581782
transform 1 0 47328 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_494
timestamp 1679581782
transform 1 0 48000 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_501
timestamp 1679581782
transform 1 0 48672 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_508
timestamp 1679581782
transform 1 0 49344 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_515
timestamp 1679581782
transform 1 0 50016 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_522
timestamp 1679581782
transform 1 0 50688 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_529
timestamp 1679581782
transform 1 0 51360 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_536
timestamp 1679581782
transform 1 0 52032 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_543
timestamp 1679581782
transform 1 0 52704 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_550
timestamp 1679581782
transform 1 0 53376 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_557
timestamp 1679581782
transform 1 0 54048 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_564
timestamp 1679581782
transform 1 0 54720 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_571
timestamp 1679581782
transform 1 0 55392 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_578
timestamp 1679581782
transform 1 0 56064 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_585
timestamp 1679581782
transform 1 0 56736 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_592
timestamp 1679581782
transform 1 0 57408 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_599
timestamp 1679581782
transform 1 0 58080 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_606
timestamp 1679581782
transform 1 0 58752 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_613
timestamp 1679581782
transform 1 0 59424 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_620
timestamp 1679581782
transform 1 0 60096 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_627
timestamp 1679581782
transform 1 0 60768 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_634
timestamp 1679581782
transform 1 0 61440 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_641
timestamp 1679581782
transform 1 0 62112 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_648
timestamp 1679581782
transform 1 0 62784 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_655
timestamp 1679581782
transform 1 0 63456 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_662
timestamp 1679581782
transform 1 0 64128 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_669
timestamp 1679581782
transform 1 0 64800 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_676
timestamp 1679581782
transform 1 0 65472 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_683
timestamp 1679581782
transform 1 0 66144 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_690
timestamp 1679581782
transform 1 0 66816 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_697
timestamp 1679581782
transform 1 0 67488 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_704
timestamp 1679581782
transform 1 0 68160 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_711
timestamp 1679581782
transform 1 0 68832 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_718
timestamp 1679581782
transform 1 0 69504 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_725
timestamp 1679581782
transform 1 0 70176 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_732
timestamp 1679581782
transform 1 0 70848 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_739
timestamp 1679581782
transform 1 0 71520 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_746
timestamp 1679581782
transform 1 0 72192 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_753
timestamp 1679581782
transform 1 0 72864 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_760
timestamp 1679581782
transform 1 0 73536 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_767
timestamp 1679581782
transform 1 0 74208 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_774
timestamp 1679581782
transform 1 0 74880 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_781
timestamp 1679581782
transform 1 0 75552 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_788
timestamp 1679581782
transform 1 0 76224 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_795
timestamp 1679581782
transform 1 0 76896 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_802
timestamp 1679581782
transform 1 0 77568 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_809
timestamp 1679581782
transform 1 0 78240 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_816
timestamp 1679581782
transform 1 0 78912 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_823
timestamp 1679581782
transform 1 0 79584 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_830
timestamp 1679581782
transform 1 0 80256 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_837
timestamp 1679581782
transform 1 0 80928 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_844
timestamp 1679581782
transform 1 0 81600 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_851
timestamp 1679581782
transform 1 0 82272 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_858
timestamp 1679581782
transform 1 0 82944 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_865
timestamp 1679581782
transform 1 0 83616 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_872
timestamp 1679581782
transform 1 0 84288 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_879
timestamp 1679581782
transform 1 0 84960 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_886
timestamp 1679581782
transform 1 0 85632 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_893
timestamp 1679581782
transform 1 0 86304 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_900
timestamp 1679581782
transform 1 0 86976 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_907
timestamp 1679581782
transform 1 0 87648 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_914
timestamp 1679581782
transform 1 0 88320 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_19_921
timestamp 1679577901
transform 1 0 88992 0 -1 15876
box -48 -56 432 834
use sg13g2_decap_8  FILLER_20_4
timestamp 1679581782
transform 1 0 960 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_11
timestamp 1679581782
transform 1 0 1632 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_18
timestamp 1679581782
transform 1 0 2304 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_25
timestamp 1679581782
transform 1 0 2976 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_32
timestamp 1679581782
transform 1 0 3648 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_39
timestamp 1679581782
transform 1 0 4320 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_46
timestamp 1679581782
transform 1 0 4992 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_53
timestamp 1679581782
transform 1 0 5664 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_60
timestamp 1679581782
transform 1 0 6336 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_67
timestamp 1679581782
transform 1 0 7008 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_74
timestamp 1679581782
transform 1 0 7680 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_81
timestamp 1679581782
transform 1 0 8352 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_88
timestamp 1679581782
transform 1 0 9024 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_95
timestamp 1679581782
transform 1 0 9696 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_102
timestamp 1679581782
transform 1 0 10368 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_109
timestamp 1679581782
transform 1 0 11040 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_116
timestamp 1679581782
transform 1 0 11712 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_123
timestamp 1679581782
transform 1 0 12384 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_130
timestamp 1679581782
transform 1 0 13056 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_137
timestamp 1679581782
transform 1 0 13728 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_144
timestamp 1679581782
transform 1 0 14400 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_151
timestamp 1679581782
transform 1 0 15072 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_158
timestamp 1679581782
transform 1 0 15744 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_165
timestamp 1679581782
transform 1 0 16416 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_172
timestamp 1679581782
transform 1 0 17088 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_179
timestamp 1679581782
transform 1 0 17760 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_186
timestamp 1679581782
transform 1 0 18432 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_193
timestamp 1679581782
transform 1 0 19104 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_200
timestamp 1679581782
transform 1 0 19776 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_207
timestamp 1679581782
transform 1 0 20448 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_214
timestamp 1679581782
transform 1 0 21120 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_221
timestamp 1679581782
transform 1 0 21792 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_228
timestamp 1679581782
transform 1 0 22464 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_235
timestamp 1679581782
transform 1 0 23136 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_242
timestamp 1679581782
transform 1 0 23808 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_249
timestamp 1679581782
transform 1 0 24480 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_256
timestamp 1679581782
transform 1 0 25152 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_263
timestamp 1679581782
transform 1 0 25824 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_270
timestamp 1679581782
transform 1 0 26496 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_277
timestamp 1679581782
transform 1 0 27168 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_284
timestamp 1679581782
transform 1 0 27840 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_291
timestamp 1679581782
transform 1 0 28512 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_298
timestamp 1679581782
transform 1 0 29184 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_305
timestamp 1679581782
transform 1 0 29856 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_312
timestamp 1679581782
transform 1 0 30528 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_319
timestamp 1679581782
transform 1 0 31200 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_326
timestamp 1679581782
transform 1 0 31872 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_333
timestamp 1679581782
transform 1 0 32544 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_340
timestamp 1679581782
transform 1 0 33216 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_347
timestamp 1679581782
transform 1 0 33888 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_354
timestamp 1679581782
transform 1 0 34560 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_361
timestamp 1679581782
transform 1 0 35232 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_368
timestamp 1679581782
transform 1 0 35904 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_375
timestamp 1679581782
transform 1 0 36576 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_382
timestamp 1679581782
transform 1 0 37248 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_389
timestamp 1679581782
transform 1 0 37920 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_396
timestamp 1679581782
transform 1 0 38592 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_403
timestamp 1679581782
transform 1 0 39264 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_410
timestamp 1679581782
transform 1 0 39936 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_417
timestamp 1679581782
transform 1 0 40608 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_424
timestamp 1679581782
transform 1 0 41280 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_431
timestamp 1679581782
transform 1 0 41952 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_438
timestamp 1679581782
transform 1 0 42624 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_445
timestamp 1679581782
transform 1 0 43296 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_452
timestamp 1679581782
transform 1 0 43968 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_459
timestamp 1679581782
transform 1 0 44640 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_466
timestamp 1679581782
transform 1 0 45312 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_473
timestamp 1679581782
transform 1 0 45984 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_480
timestamp 1679581782
transform 1 0 46656 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_487
timestamp 1679581782
transform 1 0 47328 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_494
timestamp 1679581782
transform 1 0 48000 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_501
timestamp 1679581782
transform 1 0 48672 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_508
timestamp 1679581782
transform 1 0 49344 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_515
timestamp 1679581782
transform 1 0 50016 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_522
timestamp 1679581782
transform 1 0 50688 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_529
timestamp 1679581782
transform 1 0 51360 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_536
timestamp 1679581782
transform 1 0 52032 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_543
timestamp 1679581782
transform 1 0 52704 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_550
timestamp 1679581782
transform 1 0 53376 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_557
timestamp 1679581782
transform 1 0 54048 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_564
timestamp 1679581782
transform 1 0 54720 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_571
timestamp 1679581782
transform 1 0 55392 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_578
timestamp 1679581782
transform 1 0 56064 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_585
timestamp 1679581782
transform 1 0 56736 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_592
timestamp 1679581782
transform 1 0 57408 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_599
timestamp 1679581782
transform 1 0 58080 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_606
timestamp 1679581782
transform 1 0 58752 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_613
timestamp 1679581782
transform 1 0 59424 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_620
timestamp 1679581782
transform 1 0 60096 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_627
timestamp 1679581782
transform 1 0 60768 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_634
timestamp 1679581782
transform 1 0 61440 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_641
timestamp 1679581782
transform 1 0 62112 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_648
timestamp 1679581782
transform 1 0 62784 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_655
timestamp 1679581782
transform 1 0 63456 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_662
timestamp 1679581782
transform 1 0 64128 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_669
timestamp 1679581782
transform 1 0 64800 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_676
timestamp 1679581782
transform 1 0 65472 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_683
timestamp 1679581782
transform 1 0 66144 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_690
timestamp 1679581782
transform 1 0 66816 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_697
timestamp 1679581782
transform 1 0 67488 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_704
timestamp 1679581782
transform 1 0 68160 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_711
timestamp 1679581782
transform 1 0 68832 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_718
timestamp 1679581782
transform 1 0 69504 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_725
timestamp 1679581782
transform 1 0 70176 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_732
timestamp 1679581782
transform 1 0 70848 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_739
timestamp 1679581782
transform 1 0 71520 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_746
timestamp 1679581782
transform 1 0 72192 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_753
timestamp 1679581782
transform 1 0 72864 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_760
timestamp 1679581782
transform 1 0 73536 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_767
timestamp 1679581782
transform 1 0 74208 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_774
timestamp 1679581782
transform 1 0 74880 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_781
timestamp 1679581782
transform 1 0 75552 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_788
timestamp 1679581782
transform 1 0 76224 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_795
timestamp 1679581782
transform 1 0 76896 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_802
timestamp 1679581782
transform 1 0 77568 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_809
timestamp 1679581782
transform 1 0 78240 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_816
timestamp 1679581782
transform 1 0 78912 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_823
timestamp 1679581782
transform 1 0 79584 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_830
timestamp 1679581782
transform 1 0 80256 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_837
timestamp 1679581782
transform 1 0 80928 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_844
timestamp 1679581782
transform 1 0 81600 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_851
timestamp 1679581782
transform 1 0 82272 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_858
timestamp 1679581782
transform 1 0 82944 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_865
timestamp 1679581782
transform 1 0 83616 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_872
timestamp 1679581782
transform 1 0 84288 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_879
timestamp 1679581782
transform 1 0 84960 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_886
timestamp 1679581782
transform 1 0 85632 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_893
timestamp 1679581782
transform 1 0 86304 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_900
timestamp 1679581782
transform 1 0 86976 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_907
timestamp 1679581782
transform 1 0 87648 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_914
timestamp 1679581782
transform 1 0 88320 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_921
timestamp 1679577901
transform 1 0 88992 0 1 15876
box -48 -56 432 834
use sg13g2_decap_8  FILLER_21_4
timestamp 1679581782
transform 1 0 960 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_11
timestamp 1679581782
transform 1 0 1632 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_18
timestamp 1679581782
transform 1 0 2304 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_25
timestamp 1679581782
transform 1 0 2976 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_32
timestamp 1679581782
transform 1 0 3648 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_39
timestamp 1679581782
transform 1 0 4320 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_46
timestamp 1679581782
transform 1 0 4992 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_53
timestamp 1679581782
transform 1 0 5664 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_60
timestamp 1679581782
transform 1 0 6336 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_67
timestamp 1679581782
transform 1 0 7008 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_74
timestamp 1679581782
transform 1 0 7680 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_81
timestamp 1679581782
transform 1 0 8352 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_88
timestamp 1679581782
transform 1 0 9024 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_95
timestamp 1679581782
transform 1 0 9696 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_102
timestamp 1679581782
transform 1 0 10368 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_109
timestamp 1679581782
transform 1 0 11040 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_116
timestamp 1679581782
transform 1 0 11712 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_123
timestamp 1679581782
transform 1 0 12384 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_130
timestamp 1679581782
transform 1 0 13056 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_137
timestamp 1679581782
transform 1 0 13728 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_144
timestamp 1679581782
transform 1 0 14400 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_151
timestamp 1679581782
transform 1 0 15072 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_158
timestamp 1679581782
transform 1 0 15744 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_165
timestamp 1679581782
transform 1 0 16416 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_172
timestamp 1679581782
transform 1 0 17088 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_179
timestamp 1679581782
transform 1 0 17760 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_186
timestamp 1679581782
transform 1 0 18432 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_193
timestamp 1679581782
transform 1 0 19104 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_200
timestamp 1679581782
transform 1 0 19776 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_207
timestamp 1679581782
transform 1 0 20448 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_214
timestamp 1679581782
transform 1 0 21120 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_221
timestamp 1679581782
transform 1 0 21792 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_228
timestamp 1679581782
transform 1 0 22464 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_235
timestamp 1679581782
transform 1 0 23136 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_242
timestamp 1679581782
transform 1 0 23808 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_249
timestamp 1679581782
transform 1 0 24480 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_256
timestamp 1679581782
transform 1 0 25152 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_263
timestamp 1679581782
transform 1 0 25824 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_270
timestamp 1679581782
transform 1 0 26496 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_277
timestamp 1679581782
transform 1 0 27168 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_284
timestamp 1679581782
transform 1 0 27840 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_291
timestamp 1679581782
transform 1 0 28512 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_298
timestamp 1679581782
transform 1 0 29184 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_305
timestamp 1679581782
transform 1 0 29856 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_312
timestamp 1679581782
transform 1 0 30528 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_319
timestamp 1679581782
transform 1 0 31200 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_326
timestamp 1679581782
transform 1 0 31872 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_333
timestamp 1679581782
transform 1 0 32544 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_340
timestamp 1679581782
transform 1 0 33216 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_347
timestamp 1679581782
transform 1 0 33888 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_354
timestamp 1679581782
transform 1 0 34560 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_361
timestamp 1679581782
transform 1 0 35232 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_368
timestamp 1679581782
transform 1 0 35904 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_375
timestamp 1679581782
transform 1 0 36576 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_382
timestamp 1679581782
transform 1 0 37248 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_389
timestamp 1679581782
transform 1 0 37920 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_396
timestamp 1679581782
transform 1 0 38592 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_403
timestamp 1679581782
transform 1 0 39264 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_410
timestamp 1679581782
transform 1 0 39936 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_417
timestamp 1679581782
transform 1 0 40608 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_424
timestamp 1679581782
transform 1 0 41280 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_431
timestamp 1679581782
transform 1 0 41952 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_438
timestamp 1679581782
transform 1 0 42624 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_445
timestamp 1679581782
transform 1 0 43296 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_452
timestamp 1679581782
transform 1 0 43968 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_459
timestamp 1679581782
transform 1 0 44640 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_466
timestamp 1679581782
transform 1 0 45312 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_473
timestamp 1679581782
transform 1 0 45984 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_480
timestamp 1679581782
transform 1 0 46656 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_487
timestamp 1679581782
transform 1 0 47328 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_494
timestamp 1679581782
transform 1 0 48000 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_501
timestamp 1679581782
transform 1 0 48672 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_508
timestamp 1679581782
transform 1 0 49344 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_515
timestamp 1679581782
transform 1 0 50016 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_522
timestamp 1679581782
transform 1 0 50688 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_529
timestamp 1679581782
transform 1 0 51360 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_536
timestamp 1679581782
transform 1 0 52032 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_543
timestamp 1679581782
transform 1 0 52704 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_550
timestamp 1679581782
transform 1 0 53376 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_557
timestamp 1679581782
transform 1 0 54048 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_564
timestamp 1679581782
transform 1 0 54720 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_571
timestamp 1679581782
transform 1 0 55392 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_578
timestamp 1679581782
transform 1 0 56064 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_585
timestamp 1679581782
transform 1 0 56736 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_592
timestamp 1679581782
transform 1 0 57408 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_599
timestamp 1679581782
transform 1 0 58080 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_606
timestamp 1679581782
transform 1 0 58752 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_613
timestamp 1679581782
transform 1 0 59424 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_620
timestamp 1679581782
transform 1 0 60096 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_627
timestamp 1679581782
transform 1 0 60768 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_634
timestamp 1679581782
transform 1 0 61440 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_641
timestamp 1679581782
transform 1 0 62112 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_648
timestamp 1679581782
transform 1 0 62784 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_655
timestamp 1679581782
transform 1 0 63456 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_662
timestamp 1679581782
transform 1 0 64128 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_669
timestamp 1679581782
transform 1 0 64800 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_676
timestamp 1679581782
transform 1 0 65472 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_683
timestamp 1679581782
transform 1 0 66144 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_690
timestamp 1679581782
transform 1 0 66816 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_697
timestamp 1679581782
transform 1 0 67488 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_704
timestamp 1679581782
transform 1 0 68160 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_711
timestamp 1679581782
transform 1 0 68832 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_718
timestamp 1679581782
transform 1 0 69504 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_725
timestamp 1679581782
transform 1 0 70176 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_732
timestamp 1679581782
transform 1 0 70848 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_739
timestamp 1679581782
transform 1 0 71520 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_746
timestamp 1679581782
transform 1 0 72192 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_753
timestamp 1679581782
transform 1 0 72864 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_760
timestamp 1679581782
transform 1 0 73536 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_767
timestamp 1679581782
transform 1 0 74208 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_774
timestamp 1679581782
transform 1 0 74880 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_781
timestamp 1679581782
transform 1 0 75552 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_788
timestamp 1679581782
transform 1 0 76224 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_795
timestamp 1679581782
transform 1 0 76896 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_802
timestamp 1679581782
transform 1 0 77568 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_809
timestamp 1679581782
transform 1 0 78240 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_816
timestamp 1679581782
transform 1 0 78912 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_823
timestamp 1679581782
transform 1 0 79584 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_830
timestamp 1679581782
transform 1 0 80256 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_837
timestamp 1679581782
transform 1 0 80928 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_844
timestamp 1679581782
transform 1 0 81600 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_851
timestamp 1679581782
transform 1 0 82272 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_858
timestamp 1679581782
transform 1 0 82944 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_865
timestamp 1679581782
transform 1 0 83616 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_872
timestamp 1679581782
transform 1 0 84288 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_879
timestamp 1679581782
transform 1 0 84960 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_886
timestamp 1679581782
transform 1 0 85632 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_893
timestamp 1679581782
transform 1 0 86304 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_900
timestamp 1679581782
transform 1 0 86976 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_907
timestamp 1679581782
transform 1 0 87648 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_914
timestamp 1679581782
transform 1 0 88320 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_921
timestamp 1679577901
transform 1 0 88992 0 -1 17388
box -48 -56 432 834
use sg13g2_decap_8  FILLER_22_4
timestamp 1679581782
transform 1 0 960 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_11
timestamp 1679581782
transform 1 0 1632 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_18
timestamp 1679581782
transform 1 0 2304 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_25
timestamp 1679581782
transform 1 0 2976 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_32
timestamp 1679581782
transform 1 0 3648 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_39
timestamp 1679581782
transform 1 0 4320 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_46
timestamp 1679581782
transform 1 0 4992 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_53
timestamp 1679581782
transform 1 0 5664 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_60
timestamp 1679581782
transform 1 0 6336 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_67
timestamp 1679581782
transform 1 0 7008 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_74
timestamp 1679581782
transform 1 0 7680 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_81
timestamp 1679581782
transform 1 0 8352 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_88
timestamp 1679581782
transform 1 0 9024 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_95
timestamp 1679581782
transform 1 0 9696 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_102
timestamp 1679581782
transform 1 0 10368 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_109
timestamp 1679581782
transform 1 0 11040 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_116
timestamp 1679581782
transform 1 0 11712 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_123
timestamp 1679581782
transform 1 0 12384 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_130
timestamp 1679581782
transform 1 0 13056 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_137
timestamp 1679581782
transform 1 0 13728 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_144
timestamp 1679581782
transform 1 0 14400 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_151
timestamp 1679581782
transform 1 0 15072 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_158
timestamp 1679581782
transform 1 0 15744 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_165
timestamp 1679581782
transform 1 0 16416 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_172
timestamp 1679581782
transform 1 0 17088 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_179
timestamp 1679581782
transform 1 0 17760 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_186
timestamp 1679581782
transform 1 0 18432 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_193
timestamp 1679581782
transform 1 0 19104 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_200
timestamp 1679581782
transform 1 0 19776 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_207
timestamp 1679581782
transform 1 0 20448 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_214
timestamp 1679581782
transform 1 0 21120 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_221
timestamp 1679581782
transform 1 0 21792 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_228
timestamp 1679581782
transform 1 0 22464 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_235
timestamp 1679581782
transform 1 0 23136 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_242
timestamp 1679581782
transform 1 0 23808 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_249
timestamp 1679581782
transform 1 0 24480 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_256
timestamp 1679581782
transform 1 0 25152 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_263
timestamp 1679581782
transform 1 0 25824 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_270
timestamp 1679581782
transform 1 0 26496 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_277
timestamp 1679581782
transform 1 0 27168 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_284
timestamp 1679581782
transform 1 0 27840 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_291
timestamp 1679581782
transform 1 0 28512 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_298
timestamp 1679581782
transform 1 0 29184 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_305
timestamp 1679581782
transform 1 0 29856 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_312
timestamp 1679581782
transform 1 0 30528 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_319
timestamp 1679581782
transform 1 0 31200 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_326
timestamp 1679581782
transform 1 0 31872 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_333
timestamp 1679581782
transform 1 0 32544 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_340
timestamp 1679581782
transform 1 0 33216 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_347
timestamp 1679581782
transform 1 0 33888 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_354
timestamp 1679581782
transform 1 0 34560 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_361
timestamp 1679581782
transform 1 0 35232 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_368
timestamp 1679581782
transform 1 0 35904 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_375
timestamp 1679581782
transform 1 0 36576 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_382
timestamp 1679581782
transform 1 0 37248 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_389
timestamp 1679581782
transform 1 0 37920 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_396
timestamp 1679581782
transform 1 0 38592 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_403
timestamp 1679581782
transform 1 0 39264 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_410
timestamp 1679581782
transform 1 0 39936 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_417
timestamp 1679581782
transform 1 0 40608 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_424
timestamp 1679581782
transform 1 0 41280 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_431
timestamp 1679581782
transform 1 0 41952 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_438
timestamp 1679581782
transform 1 0 42624 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_445
timestamp 1679581782
transform 1 0 43296 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_452
timestamp 1679581782
transform 1 0 43968 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_459
timestamp 1679581782
transform 1 0 44640 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_466
timestamp 1679581782
transform 1 0 45312 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_473
timestamp 1679581782
transform 1 0 45984 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_480
timestamp 1679581782
transform 1 0 46656 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_487
timestamp 1679581782
transform 1 0 47328 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_494
timestamp 1679581782
transform 1 0 48000 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_501
timestamp 1679581782
transform 1 0 48672 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_508
timestamp 1679581782
transform 1 0 49344 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_515
timestamp 1679581782
transform 1 0 50016 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_522
timestamp 1679581782
transform 1 0 50688 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_529
timestamp 1679581782
transform 1 0 51360 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_536
timestamp 1679581782
transform 1 0 52032 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_543
timestamp 1679581782
transform 1 0 52704 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_550
timestamp 1679581782
transform 1 0 53376 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_557
timestamp 1679581782
transform 1 0 54048 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_564
timestamp 1679581782
transform 1 0 54720 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_571
timestamp 1679581782
transform 1 0 55392 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_578
timestamp 1679581782
transform 1 0 56064 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_585
timestamp 1679581782
transform 1 0 56736 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_592
timestamp 1679581782
transform 1 0 57408 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_599
timestamp 1679581782
transform 1 0 58080 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_606
timestamp 1679581782
transform 1 0 58752 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_613
timestamp 1679581782
transform 1 0 59424 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_620
timestamp 1679581782
transform 1 0 60096 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_627
timestamp 1679581782
transform 1 0 60768 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_634
timestamp 1679581782
transform 1 0 61440 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_641
timestamp 1679581782
transform 1 0 62112 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_648
timestamp 1679581782
transform 1 0 62784 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_655
timestamp 1679581782
transform 1 0 63456 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_662
timestamp 1679581782
transform 1 0 64128 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_669
timestamp 1679581782
transform 1 0 64800 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_676
timestamp 1679581782
transform 1 0 65472 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_683
timestamp 1679581782
transform 1 0 66144 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_690
timestamp 1679581782
transform 1 0 66816 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_697
timestamp 1679581782
transform 1 0 67488 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_704
timestamp 1679581782
transform 1 0 68160 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_711
timestamp 1679581782
transform 1 0 68832 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_718
timestamp 1679581782
transform 1 0 69504 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_725
timestamp 1679581782
transform 1 0 70176 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_732
timestamp 1679581782
transform 1 0 70848 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_739
timestamp 1679581782
transform 1 0 71520 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_746
timestamp 1679581782
transform 1 0 72192 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_753
timestamp 1679581782
transform 1 0 72864 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_760
timestamp 1679581782
transform 1 0 73536 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_767
timestamp 1679581782
transform 1 0 74208 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_774
timestamp 1679581782
transform 1 0 74880 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_781
timestamp 1679581782
transform 1 0 75552 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_788
timestamp 1679581782
transform 1 0 76224 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_795
timestamp 1679581782
transform 1 0 76896 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_802
timestamp 1679581782
transform 1 0 77568 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_809
timestamp 1679581782
transform 1 0 78240 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_816
timestamp 1679581782
transform 1 0 78912 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_823
timestamp 1679581782
transform 1 0 79584 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_830
timestamp 1679581782
transform 1 0 80256 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_837
timestamp 1679581782
transform 1 0 80928 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_844
timestamp 1679581782
transform 1 0 81600 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_851
timestamp 1679581782
transform 1 0 82272 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_858
timestamp 1679581782
transform 1 0 82944 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_865
timestamp 1679581782
transform 1 0 83616 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_872
timestamp 1679581782
transform 1 0 84288 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_879
timestamp 1679581782
transform 1 0 84960 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_886
timestamp 1679581782
transform 1 0 85632 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_893
timestamp 1679581782
transform 1 0 86304 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_900
timestamp 1679581782
transform 1 0 86976 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_907
timestamp 1679581782
transform 1 0 87648 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_914
timestamp 1679581782
transform 1 0 88320 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_921
timestamp 1679577901
transform 1 0 88992 0 1 17388
box -48 -56 432 834
use sg13g2_decap_8  FILLER_23_4
timestamp 1679581782
transform 1 0 960 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_11
timestamp 1679581782
transform 1 0 1632 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_18
timestamp 1679581782
transform 1 0 2304 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_25
timestamp 1679581782
transform 1 0 2976 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_32
timestamp 1679581782
transform 1 0 3648 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_39
timestamp 1679581782
transform 1 0 4320 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_46
timestamp 1679581782
transform 1 0 4992 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_53
timestamp 1679581782
transform 1 0 5664 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_60
timestamp 1679581782
transform 1 0 6336 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_67
timestamp 1679581782
transform 1 0 7008 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_74
timestamp 1679581782
transform 1 0 7680 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_81
timestamp 1679581782
transform 1 0 8352 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_88
timestamp 1679581782
transform 1 0 9024 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_95
timestamp 1679581782
transform 1 0 9696 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_102
timestamp 1679581782
transform 1 0 10368 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_109
timestamp 1679581782
transform 1 0 11040 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_116
timestamp 1679581782
transform 1 0 11712 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_123
timestamp 1679581782
transform 1 0 12384 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_130
timestamp 1679581782
transform 1 0 13056 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_137
timestamp 1679581782
transform 1 0 13728 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_144
timestamp 1679581782
transform 1 0 14400 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_151
timestamp 1679581782
transform 1 0 15072 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_158
timestamp 1679581782
transform 1 0 15744 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_165
timestamp 1679581782
transform 1 0 16416 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_172
timestamp 1679581782
transform 1 0 17088 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_179
timestamp 1679581782
transform 1 0 17760 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_186
timestamp 1679581782
transform 1 0 18432 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_193
timestamp 1679581782
transform 1 0 19104 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_200
timestamp 1679581782
transform 1 0 19776 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_207
timestamp 1679581782
transform 1 0 20448 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_214
timestamp 1679581782
transform 1 0 21120 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_221
timestamp 1679581782
transform 1 0 21792 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_228
timestamp 1679581782
transform 1 0 22464 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_235
timestamp 1679581782
transform 1 0 23136 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_242
timestamp 1679581782
transform 1 0 23808 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_249
timestamp 1679581782
transform 1 0 24480 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_256
timestamp 1679581782
transform 1 0 25152 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_263
timestamp 1679581782
transform 1 0 25824 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_270
timestamp 1679581782
transform 1 0 26496 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_277
timestamp 1679581782
transform 1 0 27168 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_284
timestamp 1679581782
transform 1 0 27840 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_291
timestamp 1679581782
transform 1 0 28512 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_298
timestamp 1679581782
transform 1 0 29184 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_305
timestamp 1679581782
transform 1 0 29856 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_312
timestamp 1679581782
transform 1 0 30528 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_319
timestamp 1679581782
transform 1 0 31200 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_326
timestamp 1679581782
transform 1 0 31872 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_333
timestamp 1679581782
transform 1 0 32544 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_340
timestamp 1679581782
transform 1 0 33216 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_347
timestamp 1679581782
transform 1 0 33888 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_354
timestamp 1679581782
transform 1 0 34560 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_361
timestamp 1679581782
transform 1 0 35232 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_368
timestamp 1679581782
transform 1 0 35904 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_375
timestamp 1679581782
transform 1 0 36576 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_382
timestamp 1679581782
transform 1 0 37248 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_389
timestamp 1679581782
transform 1 0 37920 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_396
timestamp 1679581782
transform 1 0 38592 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_403
timestamp 1679581782
transform 1 0 39264 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_410
timestamp 1679581782
transform 1 0 39936 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_417
timestamp 1679581782
transform 1 0 40608 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_424
timestamp 1679581782
transform 1 0 41280 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_431
timestamp 1679581782
transform 1 0 41952 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_438
timestamp 1679581782
transform 1 0 42624 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_445
timestamp 1679581782
transform 1 0 43296 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_452
timestamp 1679581782
transform 1 0 43968 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_459
timestamp 1679581782
transform 1 0 44640 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_466
timestamp 1679581782
transform 1 0 45312 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_473
timestamp 1679581782
transform 1 0 45984 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_480
timestamp 1679581782
transform 1 0 46656 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_487
timestamp 1679581782
transform 1 0 47328 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_494
timestamp 1679581782
transform 1 0 48000 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_501
timestamp 1679581782
transform 1 0 48672 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_508
timestamp 1679581782
transform 1 0 49344 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_515
timestamp 1679581782
transform 1 0 50016 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_522
timestamp 1679581782
transform 1 0 50688 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_529
timestamp 1679581782
transform 1 0 51360 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_536
timestamp 1679581782
transform 1 0 52032 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_543
timestamp 1679581782
transform 1 0 52704 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_550
timestamp 1679581782
transform 1 0 53376 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_557
timestamp 1679581782
transform 1 0 54048 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_564
timestamp 1679581782
transform 1 0 54720 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_571
timestamp 1679581782
transform 1 0 55392 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_578
timestamp 1679581782
transform 1 0 56064 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_585
timestamp 1679581782
transform 1 0 56736 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_592
timestamp 1679581782
transform 1 0 57408 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_599
timestamp 1679581782
transform 1 0 58080 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_606
timestamp 1679581782
transform 1 0 58752 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_613
timestamp 1679581782
transform 1 0 59424 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_620
timestamp 1679581782
transform 1 0 60096 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_627
timestamp 1679581782
transform 1 0 60768 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_634
timestamp 1679581782
transform 1 0 61440 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_641
timestamp 1679581782
transform 1 0 62112 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_648
timestamp 1679581782
transform 1 0 62784 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_655
timestamp 1679581782
transform 1 0 63456 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_662
timestamp 1679581782
transform 1 0 64128 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_669
timestamp 1679581782
transform 1 0 64800 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_676
timestamp 1679581782
transform 1 0 65472 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_683
timestamp 1679581782
transform 1 0 66144 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_690
timestamp 1679581782
transform 1 0 66816 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_697
timestamp 1679581782
transform 1 0 67488 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_704
timestamp 1679581782
transform 1 0 68160 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_711
timestamp 1679581782
transform 1 0 68832 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_718
timestamp 1679581782
transform 1 0 69504 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_725
timestamp 1679581782
transform 1 0 70176 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_732
timestamp 1679581782
transform 1 0 70848 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_739
timestamp 1679581782
transform 1 0 71520 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_746
timestamp 1679581782
transform 1 0 72192 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_753
timestamp 1679581782
transform 1 0 72864 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_760
timestamp 1679581782
transform 1 0 73536 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_767
timestamp 1679581782
transform 1 0 74208 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_774
timestamp 1679581782
transform 1 0 74880 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_781
timestamp 1679581782
transform 1 0 75552 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_788
timestamp 1679581782
transform 1 0 76224 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_795
timestamp 1679581782
transform 1 0 76896 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_802
timestamp 1679581782
transform 1 0 77568 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_809
timestamp 1679581782
transform 1 0 78240 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_816
timestamp 1679581782
transform 1 0 78912 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_823
timestamp 1679581782
transform 1 0 79584 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_830
timestamp 1679581782
transform 1 0 80256 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_837
timestamp 1679581782
transform 1 0 80928 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_844
timestamp 1679581782
transform 1 0 81600 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_851
timestamp 1679581782
transform 1 0 82272 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_858
timestamp 1679581782
transform 1 0 82944 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_865
timestamp 1679581782
transform 1 0 83616 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_872
timestamp 1679581782
transform 1 0 84288 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_879
timestamp 1679581782
transform 1 0 84960 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_886
timestamp 1679581782
transform 1 0 85632 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_893
timestamp 1679581782
transform 1 0 86304 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_900
timestamp 1679581782
transform 1 0 86976 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_907
timestamp 1679581782
transform 1 0 87648 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_914
timestamp 1679581782
transform 1 0 88320 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_23_921
timestamp 1679577901
transform 1 0 88992 0 -1 18900
box -48 -56 432 834
use sg13g2_decap_8  FILLER_24_4
timestamp 1679581782
transform 1 0 960 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_11
timestamp 1679581782
transform 1 0 1632 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_18
timestamp 1679581782
transform 1 0 2304 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_25
timestamp 1679581782
transform 1 0 2976 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_32
timestamp 1679581782
transform 1 0 3648 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_39
timestamp 1679581782
transform 1 0 4320 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_46
timestamp 1679581782
transform 1 0 4992 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_53
timestamp 1679581782
transform 1 0 5664 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_60
timestamp 1679581782
transform 1 0 6336 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_67
timestamp 1679581782
transform 1 0 7008 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_24_74
timestamp 1677580104
transform 1 0 7680 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_76
timestamp 1677579658
transform 1 0 7872 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_82
timestamp 1679581782
transform 1 0 8448 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_89
timestamp 1679581782
transform 1 0 9120 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_96
timestamp 1679581782
transform 1 0 9792 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_103
timestamp 1679581782
transform 1 0 10464 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_110
timestamp 1679581782
transform 1 0 11136 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_117
timestamp 1679581782
transform 1 0 11808 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_124
timestamp 1679581782
transform 1 0 12480 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_131
timestamp 1679581782
transform 1 0 13152 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_138
timestamp 1679581782
transform 1 0 13824 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_145
timestamp 1679581782
transform 1 0 14496 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_152
timestamp 1679581782
transform 1 0 15168 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_159
timestamp 1679581782
transform 1 0 15840 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_166
timestamp 1679581782
transform 1 0 16512 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_173
timestamp 1679581782
transform 1 0 17184 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_180
timestamp 1679581782
transform 1 0 17856 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_187
timestamp 1679581782
transform 1 0 18528 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_194
timestamp 1679581782
transform 1 0 19200 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_201
timestamp 1679581782
transform 1 0 19872 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_208
timestamp 1679581782
transform 1 0 20544 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_215
timestamp 1679581782
transform 1 0 21216 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_222
timestamp 1679581782
transform 1 0 21888 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_229
timestamp 1679581782
transform 1 0 22560 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_236
timestamp 1679581782
transform 1 0 23232 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_243
timestamp 1679581782
transform 1 0 23904 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_250
timestamp 1679581782
transform 1 0 24576 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_257
timestamp 1679581782
transform 1 0 25248 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_264
timestamp 1679581782
transform 1 0 25920 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_271
timestamp 1679581782
transform 1 0 26592 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_278
timestamp 1679581782
transform 1 0 27264 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_285
timestamp 1679581782
transform 1 0 27936 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_292
timestamp 1679581782
transform 1 0 28608 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_299
timestamp 1679581782
transform 1 0 29280 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_306
timestamp 1679581782
transform 1 0 29952 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_313
timestamp 1679581782
transform 1 0 30624 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_320
timestamp 1679581782
transform 1 0 31296 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_327
timestamp 1679581782
transform 1 0 31968 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_334
timestamp 1679581782
transform 1 0 32640 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_341
timestamp 1679581782
transform 1 0 33312 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_348
timestamp 1679581782
transform 1 0 33984 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_355
timestamp 1679581782
transform 1 0 34656 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_362
timestamp 1679581782
transform 1 0 35328 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_369
timestamp 1679581782
transform 1 0 36000 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_376
timestamp 1679581782
transform 1 0 36672 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_383
timestamp 1679581782
transform 1 0 37344 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_390
timestamp 1679581782
transform 1 0 38016 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_397
timestamp 1679581782
transform 1 0 38688 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_404
timestamp 1679581782
transform 1 0 39360 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_411
timestamp 1679581782
transform 1 0 40032 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_418
timestamp 1679581782
transform 1 0 40704 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_425
timestamp 1679581782
transform 1 0 41376 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_432
timestamp 1679581782
transform 1 0 42048 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_439
timestamp 1679581782
transform 1 0 42720 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_446
timestamp 1679581782
transform 1 0 43392 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_453
timestamp 1679581782
transform 1 0 44064 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_460
timestamp 1679581782
transform 1 0 44736 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_467
timestamp 1679581782
transform 1 0 45408 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_474
timestamp 1679581782
transform 1 0 46080 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_481
timestamp 1679581782
transform 1 0 46752 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_488
timestamp 1679581782
transform 1 0 47424 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_495
timestamp 1679581782
transform 1 0 48096 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_502
timestamp 1679581782
transform 1 0 48768 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_509
timestamp 1679581782
transform 1 0 49440 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_516
timestamp 1679581782
transform 1 0 50112 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_523
timestamp 1679581782
transform 1 0 50784 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_530
timestamp 1679581782
transform 1 0 51456 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_537
timestamp 1679581782
transform 1 0 52128 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_544
timestamp 1679581782
transform 1 0 52800 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_551
timestamp 1679581782
transform 1 0 53472 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_558
timestamp 1679581782
transform 1 0 54144 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_565
timestamp 1679581782
transform 1 0 54816 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_572
timestamp 1679581782
transform 1 0 55488 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_579
timestamp 1679581782
transform 1 0 56160 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_586
timestamp 1679581782
transform 1 0 56832 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_593
timestamp 1679581782
transform 1 0 57504 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_600
timestamp 1679581782
transform 1 0 58176 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_607
timestamp 1679581782
transform 1 0 58848 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_614
timestamp 1679581782
transform 1 0 59520 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_621
timestamp 1679581782
transform 1 0 60192 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_628
timestamp 1679581782
transform 1 0 60864 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_635
timestamp 1679581782
transform 1 0 61536 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_642
timestamp 1679581782
transform 1 0 62208 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_649
timestamp 1679581782
transform 1 0 62880 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_656
timestamp 1679581782
transform 1 0 63552 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_663
timestamp 1679581782
transform 1 0 64224 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_670
timestamp 1679581782
transform 1 0 64896 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_677
timestamp 1679581782
transform 1 0 65568 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_684
timestamp 1679581782
transform 1 0 66240 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_691
timestamp 1679581782
transform 1 0 66912 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_698
timestamp 1679581782
transform 1 0 67584 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_705
timestamp 1679581782
transform 1 0 68256 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_712
timestamp 1679581782
transform 1 0 68928 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_719
timestamp 1679581782
transform 1 0 69600 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_726
timestamp 1679581782
transform 1 0 70272 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_733
timestamp 1679581782
transform 1 0 70944 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_740
timestamp 1679581782
transform 1 0 71616 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_747
timestamp 1679581782
transform 1 0 72288 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_754
timestamp 1679581782
transform 1 0 72960 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_761
timestamp 1679581782
transform 1 0 73632 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_768
timestamp 1679581782
transform 1 0 74304 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_775
timestamp 1679581782
transform 1 0 74976 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_782
timestamp 1679581782
transform 1 0 75648 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_789
timestamp 1679581782
transform 1 0 76320 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_796
timestamp 1679581782
transform 1 0 76992 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_803
timestamp 1679581782
transform 1 0 77664 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_810
timestamp 1679581782
transform 1 0 78336 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_817
timestamp 1679581782
transform 1 0 79008 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_824
timestamp 1679581782
transform 1 0 79680 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_831
timestamp 1679581782
transform 1 0 80352 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_838
timestamp 1679581782
transform 1 0 81024 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_845
timestamp 1679581782
transform 1 0 81696 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_852
timestamp 1679581782
transform 1 0 82368 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_859
timestamp 1679581782
transform 1 0 83040 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_866
timestamp 1679581782
transform 1 0 83712 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_873
timestamp 1679581782
transform 1 0 84384 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_880
timestamp 1679581782
transform 1 0 85056 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_887
timestamp 1679581782
transform 1 0 85728 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_894
timestamp 1679581782
transform 1 0 86400 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_901
timestamp 1679581782
transform 1 0 87072 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_908
timestamp 1679581782
transform 1 0 87744 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_915
timestamp 1679581782
transform 1 0 88416 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_24_922
timestamp 1677580104
transform 1 0 89088 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_924
timestamp 1677579658
transform 1 0 89280 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_4
timestamp 1679581782
transform 1 0 960 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_11
timestamp 1679581782
transform 1 0 1632 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_18
timestamp 1679581782
transform 1 0 2304 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_25
timestamp 1679581782
transform 1 0 2976 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_32
timestamp 1679581782
transform 1 0 3648 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_39
timestamp 1679581782
transform 1 0 4320 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_46
timestamp 1679581782
transform 1 0 4992 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_53
timestamp 1679581782
transform 1 0 5664 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_60
timestamp 1679581782
transform 1 0 6336 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_67
timestamp 1679581782
transform 1 0 7008 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_90
timestamp 1679581782
transform 1 0 9216 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_97
timestamp 1679581782
transform 1 0 9888 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_104
timestamp 1679581782
transform 1 0 10560 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_111
timestamp 1679581782
transform 1 0 11232 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_118
timestamp 1679581782
transform 1 0 11904 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_125
timestamp 1679581782
transform 1 0 12576 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_132
timestamp 1679581782
transform 1 0 13248 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_139
timestamp 1679581782
transform 1 0 13920 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_146
timestamp 1679581782
transform 1 0 14592 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_153
timestamp 1679581782
transform 1 0 15264 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_160
timestamp 1679581782
transform 1 0 15936 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_167
timestamp 1679581782
transform 1 0 16608 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_174
timestamp 1679581782
transform 1 0 17280 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_181
timestamp 1679581782
transform 1 0 17952 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_188
timestamp 1679581782
transform 1 0 18624 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_195
timestamp 1679581782
transform 1 0 19296 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_202
timestamp 1679581782
transform 1 0 19968 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_209
timestamp 1679581782
transform 1 0 20640 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_216
timestamp 1679581782
transform 1 0 21312 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_223
timestamp 1679581782
transform 1 0 21984 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_230
timestamp 1679581782
transform 1 0 22656 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_237
timestamp 1679581782
transform 1 0 23328 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_244
timestamp 1679581782
transform 1 0 24000 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_251
timestamp 1679581782
transform 1 0 24672 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_258
timestamp 1679581782
transform 1 0 25344 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_265
timestamp 1679581782
transform 1 0 26016 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_272
timestamp 1679581782
transform 1 0 26688 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_279
timestamp 1679581782
transform 1 0 27360 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_286
timestamp 1679581782
transform 1 0 28032 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_293
timestamp 1679581782
transform 1 0 28704 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_300
timestamp 1679581782
transform 1 0 29376 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_307
timestamp 1679581782
transform 1 0 30048 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_314
timestamp 1679581782
transform 1 0 30720 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_321
timestamp 1679581782
transform 1 0 31392 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_328
timestamp 1679581782
transform 1 0 32064 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_335
timestamp 1679581782
transform 1 0 32736 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_342
timestamp 1679581782
transform 1 0 33408 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_349
timestamp 1679581782
transform 1 0 34080 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_356
timestamp 1679581782
transform 1 0 34752 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_363
timestamp 1679581782
transform 1 0 35424 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_370
timestamp 1679581782
transform 1 0 36096 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_377
timestamp 1679581782
transform 1 0 36768 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_384
timestamp 1679581782
transform 1 0 37440 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_391
timestamp 1679581782
transform 1 0 38112 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_398
timestamp 1679581782
transform 1 0 38784 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_405
timestamp 1679581782
transform 1 0 39456 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_412
timestamp 1679581782
transform 1 0 40128 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_419
timestamp 1679581782
transform 1 0 40800 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_426
timestamp 1679581782
transform 1 0 41472 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_433
timestamp 1679581782
transform 1 0 42144 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_440
timestamp 1679581782
transform 1 0 42816 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_447
timestamp 1679581782
transform 1 0 43488 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_454
timestamp 1679581782
transform 1 0 44160 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_461
timestamp 1679581782
transform 1 0 44832 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_468
timestamp 1679581782
transform 1 0 45504 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_475
timestamp 1679581782
transform 1 0 46176 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_482
timestamp 1679581782
transform 1 0 46848 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_489
timestamp 1679581782
transform 1 0 47520 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_496
timestamp 1679581782
transform 1 0 48192 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_503
timestamp 1679581782
transform 1 0 48864 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_510
timestamp 1679581782
transform 1 0 49536 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_517
timestamp 1679581782
transform 1 0 50208 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_524
timestamp 1679581782
transform 1 0 50880 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_531
timestamp 1679581782
transform 1 0 51552 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_538
timestamp 1679581782
transform 1 0 52224 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_545
timestamp 1679581782
transform 1 0 52896 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_552
timestamp 1679581782
transform 1 0 53568 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_559
timestamp 1679581782
transform 1 0 54240 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_566
timestamp 1679581782
transform 1 0 54912 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_573
timestamp 1679581782
transform 1 0 55584 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_580
timestamp 1679581782
transform 1 0 56256 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_587
timestamp 1679581782
transform 1 0 56928 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_594
timestamp 1679581782
transform 1 0 57600 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_601
timestamp 1679581782
transform 1 0 58272 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_608
timestamp 1679581782
transform 1 0 58944 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_615
timestamp 1679581782
transform 1 0 59616 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_622
timestamp 1679581782
transform 1 0 60288 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_629
timestamp 1679581782
transform 1 0 60960 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_636
timestamp 1679581782
transform 1 0 61632 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_643
timestamp 1679581782
transform 1 0 62304 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_650
timestamp 1679581782
transform 1 0 62976 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_657
timestamp 1679581782
transform 1 0 63648 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_664
timestamp 1679581782
transform 1 0 64320 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_671
timestamp 1679581782
transform 1 0 64992 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_678
timestamp 1679581782
transform 1 0 65664 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_685
timestamp 1679581782
transform 1 0 66336 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_692
timestamp 1679581782
transform 1 0 67008 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_699
timestamp 1679581782
transform 1 0 67680 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_706
timestamp 1679581782
transform 1 0 68352 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_713
timestamp 1679581782
transform 1 0 69024 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_720
timestamp 1679581782
transform 1 0 69696 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_727
timestamp 1679581782
transform 1 0 70368 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_734
timestamp 1679581782
transform 1 0 71040 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_741
timestamp 1679581782
transform 1 0 71712 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_748
timestamp 1679581782
transform 1 0 72384 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_755
timestamp 1679581782
transform 1 0 73056 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_762
timestamp 1679581782
transform 1 0 73728 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_769
timestamp 1679581782
transform 1 0 74400 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_776
timestamp 1679581782
transform 1 0 75072 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_783
timestamp 1679581782
transform 1 0 75744 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_790
timestamp 1679581782
transform 1 0 76416 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_797
timestamp 1679581782
transform 1 0 77088 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_804
timestamp 1679581782
transform 1 0 77760 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_811
timestamp 1679581782
transform 1 0 78432 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_818
timestamp 1679581782
transform 1 0 79104 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_825
timestamp 1679581782
transform 1 0 79776 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_832
timestamp 1679581782
transform 1 0 80448 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_839
timestamp 1679581782
transform 1 0 81120 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_846
timestamp 1679581782
transform 1 0 81792 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_853
timestamp 1679581782
transform 1 0 82464 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_860
timestamp 1679581782
transform 1 0 83136 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_867
timestamp 1679581782
transform 1 0 83808 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_874
timestamp 1679581782
transform 1 0 84480 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_881
timestamp 1679581782
transform 1 0 85152 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_888
timestamp 1679581782
transform 1 0 85824 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_895
timestamp 1679581782
transform 1 0 86496 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_902
timestamp 1679581782
transform 1 0 87168 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_909
timestamp 1679581782
transform 1 0 87840 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_916
timestamp 1679581782
transform 1 0 88512 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_923
timestamp 1677580104
transform 1 0 89184 0 -1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_26_4
timestamp 1679581782
transform 1 0 960 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_11
timestamp 1679581782
transform 1 0 1632 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_18
timestamp 1679581782
transform 1 0 2304 0 1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_26_25
timestamp 1677580104
transform 1 0 2976 0 1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_26_40
timestamp 1679581782
transform 1 0 4416 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_47
timestamp 1679581782
transform 1 0 5088 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_54
timestamp 1679581782
transform 1 0 5760 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_61
timestamp 1679581782
transform 1 0 6432 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_68
timestamp 1679581782
transform 1 0 7104 0 1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_26_75
timestamp 1679577901
transform 1 0 7776 0 1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_26_79
timestamp 1677579658
transform 1 0 8160 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_88
timestamp 1679581782
transform 1 0 9024 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_95
timestamp 1679581782
transform 1 0 9696 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_102
timestamp 1679581782
transform 1 0 10368 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_109
timestamp 1679581782
transform 1 0 11040 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_116
timestamp 1679581782
transform 1 0 11712 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_123
timestamp 1679581782
transform 1 0 12384 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_130
timestamp 1679581782
transform 1 0 13056 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_137
timestamp 1679581782
transform 1 0 13728 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_144
timestamp 1679581782
transform 1 0 14400 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_151
timestamp 1679581782
transform 1 0 15072 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_158
timestamp 1679581782
transform 1 0 15744 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_165
timestamp 1679581782
transform 1 0 16416 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_172
timestamp 1679581782
transform 1 0 17088 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_179
timestamp 1679581782
transform 1 0 17760 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_186
timestamp 1679581782
transform 1 0 18432 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_193
timestamp 1679581782
transform 1 0 19104 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_200
timestamp 1679581782
transform 1 0 19776 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_207
timestamp 1679581782
transform 1 0 20448 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_214
timestamp 1679581782
transform 1 0 21120 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_221
timestamp 1679581782
transform 1 0 21792 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_228
timestamp 1679581782
transform 1 0 22464 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_235
timestamp 1679581782
transform 1 0 23136 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_242
timestamp 1679581782
transform 1 0 23808 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_249
timestamp 1679581782
transform 1 0 24480 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_256
timestamp 1679581782
transform 1 0 25152 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_263
timestamp 1679581782
transform 1 0 25824 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_270
timestamp 1679581782
transform 1 0 26496 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_277
timestamp 1679581782
transform 1 0 27168 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_284
timestamp 1679581782
transform 1 0 27840 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_291
timestamp 1679581782
transform 1 0 28512 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_298
timestamp 1679581782
transform 1 0 29184 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_305
timestamp 1679581782
transform 1 0 29856 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_312
timestamp 1679581782
transform 1 0 30528 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_319
timestamp 1679581782
transform 1 0 31200 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_326
timestamp 1679581782
transform 1 0 31872 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_333
timestamp 1679581782
transform 1 0 32544 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_340
timestamp 1679581782
transform 1 0 33216 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_347
timestamp 1679581782
transform 1 0 33888 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_354
timestamp 1679581782
transform 1 0 34560 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_361
timestamp 1679581782
transform 1 0 35232 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_368
timestamp 1679581782
transform 1 0 35904 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_375
timestamp 1679581782
transform 1 0 36576 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_382
timestamp 1679581782
transform 1 0 37248 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_389
timestamp 1679581782
transform 1 0 37920 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_396
timestamp 1679581782
transform 1 0 38592 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_403
timestamp 1679581782
transform 1 0 39264 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_410
timestamp 1679581782
transform 1 0 39936 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_417
timestamp 1679581782
transform 1 0 40608 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_424
timestamp 1679581782
transform 1 0 41280 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_431
timestamp 1679581782
transform 1 0 41952 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_438
timestamp 1679581782
transform 1 0 42624 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_445
timestamp 1679581782
transform 1 0 43296 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_452
timestamp 1679581782
transform 1 0 43968 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_459
timestamp 1679581782
transform 1 0 44640 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_466
timestamp 1679581782
transform 1 0 45312 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_473
timestamp 1679581782
transform 1 0 45984 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_480
timestamp 1679581782
transform 1 0 46656 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_487
timestamp 1679581782
transform 1 0 47328 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_494
timestamp 1679581782
transform 1 0 48000 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_501
timestamp 1679581782
transform 1 0 48672 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_508
timestamp 1679581782
transform 1 0 49344 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_515
timestamp 1679581782
transform 1 0 50016 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_522
timestamp 1679581782
transform 1 0 50688 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_529
timestamp 1679581782
transform 1 0 51360 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_536
timestamp 1679581782
transform 1 0 52032 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_543
timestamp 1679581782
transform 1 0 52704 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_550
timestamp 1679581782
transform 1 0 53376 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_557
timestamp 1679581782
transform 1 0 54048 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_564
timestamp 1679581782
transform 1 0 54720 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_571
timestamp 1679581782
transform 1 0 55392 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_578
timestamp 1679581782
transform 1 0 56064 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_585
timestamp 1679581782
transform 1 0 56736 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_592
timestamp 1679581782
transform 1 0 57408 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_599
timestamp 1679581782
transform 1 0 58080 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_606
timestamp 1679581782
transform 1 0 58752 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_613
timestamp 1679581782
transform 1 0 59424 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_620
timestamp 1679581782
transform 1 0 60096 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_627
timestamp 1679581782
transform 1 0 60768 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_634
timestamp 1679581782
transform 1 0 61440 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_641
timestamp 1679581782
transform 1 0 62112 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_648
timestamp 1679581782
transform 1 0 62784 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_655
timestamp 1679581782
transform 1 0 63456 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_662
timestamp 1679581782
transform 1 0 64128 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_669
timestamp 1679581782
transform 1 0 64800 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_676
timestamp 1679581782
transform 1 0 65472 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_683
timestamp 1679581782
transform 1 0 66144 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_690
timestamp 1679581782
transform 1 0 66816 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_697
timestamp 1679581782
transform 1 0 67488 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_704
timestamp 1679581782
transform 1 0 68160 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_711
timestamp 1679581782
transform 1 0 68832 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_718
timestamp 1679581782
transform 1 0 69504 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_725
timestamp 1679581782
transform 1 0 70176 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_732
timestamp 1679581782
transform 1 0 70848 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_739
timestamp 1679581782
transform 1 0 71520 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_746
timestamp 1679581782
transform 1 0 72192 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_753
timestamp 1679581782
transform 1 0 72864 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_760
timestamp 1679581782
transform 1 0 73536 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_767
timestamp 1679581782
transform 1 0 74208 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_774
timestamp 1679581782
transform 1 0 74880 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_781
timestamp 1679581782
transform 1 0 75552 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_788
timestamp 1679581782
transform 1 0 76224 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_795
timestamp 1679581782
transform 1 0 76896 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_802
timestamp 1679581782
transform 1 0 77568 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_809
timestamp 1679581782
transform 1 0 78240 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_816
timestamp 1679581782
transform 1 0 78912 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_823
timestamp 1679581782
transform 1 0 79584 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_830
timestamp 1679581782
transform 1 0 80256 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_837
timestamp 1679581782
transform 1 0 80928 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_844
timestamp 1679581782
transform 1 0 81600 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_851
timestamp 1679581782
transform 1 0 82272 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_858
timestamp 1679581782
transform 1 0 82944 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_865
timestamp 1679581782
transform 1 0 83616 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_872
timestamp 1679581782
transform 1 0 84288 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_879
timestamp 1679581782
transform 1 0 84960 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_886
timestamp 1679581782
transform 1 0 85632 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_893
timestamp 1679581782
transform 1 0 86304 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_900
timestamp 1679581782
transform 1 0 86976 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_907
timestamp 1679581782
transform 1 0 87648 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_914
timestamp 1679581782
transform 1 0 88320 0 1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_26_921
timestamp 1679577901
transform 1 0 88992 0 1 20412
box -48 -56 432 834
use sg13g2_decap_8  FILLER_27_0
timestamp 1679581782
transform 1 0 576 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_7
timestamp 1679581782
transform 1 0 1248 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_14
timestamp 1679581782
transform 1 0 1920 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_21
timestamp 1679581782
transform 1 0 2592 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_28
timestamp 1679581782
transform 1 0 3264 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_35
timestamp 1679581782
transform 1 0 3936 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_42
timestamp 1679581782
transform 1 0 4608 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_49
timestamp 1679581782
transform 1 0 5280 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_56
timestamp 1679581782
transform 1 0 5952 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_63
timestamp 1679581782
transform 1 0 6624 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_70
timestamp 1679581782
transform 1 0 7296 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_77
timestamp 1679581782
transform 1 0 7968 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_84
timestamp 1679581782
transform 1 0 8640 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_91
timestamp 1679581782
transform 1 0 9312 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_98
timestamp 1679581782
transform 1 0 9984 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_105
timestamp 1679581782
transform 1 0 10656 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_112
timestamp 1679581782
transform 1 0 11328 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_119
timestamp 1679581782
transform 1 0 12000 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_126
timestamp 1679581782
transform 1 0 12672 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_133
timestamp 1679581782
transform 1 0 13344 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_140
timestamp 1679581782
transform 1 0 14016 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_147
timestamp 1679581782
transform 1 0 14688 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_154
timestamp 1679581782
transform 1 0 15360 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_161
timestamp 1679581782
transform 1 0 16032 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_168
timestamp 1679581782
transform 1 0 16704 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_175
timestamp 1679581782
transform 1 0 17376 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_182
timestamp 1679581782
transform 1 0 18048 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_189
timestamp 1679581782
transform 1 0 18720 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_196
timestamp 1679581782
transform 1 0 19392 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_203
timestamp 1679581782
transform 1 0 20064 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_210
timestamp 1679581782
transform 1 0 20736 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_217
timestamp 1679581782
transform 1 0 21408 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_224
timestamp 1679581782
transform 1 0 22080 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_231
timestamp 1679581782
transform 1 0 22752 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_238
timestamp 1679581782
transform 1 0 23424 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_245
timestamp 1679581782
transform 1 0 24096 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_252
timestamp 1679581782
transform 1 0 24768 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_259
timestamp 1679581782
transform 1 0 25440 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_266
timestamp 1679581782
transform 1 0 26112 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_273
timestamp 1679581782
transform 1 0 26784 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_280
timestamp 1679581782
transform 1 0 27456 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_287
timestamp 1679581782
transform 1 0 28128 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_294
timestamp 1679581782
transform 1 0 28800 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_301
timestamp 1679581782
transform 1 0 29472 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_308
timestamp 1679581782
transform 1 0 30144 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_315
timestamp 1679581782
transform 1 0 30816 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_322
timestamp 1679581782
transform 1 0 31488 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_329
timestamp 1679581782
transform 1 0 32160 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_336
timestamp 1679581782
transform 1 0 32832 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_343
timestamp 1679581782
transform 1 0 33504 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_350
timestamp 1679581782
transform 1 0 34176 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_357
timestamp 1679581782
transform 1 0 34848 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_364
timestamp 1679581782
transform 1 0 35520 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_371
timestamp 1679581782
transform 1 0 36192 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_378
timestamp 1679581782
transform 1 0 36864 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_385
timestamp 1679581782
transform 1 0 37536 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_392
timestamp 1679581782
transform 1 0 38208 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_399
timestamp 1679581782
transform 1 0 38880 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_406
timestamp 1679581782
transform 1 0 39552 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_413
timestamp 1679581782
transform 1 0 40224 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_420
timestamp 1679581782
transform 1 0 40896 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_427
timestamp 1679581782
transform 1 0 41568 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_434
timestamp 1679581782
transform 1 0 42240 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_441
timestamp 1679581782
transform 1 0 42912 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_448
timestamp 1679581782
transform 1 0 43584 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_455
timestamp 1679581782
transform 1 0 44256 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_462
timestamp 1679581782
transform 1 0 44928 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_469
timestamp 1679581782
transform 1 0 45600 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_476
timestamp 1679581782
transform 1 0 46272 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_483
timestamp 1679581782
transform 1 0 46944 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_490
timestamp 1679581782
transform 1 0 47616 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_497
timestamp 1679581782
transform 1 0 48288 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_504
timestamp 1679581782
transform 1 0 48960 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_511
timestamp 1679581782
transform 1 0 49632 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_518
timestamp 1679581782
transform 1 0 50304 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_525
timestamp 1679581782
transform 1 0 50976 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_532
timestamp 1679581782
transform 1 0 51648 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_539
timestamp 1679581782
transform 1 0 52320 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_546
timestamp 1679581782
transform 1 0 52992 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_553
timestamp 1679581782
transform 1 0 53664 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_560
timestamp 1679581782
transform 1 0 54336 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_567
timestamp 1679581782
transform 1 0 55008 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_574
timestamp 1679581782
transform 1 0 55680 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_581
timestamp 1679581782
transform 1 0 56352 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_588
timestamp 1679581782
transform 1 0 57024 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_595
timestamp 1679581782
transform 1 0 57696 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_602
timestamp 1679581782
transform 1 0 58368 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_609
timestamp 1679581782
transform 1 0 59040 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_616
timestamp 1679581782
transform 1 0 59712 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_623
timestamp 1679581782
transform 1 0 60384 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_630
timestamp 1679581782
transform 1 0 61056 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_637
timestamp 1679581782
transform 1 0 61728 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_644
timestamp 1679581782
transform 1 0 62400 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_651
timestamp 1679581782
transform 1 0 63072 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_658
timestamp 1679581782
transform 1 0 63744 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_665
timestamp 1679581782
transform 1 0 64416 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_672
timestamp 1679581782
transform 1 0 65088 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_679
timestamp 1679581782
transform 1 0 65760 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_686
timestamp 1679581782
transform 1 0 66432 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_693
timestamp 1679581782
transform 1 0 67104 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_700
timestamp 1679581782
transform 1 0 67776 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_707
timestamp 1679581782
transform 1 0 68448 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_714
timestamp 1679581782
transform 1 0 69120 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_721
timestamp 1679581782
transform 1 0 69792 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_728
timestamp 1679581782
transform 1 0 70464 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_735
timestamp 1679581782
transform 1 0 71136 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_742
timestamp 1679581782
transform 1 0 71808 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_749
timestamp 1679581782
transform 1 0 72480 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_756
timestamp 1679581782
transform 1 0 73152 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_763
timestamp 1679581782
transform 1 0 73824 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_770
timestamp 1679581782
transform 1 0 74496 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_777
timestamp 1679581782
transform 1 0 75168 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_784
timestamp 1679581782
transform 1 0 75840 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_791
timestamp 1679581782
transform 1 0 76512 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_798
timestamp 1679581782
transform 1 0 77184 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_805
timestamp 1679581782
transform 1 0 77856 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_812
timestamp 1679581782
transform 1 0 78528 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_819
timestamp 1679581782
transform 1 0 79200 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_826
timestamp 1679581782
transform 1 0 79872 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_833
timestamp 1679581782
transform 1 0 80544 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_840
timestamp 1679581782
transform 1 0 81216 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_847
timestamp 1679581782
transform 1 0 81888 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_854
timestamp 1679581782
transform 1 0 82560 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_861
timestamp 1679581782
transform 1 0 83232 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_868
timestamp 1679581782
transform 1 0 83904 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_875
timestamp 1679581782
transform 1 0 84576 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_882
timestamp 1679581782
transform 1 0 85248 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_889
timestamp 1679581782
transform 1 0 85920 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_896
timestamp 1679581782
transform 1 0 86592 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_903
timestamp 1679581782
transform 1 0 87264 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_910
timestamp 1679581782
transform 1 0 87936 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_917
timestamp 1679581782
transform 1 0 88608 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_1  FILLER_27_924
timestamp 1677579658
transform 1 0 89280 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_4
timestamp 1679581782
transform 1 0 960 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_11
timestamp 1679581782
transform 1 0 1632 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_18
timestamp 1679581782
transform 1 0 2304 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_25
timestamp 1679581782
transform 1 0 2976 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_32
timestamp 1679581782
transform 1 0 3648 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_39
timestamp 1679581782
transform 1 0 4320 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_46
timestamp 1679581782
transform 1 0 4992 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_53
timestamp 1679581782
transform 1 0 5664 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_60
timestamp 1679581782
transform 1 0 6336 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_67
timestamp 1679581782
transform 1 0 7008 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_74
timestamp 1679581782
transform 1 0 7680 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_81
timestamp 1679581782
transform 1 0 8352 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_88
timestamp 1679581782
transform 1 0 9024 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_95
timestamp 1679581782
transform 1 0 9696 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_102
timestamp 1679577901
transform 1 0 10368 0 1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_28_106
timestamp 1677580104
transform 1 0 10752 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_116
timestamp 1677579658
transform 1 0 11712 0 1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_125
timestamp 1679581782
transform 1 0 12576 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_132
timestamp 1679581782
transform 1 0 13248 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_139
timestamp 1679581782
transform 1 0 13920 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_146
timestamp 1679581782
transform 1 0 14592 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_153
timestamp 1679581782
transform 1 0 15264 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_160
timestamp 1679581782
transform 1 0 15936 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_167
timestamp 1679581782
transform 1 0 16608 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_174
timestamp 1679581782
transform 1 0 17280 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_181
timestamp 1679581782
transform 1 0 17952 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_188
timestamp 1679581782
transform 1 0 18624 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_195
timestamp 1679581782
transform 1 0 19296 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_202
timestamp 1679581782
transform 1 0 19968 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_209
timestamp 1679581782
transform 1 0 20640 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_216
timestamp 1679581782
transform 1 0 21312 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_223
timestamp 1679581782
transform 1 0 21984 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_230
timestamp 1679581782
transform 1 0 22656 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_237
timestamp 1679581782
transform 1 0 23328 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_244
timestamp 1679581782
transform 1 0 24000 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_251
timestamp 1679581782
transform 1 0 24672 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_258
timestamp 1679581782
transform 1 0 25344 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_265
timestamp 1679581782
transform 1 0 26016 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_272
timestamp 1679581782
transform 1 0 26688 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_279
timestamp 1679581782
transform 1 0 27360 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_286
timestamp 1679581782
transform 1 0 28032 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_293
timestamp 1679581782
transform 1 0 28704 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_300
timestamp 1679581782
transform 1 0 29376 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_307
timestamp 1679581782
transform 1 0 30048 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_314
timestamp 1679581782
transform 1 0 30720 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_321
timestamp 1679581782
transform 1 0 31392 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_328
timestamp 1679581782
transform 1 0 32064 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_335
timestamp 1679581782
transform 1 0 32736 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_342
timestamp 1679581782
transform 1 0 33408 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_349
timestamp 1679581782
transform 1 0 34080 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_356
timestamp 1679581782
transform 1 0 34752 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_363
timestamp 1679581782
transform 1 0 35424 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_370
timestamp 1679581782
transform 1 0 36096 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_377
timestamp 1679581782
transform 1 0 36768 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_384
timestamp 1679581782
transform 1 0 37440 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_391
timestamp 1679581782
transform 1 0 38112 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_398
timestamp 1679581782
transform 1 0 38784 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_405
timestamp 1679581782
transform 1 0 39456 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_412
timestamp 1679581782
transform 1 0 40128 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_419
timestamp 1679581782
transform 1 0 40800 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_426
timestamp 1679581782
transform 1 0 41472 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_433
timestamp 1679581782
transform 1 0 42144 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_440
timestamp 1679581782
transform 1 0 42816 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_447
timestamp 1679581782
transform 1 0 43488 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_454
timestamp 1679581782
transform 1 0 44160 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_461
timestamp 1679581782
transform 1 0 44832 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_468
timestamp 1679581782
transform 1 0 45504 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_475
timestamp 1679581782
transform 1 0 46176 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_482
timestamp 1679581782
transform 1 0 46848 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_489
timestamp 1679581782
transform 1 0 47520 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_496
timestamp 1679581782
transform 1 0 48192 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_503
timestamp 1679581782
transform 1 0 48864 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_510
timestamp 1679581782
transform 1 0 49536 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_517
timestamp 1679581782
transform 1 0 50208 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_524
timestamp 1679581782
transform 1 0 50880 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_531
timestamp 1679581782
transform 1 0 51552 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_538
timestamp 1679581782
transform 1 0 52224 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_545
timestamp 1679581782
transform 1 0 52896 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_552
timestamp 1679581782
transform 1 0 53568 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_559
timestamp 1679581782
transform 1 0 54240 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_566
timestamp 1679581782
transform 1 0 54912 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_573
timestamp 1679581782
transform 1 0 55584 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_580
timestamp 1679581782
transform 1 0 56256 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_587
timestamp 1679581782
transform 1 0 56928 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_594
timestamp 1679581782
transform 1 0 57600 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_601
timestamp 1679581782
transform 1 0 58272 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_608
timestamp 1679581782
transform 1 0 58944 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_615
timestamp 1679581782
transform 1 0 59616 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_622
timestamp 1679581782
transform 1 0 60288 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_629
timestamp 1679581782
transform 1 0 60960 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_636
timestamp 1679581782
transform 1 0 61632 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_643
timestamp 1679581782
transform 1 0 62304 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_650
timestamp 1679581782
transform 1 0 62976 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_657
timestamp 1679581782
transform 1 0 63648 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_664
timestamp 1679581782
transform 1 0 64320 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_671
timestamp 1679581782
transform 1 0 64992 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_678
timestamp 1679581782
transform 1 0 65664 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_685
timestamp 1679581782
transform 1 0 66336 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_692
timestamp 1679581782
transform 1 0 67008 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_699
timestamp 1679581782
transform 1 0 67680 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_706
timestamp 1679581782
transform 1 0 68352 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_713
timestamp 1679581782
transform 1 0 69024 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_720
timestamp 1679581782
transform 1 0 69696 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_727
timestamp 1679581782
transform 1 0 70368 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_734
timestamp 1679581782
transform 1 0 71040 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_741
timestamp 1679581782
transform 1 0 71712 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_748
timestamp 1679581782
transform 1 0 72384 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_755
timestamp 1679581782
transform 1 0 73056 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_762
timestamp 1679581782
transform 1 0 73728 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_769
timestamp 1679581782
transform 1 0 74400 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_776
timestamp 1679581782
transform 1 0 75072 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_783
timestamp 1679581782
transform 1 0 75744 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_790
timestamp 1679581782
transform 1 0 76416 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_797
timestamp 1679581782
transform 1 0 77088 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_804
timestamp 1679581782
transform 1 0 77760 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_811
timestamp 1679581782
transform 1 0 78432 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_818
timestamp 1679581782
transform 1 0 79104 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_825
timestamp 1679581782
transform 1 0 79776 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_832
timestamp 1679581782
transform 1 0 80448 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_839
timestamp 1679581782
transform 1 0 81120 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_846
timestamp 1679581782
transform 1 0 81792 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_853
timestamp 1679581782
transform 1 0 82464 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_860
timestamp 1679581782
transform 1 0 83136 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_867
timestamp 1679581782
transform 1 0 83808 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_874
timestamp 1679581782
transform 1 0 84480 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_881
timestamp 1679581782
transform 1 0 85152 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_888
timestamp 1679581782
transform 1 0 85824 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_895
timestamp 1679581782
transform 1 0 86496 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_902
timestamp 1679581782
transform 1 0 87168 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_909
timestamp 1679581782
transform 1 0 87840 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_916
timestamp 1679581782
transform 1 0 88512 0 1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_28_923
timestamp 1677580104
transform 1 0 89184 0 1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_29_4
timestamp 1679581782
transform 1 0 960 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_11
timestamp 1679581782
transform 1 0 1632 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_18
timestamp 1679581782
transform 1 0 2304 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_25
timestamp 1679581782
transform 1 0 2976 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_32
timestamp 1679581782
transform 1 0 3648 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_39
timestamp 1679581782
transform 1 0 4320 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_46
timestamp 1679581782
transform 1 0 4992 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_53
timestamp 1679581782
transform 1 0 5664 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_60
timestamp 1679581782
transform 1 0 6336 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_67
timestamp 1679581782
transform 1 0 7008 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_74
timestamp 1679581782
transform 1 0 7680 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_81
timestamp 1679581782
transform 1 0 8352 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_88
timestamp 1679581782
transform 1 0 9024 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_95
timestamp 1679581782
transform 1 0 9696 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_102
timestamp 1679581782
transform 1 0 10368 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_109
timestamp 1679581782
transform 1 0 11040 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_29_116
timestamp 1677580104
transform 1 0 11712 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_118
timestamp 1677579658
transform 1 0 11904 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_29_124
timestamp 1679581782
transform 1 0 12480 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_131
timestamp 1679581782
transform 1 0 13152 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_138
timestamp 1679581782
transform 1 0 13824 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_145
timestamp 1679581782
transform 1 0 14496 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_152
timestamp 1679581782
transform 1 0 15168 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_159
timestamp 1679581782
transform 1 0 15840 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_166
timestamp 1679581782
transform 1 0 16512 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_173
timestamp 1679581782
transform 1 0 17184 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_180
timestamp 1679581782
transform 1 0 17856 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_187
timestamp 1679581782
transform 1 0 18528 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_194
timestamp 1679581782
transform 1 0 19200 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_201
timestamp 1679581782
transform 1 0 19872 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_208
timestamp 1679581782
transform 1 0 20544 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_215
timestamp 1679581782
transform 1 0 21216 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_222
timestamp 1679581782
transform 1 0 21888 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_229
timestamp 1679581782
transform 1 0 22560 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_236
timestamp 1679581782
transform 1 0 23232 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_243
timestamp 1679581782
transform 1 0 23904 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_250
timestamp 1679581782
transform 1 0 24576 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_257
timestamp 1679581782
transform 1 0 25248 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_264
timestamp 1679581782
transform 1 0 25920 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_271
timestamp 1679581782
transform 1 0 26592 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_278
timestamp 1679581782
transform 1 0 27264 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_285
timestamp 1679581782
transform 1 0 27936 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_292
timestamp 1679581782
transform 1 0 28608 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_299
timestamp 1679581782
transform 1 0 29280 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_306
timestamp 1679581782
transform 1 0 29952 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_313
timestamp 1679581782
transform 1 0 30624 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_320
timestamp 1679581782
transform 1 0 31296 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_327
timestamp 1679581782
transform 1 0 31968 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_334
timestamp 1679581782
transform 1 0 32640 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_341
timestamp 1679581782
transform 1 0 33312 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_348
timestamp 1679581782
transform 1 0 33984 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_355
timestamp 1679581782
transform 1 0 34656 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_362
timestamp 1679581782
transform 1 0 35328 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_369
timestamp 1679581782
transform 1 0 36000 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_376
timestamp 1679581782
transform 1 0 36672 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_383
timestamp 1679581782
transform 1 0 37344 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_390
timestamp 1679581782
transform 1 0 38016 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_397
timestamp 1679581782
transform 1 0 38688 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_404
timestamp 1679581782
transform 1 0 39360 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_411
timestamp 1679581782
transform 1 0 40032 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_418
timestamp 1679581782
transform 1 0 40704 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_425
timestamp 1679581782
transform 1 0 41376 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_432
timestamp 1679581782
transform 1 0 42048 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_439
timestamp 1679581782
transform 1 0 42720 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_446
timestamp 1679581782
transform 1 0 43392 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_453
timestamp 1679581782
transform 1 0 44064 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_460
timestamp 1679581782
transform 1 0 44736 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_467
timestamp 1679581782
transform 1 0 45408 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_474
timestamp 1679581782
transform 1 0 46080 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_481
timestamp 1679581782
transform 1 0 46752 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_488
timestamp 1679581782
transform 1 0 47424 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_495
timestamp 1679581782
transform 1 0 48096 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_502
timestamp 1679581782
transform 1 0 48768 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_509
timestamp 1679581782
transform 1 0 49440 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_516
timestamp 1679581782
transform 1 0 50112 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_523
timestamp 1679581782
transform 1 0 50784 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_530
timestamp 1679581782
transform 1 0 51456 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_537
timestamp 1679581782
transform 1 0 52128 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_544
timestamp 1679581782
transform 1 0 52800 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_551
timestamp 1679581782
transform 1 0 53472 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_558
timestamp 1679581782
transform 1 0 54144 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_565
timestamp 1679581782
transform 1 0 54816 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_572
timestamp 1679581782
transform 1 0 55488 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_579
timestamp 1679581782
transform 1 0 56160 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_586
timestamp 1679581782
transform 1 0 56832 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_593
timestamp 1679581782
transform 1 0 57504 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_600
timestamp 1679581782
transform 1 0 58176 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_607
timestamp 1679581782
transform 1 0 58848 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_614
timestamp 1679581782
transform 1 0 59520 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_621
timestamp 1679581782
transform 1 0 60192 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_628
timestamp 1679581782
transform 1 0 60864 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_635
timestamp 1679581782
transform 1 0 61536 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_642
timestamp 1679581782
transform 1 0 62208 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_649
timestamp 1679581782
transform 1 0 62880 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_656
timestamp 1679581782
transform 1 0 63552 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_663
timestamp 1679581782
transform 1 0 64224 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_670
timestamp 1679581782
transform 1 0 64896 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_677
timestamp 1679581782
transform 1 0 65568 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_684
timestamp 1679581782
transform 1 0 66240 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_691
timestamp 1679581782
transform 1 0 66912 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_698
timestamp 1679581782
transform 1 0 67584 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_705
timestamp 1679581782
transform 1 0 68256 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_712
timestamp 1679581782
transform 1 0 68928 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_719
timestamp 1679581782
transform 1 0 69600 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_726
timestamp 1679581782
transform 1 0 70272 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_733
timestamp 1679581782
transform 1 0 70944 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_740
timestamp 1679581782
transform 1 0 71616 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_747
timestamp 1679581782
transform 1 0 72288 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_754
timestamp 1679581782
transform 1 0 72960 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_761
timestamp 1679581782
transform 1 0 73632 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_768
timestamp 1679581782
transform 1 0 74304 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_775
timestamp 1679581782
transform 1 0 74976 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_782
timestamp 1679581782
transform 1 0 75648 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_789
timestamp 1679581782
transform 1 0 76320 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_796
timestamp 1679581782
transform 1 0 76992 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_803
timestamp 1679581782
transform 1 0 77664 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_810
timestamp 1679581782
transform 1 0 78336 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_817
timestamp 1679581782
transform 1 0 79008 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_824
timestamp 1679581782
transform 1 0 79680 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_831
timestamp 1679581782
transform 1 0 80352 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_838
timestamp 1679581782
transform 1 0 81024 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_845
timestamp 1679581782
transform 1 0 81696 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_852
timestamp 1679581782
transform 1 0 82368 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_859
timestamp 1679581782
transform 1 0 83040 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_866
timestamp 1679581782
transform 1 0 83712 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_873
timestamp 1679581782
transform 1 0 84384 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_880
timestamp 1679581782
transform 1 0 85056 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_887
timestamp 1679581782
transform 1 0 85728 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_894
timestamp 1679581782
transform 1 0 86400 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_901
timestamp 1679581782
transform 1 0 87072 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_908
timestamp 1679581782
transform 1 0 87744 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_915
timestamp 1679581782
transform 1 0 88416 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_29_922
timestamp 1677580104
transform 1 0 89088 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_924
timestamp 1677579658
transform 1 0 89280 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_4
timestamp 1679581782
transform 1 0 960 0 1 23436
box -48 -56 720 834
use sg13g2_fill_1  FILLER_30_11
timestamp 1677579658
transform 1 0 1632 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_24
timestamp 1679581782
transform 1 0 2880 0 1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_31
timestamp 1679577901
transform 1 0 3552 0 1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_30_35
timestamp 1677579658
transform 1 0 3936 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_40
timestamp 1679581782
transform 1 0 4416 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_47
timestamp 1679581782
transform 1 0 5088 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_54
timestamp 1679581782
transform 1 0 5760 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_61
timestamp 1679581782
transform 1 0 6432 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_68
timestamp 1679581782
transform 1 0 7104 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_75
timestamp 1679581782
transform 1 0 7776 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_82
timestamp 1679581782
transform 1 0 8448 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_89
timestamp 1679581782
transform 1 0 9120 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_96
timestamp 1679581782
transform 1 0 9792 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_103
timestamp 1679581782
transform 1 0 10464 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_114
timestamp 1679581782
transform 1 0 11520 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_121
timestamp 1679581782
transform 1 0 12192 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_128
timestamp 1679581782
transform 1 0 12864 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_135
timestamp 1679581782
transform 1 0 13536 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_142
timestamp 1679581782
transform 1 0 14208 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_149
timestamp 1679581782
transform 1 0 14880 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_156
timestamp 1679581782
transform 1 0 15552 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_163
timestamp 1679581782
transform 1 0 16224 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_170
timestamp 1679581782
transform 1 0 16896 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_177
timestamp 1679581782
transform 1 0 17568 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_184
timestamp 1679581782
transform 1 0 18240 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_191
timestamp 1679581782
transform 1 0 18912 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_198
timestamp 1679581782
transform 1 0 19584 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_205
timestamp 1679581782
transform 1 0 20256 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_212
timestamp 1679581782
transform 1 0 20928 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_219
timestamp 1679581782
transform 1 0 21600 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_226
timestamp 1679581782
transform 1 0 22272 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_233
timestamp 1679581782
transform 1 0 22944 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_240
timestamp 1679581782
transform 1 0 23616 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_247
timestamp 1679581782
transform 1 0 24288 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_254
timestamp 1679581782
transform 1 0 24960 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_261
timestamp 1679581782
transform 1 0 25632 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_268
timestamp 1679581782
transform 1 0 26304 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_275
timestamp 1679581782
transform 1 0 26976 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_282
timestamp 1679581782
transform 1 0 27648 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_289
timestamp 1679581782
transform 1 0 28320 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_296
timestamp 1679581782
transform 1 0 28992 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_303
timestamp 1679581782
transform 1 0 29664 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_310
timestamp 1679581782
transform 1 0 30336 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_317
timestamp 1679581782
transform 1 0 31008 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_324
timestamp 1679581782
transform 1 0 31680 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_331
timestamp 1679581782
transform 1 0 32352 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_338
timestamp 1679581782
transform 1 0 33024 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_345
timestamp 1679581782
transform 1 0 33696 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_352
timestamp 1679581782
transform 1 0 34368 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_359
timestamp 1679581782
transform 1 0 35040 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_366
timestamp 1679581782
transform 1 0 35712 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_373
timestamp 1679581782
transform 1 0 36384 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_380
timestamp 1679581782
transform 1 0 37056 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_387
timestamp 1679581782
transform 1 0 37728 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_394
timestamp 1679581782
transform 1 0 38400 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_401
timestamp 1679581782
transform 1 0 39072 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_408
timestamp 1679581782
transform 1 0 39744 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_415
timestamp 1679581782
transform 1 0 40416 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_422
timestamp 1679581782
transform 1 0 41088 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_429
timestamp 1679581782
transform 1 0 41760 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_436
timestamp 1679581782
transform 1 0 42432 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_443
timestamp 1679581782
transform 1 0 43104 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_450
timestamp 1679581782
transform 1 0 43776 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_457
timestamp 1679581782
transform 1 0 44448 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_464
timestamp 1679581782
transform 1 0 45120 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_471
timestamp 1679581782
transform 1 0 45792 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_478
timestamp 1679581782
transform 1 0 46464 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_485
timestamp 1679581782
transform 1 0 47136 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_492
timestamp 1679581782
transform 1 0 47808 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_499
timestamp 1679581782
transform 1 0 48480 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_506
timestamp 1679581782
transform 1 0 49152 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_513
timestamp 1679581782
transform 1 0 49824 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_520
timestamp 1679581782
transform 1 0 50496 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_527
timestamp 1679581782
transform 1 0 51168 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_534
timestamp 1679581782
transform 1 0 51840 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_541
timestamp 1679581782
transform 1 0 52512 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_548
timestamp 1679581782
transform 1 0 53184 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_555
timestamp 1679581782
transform 1 0 53856 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_562
timestamp 1679581782
transform 1 0 54528 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_569
timestamp 1679581782
transform 1 0 55200 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_576
timestamp 1679581782
transform 1 0 55872 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_583
timestamp 1679581782
transform 1 0 56544 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_590
timestamp 1679581782
transform 1 0 57216 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_597
timestamp 1679581782
transform 1 0 57888 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_604
timestamp 1679581782
transform 1 0 58560 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_611
timestamp 1679581782
transform 1 0 59232 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_618
timestamp 1679581782
transform 1 0 59904 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_625
timestamp 1679581782
transform 1 0 60576 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_632
timestamp 1679581782
transform 1 0 61248 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_639
timestamp 1679581782
transform 1 0 61920 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_646
timestamp 1679581782
transform 1 0 62592 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_653
timestamp 1679581782
transform 1 0 63264 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_660
timestamp 1679581782
transform 1 0 63936 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_667
timestamp 1679581782
transform 1 0 64608 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_674
timestamp 1679581782
transform 1 0 65280 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_681
timestamp 1679581782
transform 1 0 65952 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_688
timestamp 1679581782
transform 1 0 66624 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_695
timestamp 1679581782
transform 1 0 67296 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_702
timestamp 1679581782
transform 1 0 67968 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_709
timestamp 1679581782
transform 1 0 68640 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_716
timestamp 1679581782
transform 1 0 69312 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_723
timestamp 1679581782
transform 1 0 69984 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_730
timestamp 1679581782
transform 1 0 70656 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_737
timestamp 1679581782
transform 1 0 71328 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_744
timestamp 1679581782
transform 1 0 72000 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_751
timestamp 1679581782
transform 1 0 72672 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_758
timestamp 1679581782
transform 1 0 73344 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_765
timestamp 1679581782
transform 1 0 74016 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_772
timestamp 1679581782
transform 1 0 74688 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_779
timestamp 1679581782
transform 1 0 75360 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_786
timestamp 1679581782
transform 1 0 76032 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_793
timestamp 1679581782
transform 1 0 76704 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_800
timestamp 1679581782
transform 1 0 77376 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_807
timestamp 1679581782
transform 1 0 78048 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_814
timestamp 1679581782
transform 1 0 78720 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_821
timestamp 1679581782
transform 1 0 79392 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_828
timestamp 1679581782
transform 1 0 80064 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_835
timestamp 1679581782
transform 1 0 80736 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_842
timestamp 1679581782
transform 1 0 81408 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_849
timestamp 1679581782
transform 1 0 82080 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_856
timestamp 1679581782
transform 1 0 82752 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_863
timestamp 1679581782
transform 1 0 83424 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_870
timestamp 1679581782
transform 1 0 84096 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_877
timestamp 1679581782
transform 1 0 84768 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_884
timestamp 1679581782
transform 1 0 85440 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_891
timestamp 1679581782
transform 1 0 86112 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_898
timestamp 1679581782
transform 1 0 86784 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_905
timestamp 1679581782
transform 1 0 87456 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_912
timestamp 1679581782
transform 1 0 88128 0 1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_919
timestamp 1679577901
transform 1 0 88800 0 1 23436
box -48 -56 432 834
use sg13g2_fill_2  FILLER_30_923
timestamp 1677580104
transform 1 0 89184 0 1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_31_4
timestamp 1679581782
transform 1 0 960 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_11
timestamp 1679581782
transform 1 0 1632 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_18
timestamp 1679581782
transform 1 0 2304 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_25
timestamp 1679581782
transform 1 0 2976 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_31_32
timestamp 1679577901
transform 1 0 3648 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_40
timestamp 1677580104
transform 1 0 4416 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_31_45
timestamp 1677580104
transform 1 0 4896 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_47
timestamp 1677579658
transform 1 0 5088 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_31_56
timestamp 1677580104
transform 1 0 5952 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_58
timestamp 1677579658
transform 1 0 6144 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_67
timestamp 1679581782
transform 1 0 7008 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_74
timestamp 1679581782
transform 1 0 7680 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_81
timestamp 1679581782
transform 1 0 8352 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_88
timestamp 1679581782
transform 1 0 9024 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_31_100
timestamp 1679577901
transform 1 0 10176 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_104
timestamp 1677580104
transform 1 0 10560 0 -1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_31_111
timestamp 1679581782
transform 1 0 11232 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_122
timestamp 1679581782
transform 1 0 12288 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_129
timestamp 1679581782
transform 1 0 12960 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_136
timestamp 1679581782
transform 1 0 13632 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_143
timestamp 1679581782
transform 1 0 14304 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_150
timestamp 1679581782
transform 1 0 14976 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_157
timestamp 1679581782
transform 1 0 15648 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_164
timestamp 1679581782
transform 1 0 16320 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_171
timestamp 1679581782
transform 1 0 16992 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_178
timestamp 1679581782
transform 1 0 17664 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_185
timestamp 1679581782
transform 1 0 18336 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_192
timestamp 1679581782
transform 1 0 19008 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_199
timestamp 1679581782
transform 1 0 19680 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_206
timestamp 1679581782
transform 1 0 20352 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_213
timestamp 1679581782
transform 1 0 21024 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_220
timestamp 1679581782
transform 1 0 21696 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_227
timestamp 1679581782
transform 1 0 22368 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_234
timestamp 1679581782
transform 1 0 23040 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_241
timestamp 1679581782
transform 1 0 23712 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_248
timestamp 1679581782
transform 1 0 24384 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_255
timestamp 1679581782
transform 1 0 25056 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_262
timestamp 1679581782
transform 1 0 25728 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_269
timestamp 1679581782
transform 1 0 26400 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_276
timestamp 1679581782
transform 1 0 27072 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_283
timestamp 1679581782
transform 1 0 27744 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_290
timestamp 1679581782
transform 1 0 28416 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_297
timestamp 1679581782
transform 1 0 29088 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_304
timestamp 1679581782
transform 1 0 29760 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_311
timestamp 1679581782
transform 1 0 30432 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_318
timestamp 1679581782
transform 1 0 31104 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_325
timestamp 1679581782
transform 1 0 31776 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_332
timestamp 1679581782
transform 1 0 32448 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_339
timestamp 1679581782
transform 1 0 33120 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_346
timestamp 1679581782
transform 1 0 33792 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_353
timestamp 1679581782
transform 1 0 34464 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_360
timestamp 1679581782
transform 1 0 35136 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_367
timestamp 1679581782
transform 1 0 35808 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_374
timestamp 1679581782
transform 1 0 36480 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_381
timestamp 1679581782
transform 1 0 37152 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_388
timestamp 1679581782
transform 1 0 37824 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_395
timestamp 1679581782
transform 1 0 38496 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_402
timestamp 1679581782
transform 1 0 39168 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_409
timestamp 1679581782
transform 1 0 39840 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_416
timestamp 1679581782
transform 1 0 40512 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_423
timestamp 1679581782
transform 1 0 41184 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_430
timestamp 1679581782
transform 1 0 41856 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_437
timestamp 1679581782
transform 1 0 42528 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_444
timestamp 1679581782
transform 1 0 43200 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_451
timestamp 1679581782
transform 1 0 43872 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_458
timestamp 1679581782
transform 1 0 44544 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_465
timestamp 1679581782
transform 1 0 45216 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_472
timestamp 1679581782
transform 1 0 45888 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_479
timestamp 1679581782
transform 1 0 46560 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_486
timestamp 1679581782
transform 1 0 47232 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_493
timestamp 1679581782
transform 1 0 47904 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_500
timestamp 1679581782
transform 1 0 48576 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_507
timestamp 1679581782
transform 1 0 49248 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_514
timestamp 1679581782
transform 1 0 49920 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_521
timestamp 1679581782
transform 1 0 50592 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_528
timestamp 1679581782
transform 1 0 51264 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_535
timestamp 1679581782
transform 1 0 51936 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_542
timestamp 1679581782
transform 1 0 52608 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_549
timestamp 1679581782
transform 1 0 53280 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_556
timestamp 1679581782
transform 1 0 53952 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_563
timestamp 1679581782
transform 1 0 54624 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_570
timestamp 1679581782
transform 1 0 55296 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_577
timestamp 1679581782
transform 1 0 55968 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_584
timestamp 1679581782
transform 1 0 56640 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_591
timestamp 1679581782
transform 1 0 57312 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_598
timestamp 1679581782
transform 1 0 57984 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_605
timestamp 1679581782
transform 1 0 58656 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_612
timestamp 1679581782
transform 1 0 59328 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_619
timestamp 1679581782
transform 1 0 60000 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_626
timestamp 1679581782
transform 1 0 60672 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_633
timestamp 1679581782
transform 1 0 61344 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_640
timestamp 1679581782
transform 1 0 62016 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_647
timestamp 1679581782
transform 1 0 62688 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_654
timestamp 1679581782
transform 1 0 63360 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_661
timestamp 1679581782
transform 1 0 64032 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_668
timestamp 1679581782
transform 1 0 64704 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_675
timestamp 1679581782
transform 1 0 65376 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_682
timestamp 1679581782
transform 1 0 66048 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_689
timestamp 1679581782
transform 1 0 66720 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_696
timestamp 1679581782
transform 1 0 67392 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_703
timestamp 1679581782
transform 1 0 68064 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_710
timestamp 1679581782
transform 1 0 68736 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_717
timestamp 1679581782
transform 1 0 69408 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_724
timestamp 1679581782
transform 1 0 70080 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_731
timestamp 1679581782
transform 1 0 70752 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_738
timestamp 1679581782
transform 1 0 71424 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_745
timestamp 1679581782
transform 1 0 72096 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_752
timestamp 1679581782
transform 1 0 72768 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_759
timestamp 1679581782
transform 1 0 73440 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_766
timestamp 1679581782
transform 1 0 74112 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_773
timestamp 1679581782
transform 1 0 74784 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_780
timestamp 1679581782
transform 1 0 75456 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_787
timestamp 1679581782
transform 1 0 76128 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_794
timestamp 1679581782
transform 1 0 76800 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_801
timestamp 1679581782
transform 1 0 77472 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_808
timestamp 1679581782
transform 1 0 78144 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_815
timestamp 1679581782
transform 1 0 78816 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_822
timestamp 1679581782
transform 1 0 79488 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_829
timestamp 1679581782
transform 1 0 80160 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_836
timestamp 1679581782
transform 1 0 80832 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_843
timestamp 1679581782
transform 1 0 81504 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_850
timestamp 1679581782
transform 1 0 82176 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_857
timestamp 1679581782
transform 1 0 82848 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_864
timestamp 1679581782
transform 1 0 83520 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_871
timestamp 1679581782
transform 1 0 84192 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_878
timestamp 1679581782
transform 1 0 84864 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_885
timestamp 1679581782
transform 1 0 85536 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_892
timestamp 1679581782
transform 1 0 86208 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_899
timestamp 1679581782
transform 1 0 86880 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_906
timestamp 1679581782
transform 1 0 87552 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_913
timestamp 1679581782
transform 1 0 88224 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_31_920
timestamp 1679577901
transform 1 0 88896 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_31_924
timestamp 1677579658
transform 1 0 89280 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_4
timestamp 1679581782
transform 1 0 960 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_11
timestamp 1679581782
transform 1 0 1632 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_18
timestamp 1679581782
transform 1 0 2304 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_25
timestamp 1679581782
transform 1 0 2976 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_32
timestamp 1679581782
transform 1 0 3648 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_39
timestamp 1679581782
transform 1 0 4320 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_46
timestamp 1679581782
transform 1 0 4992 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_53
timestamp 1679581782
transform 1 0 5664 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_60
timestamp 1679581782
transform 1 0 6336 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_67
timestamp 1679581782
transform 1 0 7008 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_74
timestamp 1679581782
transform 1 0 7680 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_81
timestamp 1679581782
transform 1 0 8352 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_88
timestamp 1679581782
transform 1 0 9024 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_95
timestamp 1679581782
transform 1 0 9696 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_102
timestamp 1679581782
transform 1 0 10368 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_109
timestamp 1679581782
transform 1 0 11040 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_116
timestamp 1679577901
transform 1 0 11712 0 1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_32_120
timestamp 1677580104
transform 1 0 12096 0 1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_32_130
timestamp 1679581782
transform 1 0 13056 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_137
timestamp 1679581782
transform 1 0 13728 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_144
timestamp 1679581782
transform 1 0 14400 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_151
timestamp 1679581782
transform 1 0 15072 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_158
timestamp 1679581782
transform 1 0 15744 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_165
timestamp 1679581782
transform 1 0 16416 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_172
timestamp 1679581782
transform 1 0 17088 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_179
timestamp 1679581782
transform 1 0 17760 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_186
timestamp 1679581782
transform 1 0 18432 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_193
timestamp 1679581782
transform 1 0 19104 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_200
timestamp 1679581782
transform 1 0 19776 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_207
timestamp 1679581782
transform 1 0 20448 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_214
timestamp 1679581782
transform 1 0 21120 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_221
timestamp 1679581782
transform 1 0 21792 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_228
timestamp 1679581782
transform 1 0 22464 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_235
timestamp 1679581782
transform 1 0 23136 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_242
timestamp 1679581782
transform 1 0 23808 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_249
timestamp 1679581782
transform 1 0 24480 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_256
timestamp 1679581782
transform 1 0 25152 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_263
timestamp 1679581782
transform 1 0 25824 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_270
timestamp 1679581782
transform 1 0 26496 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_277
timestamp 1679581782
transform 1 0 27168 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_284
timestamp 1679581782
transform 1 0 27840 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_291
timestamp 1679581782
transform 1 0 28512 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_298
timestamp 1679581782
transform 1 0 29184 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_305
timestamp 1679581782
transform 1 0 29856 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_312
timestamp 1679581782
transform 1 0 30528 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_319
timestamp 1679581782
transform 1 0 31200 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_326
timestamp 1679581782
transform 1 0 31872 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_333
timestamp 1679581782
transform 1 0 32544 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_340
timestamp 1679581782
transform 1 0 33216 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_347
timestamp 1679581782
transform 1 0 33888 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_354
timestamp 1679581782
transform 1 0 34560 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_361
timestamp 1679581782
transform 1 0 35232 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_368
timestamp 1679581782
transform 1 0 35904 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_375
timestamp 1679581782
transform 1 0 36576 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_382
timestamp 1679581782
transform 1 0 37248 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_389
timestamp 1679581782
transform 1 0 37920 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_396
timestamp 1679581782
transform 1 0 38592 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_403
timestamp 1679581782
transform 1 0 39264 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_410
timestamp 1679581782
transform 1 0 39936 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_417
timestamp 1679581782
transform 1 0 40608 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_424
timestamp 1679581782
transform 1 0 41280 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_431
timestamp 1679581782
transform 1 0 41952 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_438
timestamp 1679581782
transform 1 0 42624 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_445
timestamp 1679581782
transform 1 0 43296 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_452
timestamp 1679581782
transform 1 0 43968 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_459
timestamp 1679581782
transform 1 0 44640 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_466
timestamp 1679581782
transform 1 0 45312 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_473
timestamp 1679581782
transform 1 0 45984 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_480
timestamp 1679581782
transform 1 0 46656 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_487
timestamp 1679581782
transform 1 0 47328 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_494
timestamp 1679581782
transform 1 0 48000 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_501
timestamp 1679581782
transform 1 0 48672 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_508
timestamp 1679581782
transform 1 0 49344 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_515
timestamp 1679581782
transform 1 0 50016 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_522
timestamp 1679581782
transform 1 0 50688 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_529
timestamp 1679581782
transform 1 0 51360 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_536
timestamp 1679581782
transform 1 0 52032 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_543
timestamp 1679581782
transform 1 0 52704 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_550
timestamp 1679581782
transform 1 0 53376 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_557
timestamp 1679581782
transform 1 0 54048 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_564
timestamp 1679581782
transform 1 0 54720 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_571
timestamp 1679581782
transform 1 0 55392 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_578
timestamp 1679581782
transform 1 0 56064 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_585
timestamp 1679581782
transform 1 0 56736 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_592
timestamp 1679581782
transform 1 0 57408 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_599
timestamp 1679581782
transform 1 0 58080 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_606
timestamp 1679581782
transform 1 0 58752 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_613
timestamp 1679581782
transform 1 0 59424 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_620
timestamp 1679581782
transform 1 0 60096 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_627
timestamp 1679581782
transform 1 0 60768 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_634
timestamp 1679581782
transform 1 0 61440 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_641
timestamp 1679581782
transform 1 0 62112 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_648
timestamp 1679581782
transform 1 0 62784 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_655
timestamp 1679581782
transform 1 0 63456 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_662
timestamp 1679581782
transform 1 0 64128 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_669
timestamp 1679581782
transform 1 0 64800 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_676
timestamp 1679581782
transform 1 0 65472 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_683
timestamp 1679581782
transform 1 0 66144 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_690
timestamp 1679581782
transform 1 0 66816 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_697
timestamp 1679581782
transform 1 0 67488 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_704
timestamp 1679581782
transform 1 0 68160 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_711
timestamp 1679581782
transform 1 0 68832 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_718
timestamp 1679581782
transform 1 0 69504 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_725
timestamp 1679581782
transform 1 0 70176 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_732
timestamp 1679581782
transform 1 0 70848 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_739
timestamp 1679581782
transform 1 0 71520 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_746
timestamp 1679581782
transform 1 0 72192 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_753
timestamp 1679581782
transform 1 0 72864 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_760
timestamp 1679581782
transform 1 0 73536 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_767
timestamp 1679581782
transform 1 0 74208 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_774
timestamp 1679581782
transform 1 0 74880 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_781
timestamp 1679581782
transform 1 0 75552 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_788
timestamp 1679581782
transform 1 0 76224 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_795
timestamp 1679581782
transform 1 0 76896 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_802
timestamp 1679581782
transform 1 0 77568 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_809
timestamp 1679581782
transform 1 0 78240 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_816
timestamp 1679581782
transform 1 0 78912 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_823
timestamp 1679581782
transform 1 0 79584 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_830
timestamp 1679581782
transform 1 0 80256 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_837
timestamp 1679581782
transform 1 0 80928 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_844
timestamp 1679581782
transform 1 0 81600 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_851
timestamp 1679581782
transform 1 0 82272 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_858
timestamp 1679581782
transform 1 0 82944 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_865
timestamp 1679581782
transform 1 0 83616 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_872
timestamp 1679581782
transform 1 0 84288 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_879
timestamp 1679581782
transform 1 0 84960 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_886
timestamp 1679581782
transform 1 0 85632 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_893
timestamp 1679581782
transform 1 0 86304 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_900
timestamp 1679581782
transform 1 0 86976 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_907
timestamp 1679581782
transform 1 0 87648 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_914
timestamp 1679581782
transform 1 0 88320 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_921
timestamp 1679577901
transform 1 0 88992 0 1 24948
box -48 -56 432 834
use sg13g2_decap_8  FILLER_33_4
timestamp 1679581782
transform 1 0 960 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_11
timestamp 1679581782
transform 1 0 1632 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_18
timestamp 1679581782
transform 1 0 2304 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_25
timestamp 1679577901
transform 1 0 2976 0 -1 26460
box -48 -56 432 834
use sg13g2_decap_8  FILLER_33_33
timestamp 1679581782
transform 1 0 3744 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_40
timestamp 1679581782
transform 1 0 4416 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_51
timestamp 1679581782
transform 1 0 5472 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_58
timestamp 1679581782
transform 1 0 6144 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_65
timestamp 1679581782
transform 1 0 6816 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_72
timestamp 1679581782
transform 1 0 7488 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_79
timestamp 1679581782
transform 1 0 8160 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_86
timestamp 1679581782
transform 1 0 8832 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_93
timestamp 1679581782
transform 1 0 9504 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_100
timestamp 1679581782
transform 1 0 10176 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_33_107
timestamp 1677580104
transform 1 0 10848 0 -1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_33_114
timestamp 1679581782
transform 1 0 11520 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_121
timestamp 1679581782
transform 1 0 12192 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_128
timestamp 1679581782
transform 1 0 12864 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_135
timestamp 1679581782
transform 1 0 13536 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_142
timestamp 1679581782
transform 1 0 14208 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_149
timestamp 1679581782
transform 1 0 14880 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_156
timestamp 1679581782
transform 1 0 15552 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_163
timestamp 1679581782
transform 1 0 16224 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_170
timestamp 1679581782
transform 1 0 16896 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_177
timestamp 1679581782
transform 1 0 17568 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_184
timestamp 1679581782
transform 1 0 18240 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_191
timestamp 1679581782
transform 1 0 18912 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_198
timestamp 1679581782
transform 1 0 19584 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_205
timestamp 1679581782
transform 1 0 20256 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_212
timestamp 1679581782
transform 1 0 20928 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_219
timestamp 1679581782
transform 1 0 21600 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_226
timestamp 1679581782
transform 1 0 22272 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_233
timestamp 1679581782
transform 1 0 22944 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_240
timestamp 1679581782
transform 1 0 23616 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_247
timestamp 1679581782
transform 1 0 24288 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_254
timestamp 1679581782
transform 1 0 24960 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_261
timestamp 1679581782
transform 1 0 25632 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_268
timestamp 1679581782
transform 1 0 26304 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_275
timestamp 1679581782
transform 1 0 26976 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_282
timestamp 1679581782
transform 1 0 27648 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_289
timestamp 1679581782
transform 1 0 28320 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_296
timestamp 1679581782
transform 1 0 28992 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_303
timestamp 1679581782
transform 1 0 29664 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_310
timestamp 1679581782
transform 1 0 30336 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_317
timestamp 1679581782
transform 1 0 31008 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_324
timestamp 1679581782
transform 1 0 31680 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_331
timestamp 1679581782
transform 1 0 32352 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_338
timestamp 1679581782
transform 1 0 33024 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_345
timestamp 1679581782
transform 1 0 33696 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_352
timestamp 1679581782
transform 1 0 34368 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_359
timestamp 1679581782
transform 1 0 35040 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_366
timestamp 1679581782
transform 1 0 35712 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_373
timestamp 1679581782
transform 1 0 36384 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_380
timestamp 1679581782
transform 1 0 37056 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_387
timestamp 1679581782
transform 1 0 37728 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_394
timestamp 1679581782
transform 1 0 38400 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_401
timestamp 1679581782
transform 1 0 39072 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_408
timestamp 1679581782
transform 1 0 39744 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_415
timestamp 1679581782
transform 1 0 40416 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_422
timestamp 1679581782
transform 1 0 41088 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_429
timestamp 1679581782
transform 1 0 41760 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_436
timestamp 1679581782
transform 1 0 42432 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_443
timestamp 1679581782
transform 1 0 43104 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_450
timestamp 1679581782
transform 1 0 43776 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_457
timestamp 1679581782
transform 1 0 44448 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_464
timestamp 1679581782
transform 1 0 45120 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_471
timestamp 1679581782
transform 1 0 45792 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_478
timestamp 1679581782
transform 1 0 46464 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_485
timestamp 1679581782
transform 1 0 47136 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_492
timestamp 1679581782
transform 1 0 47808 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_499
timestamp 1679581782
transform 1 0 48480 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_506
timestamp 1679581782
transform 1 0 49152 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_513
timestamp 1679581782
transform 1 0 49824 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_520
timestamp 1679581782
transform 1 0 50496 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_527
timestamp 1679581782
transform 1 0 51168 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_534
timestamp 1679581782
transform 1 0 51840 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_541
timestamp 1679581782
transform 1 0 52512 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_548
timestamp 1679581782
transform 1 0 53184 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_555
timestamp 1679581782
transform 1 0 53856 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_562
timestamp 1679581782
transform 1 0 54528 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_569
timestamp 1679581782
transform 1 0 55200 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_576
timestamp 1679581782
transform 1 0 55872 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_583
timestamp 1679581782
transform 1 0 56544 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_590
timestamp 1679581782
transform 1 0 57216 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_597
timestamp 1679581782
transform 1 0 57888 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_604
timestamp 1679581782
transform 1 0 58560 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_611
timestamp 1679581782
transform 1 0 59232 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_618
timestamp 1679581782
transform 1 0 59904 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_625
timestamp 1679581782
transform 1 0 60576 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_632
timestamp 1679581782
transform 1 0 61248 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_639
timestamp 1679581782
transform 1 0 61920 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_646
timestamp 1679581782
transform 1 0 62592 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_653
timestamp 1679581782
transform 1 0 63264 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_660
timestamp 1679581782
transform 1 0 63936 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_667
timestamp 1679581782
transform 1 0 64608 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_674
timestamp 1679581782
transform 1 0 65280 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_681
timestamp 1679581782
transform 1 0 65952 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_688
timestamp 1679581782
transform 1 0 66624 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_695
timestamp 1679581782
transform 1 0 67296 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_702
timestamp 1679581782
transform 1 0 67968 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_709
timestamp 1679581782
transform 1 0 68640 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_716
timestamp 1679581782
transform 1 0 69312 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_723
timestamp 1679581782
transform 1 0 69984 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_730
timestamp 1679581782
transform 1 0 70656 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_737
timestamp 1679581782
transform 1 0 71328 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_744
timestamp 1679581782
transform 1 0 72000 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_751
timestamp 1679581782
transform 1 0 72672 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_758
timestamp 1679581782
transform 1 0 73344 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_765
timestamp 1679581782
transform 1 0 74016 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_772
timestamp 1679581782
transform 1 0 74688 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_779
timestamp 1679581782
transform 1 0 75360 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_786
timestamp 1679581782
transform 1 0 76032 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_793
timestamp 1679581782
transform 1 0 76704 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_800
timestamp 1679581782
transform 1 0 77376 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_807
timestamp 1679581782
transform 1 0 78048 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_814
timestamp 1679581782
transform 1 0 78720 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_821
timestamp 1679581782
transform 1 0 79392 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_828
timestamp 1679581782
transform 1 0 80064 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_835
timestamp 1679581782
transform 1 0 80736 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_842
timestamp 1679581782
transform 1 0 81408 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_849
timestamp 1679581782
transform 1 0 82080 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_856
timestamp 1679581782
transform 1 0 82752 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_863
timestamp 1679581782
transform 1 0 83424 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_870
timestamp 1679581782
transform 1 0 84096 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_877
timestamp 1679581782
transform 1 0 84768 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_884
timestamp 1679581782
transform 1 0 85440 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_891
timestamp 1679581782
transform 1 0 86112 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_898
timestamp 1679581782
transform 1 0 86784 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_905
timestamp 1679581782
transform 1 0 87456 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_912
timestamp 1679581782
transform 1 0 88128 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_919
timestamp 1679577901
transform 1 0 88800 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_33_923
timestamp 1677580104
transform 1 0 89184 0 -1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_34_4
timestamp 1679581782
transform 1 0 960 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_11
timestamp 1679581782
transform 1 0 1632 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_18
timestamp 1679581782
transform 1 0 2304 0 1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_34_25
timestamp 1679577901
transform 1 0 2976 0 1 26460
box -48 -56 432 834
use sg13g2_decap_8  FILLER_34_49
timestamp 1679581782
transform 1 0 5280 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_56
timestamp 1679581782
transform 1 0 5952 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_63
timestamp 1679581782
transform 1 0 6624 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_70
timestamp 1679581782
transform 1 0 7296 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_77
timestamp 1679581782
transform 1 0 7968 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_84
timestamp 1679581782
transform 1 0 8640 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_91
timestamp 1679581782
transform 1 0 9312 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_98
timestamp 1679581782
transform 1 0 9984 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_118
timestamp 1679581782
transform 1 0 11904 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_125
timestamp 1679581782
transform 1 0 12576 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_132
timestamp 1679581782
transform 1 0 13248 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_139
timestamp 1679581782
transform 1 0 13920 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_146
timestamp 1679581782
transform 1 0 14592 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_153
timestamp 1679581782
transform 1 0 15264 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_160
timestamp 1679581782
transform 1 0 15936 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_167
timestamp 1679581782
transform 1 0 16608 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_174
timestamp 1679581782
transform 1 0 17280 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_181
timestamp 1679581782
transform 1 0 17952 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_188
timestamp 1679581782
transform 1 0 18624 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_195
timestamp 1679581782
transform 1 0 19296 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_202
timestamp 1679581782
transform 1 0 19968 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_209
timestamp 1679581782
transform 1 0 20640 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_216
timestamp 1679581782
transform 1 0 21312 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_223
timestamp 1679581782
transform 1 0 21984 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_230
timestamp 1679581782
transform 1 0 22656 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_237
timestamp 1679581782
transform 1 0 23328 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_244
timestamp 1679581782
transform 1 0 24000 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_251
timestamp 1679581782
transform 1 0 24672 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_258
timestamp 1679581782
transform 1 0 25344 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_265
timestamp 1679581782
transform 1 0 26016 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_272
timestamp 1679581782
transform 1 0 26688 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_279
timestamp 1679581782
transform 1 0 27360 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_286
timestamp 1679581782
transform 1 0 28032 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_293
timestamp 1679581782
transform 1 0 28704 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_300
timestamp 1679581782
transform 1 0 29376 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_307
timestamp 1679581782
transform 1 0 30048 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_314
timestamp 1679581782
transform 1 0 30720 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_321
timestamp 1679581782
transform 1 0 31392 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_328
timestamp 1679581782
transform 1 0 32064 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_335
timestamp 1679581782
transform 1 0 32736 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_342
timestamp 1679581782
transform 1 0 33408 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_349
timestamp 1679581782
transform 1 0 34080 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_356
timestamp 1679581782
transform 1 0 34752 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_363
timestamp 1679581782
transform 1 0 35424 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_370
timestamp 1679581782
transform 1 0 36096 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_377
timestamp 1679581782
transform 1 0 36768 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_384
timestamp 1679581782
transform 1 0 37440 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_391
timestamp 1679581782
transform 1 0 38112 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_398
timestamp 1679581782
transform 1 0 38784 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_405
timestamp 1679581782
transform 1 0 39456 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_412
timestamp 1679581782
transform 1 0 40128 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_419
timestamp 1679581782
transform 1 0 40800 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_426
timestamp 1679581782
transform 1 0 41472 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_433
timestamp 1679581782
transform 1 0 42144 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_440
timestamp 1679581782
transform 1 0 42816 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_447
timestamp 1679581782
transform 1 0 43488 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_454
timestamp 1679581782
transform 1 0 44160 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_461
timestamp 1679581782
transform 1 0 44832 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_468
timestamp 1679581782
transform 1 0 45504 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_475
timestamp 1679581782
transform 1 0 46176 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_482
timestamp 1679581782
transform 1 0 46848 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_489
timestamp 1679581782
transform 1 0 47520 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_496
timestamp 1679581782
transform 1 0 48192 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_503
timestamp 1679581782
transform 1 0 48864 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_510
timestamp 1679581782
transform 1 0 49536 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_517
timestamp 1679581782
transform 1 0 50208 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_524
timestamp 1679581782
transform 1 0 50880 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_531
timestamp 1679581782
transform 1 0 51552 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_538
timestamp 1679581782
transform 1 0 52224 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_545
timestamp 1679581782
transform 1 0 52896 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_552
timestamp 1679581782
transform 1 0 53568 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_559
timestamp 1679581782
transform 1 0 54240 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_566
timestamp 1679581782
transform 1 0 54912 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_573
timestamp 1679581782
transform 1 0 55584 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_580
timestamp 1679581782
transform 1 0 56256 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_587
timestamp 1679581782
transform 1 0 56928 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_594
timestamp 1679581782
transform 1 0 57600 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_601
timestamp 1679581782
transform 1 0 58272 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_608
timestamp 1679581782
transform 1 0 58944 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_615
timestamp 1679581782
transform 1 0 59616 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_622
timestamp 1679581782
transform 1 0 60288 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_629
timestamp 1679581782
transform 1 0 60960 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_636
timestamp 1679581782
transform 1 0 61632 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_643
timestamp 1679581782
transform 1 0 62304 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_650
timestamp 1679581782
transform 1 0 62976 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_657
timestamp 1679581782
transform 1 0 63648 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_664
timestamp 1679581782
transform 1 0 64320 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_671
timestamp 1679581782
transform 1 0 64992 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_678
timestamp 1679581782
transform 1 0 65664 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_685
timestamp 1679581782
transform 1 0 66336 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_692
timestamp 1679581782
transform 1 0 67008 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_699
timestamp 1679581782
transform 1 0 67680 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_706
timestamp 1679581782
transform 1 0 68352 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_713
timestamp 1679581782
transform 1 0 69024 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_720
timestamp 1679581782
transform 1 0 69696 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_727
timestamp 1679581782
transform 1 0 70368 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_734
timestamp 1679581782
transform 1 0 71040 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_741
timestamp 1679581782
transform 1 0 71712 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_748
timestamp 1679581782
transform 1 0 72384 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_755
timestamp 1679581782
transform 1 0 73056 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_762
timestamp 1679581782
transform 1 0 73728 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_769
timestamp 1679581782
transform 1 0 74400 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_776
timestamp 1679581782
transform 1 0 75072 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_783
timestamp 1679581782
transform 1 0 75744 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_790
timestamp 1679581782
transform 1 0 76416 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_797
timestamp 1679581782
transform 1 0 77088 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_804
timestamp 1679581782
transform 1 0 77760 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_811
timestamp 1679581782
transform 1 0 78432 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_818
timestamp 1679581782
transform 1 0 79104 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_825
timestamp 1679581782
transform 1 0 79776 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_832
timestamp 1679581782
transform 1 0 80448 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_839
timestamp 1679581782
transform 1 0 81120 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_846
timestamp 1679581782
transform 1 0 81792 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_853
timestamp 1679581782
transform 1 0 82464 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_860
timestamp 1679581782
transform 1 0 83136 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_867
timestamp 1679581782
transform 1 0 83808 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_874
timestamp 1679581782
transform 1 0 84480 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_881
timestamp 1679581782
transform 1 0 85152 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_888
timestamp 1679581782
transform 1 0 85824 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_895
timestamp 1679581782
transform 1 0 86496 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_902
timestamp 1679581782
transform 1 0 87168 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_909
timestamp 1679581782
transform 1 0 87840 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_916
timestamp 1679581782
transform 1 0 88512 0 1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_34_923
timestamp 1677580104
transform 1 0 89184 0 1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_35_4
timestamp 1679581782
transform 1 0 960 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_11
timestamp 1679581782
transform 1 0 1632 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_18
timestamp 1679581782
transform 1 0 2304 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_25
timestamp 1679581782
transform 1 0 2976 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_32
timestamp 1679581782
transform 1 0 3648 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_39
timestamp 1679581782
transform 1 0 4320 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_46
timestamp 1679581782
transform 1 0 4992 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_53
timestamp 1679581782
transform 1 0 5664 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_60
timestamp 1679581782
transform 1 0 6336 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_67
timestamp 1679581782
transform 1 0 7008 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_74
timestamp 1679581782
transform 1 0 7680 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_81
timestamp 1679581782
transform 1 0 8352 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_88
timestamp 1679581782
transform 1 0 9024 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_95
timestamp 1679581782
transform 1 0 9696 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_102
timestamp 1679581782
transform 1 0 10368 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_114
timestamp 1679581782
transform 1 0 11520 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_121
timestamp 1679581782
transform 1 0 12192 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_128
timestamp 1679581782
transform 1 0 12864 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_135
timestamp 1679581782
transform 1 0 13536 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_142
timestamp 1679581782
transform 1 0 14208 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_149
timestamp 1679581782
transform 1 0 14880 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_156
timestamp 1679581782
transform 1 0 15552 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_163
timestamp 1679581782
transform 1 0 16224 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_170
timestamp 1679581782
transform 1 0 16896 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_177
timestamp 1679581782
transform 1 0 17568 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_184
timestamp 1679581782
transform 1 0 18240 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_191
timestamp 1679581782
transform 1 0 18912 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_198
timestamp 1679581782
transform 1 0 19584 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_205
timestamp 1679581782
transform 1 0 20256 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_212
timestamp 1679581782
transform 1 0 20928 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_219
timestamp 1679581782
transform 1 0 21600 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_226
timestamp 1679581782
transform 1 0 22272 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_233
timestamp 1679581782
transform 1 0 22944 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_240
timestamp 1679581782
transform 1 0 23616 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_247
timestamp 1679581782
transform 1 0 24288 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_254
timestamp 1679581782
transform 1 0 24960 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_261
timestamp 1679581782
transform 1 0 25632 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_268
timestamp 1679581782
transform 1 0 26304 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_275
timestamp 1679581782
transform 1 0 26976 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_282
timestamp 1679581782
transform 1 0 27648 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_289
timestamp 1679581782
transform 1 0 28320 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_296
timestamp 1679581782
transform 1 0 28992 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_303
timestamp 1679581782
transform 1 0 29664 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_310
timestamp 1679581782
transform 1 0 30336 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_317
timestamp 1679581782
transform 1 0 31008 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_324
timestamp 1679581782
transform 1 0 31680 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_331
timestamp 1679581782
transform 1 0 32352 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_338
timestamp 1679581782
transform 1 0 33024 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_345
timestamp 1679581782
transform 1 0 33696 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_352
timestamp 1679581782
transform 1 0 34368 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_359
timestamp 1679581782
transform 1 0 35040 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_366
timestamp 1679581782
transform 1 0 35712 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_373
timestamp 1679581782
transform 1 0 36384 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_380
timestamp 1679581782
transform 1 0 37056 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_387
timestamp 1679581782
transform 1 0 37728 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_394
timestamp 1679581782
transform 1 0 38400 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_401
timestamp 1679581782
transform 1 0 39072 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_408
timestamp 1679581782
transform 1 0 39744 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_415
timestamp 1679581782
transform 1 0 40416 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_422
timestamp 1679581782
transform 1 0 41088 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_429
timestamp 1679581782
transform 1 0 41760 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_436
timestamp 1679581782
transform 1 0 42432 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_443
timestamp 1679581782
transform 1 0 43104 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_450
timestamp 1679581782
transform 1 0 43776 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_457
timestamp 1679581782
transform 1 0 44448 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_464
timestamp 1679581782
transform 1 0 45120 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_471
timestamp 1679581782
transform 1 0 45792 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_478
timestamp 1679581782
transform 1 0 46464 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_485
timestamp 1679581782
transform 1 0 47136 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_492
timestamp 1679581782
transform 1 0 47808 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_499
timestamp 1679581782
transform 1 0 48480 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_506
timestamp 1679581782
transform 1 0 49152 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_513
timestamp 1679581782
transform 1 0 49824 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_520
timestamp 1679581782
transform 1 0 50496 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_527
timestamp 1679581782
transform 1 0 51168 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_534
timestamp 1679581782
transform 1 0 51840 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_541
timestamp 1679581782
transform 1 0 52512 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_548
timestamp 1679581782
transform 1 0 53184 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_555
timestamp 1679581782
transform 1 0 53856 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_562
timestamp 1679581782
transform 1 0 54528 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_569
timestamp 1679581782
transform 1 0 55200 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_576
timestamp 1679581782
transform 1 0 55872 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_583
timestamp 1679581782
transform 1 0 56544 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_590
timestamp 1679581782
transform 1 0 57216 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_597
timestamp 1679581782
transform 1 0 57888 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_604
timestamp 1679581782
transform 1 0 58560 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_611
timestamp 1679581782
transform 1 0 59232 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_618
timestamp 1679581782
transform 1 0 59904 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_625
timestamp 1679581782
transform 1 0 60576 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_632
timestamp 1679581782
transform 1 0 61248 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_639
timestamp 1679581782
transform 1 0 61920 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_646
timestamp 1679581782
transform 1 0 62592 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_653
timestamp 1679581782
transform 1 0 63264 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_660
timestamp 1679581782
transform 1 0 63936 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_667
timestamp 1679581782
transform 1 0 64608 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_674
timestamp 1679581782
transform 1 0 65280 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_681
timestamp 1679581782
transform 1 0 65952 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_688
timestamp 1679581782
transform 1 0 66624 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_695
timestamp 1679581782
transform 1 0 67296 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_702
timestamp 1679581782
transform 1 0 67968 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_709
timestamp 1679581782
transform 1 0 68640 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_716
timestamp 1679581782
transform 1 0 69312 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_723
timestamp 1679581782
transform 1 0 69984 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_730
timestamp 1679581782
transform 1 0 70656 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_737
timestamp 1679581782
transform 1 0 71328 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_744
timestamp 1679581782
transform 1 0 72000 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_751
timestamp 1679581782
transform 1 0 72672 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_758
timestamp 1679581782
transform 1 0 73344 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_765
timestamp 1679581782
transform 1 0 74016 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_772
timestamp 1679581782
transform 1 0 74688 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_779
timestamp 1679581782
transform 1 0 75360 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_786
timestamp 1679581782
transform 1 0 76032 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_793
timestamp 1679581782
transform 1 0 76704 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_800
timestamp 1679581782
transform 1 0 77376 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_807
timestamp 1679581782
transform 1 0 78048 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_814
timestamp 1679581782
transform 1 0 78720 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_821
timestamp 1679581782
transform 1 0 79392 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_828
timestamp 1679581782
transform 1 0 80064 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_835
timestamp 1679581782
transform 1 0 80736 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_842
timestamp 1679581782
transform 1 0 81408 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_849
timestamp 1679581782
transform 1 0 82080 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_856
timestamp 1679581782
transform 1 0 82752 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_863
timestamp 1679581782
transform 1 0 83424 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_870
timestamp 1679581782
transform 1 0 84096 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_877
timestamp 1679581782
transform 1 0 84768 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_884
timestamp 1679581782
transform 1 0 85440 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_891
timestamp 1679581782
transform 1 0 86112 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_898
timestamp 1679581782
transform 1 0 86784 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_905
timestamp 1679581782
transform 1 0 87456 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_912
timestamp 1679581782
transform 1 0 88128 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_35_919
timestamp 1679577901
transform 1 0 88800 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_35_923
timestamp 1677580104
transform 1 0 89184 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_36_4
timestamp 1679581782
transform 1 0 960 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_11
timestamp 1679581782
transform 1 0 1632 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_18
timestamp 1679581782
transform 1 0 2304 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_25
timestamp 1679581782
transform 1 0 2976 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_32
timestamp 1679581782
transform 1 0 3648 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_39
timestamp 1679581782
transform 1 0 4320 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_46
timestamp 1679581782
transform 1 0 4992 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_53
timestamp 1679581782
transform 1 0 5664 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_60
timestamp 1679581782
transform 1 0 6336 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_67
timestamp 1679581782
transform 1 0 7008 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_74
timestamp 1679581782
transform 1 0 7680 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_81
timestamp 1679581782
transform 1 0 8352 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_88
timestamp 1679581782
transform 1 0 9024 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_95
timestamp 1679581782
transform 1 0 9696 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_102
timestamp 1679581782
transform 1 0 10368 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_109
timestamp 1679581782
transform 1 0 11040 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_116
timestamp 1679581782
transform 1 0 11712 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_123
timestamp 1679581782
transform 1 0 12384 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_130
timestamp 1679581782
transform 1 0 13056 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_137
timestamp 1679581782
transform 1 0 13728 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_144
timestamp 1679581782
transform 1 0 14400 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_151
timestamp 1679581782
transform 1 0 15072 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_158
timestamp 1679581782
transform 1 0 15744 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_165
timestamp 1679581782
transform 1 0 16416 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_172
timestamp 1679581782
transform 1 0 17088 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_179
timestamp 1679581782
transform 1 0 17760 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_186
timestamp 1679581782
transform 1 0 18432 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_193
timestamp 1679581782
transform 1 0 19104 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_200
timestamp 1679581782
transform 1 0 19776 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_207
timestamp 1679581782
transform 1 0 20448 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_214
timestamp 1679581782
transform 1 0 21120 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_221
timestamp 1679581782
transform 1 0 21792 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_228
timestamp 1679581782
transform 1 0 22464 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_235
timestamp 1679581782
transform 1 0 23136 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_242
timestamp 1679581782
transform 1 0 23808 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_249
timestamp 1679581782
transform 1 0 24480 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_256
timestamp 1679581782
transform 1 0 25152 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_263
timestamp 1679581782
transform 1 0 25824 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_270
timestamp 1679581782
transform 1 0 26496 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_277
timestamp 1679581782
transform 1 0 27168 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_284
timestamp 1679581782
transform 1 0 27840 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_291
timestamp 1679581782
transform 1 0 28512 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_298
timestamp 1679581782
transform 1 0 29184 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_305
timestamp 1679581782
transform 1 0 29856 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_312
timestamp 1679581782
transform 1 0 30528 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_319
timestamp 1679581782
transform 1 0 31200 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_326
timestamp 1679581782
transform 1 0 31872 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_333
timestamp 1679581782
transform 1 0 32544 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_340
timestamp 1679581782
transform 1 0 33216 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_347
timestamp 1679581782
transform 1 0 33888 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_354
timestamp 1679581782
transform 1 0 34560 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_361
timestamp 1679581782
transform 1 0 35232 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_368
timestamp 1679581782
transform 1 0 35904 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_375
timestamp 1679581782
transform 1 0 36576 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_382
timestamp 1679581782
transform 1 0 37248 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_389
timestamp 1679581782
transform 1 0 37920 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_396
timestamp 1679581782
transform 1 0 38592 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_403
timestamp 1679581782
transform 1 0 39264 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_410
timestamp 1679581782
transform 1 0 39936 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_417
timestamp 1679581782
transform 1 0 40608 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_424
timestamp 1679581782
transform 1 0 41280 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_431
timestamp 1679581782
transform 1 0 41952 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_438
timestamp 1679581782
transform 1 0 42624 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_445
timestamp 1679581782
transform 1 0 43296 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_452
timestamp 1679581782
transform 1 0 43968 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_459
timestamp 1679581782
transform 1 0 44640 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_466
timestamp 1679581782
transform 1 0 45312 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_473
timestamp 1679581782
transform 1 0 45984 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_480
timestamp 1679581782
transform 1 0 46656 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_487
timestamp 1679581782
transform 1 0 47328 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_494
timestamp 1679581782
transform 1 0 48000 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_501
timestamp 1679581782
transform 1 0 48672 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_508
timestamp 1679581782
transform 1 0 49344 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_515
timestamp 1679581782
transform 1 0 50016 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_522
timestamp 1679581782
transform 1 0 50688 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_529
timestamp 1679581782
transform 1 0 51360 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_536
timestamp 1679581782
transform 1 0 52032 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_543
timestamp 1679581782
transform 1 0 52704 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_550
timestamp 1679581782
transform 1 0 53376 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_557
timestamp 1679581782
transform 1 0 54048 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_564
timestamp 1679581782
transform 1 0 54720 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_571
timestamp 1679581782
transform 1 0 55392 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_578
timestamp 1679581782
transform 1 0 56064 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_585
timestamp 1679581782
transform 1 0 56736 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_592
timestamp 1679581782
transform 1 0 57408 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_599
timestamp 1679581782
transform 1 0 58080 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_606
timestamp 1679581782
transform 1 0 58752 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_613
timestamp 1679581782
transform 1 0 59424 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_620
timestamp 1679581782
transform 1 0 60096 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_627
timestamp 1679581782
transform 1 0 60768 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_634
timestamp 1679581782
transform 1 0 61440 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_641
timestamp 1679581782
transform 1 0 62112 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_648
timestamp 1679581782
transform 1 0 62784 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_655
timestamp 1679581782
transform 1 0 63456 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_662
timestamp 1679581782
transform 1 0 64128 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_669
timestamp 1679581782
transform 1 0 64800 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_676
timestamp 1679581782
transform 1 0 65472 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_683
timestamp 1679581782
transform 1 0 66144 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_690
timestamp 1679581782
transform 1 0 66816 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_697
timestamp 1679581782
transform 1 0 67488 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_704
timestamp 1679581782
transform 1 0 68160 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_711
timestamp 1679581782
transform 1 0 68832 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_718
timestamp 1679581782
transform 1 0 69504 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_725
timestamp 1679581782
transform 1 0 70176 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_732
timestamp 1679581782
transform 1 0 70848 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_739
timestamp 1679581782
transform 1 0 71520 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_746
timestamp 1679581782
transform 1 0 72192 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_753
timestamp 1679581782
transform 1 0 72864 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_760
timestamp 1679581782
transform 1 0 73536 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_767
timestamp 1679581782
transform 1 0 74208 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_774
timestamp 1679581782
transform 1 0 74880 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_781
timestamp 1679581782
transform 1 0 75552 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_788
timestamp 1679581782
transform 1 0 76224 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_795
timestamp 1679581782
transform 1 0 76896 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_802
timestamp 1679581782
transform 1 0 77568 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_809
timestamp 1679581782
transform 1 0 78240 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_816
timestamp 1679581782
transform 1 0 78912 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_823
timestamp 1679581782
transform 1 0 79584 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_830
timestamp 1679581782
transform 1 0 80256 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_837
timestamp 1679581782
transform 1 0 80928 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_844
timestamp 1679581782
transform 1 0 81600 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_851
timestamp 1679581782
transform 1 0 82272 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_858
timestamp 1679581782
transform 1 0 82944 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_865
timestamp 1679581782
transform 1 0 83616 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_872
timestamp 1679581782
transform 1 0 84288 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_879
timestamp 1679581782
transform 1 0 84960 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_886
timestamp 1679581782
transform 1 0 85632 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_893
timestamp 1679581782
transform 1 0 86304 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_900
timestamp 1679581782
transform 1 0 86976 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_907
timestamp 1679581782
transform 1 0 87648 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_914
timestamp 1679581782
transform 1 0 88320 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_921
timestamp 1679577901
transform 1 0 88992 0 1 27972
box -48 -56 432 834
use sg13g2_decap_8  FILLER_37_0
timestamp 1679581782
transform 1 0 576 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_7
timestamp 1679581782
transform 1 0 1248 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_14
timestamp 1679581782
transform 1 0 1920 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_21
timestamp 1679581782
transform 1 0 2592 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_28
timestamp 1679581782
transform 1 0 3264 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_35
timestamp 1679581782
transform 1 0 3936 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_42
timestamp 1679581782
transform 1 0 4608 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_49
timestamp 1679581782
transform 1 0 5280 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_56
timestamp 1679581782
transform 1 0 5952 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_63
timestamp 1679581782
transform 1 0 6624 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_70
timestamp 1679581782
transform 1 0 7296 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_77
timestamp 1679581782
transform 1 0 7968 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_84
timestamp 1679581782
transform 1 0 8640 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_91
timestamp 1679581782
transform 1 0 9312 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_98
timestamp 1679581782
transform 1 0 9984 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_105
timestamp 1679581782
transform 1 0 10656 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_112
timestamp 1679581782
transform 1 0 11328 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_119
timestamp 1679581782
transform 1 0 12000 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_126
timestamp 1679581782
transform 1 0 12672 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_133
timestamp 1679581782
transform 1 0 13344 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_140
timestamp 1679581782
transform 1 0 14016 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_147
timestamp 1679581782
transform 1 0 14688 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_154
timestamp 1679581782
transform 1 0 15360 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_161
timestamp 1679581782
transform 1 0 16032 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_168
timestamp 1679581782
transform 1 0 16704 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_175
timestamp 1679581782
transform 1 0 17376 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_182
timestamp 1679581782
transform 1 0 18048 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_189
timestamp 1679581782
transform 1 0 18720 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_196
timestamp 1679581782
transform 1 0 19392 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_203
timestamp 1679581782
transform 1 0 20064 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_210
timestamp 1679581782
transform 1 0 20736 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_217
timestamp 1679581782
transform 1 0 21408 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_224
timestamp 1679581782
transform 1 0 22080 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_231
timestamp 1679581782
transform 1 0 22752 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_238
timestamp 1679581782
transform 1 0 23424 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_245
timestamp 1679581782
transform 1 0 24096 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_252
timestamp 1679581782
transform 1 0 24768 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_259
timestamp 1679581782
transform 1 0 25440 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_266
timestamp 1679581782
transform 1 0 26112 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_273
timestamp 1679581782
transform 1 0 26784 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_280
timestamp 1679581782
transform 1 0 27456 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_287
timestamp 1679581782
transform 1 0 28128 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_294
timestamp 1679581782
transform 1 0 28800 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_301
timestamp 1679581782
transform 1 0 29472 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_308
timestamp 1679581782
transform 1 0 30144 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_315
timestamp 1679581782
transform 1 0 30816 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_322
timestamp 1679581782
transform 1 0 31488 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_329
timestamp 1679581782
transform 1 0 32160 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_336
timestamp 1679581782
transform 1 0 32832 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_343
timestamp 1679581782
transform 1 0 33504 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_350
timestamp 1679581782
transform 1 0 34176 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_357
timestamp 1679581782
transform 1 0 34848 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_364
timestamp 1679581782
transform 1 0 35520 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_371
timestamp 1679581782
transform 1 0 36192 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_378
timestamp 1679581782
transform 1 0 36864 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_385
timestamp 1679581782
transform 1 0 37536 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_392
timestamp 1679581782
transform 1 0 38208 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_399
timestamp 1679581782
transform 1 0 38880 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_406
timestamp 1679581782
transform 1 0 39552 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_413
timestamp 1679581782
transform 1 0 40224 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_420
timestamp 1679581782
transform 1 0 40896 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_427
timestamp 1679581782
transform 1 0 41568 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_434
timestamp 1679581782
transform 1 0 42240 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_441
timestamp 1679581782
transform 1 0 42912 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_448
timestamp 1679581782
transform 1 0 43584 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_455
timestamp 1679581782
transform 1 0 44256 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_462
timestamp 1679581782
transform 1 0 44928 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_469
timestamp 1679581782
transform 1 0 45600 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_476
timestamp 1679581782
transform 1 0 46272 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_483
timestamp 1679581782
transform 1 0 46944 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_490
timestamp 1679581782
transform 1 0 47616 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_497
timestamp 1679581782
transform 1 0 48288 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_504
timestamp 1679581782
transform 1 0 48960 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_511
timestamp 1679581782
transform 1 0 49632 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_518
timestamp 1679581782
transform 1 0 50304 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_525
timestamp 1679581782
transform 1 0 50976 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_532
timestamp 1679581782
transform 1 0 51648 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_539
timestamp 1679581782
transform 1 0 52320 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_546
timestamp 1679581782
transform 1 0 52992 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_553
timestamp 1679581782
transform 1 0 53664 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_560
timestamp 1679581782
transform 1 0 54336 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_567
timestamp 1679581782
transform 1 0 55008 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_574
timestamp 1679581782
transform 1 0 55680 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_581
timestamp 1679581782
transform 1 0 56352 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_588
timestamp 1679581782
transform 1 0 57024 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_595
timestamp 1679581782
transform 1 0 57696 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_602
timestamp 1679581782
transform 1 0 58368 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_609
timestamp 1679581782
transform 1 0 59040 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_616
timestamp 1679581782
transform 1 0 59712 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_623
timestamp 1679581782
transform 1 0 60384 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_630
timestamp 1679581782
transform 1 0 61056 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_637
timestamp 1679581782
transform 1 0 61728 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_644
timestamp 1679581782
transform 1 0 62400 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_651
timestamp 1679581782
transform 1 0 63072 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_658
timestamp 1679581782
transform 1 0 63744 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_665
timestamp 1679581782
transform 1 0 64416 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_672
timestamp 1679581782
transform 1 0 65088 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_679
timestamp 1679581782
transform 1 0 65760 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_686
timestamp 1679581782
transform 1 0 66432 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_693
timestamp 1679581782
transform 1 0 67104 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_700
timestamp 1679581782
transform 1 0 67776 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_707
timestamp 1679581782
transform 1 0 68448 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_714
timestamp 1679581782
transform 1 0 69120 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_721
timestamp 1679581782
transform 1 0 69792 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_728
timestamp 1679581782
transform 1 0 70464 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_735
timestamp 1679581782
transform 1 0 71136 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_742
timestamp 1679581782
transform 1 0 71808 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_749
timestamp 1679581782
transform 1 0 72480 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_756
timestamp 1679581782
transform 1 0 73152 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_763
timestamp 1679581782
transform 1 0 73824 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_770
timestamp 1679581782
transform 1 0 74496 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_777
timestamp 1679581782
transform 1 0 75168 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_784
timestamp 1679581782
transform 1 0 75840 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_791
timestamp 1679581782
transform 1 0 76512 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_798
timestamp 1679581782
transform 1 0 77184 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_805
timestamp 1679581782
transform 1 0 77856 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_812
timestamp 1679581782
transform 1 0 78528 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_819
timestamp 1679581782
transform 1 0 79200 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_826
timestamp 1679581782
transform 1 0 79872 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_833
timestamp 1679581782
transform 1 0 80544 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_840
timestamp 1679581782
transform 1 0 81216 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_847
timestamp 1679581782
transform 1 0 81888 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_854
timestamp 1679581782
transform 1 0 82560 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_861
timestamp 1679581782
transform 1 0 83232 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_868
timestamp 1679581782
transform 1 0 83904 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_875
timestamp 1679581782
transform 1 0 84576 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_882
timestamp 1679581782
transform 1 0 85248 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_889
timestamp 1679581782
transform 1 0 85920 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_896
timestamp 1679581782
transform 1 0 86592 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_903
timestamp 1679581782
transform 1 0 87264 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_910
timestamp 1679581782
transform 1 0 87936 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_917
timestamp 1679581782
transform 1 0 88608 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_1  FILLER_37_924
timestamp 1677579658
transform 1 0 89280 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_4
timestamp 1679581782
transform 1 0 960 0 1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_38_11
timestamp 1679577901
transform 1 0 1632 0 1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_38_15
timestamp 1677580104
transform 1 0 2016 0 1 29484
box -48 -56 240 834
use sg13g2_decap_8  FILLER_38_33
timestamp 1679581782
transform 1 0 3744 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_40
timestamp 1679581782
transform 1 0 4416 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_47
timestamp 1679581782
transform 1 0 5088 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_54
timestamp 1679581782
transform 1 0 5760 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_61
timestamp 1679581782
transform 1 0 6432 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_68
timestamp 1679581782
transform 1 0 7104 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_75
timestamp 1679581782
transform 1 0 7776 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_82
timestamp 1679581782
transform 1 0 8448 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_89
timestamp 1679581782
transform 1 0 9120 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_96
timestamp 1679581782
transform 1 0 9792 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_103
timestamp 1679581782
transform 1 0 10464 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_110
timestamp 1679581782
transform 1 0 11136 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_117
timestamp 1679581782
transform 1 0 11808 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_124
timestamp 1679581782
transform 1 0 12480 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_131
timestamp 1679581782
transform 1 0 13152 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_138
timestamp 1679581782
transform 1 0 13824 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_145
timestamp 1679581782
transform 1 0 14496 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_152
timestamp 1679581782
transform 1 0 15168 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_159
timestamp 1679581782
transform 1 0 15840 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_166
timestamp 1679581782
transform 1 0 16512 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_173
timestamp 1679581782
transform 1 0 17184 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_180
timestamp 1679581782
transform 1 0 17856 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_187
timestamp 1679581782
transform 1 0 18528 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_194
timestamp 1679581782
transform 1 0 19200 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_201
timestamp 1679581782
transform 1 0 19872 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_208
timestamp 1679581782
transform 1 0 20544 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_215
timestamp 1679581782
transform 1 0 21216 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_222
timestamp 1679581782
transform 1 0 21888 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_229
timestamp 1679581782
transform 1 0 22560 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_236
timestamp 1679581782
transform 1 0 23232 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_243
timestamp 1679581782
transform 1 0 23904 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_250
timestamp 1679581782
transform 1 0 24576 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_257
timestamp 1679581782
transform 1 0 25248 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_264
timestamp 1679581782
transform 1 0 25920 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_271
timestamp 1679581782
transform 1 0 26592 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_278
timestamp 1679581782
transform 1 0 27264 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_285
timestamp 1679581782
transform 1 0 27936 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_292
timestamp 1679581782
transform 1 0 28608 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_299
timestamp 1679581782
transform 1 0 29280 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_306
timestamp 1679581782
transform 1 0 29952 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_313
timestamp 1679581782
transform 1 0 30624 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_320
timestamp 1679581782
transform 1 0 31296 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_327
timestamp 1679581782
transform 1 0 31968 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_334
timestamp 1679581782
transform 1 0 32640 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_341
timestamp 1679581782
transform 1 0 33312 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_348
timestamp 1679581782
transform 1 0 33984 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_355
timestamp 1679581782
transform 1 0 34656 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_362
timestamp 1679581782
transform 1 0 35328 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_369
timestamp 1679581782
transform 1 0 36000 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_376
timestamp 1679581782
transform 1 0 36672 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_383
timestamp 1679581782
transform 1 0 37344 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_390
timestamp 1679581782
transform 1 0 38016 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_397
timestamp 1679581782
transform 1 0 38688 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_404
timestamp 1679581782
transform 1 0 39360 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_411
timestamp 1679581782
transform 1 0 40032 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_418
timestamp 1679581782
transform 1 0 40704 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_425
timestamp 1679581782
transform 1 0 41376 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_432
timestamp 1679581782
transform 1 0 42048 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_439
timestamp 1679581782
transform 1 0 42720 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_446
timestamp 1679581782
transform 1 0 43392 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_453
timestamp 1679581782
transform 1 0 44064 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_460
timestamp 1679581782
transform 1 0 44736 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_467
timestamp 1679581782
transform 1 0 45408 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_474
timestamp 1679581782
transform 1 0 46080 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_481
timestamp 1679581782
transform 1 0 46752 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_488
timestamp 1679581782
transform 1 0 47424 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_495
timestamp 1679581782
transform 1 0 48096 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_502
timestamp 1679581782
transform 1 0 48768 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_509
timestamp 1679581782
transform 1 0 49440 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_516
timestamp 1679581782
transform 1 0 50112 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_523
timestamp 1679581782
transform 1 0 50784 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_530
timestamp 1679581782
transform 1 0 51456 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_537
timestamp 1679581782
transform 1 0 52128 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_544
timestamp 1679581782
transform 1 0 52800 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_551
timestamp 1679581782
transform 1 0 53472 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_558
timestamp 1679581782
transform 1 0 54144 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_565
timestamp 1679581782
transform 1 0 54816 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_572
timestamp 1679581782
transform 1 0 55488 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_579
timestamp 1679581782
transform 1 0 56160 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_586
timestamp 1679581782
transform 1 0 56832 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_593
timestamp 1679581782
transform 1 0 57504 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_600
timestamp 1679581782
transform 1 0 58176 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_607
timestamp 1679581782
transform 1 0 58848 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_614
timestamp 1679581782
transform 1 0 59520 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_621
timestamp 1679581782
transform 1 0 60192 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_628
timestamp 1679581782
transform 1 0 60864 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_635
timestamp 1679581782
transform 1 0 61536 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_642
timestamp 1679581782
transform 1 0 62208 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_649
timestamp 1679581782
transform 1 0 62880 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_656
timestamp 1679581782
transform 1 0 63552 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_663
timestamp 1679581782
transform 1 0 64224 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_670
timestamp 1679581782
transform 1 0 64896 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_677
timestamp 1679581782
transform 1 0 65568 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_684
timestamp 1679581782
transform 1 0 66240 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_691
timestamp 1679581782
transform 1 0 66912 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_698
timestamp 1679581782
transform 1 0 67584 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_705
timestamp 1679581782
transform 1 0 68256 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_712
timestamp 1679581782
transform 1 0 68928 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_719
timestamp 1679581782
transform 1 0 69600 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_726
timestamp 1679581782
transform 1 0 70272 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_733
timestamp 1679581782
transform 1 0 70944 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_740
timestamp 1679581782
transform 1 0 71616 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_747
timestamp 1679581782
transform 1 0 72288 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_754
timestamp 1679581782
transform 1 0 72960 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_761
timestamp 1679581782
transform 1 0 73632 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_768
timestamp 1679581782
transform 1 0 74304 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_775
timestamp 1679581782
transform 1 0 74976 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_782
timestamp 1679581782
transform 1 0 75648 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_789
timestamp 1679581782
transform 1 0 76320 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_796
timestamp 1679581782
transform 1 0 76992 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_803
timestamp 1679581782
transform 1 0 77664 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_810
timestamp 1679581782
transform 1 0 78336 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_817
timestamp 1679581782
transform 1 0 79008 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_824
timestamp 1679581782
transform 1 0 79680 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_831
timestamp 1679581782
transform 1 0 80352 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_838
timestamp 1679581782
transform 1 0 81024 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_845
timestamp 1679581782
transform 1 0 81696 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_852
timestamp 1679581782
transform 1 0 82368 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_859
timestamp 1679581782
transform 1 0 83040 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_866
timestamp 1679581782
transform 1 0 83712 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_873
timestamp 1679581782
transform 1 0 84384 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_880
timestamp 1679581782
transform 1 0 85056 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_887
timestamp 1679581782
transform 1 0 85728 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_894
timestamp 1679581782
transform 1 0 86400 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_901
timestamp 1679581782
transform 1 0 87072 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_908
timestamp 1679581782
transform 1 0 87744 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_915
timestamp 1679581782
transform 1 0 88416 0 1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_38_922
timestamp 1677580104
transform 1 0 89088 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_924
timestamp 1677579658
transform 1 0 89280 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_4
timestamp 1679581782
transform 1 0 960 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_11
timestamp 1679581782
transform 1 0 1632 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_39_18
timestamp 1677580104
transform 1 0 2304 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_20
timestamp 1677579658
transform 1 0 2496 0 -1 30996
box -48 -56 144 834
use sg13g2_fill_1  FILLER_39_29
timestamp 1677579658
transform 1 0 3360 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_35
timestamp 1679581782
transform 1 0 3936 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_42
timestamp 1679581782
transform 1 0 4608 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_49
timestamp 1679581782
transform 1 0 5280 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_56
timestamp 1679581782
transform 1 0 5952 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_63
timestamp 1679581782
transform 1 0 6624 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_70
timestamp 1679581782
transform 1 0 7296 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_77
timestamp 1679581782
transform 1 0 7968 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_84
timestamp 1679581782
transform 1 0 8640 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_91
timestamp 1679581782
transform 1 0 9312 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_98
timestamp 1679581782
transform 1 0 9984 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_105
timestamp 1679581782
transform 1 0 10656 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_112
timestamp 1679581782
transform 1 0 11328 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_119
timestamp 1679581782
transform 1 0 12000 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_126
timestamp 1679581782
transform 1 0 12672 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_133
timestamp 1679581782
transform 1 0 13344 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_140
timestamp 1679581782
transform 1 0 14016 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_147
timestamp 1679581782
transform 1 0 14688 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_154
timestamp 1679581782
transform 1 0 15360 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_161
timestamp 1679581782
transform 1 0 16032 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_168
timestamp 1679581782
transform 1 0 16704 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_175
timestamp 1679581782
transform 1 0 17376 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_182
timestamp 1679581782
transform 1 0 18048 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_189
timestamp 1679581782
transform 1 0 18720 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_196
timestamp 1679581782
transform 1 0 19392 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_203
timestamp 1679581782
transform 1 0 20064 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_210
timestamp 1679581782
transform 1 0 20736 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_217
timestamp 1679581782
transform 1 0 21408 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_224
timestamp 1679581782
transform 1 0 22080 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_231
timestamp 1679581782
transform 1 0 22752 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_238
timestamp 1679581782
transform 1 0 23424 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_245
timestamp 1679581782
transform 1 0 24096 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_252
timestamp 1679581782
transform 1 0 24768 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_259
timestamp 1679581782
transform 1 0 25440 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_266
timestamp 1679581782
transform 1 0 26112 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_273
timestamp 1679581782
transform 1 0 26784 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_280
timestamp 1679581782
transform 1 0 27456 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_287
timestamp 1679581782
transform 1 0 28128 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_294
timestamp 1679581782
transform 1 0 28800 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_301
timestamp 1679581782
transform 1 0 29472 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_308
timestamp 1679581782
transform 1 0 30144 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_315
timestamp 1679581782
transform 1 0 30816 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_322
timestamp 1679581782
transform 1 0 31488 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_329
timestamp 1679581782
transform 1 0 32160 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_336
timestamp 1679581782
transform 1 0 32832 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_343
timestamp 1679581782
transform 1 0 33504 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_350
timestamp 1679581782
transform 1 0 34176 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_357
timestamp 1679581782
transform 1 0 34848 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_364
timestamp 1679581782
transform 1 0 35520 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_371
timestamp 1679581782
transform 1 0 36192 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_378
timestamp 1679581782
transform 1 0 36864 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_385
timestamp 1679581782
transform 1 0 37536 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_392
timestamp 1679581782
transform 1 0 38208 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_399
timestamp 1679581782
transform 1 0 38880 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_406
timestamp 1679581782
transform 1 0 39552 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_413
timestamp 1679581782
transform 1 0 40224 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_420
timestamp 1679581782
transform 1 0 40896 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_427
timestamp 1679581782
transform 1 0 41568 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_434
timestamp 1679581782
transform 1 0 42240 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_441
timestamp 1679581782
transform 1 0 42912 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_448
timestamp 1679581782
transform 1 0 43584 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_455
timestamp 1679581782
transform 1 0 44256 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_462
timestamp 1679581782
transform 1 0 44928 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_469
timestamp 1679581782
transform 1 0 45600 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_476
timestamp 1679581782
transform 1 0 46272 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_483
timestamp 1679581782
transform 1 0 46944 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_490
timestamp 1679581782
transform 1 0 47616 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_497
timestamp 1679581782
transform 1 0 48288 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_504
timestamp 1679581782
transform 1 0 48960 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_511
timestamp 1679581782
transform 1 0 49632 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_518
timestamp 1679581782
transform 1 0 50304 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_525
timestamp 1679581782
transform 1 0 50976 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_532
timestamp 1679581782
transform 1 0 51648 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_539
timestamp 1679581782
transform 1 0 52320 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_546
timestamp 1679581782
transform 1 0 52992 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_553
timestamp 1679581782
transform 1 0 53664 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_560
timestamp 1679581782
transform 1 0 54336 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_567
timestamp 1679581782
transform 1 0 55008 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_574
timestamp 1679581782
transform 1 0 55680 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_581
timestamp 1679581782
transform 1 0 56352 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_588
timestamp 1679581782
transform 1 0 57024 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_595
timestamp 1679581782
transform 1 0 57696 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_602
timestamp 1679581782
transform 1 0 58368 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_609
timestamp 1679581782
transform 1 0 59040 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_616
timestamp 1679581782
transform 1 0 59712 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_623
timestamp 1679581782
transform 1 0 60384 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_630
timestamp 1679581782
transform 1 0 61056 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_637
timestamp 1679581782
transform 1 0 61728 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_644
timestamp 1679581782
transform 1 0 62400 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_651
timestamp 1679581782
transform 1 0 63072 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_658
timestamp 1679581782
transform 1 0 63744 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_665
timestamp 1679581782
transform 1 0 64416 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_672
timestamp 1679581782
transform 1 0 65088 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_679
timestamp 1679581782
transform 1 0 65760 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_686
timestamp 1679581782
transform 1 0 66432 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_693
timestamp 1679581782
transform 1 0 67104 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_700
timestamp 1679581782
transform 1 0 67776 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_707
timestamp 1679581782
transform 1 0 68448 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_714
timestamp 1679581782
transform 1 0 69120 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_721
timestamp 1679581782
transform 1 0 69792 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_728
timestamp 1679581782
transform 1 0 70464 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_735
timestamp 1679581782
transform 1 0 71136 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_742
timestamp 1679581782
transform 1 0 71808 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_749
timestamp 1679581782
transform 1 0 72480 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_756
timestamp 1679581782
transform 1 0 73152 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_763
timestamp 1679581782
transform 1 0 73824 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_770
timestamp 1679581782
transform 1 0 74496 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_777
timestamp 1679581782
transform 1 0 75168 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_784
timestamp 1679581782
transform 1 0 75840 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_791
timestamp 1679581782
transform 1 0 76512 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_798
timestamp 1679581782
transform 1 0 77184 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_805
timestamp 1679581782
transform 1 0 77856 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_812
timestamp 1679581782
transform 1 0 78528 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_819
timestamp 1679581782
transform 1 0 79200 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_826
timestamp 1679581782
transform 1 0 79872 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_833
timestamp 1679581782
transform 1 0 80544 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_840
timestamp 1679581782
transform 1 0 81216 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_847
timestamp 1679581782
transform 1 0 81888 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_854
timestamp 1679581782
transform 1 0 82560 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_861
timestamp 1679581782
transform 1 0 83232 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_868
timestamp 1679581782
transform 1 0 83904 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_875
timestamp 1679581782
transform 1 0 84576 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_882
timestamp 1679581782
transform 1 0 85248 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_889
timestamp 1679581782
transform 1 0 85920 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_896
timestamp 1679581782
transform 1 0 86592 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_903
timestamp 1679581782
transform 1 0 87264 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_910
timestamp 1679581782
transform 1 0 87936 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_917
timestamp 1679581782
transform 1 0 88608 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_1  FILLER_39_924
timestamp 1677579658
transform 1 0 89280 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_4
timestamp 1679581782
transform 1 0 960 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_11
timestamp 1679581782
transform 1 0 1632 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_18
timestamp 1679581782
transform 1 0 2304 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_25
timestamp 1679581782
transform 1 0 2976 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_32
timestamp 1679581782
transform 1 0 3648 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_39
timestamp 1679581782
transform 1 0 4320 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_46
timestamp 1679581782
transform 1 0 4992 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_53
timestamp 1679581782
transform 1 0 5664 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_60
timestamp 1679581782
transform 1 0 6336 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_67
timestamp 1679581782
transform 1 0 7008 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_74
timestamp 1679581782
transform 1 0 7680 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_81
timestamp 1679581782
transform 1 0 8352 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_88
timestamp 1679581782
transform 1 0 9024 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_95
timestamp 1679581782
transform 1 0 9696 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_102
timestamp 1679581782
transform 1 0 10368 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_109
timestamp 1679581782
transform 1 0 11040 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_116
timestamp 1679581782
transform 1 0 11712 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_123
timestamp 1679581782
transform 1 0 12384 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_130
timestamp 1679581782
transform 1 0 13056 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_137
timestamp 1679581782
transform 1 0 13728 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_144
timestamp 1679581782
transform 1 0 14400 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_151
timestamp 1679581782
transform 1 0 15072 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_158
timestamp 1679581782
transform 1 0 15744 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_165
timestamp 1679581782
transform 1 0 16416 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_172
timestamp 1679581782
transform 1 0 17088 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_179
timestamp 1679581782
transform 1 0 17760 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_186
timestamp 1679581782
transform 1 0 18432 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_193
timestamp 1679581782
transform 1 0 19104 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_200
timestamp 1679581782
transform 1 0 19776 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_207
timestamp 1679581782
transform 1 0 20448 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_214
timestamp 1679581782
transform 1 0 21120 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_221
timestamp 1679581782
transform 1 0 21792 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_228
timestamp 1679581782
transform 1 0 22464 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_235
timestamp 1679581782
transform 1 0 23136 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_242
timestamp 1679581782
transform 1 0 23808 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_249
timestamp 1679581782
transform 1 0 24480 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_256
timestamp 1679581782
transform 1 0 25152 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_263
timestamp 1679581782
transform 1 0 25824 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_270
timestamp 1679581782
transform 1 0 26496 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_277
timestamp 1679581782
transform 1 0 27168 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_284
timestamp 1679581782
transform 1 0 27840 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_291
timestamp 1679581782
transform 1 0 28512 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_298
timestamp 1679581782
transform 1 0 29184 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_305
timestamp 1679581782
transform 1 0 29856 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_312
timestamp 1679581782
transform 1 0 30528 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_319
timestamp 1679581782
transform 1 0 31200 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_326
timestamp 1679581782
transform 1 0 31872 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_333
timestamp 1679581782
transform 1 0 32544 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_340
timestamp 1679581782
transform 1 0 33216 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_347
timestamp 1679581782
transform 1 0 33888 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_354
timestamp 1679581782
transform 1 0 34560 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_361
timestamp 1679581782
transform 1 0 35232 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_368
timestamp 1679581782
transform 1 0 35904 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_375
timestamp 1679581782
transform 1 0 36576 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_382
timestamp 1679581782
transform 1 0 37248 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_389
timestamp 1679581782
transform 1 0 37920 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_396
timestamp 1679581782
transform 1 0 38592 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_403
timestamp 1679581782
transform 1 0 39264 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_410
timestamp 1679581782
transform 1 0 39936 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_417
timestamp 1679581782
transform 1 0 40608 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_424
timestamp 1679581782
transform 1 0 41280 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_431
timestamp 1679581782
transform 1 0 41952 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_438
timestamp 1679581782
transform 1 0 42624 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_445
timestamp 1679581782
transform 1 0 43296 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_452
timestamp 1679581782
transform 1 0 43968 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_459
timestamp 1679581782
transform 1 0 44640 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_466
timestamp 1679581782
transform 1 0 45312 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_473
timestamp 1679581782
transform 1 0 45984 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_480
timestamp 1679581782
transform 1 0 46656 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_487
timestamp 1679581782
transform 1 0 47328 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_494
timestamp 1679581782
transform 1 0 48000 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_501
timestamp 1679581782
transform 1 0 48672 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_508
timestamp 1679581782
transform 1 0 49344 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_515
timestamp 1679581782
transform 1 0 50016 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_522
timestamp 1679581782
transform 1 0 50688 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_529
timestamp 1679581782
transform 1 0 51360 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_536
timestamp 1679581782
transform 1 0 52032 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_543
timestamp 1679581782
transform 1 0 52704 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_550
timestamp 1679581782
transform 1 0 53376 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_557
timestamp 1679581782
transform 1 0 54048 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_564
timestamp 1679581782
transform 1 0 54720 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_571
timestamp 1679581782
transform 1 0 55392 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_578
timestamp 1679581782
transform 1 0 56064 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_585
timestamp 1679581782
transform 1 0 56736 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_592
timestamp 1679581782
transform 1 0 57408 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_599
timestamp 1679581782
transform 1 0 58080 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_606
timestamp 1679581782
transform 1 0 58752 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_613
timestamp 1679581782
transform 1 0 59424 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_620
timestamp 1679581782
transform 1 0 60096 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_627
timestamp 1679581782
transform 1 0 60768 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_634
timestamp 1679581782
transform 1 0 61440 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_641
timestamp 1679581782
transform 1 0 62112 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_648
timestamp 1679581782
transform 1 0 62784 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_655
timestamp 1679581782
transform 1 0 63456 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_662
timestamp 1679581782
transform 1 0 64128 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_669
timestamp 1679581782
transform 1 0 64800 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_676
timestamp 1679581782
transform 1 0 65472 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_683
timestamp 1679581782
transform 1 0 66144 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_690
timestamp 1679581782
transform 1 0 66816 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_697
timestamp 1679581782
transform 1 0 67488 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_704
timestamp 1679581782
transform 1 0 68160 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_711
timestamp 1679581782
transform 1 0 68832 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_718
timestamp 1679581782
transform 1 0 69504 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_725
timestamp 1679581782
transform 1 0 70176 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_732
timestamp 1679581782
transform 1 0 70848 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_739
timestamp 1679581782
transform 1 0 71520 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_746
timestamp 1679581782
transform 1 0 72192 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_753
timestamp 1679581782
transform 1 0 72864 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_760
timestamp 1679581782
transform 1 0 73536 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_767
timestamp 1679581782
transform 1 0 74208 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_774
timestamp 1679581782
transform 1 0 74880 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_781
timestamp 1679581782
transform 1 0 75552 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_788
timestamp 1679581782
transform 1 0 76224 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_795
timestamp 1679581782
transform 1 0 76896 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_802
timestamp 1679581782
transform 1 0 77568 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_809
timestamp 1679581782
transform 1 0 78240 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_816
timestamp 1679581782
transform 1 0 78912 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_823
timestamp 1679581782
transform 1 0 79584 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_830
timestamp 1679581782
transform 1 0 80256 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_837
timestamp 1679581782
transform 1 0 80928 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_844
timestamp 1679581782
transform 1 0 81600 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_851
timestamp 1679581782
transform 1 0 82272 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_858
timestamp 1679581782
transform 1 0 82944 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_865
timestamp 1679581782
transform 1 0 83616 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_872
timestamp 1679581782
transform 1 0 84288 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_879
timestamp 1679581782
transform 1 0 84960 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_886
timestamp 1679581782
transform 1 0 85632 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_893
timestamp 1679581782
transform 1 0 86304 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_900
timestamp 1679581782
transform 1 0 86976 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_907
timestamp 1679581782
transform 1 0 87648 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_914
timestamp 1679581782
transform 1 0 88320 0 1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_921
timestamp 1679577901
transform 1 0 88992 0 1 30996
box -48 -56 432 834
use sg13g2_decap_8  FILLER_41_4
timestamp 1679581782
transform 1 0 960 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_11
timestamp 1679581782
transform 1 0 1632 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_18
timestamp 1679581782
transform 1 0 2304 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_25
timestamp 1679581782
transform 1 0 2976 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_41_32
timestamp 1679577901
transform 1 0 3648 0 -1 32508
box -48 -56 432 834
use sg13g2_decap_8  FILLER_41_44
timestamp 1679581782
transform 1 0 4800 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_51
timestamp 1679581782
transform 1 0 5472 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_58
timestamp 1679581782
transform 1 0 6144 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_65
timestamp 1679581782
transform 1 0 6816 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_72
timestamp 1679581782
transform 1 0 7488 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_79
timestamp 1679581782
transform 1 0 8160 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_86
timestamp 1679581782
transform 1 0 8832 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_93
timestamp 1679581782
transform 1 0 9504 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_100
timestamp 1679581782
transform 1 0 10176 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_107
timestamp 1679581782
transform 1 0 10848 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_114
timestamp 1679581782
transform 1 0 11520 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_121
timestamp 1679581782
transform 1 0 12192 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_128
timestamp 1679581782
transform 1 0 12864 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_135
timestamp 1679581782
transform 1 0 13536 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_142
timestamp 1679581782
transform 1 0 14208 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_149
timestamp 1679581782
transform 1 0 14880 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_156
timestamp 1679581782
transform 1 0 15552 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_163
timestamp 1679581782
transform 1 0 16224 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_170
timestamp 1679581782
transform 1 0 16896 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_177
timestamp 1679581782
transform 1 0 17568 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_184
timestamp 1679581782
transform 1 0 18240 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_191
timestamp 1679581782
transform 1 0 18912 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_198
timestamp 1679581782
transform 1 0 19584 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_205
timestamp 1679581782
transform 1 0 20256 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_212
timestamp 1679581782
transform 1 0 20928 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_219
timestamp 1679581782
transform 1 0 21600 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_226
timestamp 1679581782
transform 1 0 22272 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_233
timestamp 1679581782
transform 1 0 22944 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_240
timestamp 1679581782
transform 1 0 23616 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_247
timestamp 1679581782
transform 1 0 24288 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_254
timestamp 1679581782
transform 1 0 24960 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_261
timestamp 1679581782
transform 1 0 25632 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_268
timestamp 1679581782
transform 1 0 26304 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_275
timestamp 1679581782
transform 1 0 26976 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_282
timestamp 1679581782
transform 1 0 27648 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_289
timestamp 1679581782
transform 1 0 28320 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_296
timestamp 1679581782
transform 1 0 28992 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_303
timestamp 1679581782
transform 1 0 29664 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_310
timestamp 1679581782
transform 1 0 30336 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_317
timestamp 1679581782
transform 1 0 31008 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_324
timestamp 1679581782
transform 1 0 31680 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_331
timestamp 1679581782
transform 1 0 32352 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_338
timestamp 1679581782
transform 1 0 33024 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_345
timestamp 1679581782
transform 1 0 33696 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_352
timestamp 1679581782
transform 1 0 34368 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_359
timestamp 1679581782
transform 1 0 35040 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_366
timestamp 1679581782
transform 1 0 35712 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_373
timestamp 1679581782
transform 1 0 36384 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_380
timestamp 1679581782
transform 1 0 37056 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_387
timestamp 1679581782
transform 1 0 37728 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_394
timestamp 1679581782
transform 1 0 38400 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_401
timestamp 1679581782
transform 1 0 39072 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_408
timestamp 1679581782
transform 1 0 39744 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_415
timestamp 1679581782
transform 1 0 40416 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_422
timestamp 1679581782
transform 1 0 41088 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_429
timestamp 1679581782
transform 1 0 41760 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_436
timestamp 1679581782
transform 1 0 42432 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_443
timestamp 1679581782
transform 1 0 43104 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_450
timestamp 1679581782
transform 1 0 43776 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_457
timestamp 1679581782
transform 1 0 44448 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_464
timestamp 1679581782
transform 1 0 45120 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_471
timestamp 1679581782
transform 1 0 45792 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_478
timestamp 1679581782
transform 1 0 46464 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_485
timestamp 1679581782
transform 1 0 47136 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_492
timestamp 1679581782
transform 1 0 47808 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_499
timestamp 1679581782
transform 1 0 48480 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_506
timestamp 1679581782
transform 1 0 49152 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_513
timestamp 1679581782
transform 1 0 49824 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_520
timestamp 1679581782
transform 1 0 50496 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_527
timestamp 1679581782
transform 1 0 51168 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_534
timestamp 1679581782
transform 1 0 51840 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_541
timestamp 1679581782
transform 1 0 52512 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_548
timestamp 1679581782
transform 1 0 53184 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_555
timestamp 1679581782
transform 1 0 53856 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_562
timestamp 1679581782
transform 1 0 54528 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_569
timestamp 1679581782
transform 1 0 55200 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_576
timestamp 1679581782
transform 1 0 55872 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_583
timestamp 1679581782
transform 1 0 56544 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_590
timestamp 1679581782
transform 1 0 57216 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_597
timestamp 1679581782
transform 1 0 57888 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_604
timestamp 1679581782
transform 1 0 58560 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_611
timestamp 1679581782
transform 1 0 59232 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_618
timestamp 1679581782
transform 1 0 59904 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_625
timestamp 1679581782
transform 1 0 60576 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_632
timestamp 1679581782
transform 1 0 61248 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_639
timestamp 1679581782
transform 1 0 61920 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_646
timestamp 1679581782
transform 1 0 62592 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_653
timestamp 1679581782
transform 1 0 63264 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_660
timestamp 1679581782
transform 1 0 63936 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_667
timestamp 1679581782
transform 1 0 64608 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_674
timestamp 1679581782
transform 1 0 65280 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_681
timestamp 1679581782
transform 1 0 65952 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_688
timestamp 1679581782
transform 1 0 66624 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_695
timestamp 1679581782
transform 1 0 67296 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_702
timestamp 1679581782
transform 1 0 67968 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_709
timestamp 1679581782
transform 1 0 68640 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_716
timestamp 1679581782
transform 1 0 69312 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_723
timestamp 1679581782
transform 1 0 69984 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_730
timestamp 1679581782
transform 1 0 70656 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_737
timestamp 1679581782
transform 1 0 71328 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_744
timestamp 1679581782
transform 1 0 72000 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_751
timestamp 1679581782
transform 1 0 72672 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_758
timestamp 1679581782
transform 1 0 73344 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_765
timestamp 1679581782
transform 1 0 74016 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_772
timestamp 1679581782
transform 1 0 74688 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_779
timestamp 1679581782
transform 1 0 75360 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_786
timestamp 1679581782
transform 1 0 76032 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_793
timestamp 1679581782
transform 1 0 76704 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_800
timestamp 1679581782
transform 1 0 77376 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_807
timestamp 1679581782
transform 1 0 78048 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_814
timestamp 1679581782
transform 1 0 78720 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_821
timestamp 1679581782
transform 1 0 79392 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_828
timestamp 1679581782
transform 1 0 80064 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_835
timestamp 1679581782
transform 1 0 80736 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_842
timestamp 1679581782
transform 1 0 81408 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_849
timestamp 1679581782
transform 1 0 82080 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_856
timestamp 1679581782
transform 1 0 82752 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_863
timestamp 1679581782
transform 1 0 83424 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_870
timestamp 1679581782
transform 1 0 84096 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_877
timestamp 1679581782
transform 1 0 84768 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_884
timestamp 1679581782
transform 1 0 85440 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_891
timestamp 1679581782
transform 1 0 86112 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_898
timestamp 1679581782
transform 1 0 86784 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_905
timestamp 1679581782
transform 1 0 87456 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_912
timestamp 1679581782
transform 1 0 88128 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_41_919
timestamp 1679577901
transform 1 0 88800 0 -1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_41_923
timestamp 1677580104
transform 1 0 89184 0 -1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_42_4
timestamp 1679581782
transform 1 0 960 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_11
timestamp 1679581782
transform 1 0 1632 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_18
timestamp 1679581782
transform 1 0 2304 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_25
timestamp 1679581782
transform 1 0 2976 0 1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_42_32
timestamp 1677580104
transform 1 0 3648 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_34
timestamp 1677579658
transform 1 0 3840 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_43
timestamp 1679581782
transform 1 0 4704 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_50
timestamp 1679581782
transform 1 0 5376 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_57
timestamp 1679581782
transform 1 0 6048 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_64
timestamp 1679581782
transform 1 0 6720 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_71
timestamp 1679581782
transform 1 0 7392 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_78
timestamp 1679581782
transform 1 0 8064 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_85
timestamp 1679581782
transform 1 0 8736 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_92
timestamp 1679581782
transform 1 0 9408 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_99
timestamp 1679581782
transform 1 0 10080 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_106
timestamp 1679581782
transform 1 0 10752 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_113
timestamp 1679581782
transform 1 0 11424 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_120
timestamp 1679581782
transform 1 0 12096 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_127
timestamp 1679581782
transform 1 0 12768 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_134
timestamp 1679581782
transform 1 0 13440 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_141
timestamp 1679581782
transform 1 0 14112 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_148
timestamp 1679581782
transform 1 0 14784 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_155
timestamp 1679581782
transform 1 0 15456 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_162
timestamp 1679581782
transform 1 0 16128 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_169
timestamp 1679581782
transform 1 0 16800 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_176
timestamp 1679581782
transform 1 0 17472 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_183
timestamp 1679581782
transform 1 0 18144 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_190
timestamp 1679581782
transform 1 0 18816 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_197
timestamp 1679581782
transform 1 0 19488 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_204
timestamp 1679581782
transform 1 0 20160 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_211
timestamp 1679581782
transform 1 0 20832 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_218
timestamp 1679581782
transform 1 0 21504 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_225
timestamp 1679581782
transform 1 0 22176 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_232
timestamp 1679581782
transform 1 0 22848 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_239
timestamp 1679581782
transform 1 0 23520 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_246
timestamp 1679581782
transform 1 0 24192 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_253
timestamp 1679581782
transform 1 0 24864 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_260
timestamp 1679581782
transform 1 0 25536 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_267
timestamp 1679581782
transform 1 0 26208 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_274
timestamp 1679581782
transform 1 0 26880 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_281
timestamp 1679581782
transform 1 0 27552 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_288
timestamp 1679581782
transform 1 0 28224 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_295
timestamp 1679581782
transform 1 0 28896 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_302
timestamp 1679581782
transform 1 0 29568 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_309
timestamp 1679581782
transform 1 0 30240 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_316
timestamp 1679581782
transform 1 0 30912 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_323
timestamp 1679581782
transform 1 0 31584 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_330
timestamp 1679581782
transform 1 0 32256 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_337
timestamp 1679581782
transform 1 0 32928 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_344
timestamp 1679581782
transform 1 0 33600 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_351
timestamp 1679581782
transform 1 0 34272 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_358
timestamp 1679581782
transform 1 0 34944 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_365
timestamp 1679581782
transform 1 0 35616 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_372
timestamp 1679581782
transform 1 0 36288 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_379
timestamp 1679581782
transform 1 0 36960 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_386
timestamp 1679581782
transform 1 0 37632 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_393
timestamp 1679581782
transform 1 0 38304 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_400
timestamp 1679581782
transform 1 0 38976 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_407
timestamp 1679581782
transform 1 0 39648 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_414
timestamp 1679581782
transform 1 0 40320 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_421
timestamp 1679581782
transform 1 0 40992 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_428
timestamp 1679581782
transform 1 0 41664 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_435
timestamp 1679581782
transform 1 0 42336 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_442
timestamp 1679581782
transform 1 0 43008 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_449
timestamp 1679581782
transform 1 0 43680 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_456
timestamp 1679581782
transform 1 0 44352 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_463
timestamp 1679581782
transform 1 0 45024 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_470
timestamp 1679581782
transform 1 0 45696 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_477
timestamp 1679581782
transform 1 0 46368 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_484
timestamp 1679581782
transform 1 0 47040 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_491
timestamp 1679581782
transform 1 0 47712 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_498
timestamp 1679581782
transform 1 0 48384 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_505
timestamp 1679581782
transform 1 0 49056 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_512
timestamp 1679581782
transform 1 0 49728 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_519
timestamp 1679581782
transform 1 0 50400 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_526
timestamp 1679581782
transform 1 0 51072 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_533
timestamp 1679581782
transform 1 0 51744 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_540
timestamp 1679581782
transform 1 0 52416 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_547
timestamp 1679581782
transform 1 0 53088 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_554
timestamp 1679581782
transform 1 0 53760 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_561
timestamp 1679581782
transform 1 0 54432 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_568
timestamp 1679581782
transform 1 0 55104 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_575
timestamp 1679581782
transform 1 0 55776 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_582
timestamp 1679581782
transform 1 0 56448 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_589
timestamp 1679581782
transform 1 0 57120 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_596
timestamp 1679581782
transform 1 0 57792 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_603
timestamp 1679581782
transform 1 0 58464 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_610
timestamp 1679581782
transform 1 0 59136 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_617
timestamp 1679581782
transform 1 0 59808 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_624
timestamp 1679581782
transform 1 0 60480 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_631
timestamp 1679581782
transform 1 0 61152 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_638
timestamp 1679581782
transform 1 0 61824 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_645
timestamp 1679581782
transform 1 0 62496 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_652
timestamp 1679581782
transform 1 0 63168 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_659
timestamp 1679581782
transform 1 0 63840 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_666
timestamp 1679581782
transform 1 0 64512 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_673
timestamp 1679581782
transform 1 0 65184 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_680
timestamp 1679581782
transform 1 0 65856 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_687
timestamp 1679581782
transform 1 0 66528 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_694
timestamp 1679581782
transform 1 0 67200 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_701
timestamp 1679581782
transform 1 0 67872 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_708
timestamp 1679581782
transform 1 0 68544 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_715
timestamp 1679581782
transform 1 0 69216 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_722
timestamp 1679581782
transform 1 0 69888 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_729
timestamp 1679581782
transform 1 0 70560 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_736
timestamp 1679581782
transform 1 0 71232 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_743
timestamp 1679581782
transform 1 0 71904 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_750
timestamp 1679581782
transform 1 0 72576 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_757
timestamp 1679581782
transform 1 0 73248 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_764
timestamp 1679581782
transform 1 0 73920 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_771
timestamp 1679581782
transform 1 0 74592 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_778
timestamp 1679581782
transform 1 0 75264 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_785
timestamp 1679581782
transform 1 0 75936 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_792
timestamp 1679581782
transform 1 0 76608 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_799
timestamp 1679581782
transform 1 0 77280 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_806
timestamp 1679581782
transform 1 0 77952 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_813
timestamp 1679581782
transform 1 0 78624 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_820
timestamp 1679581782
transform 1 0 79296 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_827
timestamp 1679581782
transform 1 0 79968 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_834
timestamp 1679581782
transform 1 0 80640 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_841
timestamp 1679581782
transform 1 0 81312 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_848
timestamp 1679581782
transform 1 0 81984 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_855
timestamp 1679581782
transform 1 0 82656 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_862
timestamp 1679581782
transform 1 0 83328 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_869
timestamp 1679581782
transform 1 0 84000 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_876
timestamp 1679581782
transform 1 0 84672 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_883
timestamp 1679581782
transform 1 0 85344 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_890
timestamp 1679581782
transform 1 0 86016 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_897
timestamp 1679581782
transform 1 0 86688 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_904
timestamp 1679581782
transform 1 0 87360 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_911
timestamp 1679581782
transform 1 0 88032 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_918
timestamp 1679581782
transform 1 0 88704 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_4
timestamp 1679581782
transform 1 0 960 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_11
timestamp 1679581782
transform 1 0 1632 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_18
timestamp 1679581782
transform 1 0 2304 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_25
timestamp 1679581782
transform 1 0 2976 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_32
timestamp 1679581782
transform 1 0 3648 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_39
timestamp 1679581782
transform 1 0 4320 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_46
timestamp 1679581782
transform 1 0 4992 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_53
timestamp 1679581782
transform 1 0 5664 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_60
timestamp 1679581782
transform 1 0 6336 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_67
timestamp 1679581782
transform 1 0 7008 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_74
timestamp 1679581782
transform 1 0 7680 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_81
timestamp 1679581782
transform 1 0 8352 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_88
timestamp 1679581782
transform 1 0 9024 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_95
timestamp 1679581782
transform 1 0 9696 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_102
timestamp 1679581782
transform 1 0 10368 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_109
timestamp 1679581782
transform 1 0 11040 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_116
timestamp 1679581782
transform 1 0 11712 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_123
timestamp 1679581782
transform 1 0 12384 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_130
timestamp 1679581782
transform 1 0 13056 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_137
timestamp 1679581782
transform 1 0 13728 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_144
timestamp 1679581782
transform 1 0 14400 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_151
timestamp 1679581782
transform 1 0 15072 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_158
timestamp 1679581782
transform 1 0 15744 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_165
timestamp 1679581782
transform 1 0 16416 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_172
timestamp 1679581782
transform 1 0 17088 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_179
timestamp 1679581782
transform 1 0 17760 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_186
timestamp 1679581782
transform 1 0 18432 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_193
timestamp 1679581782
transform 1 0 19104 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_200
timestamp 1679581782
transform 1 0 19776 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_207
timestamp 1679581782
transform 1 0 20448 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_214
timestamp 1679581782
transform 1 0 21120 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_221
timestamp 1679581782
transform 1 0 21792 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_228
timestamp 1679581782
transform 1 0 22464 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_235
timestamp 1679581782
transform 1 0 23136 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_242
timestamp 1679581782
transform 1 0 23808 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_249
timestamp 1679581782
transform 1 0 24480 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_256
timestamp 1679581782
transform 1 0 25152 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_263
timestamp 1679581782
transform 1 0 25824 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_270
timestamp 1679581782
transform 1 0 26496 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_277
timestamp 1679581782
transform 1 0 27168 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_284
timestamp 1679581782
transform 1 0 27840 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_291
timestamp 1679581782
transform 1 0 28512 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_298
timestamp 1679581782
transform 1 0 29184 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_305
timestamp 1679581782
transform 1 0 29856 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_312
timestamp 1679581782
transform 1 0 30528 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_319
timestamp 1679581782
transform 1 0 31200 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_326
timestamp 1679581782
transform 1 0 31872 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_333
timestamp 1679581782
transform 1 0 32544 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_340
timestamp 1679581782
transform 1 0 33216 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_347
timestamp 1679581782
transform 1 0 33888 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_354
timestamp 1679581782
transform 1 0 34560 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_361
timestamp 1679581782
transform 1 0 35232 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_368
timestamp 1679581782
transform 1 0 35904 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_375
timestamp 1679581782
transform 1 0 36576 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_382
timestamp 1679581782
transform 1 0 37248 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_389
timestamp 1679581782
transform 1 0 37920 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_396
timestamp 1679581782
transform 1 0 38592 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_403
timestamp 1679581782
transform 1 0 39264 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_410
timestamp 1679581782
transform 1 0 39936 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_417
timestamp 1679581782
transform 1 0 40608 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_424
timestamp 1679581782
transform 1 0 41280 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_431
timestamp 1679581782
transform 1 0 41952 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_438
timestamp 1679581782
transform 1 0 42624 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_445
timestamp 1679581782
transform 1 0 43296 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_452
timestamp 1679581782
transform 1 0 43968 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_459
timestamp 1679581782
transform 1 0 44640 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_466
timestamp 1679581782
transform 1 0 45312 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_473
timestamp 1679581782
transform 1 0 45984 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_480
timestamp 1679581782
transform 1 0 46656 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_487
timestamp 1679581782
transform 1 0 47328 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_494
timestamp 1679581782
transform 1 0 48000 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_501
timestamp 1679581782
transform 1 0 48672 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_508
timestamp 1679581782
transform 1 0 49344 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_515
timestamp 1679581782
transform 1 0 50016 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_522
timestamp 1679581782
transform 1 0 50688 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_529
timestamp 1679581782
transform 1 0 51360 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_536
timestamp 1679581782
transform 1 0 52032 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_543
timestamp 1679581782
transform 1 0 52704 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_550
timestamp 1679581782
transform 1 0 53376 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_557
timestamp 1679581782
transform 1 0 54048 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_564
timestamp 1679581782
transform 1 0 54720 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_571
timestamp 1679581782
transform 1 0 55392 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_578
timestamp 1679581782
transform 1 0 56064 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_585
timestamp 1679581782
transform 1 0 56736 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_592
timestamp 1679581782
transform 1 0 57408 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_599
timestamp 1679581782
transform 1 0 58080 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_606
timestamp 1679581782
transform 1 0 58752 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_613
timestamp 1679581782
transform 1 0 59424 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_620
timestamp 1679581782
transform 1 0 60096 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_627
timestamp 1679581782
transform 1 0 60768 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_634
timestamp 1679581782
transform 1 0 61440 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_641
timestamp 1679581782
transform 1 0 62112 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_648
timestamp 1679581782
transform 1 0 62784 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_655
timestamp 1679581782
transform 1 0 63456 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_662
timestamp 1679581782
transform 1 0 64128 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_669
timestamp 1679581782
transform 1 0 64800 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_676
timestamp 1679581782
transform 1 0 65472 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_683
timestamp 1679581782
transform 1 0 66144 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_690
timestamp 1679581782
transform 1 0 66816 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_697
timestamp 1679581782
transform 1 0 67488 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_704
timestamp 1679581782
transform 1 0 68160 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_711
timestamp 1679581782
transform 1 0 68832 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_718
timestamp 1679581782
transform 1 0 69504 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_725
timestamp 1679581782
transform 1 0 70176 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_732
timestamp 1679581782
transform 1 0 70848 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_739
timestamp 1679581782
transform 1 0 71520 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_746
timestamp 1679581782
transform 1 0 72192 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_753
timestamp 1679581782
transform 1 0 72864 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_760
timestamp 1679581782
transform 1 0 73536 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_767
timestamp 1679581782
transform 1 0 74208 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_774
timestamp 1679581782
transform 1 0 74880 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_781
timestamp 1679581782
transform 1 0 75552 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_788
timestamp 1679581782
transform 1 0 76224 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_795
timestamp 1679581782
transform 1 0 76896 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_802
timestamp 1679581782
transform 1 0 77568 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_809
timestamp 1679581782
transform 1 0 78240 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_816
timestamp 1679581782
transform 1 0 78912 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_823
timestamp 1679581782
transform 1 0 79584 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_830
timestamp 1679581782
transform 1 0 80256 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_837
timestamp 1679581782
transform 1 0 80928 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_844
timestamp 1679581782
transform 1 0 81600 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_851
timestamp 1679581782
transform 1 0 82272 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_858
timestamp 1679581782
transform 1 0 82944 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_865
timestamp 1679581782
transform 1 0 83616 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_872
timestamp 1679581782
transform 1 0 84288 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_879
timestamp 1679581782
transform 1 0 84960 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_886
timestamp 1679581782
transform 1 0 85632 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_893
timestamp 1679581782
transform 1 0 86304 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_900
timestamp 1679581782
transform 1 0 86976 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_907
timestamp 1679581782
transform 1 0 87648 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_914
timestamp 1679581782
transform 1 0 88320 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_43_921
timestamp 1679577901
transform 1 0 88992 0 -1 34020
box -48 -56 432 834
use sg13g2_decap_8  FILLER_44_4
timestamp 1679581782
transform 1 0 960 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_11
timestamp 1679581782
transform 1 0 1632 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_18
timestamp 1679581782
transform 1 0 2304 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_25
timestamp 1679581782
transform 1 0 2976 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_32
timestamp 1679581782
transform 1 0 3648 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_39
timestamp 1679581782
transform 1 0 4320 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_46
timestamp 1679581782
transform 1 0 4992 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_53
timestamp 1679581782
transform 1 0 5664 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_60
timestamp 1679581782
transform 1 0 6336 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_67
timestamp 1679581782
transform 1 0 7008 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_74
timestamp 1679581782
transform 1 0 7680 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_81
timestamp 1679581782
transform 1 0 8352 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_88
timestamp 1679581782
transform 1 0 9024 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_95
timestamp 1679581782
transform 1 0 9696 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_102
timestamp 1679581782
transform 1 0 10368 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_109
timestamp 1679581782
transform 1 0 11040 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_116
timestamp 1679581782
transform 1 0 11712 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_123
timestamp 1679581782
transform 1 0 12384 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_130
timestamp 1679581782
transform 1 0 13056 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_137
timestamp 1679581782
transform 1 0 13728 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_144
timestamp 1679581782
transform 1 0 14400 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_151
timestamp 1679581782
transform 1 0 15072 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_158
timestamp 1679581782
transform 1 0 15744 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_165
timestamp 1679581782
transform 1 0 16416 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_172
timestamp 1679581782
transform 1 0 17088 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_179
timestamp 1679581782
transform 1 0 17760 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_186
timestamp 1679581782
transform 1 0 18432 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_193
timestamp 1679581782
transform 1 0 19104 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_200
timestamp 1679581782
transform 1 0 19776 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_207
timestamp 1679581782
transform 1 0 20448 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_214
timestamp 1679581782
transform 1 0 21120 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_221
timestamp 1679581782
transform 1 0 21792 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_228
timestamp 1679581782
transform 1 0 22464 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_235
timestamp 1679581782
transform 1 0 23136 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_242
timestamp 1679581782
transform 1 0 23808 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_249
timestamp 1679581782
transform 1 0 24480 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_256
timestamp 1679581782
transform 1 0 25152 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_263
timestamp 1679581782
transform 1 0 25824 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_270
timestamp 1679581782
transform 1 0 26496 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_277
timestamp 1679581782
transform 1 0 27168 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_284
timestamp 1679581782
transform 1 0 27840 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_291
timestamp 1679581782
transform 1 0 28512 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_298
timestamp 1679581782
transform 1 0 29184 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_305
timestamp 1679581782
transform 1 0 29856 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_312
timestamp 1679581782
transform 1 0 30528 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_319
timestamp 1679581782
transform 1 0 31200 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_326
timestamp 1679581782
transform 1 0 31872 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_333
timestamp 1679581782
transform 1 0 32544 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_340
timestamp 1679581782
transform 1 0 33216 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_347
timestamp 1679581782
transform 1 0 33888 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_354
timestamp 1679581782
transform 1 0 34560 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_361
timestamp 1679581782
transform 1 0 35232 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_368
timestamp 1679581782
transform 1 0 35904 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_375
timestamp 1679581782
transform 1 0 36576 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_382
timestamp 1679581782
transform 1 0 37248 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_389
timestamp 1679581782
transform 1 0 37920 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_396
timestamp 1679581782
transform 1 0 38592 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_403
timestamp 1679581782
transform 1 0 39264 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_410
timestamp 1679581782
transform 1 0 39936 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_417
timestamp 1679581782
transform 1 0 40608 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_424
timestamp 1679581782
transform 1 0 41280 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_431
timestamp 1679581782
transform 1 0 41952 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_438
timestamp 1679581782
transform 1 0 42624 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_445
timestamp 1679581782
transform 1 0 43296 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_452
timestamp 1679581782
transform 1 0 43968 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_459
timestamp 1679581782
transform 1 0 44640 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_466
timestamp 1679581782
transform 1 0 45312 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_473
timestamp 1679581782
transform 1 0 45984 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_480
timestamp 1679581782
transform 1 0 46656 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_487
timestamp 1679581782
transform 1 0 47328 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_494
timestamp 1679581782
transform 1 0 48000 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_501
timestamp 1679581782
transform 1 0 48672 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_508
timestamp 1679581782
transform 1 0 49344 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_515
timestamp 1679581782
transform 1 0 50016 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_522
timestamp 1679581782
transform 1 0 50688 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_529
timestamp 1679581782
transform 1 0 51360 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_536
timestamp 1679581782
transform 1 0 52032 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_543
timestamp 1679581782
transform 1 0 52704 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_550
timestamp 1679581782
transform 1 0 53376 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_557
timestamp 1679581782
transform 1 0 54048 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_564
timestamp 1679581782
transform 1 0 54720 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_571
timestamp 1679581782
transform 1 0 55392 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_578
timestamp 1679581782
transform 1 0 56064 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_585
timestamp 1679581782
transform 1 0 56736 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_592
timestamp 1679581782
transform 1 0 57408 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_599
timestamp 1679581782
transform 1 0 58080 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_606
timestamp 1679581782
transform 1 0 58752 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_613
timestamp 1679581782
transform 1 0 59424 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_620
timestamp 1679581782
transform 1 0 60096 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_627
timestamp 1679581782
transform 1 0 60768 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_634
timestamp 1679581782
transform 1 0 61440 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_641
timestamp 1679581782
transform 1 0 62112 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_648
timestamp 1679581782
transform 1 0 62784 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_655
timestamp 1679581782
transform 1 0 63456 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_662
timestamp 1679581782
transform 1 0 64128 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_669
timestamp 1679581782
transform 1 0 64800 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_676
timestamp 1679581782
transform 1 0 65472 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_683
timestamp 1679581782
transform 1 0 66144 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_690
timestamp 1679581782
transform 1 0 66816 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_697
timestamp 1679581782
transform 1 0 67488 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_704
timestamp 1679581782
transform 1 0 68160 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_711
timestamp 1679581782
transform 1 0 68832 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_718
timestamp 1679581782
transform 1 0 69504 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_725
timestamp 1679581782
transform 1 0 70176 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_732
timestamp 1679581782
transform 1 0 70848 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_739
timestamp 1679581782
transform 1 0 71520 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_746
timestamp 1679581782
transform 1 0 72192 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_753
timestamp 1679581782
transform 1 0 72864 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_760
timestamp 1679581782
transform 1 0 73536 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_767
timestamp 1679581782
transform 1 0 74208 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_774
timestamp 1679581782
transform 1 0 74880 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_781
timestamp 1679581782
transform 1 0 75552 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_788
timestamp 1679581782
transform 1 0 76224 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_795
timestamp 1679581782
transform 1 0 76896 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_802
timestamp 1679581782
transform 1 0 77568 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_809
timestamp 1679581782
transform 1 0 78240 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_816
timestamp 1679581782
transform 1 0 78912 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_823
timestamp 1679581782
transform 1 0 79584 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_830
timestamp 1679581782
transform 1 0 80256 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_837
timestamp 1679581782
transform 1 0 80928 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_844
timestamp 1679581782
transform 1 0 81600 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_851
timestamp 1679581782
transform 1 0 82272 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_858
timestamp 1679581782
transform 1 0 82944 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_865
timestamp 1679581782
transform 1 0 83616 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_872
timestamp 1679581782
transform 1 0 84288 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_879
timestamp 1679581782
transform 1 0 84960 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_886
timestamp 1679581782
transform 1 0 85632 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_893
timestamp 1679581782
transform 1 0 86304 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_900
timestamp 1679581782
transform 1 0 86976 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_907
timestamp 1679581782
transform 1 0 87648 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_914
timestamp 1679581782
transform 1 0 88320 0 1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_44_921
timestamp 1679577901
transform 1 0 88992 0 1 34020
box -48 -56 432 834
use sg13g2_decap_8  FILLER_45_4
timestamp 1679581782
transform 1 0 960 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_11
timestamp 1679581782
transform 1 0 1632 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_18
timestamp 1679581782
transform 1 0 2304 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_25
timestamp 1679581782
transform 1 0 2976 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_32
timestamp 1679581782
transform 1 0 3648 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_39
timestamp 1679581782
transform 1 0 4320 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_46
timestamp 1679581782
transform 1 0 4992 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_53
timestamp 1679581782
transform 1 0 5664 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_60
timestamp 1679581782
transform 1 0 6336 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_67
timestamp 1679581782
transform 1 0 7008 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_74
timestamp 1679581782
transform 1 0 7680 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_81
timestamp 1679581782
transform 1 0 8352 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_88
timestamp 1679581782
transform 1 0 9024 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_95
timestamp 1679581782
transform 1 0 9696 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_102
timestamp 1679581782
transform 1 0 10368 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_109
timestamp 1679581782
transform 1 0 11040 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_116
timestamp 1679581782
transform 1 0 11712 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_123
timestamp 1679581782
transform 1 0 12384 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_130
timestamp 1679581782
transform 1 0 13056 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_137
timestamp 1679581782
transform 1 0 13728 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_144
timestamp 1679581782
transform 1 0 14400 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_151
timestamp 1679581782
transform 1 0 15072 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_158
timestamp 1679581782
transform 1 0 15744 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_165
timestamp 1679581782
transform 1 0 16416 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_172
timestamp 1679581782
transform 1 0 17088 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_179
timestamp 1679581782
transform 1 0 17760 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_186
timestamp 1679581782
transform 1 0 18432 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_193
timestamp 1679581782
transform 1 0 19104 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_200
timestamp 1679581782
transform 1 0 19776 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_207
timestamp 1679581782
transform 1 0 20448 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_214
timestamp 1679581782
transform 1 0 21120 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_221
timestamp 1679581782
transform 1 0 21792 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_228
timestamp 1679581782
transform 1 0 22464 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_235
timestamp 1679581782
transform 1 0 23136 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_242
timestamp 1679581782
transform 1 0 23808 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_249
timestamp 1679581782
transform 1 0 24480 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_256
timestamp 1679581782
transform 1 0 25152 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_263
timestamp 1679581782
transform 1 0 25824 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_270
timestamp 1679581782
transform 1 0 26496 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_277
timestamp 1679581782
transform 1 0 27168 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_284
timestamp 1679581782
transform 1 0 27840 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_291
timestamp 1679581782
transform 1 0 28512 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_298
timestamp 1679581782
transform 1 0 29184 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_305
timestamp 1679581782
transform 1 0 29856 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_312
timestamp 1679581782
transform 1 0 30528 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_319
timestamp 1679581782
transform 1 0 31200 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_326
timestamp 1679581782
transform 1 0 31872 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_333
timestamp 1679581782
transform 1 0 32544 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_340
timestamp 1679581782
transform 1 0 33216 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_347
timestamp 1679581782
transform 1 0 33888 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_354
timestamp 1679581782
transform 1 0 34560 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_361
timestamp 1679581782
transform 1 0 35232 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_368
timestamp 1679581782
transform 1 0 35904 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_375
timestamp 1679581782
transform 1 0 36576 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_382
timestamp 1679581782
transform 1 0 37248 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_389
timestamp 1679581782
transform 1 0 37920 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_396
timestamp 1679581782
transform 1 0 38592 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_403
timestamp 1679581782
transform 1 0 39264 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_410
timestamp 1679581782
transform 1 0 39936 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_417
timestamp 1679581782
transform 1 0 40608 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_424
timestamp 1679581782
transform 1 0 41280 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_431
timestamp 1679581782
transform 1 0 41952 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_438
timestamp 1679581782
transform 1 0 42624 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_445
timestamp 1679581782
transform 1 0 43296 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_452
timestamp 1679581782
transform 1 0 43968 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_459
timestamp 1679581782
transform 1 0 44640 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_466
timestamp 1679581782
transform 1 0 45312 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_473
timestamp 1679581782
transform 1 0 45984 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_480
timestamp 1679581782
transform 1 0 46656 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_487
timestamp 1679581782
transform 1 0 47328 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_494
timestamp 1679581782
transform 1 0 48000 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_501
timestamp 1679581782
transform 1 0 48672 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_508
timestamp 1679581782
transform 1 0 49344 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_515
timestamp 1679581782
transform 1 0 50016 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_522
timestamp 1679581782
transform 1 0 50688 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_529
timestamp 1679581782
transform 1 0 51360 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_536
timestamp 1679581782
transform 1 0 52032 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_543
timestamp 1679581782
transform 1 0 52704 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_550
timestamp 1679581782
transform 1 0 53376 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_557
timestamp 1679581782
transform 1 0 54048 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_564
timestamp 1679581782
transform 1 0 54720 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_571
timestamp 1679581782
transform 1 0 55392 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_578
timestamp 1679581782
transform 1 0 56064 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_585
timestamp 1679581782
transform 1 0 56736 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_592
timestamp 1679581782
transform 1 0 57408 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_599
timestamp 1679581782
transform 1 0 58080 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_606
timestamp 1679581782
transform 1 0 58752 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_613
timestamp 1679581782
transform 1 0 59424 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_620
timestamp 1679581782
transform 1 0 60096 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_627
timestamp 1679581782
transform 1 0 60768 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_634
timestamp 1679581782
transform 1 0 61440 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_641
timestamp 1679581782
transform 1 0 62112 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_648
timestamp 1679581782
transform 1 0 62784 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_655
timestamp 1679581782
transform 1 0 63456 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_662
timestamp 1679581782
transform 1 0 64128 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_669
timestamp 1679581782
transform 1 0 64800 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_676
timestamp 1679581782
transform 1 0 65472 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_683
timestamp 1679581782
transform 1 0 66144 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_690
timestamp 1679581782
transform 1 0 66816 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_697
timestamp 1679581782
transform 1 0 67488 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_704
timestamp 1679581782
transform 1 0 68160 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_711
timestamp 1679581782
transform 1 0 68832 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_718
timestamp 1679581782
transform 1 0 69504 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_725
timestamp 1679581782
transform 1 0 70176 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_732
timestamp 1679581782
transform 1 0 70848 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_739
timestamp 1679581782
transform 1 0 71520 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_746
timestamp 1679581782
transform 1 0 72192 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_753
timestamp 1679581782
transform 1 0 72864 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_760
timestamp 1679581782
transform 1 0 73536 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_767
timestamp 1679581782
transform 1 0 74208 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_774
timestamp 1679581782
transform 1 0 74880 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_781
timestamp 1679581782
transform 1 0 75552 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_788
timestamp 1679581782
transform 1 0 76224 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_795
timestamp 1679581782
transform 1 0 76896 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_802
timestamp 1679581782
transform 1 0 77568 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_809
timestamp 1679581782
transform 1 0 78240 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_816
timestamp 1679581782
transform 1 0 78912 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_823
timestamp 1679581782
transform 1 0 79584 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_830
timestamp 1679581782
transform 1 0 80256 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_837
timestamp 1679581782
transform 1 0 80928 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_844
timestamp 1679581782
transform 1 0 81600 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_851
timestamp 1679581782
transform 1 0 82272 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_858
timestamp 1679581782
transform 1 0 82944 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_865
timestamp 1679581782
transform 1 0 83616 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_872
timestamp 1679581782
transform 1 0 84288 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_879
timestamp 1679581782
transform 1 0 84960 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_886
timestamp 1679581782
transform 1 0 85632 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_893
timestamp 1679581782
transform 1 0 86304 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_900
timestamp 1679581782
transform 1 0 86976 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_907
timestamp 1679581782
transform 1 0 87648 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_914
timestamp 1679581782
transform 1 0 88320 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_45_921
timestamp 1679577901
transform 1 0 88992 0 -1 35532
box -48 -56 432 834
use sg13g2_decap_8  FILLER_46_0
timestamp 1679581782
transform 1 0 576 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_7
timestamp 1679581782
transform 1 0 1248 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_14
timestamp 1679581782
transform 1 0 1920 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_21
timestamp 1679581782
transform 1 0 2592 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_28
timestamp 1679581782
transform 1 0 3264 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_35
timestamp 1679581782
transform 1 0 3936 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_42
timestamp 1679581782
transform 1 0 4608 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_49
timestamp 1679581782
transform 1 0 5280 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_56
timestamp 1679581782
transform 1 0 5952 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_63
timestamp 1679581782
transform 1 0 6624 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_70
timestamp 1679581782
transform 1 0 7296 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_77
timestamp 1679581782
transform 1 0 7968 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_84
timestamp 1679581782
transform 1 0 8640 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_91
timestamp 1679581782
transform 1 0 9312 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_98
timestamp 1679581782
transform 1 0 9984 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_105
timestamp 1679581782
transform 1 0 10656 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_112
timestamp 1679581782
transform 1 0 11328 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_119
timestamp 1679581782
transform 1 0 12000 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_126
timestamp 1679581782
transform 1 0 12672 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_133
timestamp 1679581782
transform 1 0 13344 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_140
timestamp 1679581782
transform 1 0 14016 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_147
timestamp 1679581782
transform 1 0 14688 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_154
timestamp 1679581782
transform 1 0 15360 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_161
timestamp 1679581782
transform 1 0 16032 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_168
timestamp 1679581782
transform 1 0 16704 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_175
timestamp 1679581782
transform 1 0 17376 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_182
timestamp 1679581782
transform 1 0 18048 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_189
timestamp 1679581782
transform 1 0 18720 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_196
timestamp 1679581782
transform 1 0 19392 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_203
timestamp 1679581782
transform 1 0 20064 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_210
timestamp 1679581782
transform 1 0 20736 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_217
timestamp 1679581782
transform 1 0 21408 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_224
timestamp 1679581782
transform 1 0 22080 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_231
timestamp 1679581782
transform 1 0 22752 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_238
timestamp 1679581782
transform 1 0 23424 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_245
timestamp 1679581782
transform 1 0 24096 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_252
timestamp 1679581782
transform 1 0 24768 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_259
timestamp 1679581782
transform 1 0 25440 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_266
timestamp 1679581782
transform 1 0 26112 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_273
timestamp 1679581782
transform 1 0 26784 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_280
timestamp 1679581782
transform 1 0 27456 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_287
timestamp 1679581782
transform 1 0 28128 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_294
timestamp 1679581782
transform 1 0 28800 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_301
timestamp 1679581782
transform 1 0 29472 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_308
timestamp 1679581782
transform 1 0 30144 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_315
timestamp 1679581782
transform 1 0 30816 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_322
timestamp 1679581782
transform 1 0 31488 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_329
timestamp 1679581782
transform 1 0 32160 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_336
timestamp 1679581782
transform 1 0 32832 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_343
timestamp 1679581782
transform 1 0 33504 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_350
timestamp 1679581782
transform 1 0 34176 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_357
timestamp 1679581782
transform 1 0 34848 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_364
timestamp 1679581782
transform 1 0 35520 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_371
timestamp 1679581782
transform 1 0 36192 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_378
timestamp 1679581782
transform 1 0 36864 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_385
timestamp 1679581782
transform 1 0 37536 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_392
timestamp 1679581782
transform 1 0 38208 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_399
timestamp 1679581782
transform 1 0 38880 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_406
timestamp 1679581782
transform 1 0 39552 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_413
timestamp 1679581782
transform 1 0 40224 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_420
timestamp 1679581782
transform 1 0 40896 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_427
timestamp 1679581782
transform 1 0 41568 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_434
timestamp 1679581782
transform 1 0 42240 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_441
timestamp 1679581782
transform 1 0 42912 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_448
timestamp 1679581782
transform 1 0 43584 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_455
timestamp 1679581782
transform 1 0 44256 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_462
timestamp 1679581782
transform 1 0 44928 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_469
timestamp 1679581782
transform 1 0 45600 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_476
timestamp 1679581782
transform 1 0 46272 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_483
timestamp 1679581782
transform 1 0 46944 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_490
timestamp 1679581782
transform 1 0 47616 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_497
timestamp 1679581782
transform 1 0 48288 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_504
timestamp 1679581782
transform 1 0 48960 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_511
timestamp 1679581782
transform 1 0 49632 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_518
timestamp 1679581782
transform 1 0 50304 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_525
timestamp 1679581782
transform 1 0 50976 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_532
timestamp 1679581782
transform 1 0 51648 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_539
timestamp 1679581782
transform 1 0 52320 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_546
timestamp 1679581782
transform 1 0 52992 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_553
timestamp 1679581782
transform 1 0 53664 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_560
timestamp 1679581782
transform 1 0 54336 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_567
timestamp 1679581782
transform 1 0 55008 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_574
timestamp 1679581782
transform 1 0 55680 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_581
timestamp 1679581782
transform 1 0 56352 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_588
timestamp 1679581782
transform 1 0 57024 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_595
timestamp 1679581782
transform 1 0 57696 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_602
timestamp 1679581782
transform 1 0 58368 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_609
timestamp 1679581782
transform 1 0 59040 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_616
timestamp 1679581782
transform 1 0 59712 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_623
timestamp 1679581782
transform 1 0 60384 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_630
timestamp 1679581782
transform 1 0 61056 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_637
timestamp 1679581782
transform 1 0 61728 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_644
timestamp 1679581782
transform 1 0 62400 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_651
timestamp 1679581782
transform 1 0 63072 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_658
timestamp 1679581782
transform 1 0 63744 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_665
timestamp 1679581782
transform 1 0 64416 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_672
timestamp 1679581782
transform 1 0 65088 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_679
timestamp 1679581782
transform 1 0 65760 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_686
timestamp 1679581782
transform 1 0 66432 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_693
timestamp 1679581782
transform 1 0 67104 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_700
timestamp 1679581782
transform 1 0 67776 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_707
timestamp 1679581782
transform 1 0 68448 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_714
timestamp 1679581782
transform 1 0 69120 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_721
timestamp 1679581782
transform 1 0 69792 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_728
timestamp 1679581782
transform 1 0 70464 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_735
timestamp 1679581782
transform 1 0 71136 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_742
timestamp 1679581782
transform 1 0 71808 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_749
timestamp 1679581782
transform 1 0 72480 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_756
timestamp 1679581782
transform 1 0 73152 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_763
timestamp 1679581782
transform 1 0 73824 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_770
timestamp 1679581782
transform 1 0 74496 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_777
timestamp 1679581782
transform 1 0 75168 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_784
timestamp 1679581782
transform 1 0 75840 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_791
timestamp 1679581782
transform 1 0 76512 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_798
timestamp 1679581782
transform 1 0 77184 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_805
timestamp 1679581782
transform 1 0 77856 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_812
timestamp 1679581782
transform 1 0 78528 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_819
timestamp 1679581782
transform 1 0 79200 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_826
timestamp 1679581782
transform 1 0 79872 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_833
timestamp 1679581782
transform 1 0 80544 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_840
timestamp 1679581782
transform 1 0 81216 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_847
timestamp 1679581782
transform 1 0 81888 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_854
timestamp 1679581782
transform 1 0 82560 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_861
timestamp 1679581782
transform 1 0 83232 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_868
timestamp 1679581782
transform 1 0 83904 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_875
timestamp 1679581782
transform 1 0 84576 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_882
timestamp 1679581782
transform 1 0 85248 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_889
timestamp 1679581782
transform 1 0 85920 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_896
timestamp 1679581782
transform 1 0 86592 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_903
timestamp 1679581782
transform 1 0 87264 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_910
timestamp 1679581782
transform 1 0 87936 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_917
timestamp 1679581782
transform 1 0 88608 0 1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_46_924
timestamp 1677579658
transform 1 0 89280 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_47_0
timestamp 1679581782
transform 1 0 576 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_7
timestamp 1679581782
transform 1 0 1248 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_14
timestamp 1679581782
transform 1 0 1920 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_21
timestamp 1679581782
transform 1 0 2592 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_28
timestamp 1679581782
transform 1 0 3264 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_35
timestamp 1679581782
transform 1 0 3936 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_42
timestamp 1679581782
transform 1 0 4608 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_49
timestamp 1679581782
transform 1 0 5280 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_56
timestamp 1679581782
transform 1 0 5952 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_63
timestamp 1679581782
transform 1 0 6624 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_70
timestamp 1679581782
transform 1 0 7296 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_77
timestamp 1679581782
transform 1 0 7968 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_84
timestamp 1679581782
transform 1 0 8640 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_91
timestamp 1679581782
transform 1 0 9312 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_98
timestamp 1679581782
transform 1 0 9984 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_105
timestamp 1679581782
transform 1 0 10656 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_112
timestamp 1679581782
transform 1 0 11328 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_119
timestamp 1679581782
transform 1 0 12000 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_126
timestamp 1679581782
transform 1 0 12672 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_133
timestamp 1679581782
transform 1 0 13344 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_140
timestamp 1679581782
transform 1 0 14016 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_147
timestamp 1679581782
transform 1 0 14688 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_154
timestamp 1679581782
transform 1 0 15360 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_161
timestamp 1679581782
transform 1 0 16032 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_168
timestamp 1679581782
transform 1 0 16704 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_175
timestamp 1679581782
transform 1 0 17376 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_182
timestamp 1679581782
transform 1 0 18048 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_189
timestamp 1679581782
transform 1 0 18720 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_196
timestamp 1679581782
transform 1 0 19392 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_203
timestamp 1679581782
transform 1 0 20064 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_210
timestamp 1679581782
transform 1 0 20736 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_217
timestamp 1679581782
transform 1 0 21408 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_224
timestamp 1679581782
transform 1 0 22080 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_231
timestamp 1679581782
transform 1 0 22752 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_238
timestamp 1679581782
transform 1 0 23424 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_245
timestamp 1679581782
transform 1 0 24096 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_252
timestamp 1679581782
transform 1 0 24768 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_259
timestamp 1679581782
transform 1 0 25440 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_266
timestamp 1679581782
transform 1 0 26112 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_273
timestamp 1679581782
transform 1 0 26784 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_280
timestamp 1679581782
transform 1 0 27456 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_287
timestamp 1679581782
transform 1 0 28128 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_294
timestamp 1679581782
transform 1 0 28800 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_301
timestamp 1679581782
transform 1 0 29472 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_308
timestamp 1679581782
transform 1 0 30144 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_315
timestamp 1679581782
transform 1 0 30816 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_322
timestamp 1679581782
transform 1 0 31488 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_329
timestamp 1679581782
transform 1 0 32160 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_336
timestamp 1679581782
transform 1 0 32832 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_343
timestamp 1679581782
transform 1 0 33504 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_350
timestamp 1679581782
transform 1 0 34176 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_357
timestamp 1679581782
transform 1 0 34848 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_364
timestamp 1679581782
transform 1 0 35520 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_371
timestamp 1679581782
transform 1 0 36192 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_378
timestamp 1679581782
transform 1 0 36864 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_385
timestamp 1679581782
transform 1 0 37536 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_392
timestamp 1679581782
transform 1 0 38208 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_399
timestamp 1679581782
transform 1 0 38880 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_406
timestamp 1679581782
transform 1 0 39552 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_413
timestamp 1679581782
transform 1 0 40224 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_420
timestamp 1679581782
transform 1 0 40896 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_427
timestamp 1679581782
transform 1 0 41568 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_434
timestamp 1679581782
transform 1 0 42240 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_441
timestamp 1679581782
transform 1 0 42912 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_448
timestamp 1679581782
transform 1 0 43584 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_455
timestamp 1679581782
transform 1 0 44256 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_462
timestamp 1679581782
transform 1 0 44928 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_469
timestamp 1679581782
transform 1 0 45600 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_476
timestamp 1679581782
transform 1 0 46272 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_483
timestamp 1679581782
transform 1 0 46944 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_490
timestamp 1679581782
transform 1 0 47616 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_497
timestamp 1679581782
transform 1 0 48288 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_504
timestamp 1679581782
transform 1 0 48960 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_511
timestamp 1679581782
transform 1 0 49632 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_518
timestamp 1679581782
transform 1 0 50304 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_525
timestamp 1679581782
transform 1 0 50976 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_532
timestamp 1679581782
transform 1 0 51648 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_539
timestamp 1679581782
transform 1 0 52320 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_546
timestamp 1679581782
transform 1 0 52992 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_553
timestamp 1679581782
transform 1 0 53664 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_560
timestamp 1679581782
transform 1 0 54336 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_567
timestamp 1679581782
transform 1 0 55008 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_574
timestamp 1679581782
transform 1 0 55680 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_581
timestamp 1679581782
transform 1 0 56352 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_588
timestamp 1679581782
transform 1 0 57024 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_595
timestamp 1679581782
transform 1 0 57696 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_602
timestamp 1679581782
transform 1 0 58368 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_609
timestamp 1679581782
transform 1 0 59040 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_616
timestamp 1679581782
transform 1 0 59712 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_623
timestamp 1679581782
transform 1 0 60384 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_630
timestamp 1679581782
transform 1 0 61056 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_637
timestamp 1679581782
transform 1 0 61728 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_644
timestamp 1679581782
transform 1 0 62400 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_651
timestamp 1679581782
transform 1 0 63072 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_658
timestamp 1679581782
transform 1 0 63744 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_665
timestamp 1679581782
transform 1 0 64416 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_672
timestamp 1679581782
transform 1 0 65088 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_679
timestamp 1679581782
transform 1 0 65760 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_686
timestamp 1679581782
transform 1 0 66432 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_693
timestamp 1679581782
transform 1 0 67104 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_700
timestamp 1679581782
transform 1 0 67776 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_707
timestamp 1679581782
transform 1 0 68448 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_714
timestamp 1679581782
transform 1 0 69120 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_721
timestamp 1679581782
transform 1 0 69792 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_728
timestamp 1679581782
transform 1 0 70464 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_735
timestamp 1679581782
transform 1 0 71136 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_742
timestamp 1679581782
transform 1 0 71808 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_749
timestamp 1679581782
transform 1 0 72480 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_756
timestamp 1679581782
transform 1 0 73152 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_763
timestamp 1679581782
transform 1 0 73824 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_770
timestamp 1679581782
transform 1 0 74496 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_777
timestamp 1679581782
transform 1 0 75168 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_784
timestamp 1679581782
transform 1 0 75840 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_791
timestamp 1679581782
transform 1 0 76512 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_798
timestamp 1679581782
transform 1 0 77184 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_805
timestamp 1679581782
transform 1 0 77856 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_812
timestamp 1679581782
transform 1 0 78528 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_819
timestamp 1679581782
transform 1 0 79200 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_826
timestamp 1679581782
transform 1 0 79872 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_833
timestamp 1679581782
transform 1 0 80544 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_840
timestamp 1679581782
transform 1 0 81216 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_847
timestamp 1679581782
transform 1 0 81888 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_854
timestamp 1679581782
transform 1 0 82560 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_861
timestamp 1679581782
transform 1 0 83232 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_868
timestamp 1679581782
transform 1 0 83904 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_875
timestamp 1679581782
transform 1 0 84576 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_882
timestamp 1679581782
transform 1 0 85248 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_889
timestamp 1679581782
transform 1 0 85920 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_896
timestamp 1679581782
transform 1 0 86592 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_903
timestamp 1679581782
transform 1 0 87264 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_910
timestamp 1679581782
transform 1 0 87936 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_917
timestamp 1679581782
transform 1 0 88608 0 -1 37044
box -48 -56 720 834
use sg13g2_fill_1  FILLER_47_924
timestamp 1677579658
transform 1 0 89280 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_48_0
timestamp 1679581782
transform 1 0 576 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_7
timestamp 1679581782
transform 1 0 1248 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_14
timestamp 1679581782
transform 1 0 1920 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_21
timestamp 1679581782
transform 1 0 2592 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_28
timestamp 1679581782
transform 1 0 3264 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_35
timestamp 1679581782
transform 1 0 3936 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_42
timestamp 1679581782
transform 1 0 4608 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_49
timestamp 1679581782
transform 1 0 5280 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_56
timestamp 1679581782
transform 1 0 5952 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_63
timestamp 1679581782
transform 1 0 6624 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_70
timestamp 1679581782
transform 1 0 7296 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_77
timestamp 1679581782
transform 1 0 7968 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_84
timestamp 1679581782
transform 1 0 8640 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_91
timestamp 1679581782
transform 1 0 9312 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_98
timestamp 1679581782
transform 1 0 9984 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_105
timestamp 1679581782
transform 1 0 10656 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_112
timestamp 1679581782
transform 1 0 11328 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_119
timestamp 1679581782
transform 1 0 12000 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_126
timestamp 1679581782
transform 1 0 12672 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_133
timestamp 1679581782
transform 1 0 13344 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_140
timestamp 1679581782
transform 1 0 14016 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_147
timestamp 1679581782
transform 1 0 14688 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_154
timestamp 1679581782
transform 1 0 15360 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_161
timestamp 1679581782
transform 1 0 16032 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_168
timestamp 1679581782
transform 1 0 16704 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_175
timestamp 1679581782
transform 1 0 17376 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_182
timestamp 1679581782
transform 1 0 18048 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_189
timestamp 1679581782
transform 1 0 18720 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_196
timestamp 1679581782
transform 1 0 19392 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_203
timestamp 1679581782
transform 1 0 20064 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_210
timestamp 1679581782
transform 1 0 20736 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_217
timestamp 1679581782
transform 1 0 21408 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_224
timestamp 1679581782
transform 1 0 22080 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_231
timestamp 1679581782
transform 1 0 22752 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_238
timestamp 1679581782
transform 1 0 23424 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_245
timestamp 1679581782
transform 1 0 24096 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_252
timestamp 1679581782
transform 1 0 24768 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_259
timestamp 1679581782
transform 1 0 25440 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_266
timestamp 1679581782
transform 1 0 26112 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_273
timestamp 1679581782
transform 1 0 26784 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_280
timestamp 1679581782
transform 1 0 27456 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_287
timestamp 1679581782
transform 1 0 28128 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_294
timestamp 1679581782
transform 1 0 28800 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_301
timestamp 1679581782
transform 1 0 29472 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_308
timestamp 1679581782
transform 1 0 30144 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_315
timestamp 1679581782
transform 1 0 30816 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_322
timestamp 1679581782
transform 1 0 31488 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_329
timestamp 1679581782
transform 1 0 32160 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_336
timestamp 1679581782
transform 1 0 32832 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_343
timestamp 1679581782
transform 1 0 33504 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_350
timestamp 1679581782
transform 1 0 34176 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_357
timestamp 1679581782
transform 1 0 34848 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_364
timestamp 1679581782
transform 1 0 35520 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_371
timestamp 1679581782
transform 1 0 36192 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_378
timestamp 1679581782
transform 1 0 36864 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_385
timestamp 1679581782
transform 1 0 37536 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_392
timestamp 1679581782
transform 1 0 38208 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_399
timestamp 1679581782
transform 1 0 38880 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_406
timestamp 1679581782
transform 1 0 39552 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_413
timestamp 1679581782
transform 1 0 40224 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_420
timestamp 1679581782
transform 1 0 40896 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_427
timestamp 1679581782
transform 1 0 41568 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_434
timestamp 1679581782
transform 1 0 42240 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_441
timestamp 1679581782
transform 1 0 42912 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_448
timestamp 1679581782
transform 1 0 43584 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_455
timestamp 1679581782
transform 1 0 44256 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_462
timestamp 1679581782
transform 1 0 44928 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_469
timestamp 1679581782
transform 1 0 45600 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_476
timestamp 1679581782
transform 1 0 46272 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_483
timestamp 1679581782
transform 1 0 46944 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_490
timestamp 1679581782
transform 1 0 47616 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_497
timestamp 1679581782
transform 1 0 48288 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_504
timestamp 1679581782
transform 1 0 48960 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_511
timestamp 1679581782
transform 1 0 49632 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_518
timestamp 1679581782
transform 1 0 50304 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_525
timestamp 1679581782
transform 1 0 50976 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_532
timestamp 1679581782
transform 1 0 51648 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_539
timestamp 1679581782
transform 1 0 52320 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_546
timestamp 1679581782
transform 1 0 52992 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_553
timestamp 1679581782
transform 1 0 53664 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_560
timestamp 1679581782
transform 1 0 54336 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_567
timestamp 1679581782
transform 1 0 55008 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_574
timestamp 1679581782
transform 1 0 55680 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_581
timestamp 1679581782
transform 1 0 56352 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_588
timestamp 1679581782
transform 1 0 57024 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_595
timestamp 1679581782
transform 1 0 57696 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_602
timestamp 1679581782
transform 1 0 58368 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_609
timestamp 1679581782
transform 1 0 59040 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_616
timestamp 1679581782
transform 1 0 59712 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_623
timestamp 1679581782
transform 1 0 60384 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_630
timestamp 1679581782
transform 1 0 61056 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_637
timestamp 1679581782
transform 1 0 61728 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_644
timestamp 1679581782
transform 1 0 62400 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_651
timestamp 1679581782
transform 1 0 63072 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_658
timestamp 1679581782
transform 1 0 63744 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_665
timestamp 1679581782
transform 1 0 64416 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_672
timestamp 1679581782
transform 1 0 65088 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_679
timestamp 1679581782
transform 1 0 65760 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_686
timestamp 1679581782
transform 1 0 66432 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_693
timestamp 1679581782
transform 1 0 67104 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_700
timestamp 1679581782
transform 1 0 67776 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_707
timestamp 1679581782
transform 1 0 68448 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_714
timestamp 1679581782
transform 1 0 69120 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_721
timestamp 1679581782
transform 1 0 69792 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_728
timestamp 1679581782
transform 1 0 70464 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_735
timestamp 1679581782
transform 1 0 71136 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_742
timestamp 1679581782
transform 1 0 71808 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_749
timestamp 1679581782
transform 1 0 72480 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_756
timestamp 1679581782
transform 1 0 73152 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_763
timestamp 1679581782
transform 1 0 73824 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_770
timestamp 1679581782
transform 1 0 74496 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_777
timestamp 1679581782
transform 1 0 75168 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_784
timestamp 1679581782
transform 1 0 75840 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_791
timestamp 1679581782
transform 1 0 76512 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_798
timestamp 1679581782
transform 1 0 77184 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_805
timestamp 1679581782
transform 1 0 77856 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_812
timestamp 1679581782
transform 1 0 78528 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_819
timestamp 1679581782
transform 1 0 79200 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_826
timestamp 1679581782
transform 1 0 79872 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_833
timestamp 1679581782
transform 1 0 80544 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_840
timestamp 1679581782
transform 1 0 81216 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_847
timestamp 1679581782
transform 1 0 81888 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_854
timestamp 1679581782
transform 1 0 82560 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_861
timestamp 1679581782
transform 1 0 83232 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_868
timestamp 1679581782
transform 1 0 83904 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_875
timestamp 1679581782
transform 1 0 84576 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_882
timestamp 1679581782
transform 1 0 85248 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_889
timestamp 1679581782
transform 1 0 85920 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_896
timestamp 1679581782
transform 1 0 86592 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_903
timestamp 1679581782
transform 1 0 87264 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_910
timestamp 1679581782
transform 1 0 87936 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_917
timestamp 1679581782
transform 1 0 88608 0 1 37044
box -48 -56 720 834
use sg13g2_fill_1  FILLER_48_924
timestamp 1677579658
transform 1 0 89280 0 1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_49_0
timestamp 1679581782
transform 1 0 576 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_7
timestamp 1679581782
transform 1 0 1248 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_14
timestamp 1679581782
transform 1 0 1920 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_21
timestamp 1679581782
transform 1 0 2592 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_28
timestamp 1679581782
transform 1 0 3264 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_35
timestamp 1679581782
transform 1 0 3936 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_42
timestamp 1679581782
transform 1 0 4608 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_49
timestamp 1679581782
transform 1 0 5280 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_56
timestamp 1679581782
transform 1 0 5952 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_63
timestamp 1679581782
transform 1 0 6624 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_70
timestamp 1679581782
transform 1 0 7296 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_77
timestamp 1679581782
transform 1 0 7968 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_84
timestamp 1679581782
transform 1 0 8640 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_91
timestamp 1679581782
transform 1 0 9312 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_98
timestamp 1679581782
transform 1 0 9984 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_105
timestamp 1679581782
transform 1 0 10656 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_112
timestamp 1679581782
transform 1 0 11328 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_119
timestamp 1679581782
transform 1 0 12000 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_126
timestamp 1679581782
transform 1 0 12672 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_133
timestamp 1679581782
transform 1 0 13344 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_140
timestamp 1679581782
transform 1 0 14016 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_147
timestamp 1679581782
transform 1 0 14688 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_154
timestamp 1679581782
transform 1 0 15360 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_161
timestamp 1679581782
transform 1 0 16032 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_168
timestamp 1679581782
transform 1 0 16704 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_175
timestamp 1679581782
transform 1 0 17376 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_182
timestamp 1679581782
transform 1 0 18048 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_189
timestamp 1679581782
transform 1 0 18720 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_196
timestamp 1679581782
transform 1 0 19392 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_203
timestamp 1679581782
transform 1 0 20064 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_210
timestamp 1679581782
transform 1 0 20736 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_217
timestamp 1679581782
transform 1 0 21408 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_224
timestamp 1679581782
transform 1 0 22080 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_231
timestamp 1679581782
transform 1 0 22752 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_238
timestamp 1679581782
transform 1 0 23424 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_245
timestamp 1679581782
transform 1 0 24096 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_252
timestamp 1679581782
transform 1 0 24768 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_259
timestamp 1679581782
transform 1 0 25440 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_266
timestamp 1679581782
transform 1 0 26112 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_273
timestamp 1679581782
transform 1 0 26784 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_280
timestamp 1679581782
transform 1 0 27456 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_287
timestamp 1679581782
transform 1 0 28128 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_294
timestamp 1679581782
transform 1 0 28800 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_301
timestamp 1679581782
transform 1 0 29472 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_308
timestamp 1679581782
transform 1 0 30144 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_315
timestamp 1679581782
transform 1 0 30816 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_322
timestamp 1679581782
transform 1 0 31488 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_329
timestamp 1679581782
transform 1 0 32160 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_336
timestamp 1679581782
transform 1 0 32832 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_343
timestamp 1679581782
transform 1 0 33504 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_350
timestamp 1679581782
transform 1 0 34176 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_357
timestamp 1679581782
transform 1 0 34848 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_364
timestamp 1679581782
transform 1 0 35520 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_371
timestamp 1679581782
transform 1 0 36192 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_378
timestamp 1679581782
transform 1 0 36864 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_385
timestamp 1679581782
transform 1 0 37536 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_392
timestamp 1679581782
transform 1 0 38208 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_399
timestamp 1679581782
transform 1 0 38880 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_406
timestamp 1679581782
transform 1 0 39552 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_413
timestamp 1679581782
transform 1 0 40224 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_420
timestamp 1679581782
transform 1 0 40896 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_427
timestamp 1679581782
transform 1 0 41568 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_434
timestamp 1679581782
transform 1 0 42240 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_441
timestamp 1679581782
transform 1 0 42912 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_448
timestamp 1679581782
transform 1 0 43584 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_455
timestamp 1679581782
transform 1 0 44256 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_462
timestamp 1679581782
transform 1 0 44928 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_469
timestamp 1679581782
transform 1 0 45600 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_476
timestamp 1679581782
transform 1 0 46272 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_483
timestamp 1679581782
transform 1 0 46944 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_490
timestamp 1679581782
transform 1 0 47616 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_497
timestamp 1679581782
transform 1 0 48288 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_504
timestamp 1679581782
transform 1 0 48960 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_511
timestamp 1679581782
transform 1 0 49632 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_518
timestamp 1679581782
transform 1 0 50304 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_525
timestamp 1679581782
transform 1 0 50976 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_532
timestamp 1679581782
transform 1 0 51648 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_539
timestamp 1679581782
transform 1 0 52320 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_546
timestamp 1679581782
transform 1 0 52992 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_553
timestamp 1679581782
transform 1 0 53664 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_560
timestamp 1679581782
transform 1 0 54336 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_567
timestamp 1679581782
transform 1 0 55008 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_574
timestamp 1679581782
transform 1 0 55680 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_581
timestamp 1679581782
transform 1 0 56352 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_588
timestamp 1679581782
transform 1 0 57024 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_595
timestamp 1679581782
transform 1 0 57696 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_602
timestamp 1679581782
transform 1 0 58368 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_609
timestamp 1679581782
transform 1 0 59040 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_616
timestamp 1679581782
transform 1 0 59712 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_623
timestamp 1679581782
transform 1 0 60384 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_630
timestamp 1679581782
transform 1 0 61056 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_637
timestamp 1679581782
transform 1 0 61728 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_644
timestamp 1679581782
transform 1 0 62400 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_651
timestamp 1679581782
transform 1 0 63072 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_658
timestamp 1679581782
transform 1 0 63744 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_665
timestamp 1679581782
transform 1 0 64416 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_672
timestamp 1679581782
transform 1 0 65088 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_679
timestamp 1679581782
transform 1 0 65760 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_686
timestamp 1679581782
transform 1 0 66432 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_693
timestamp 1679581782
transform 1 0 67104 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_700
timestamp 1679581782
transform 1 0 67776 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_707
timestamp 1679581782
transform 1 0 68448 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_714
timestamp 1679581782
transform 1 0 69120 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_721
timestamp 1679581782
transform 1 0 69792 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_728
timestamp 1679581782
transform 1 0 70464 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_735
timestamp 1679581782
transform 1 0 71136 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_742
timestamp 1679581782
transform 1 0 71808 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_749
timestamp 1679581782
transform 1 0 72480 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_756
timestamp 1679581782
transform 1 0 73152 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_763
timestamp 1679581782
transform 1 0 73824 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_770
timestamp 1679581782
transform 1 0 74496 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_777
timestamp 1679581782
transform 1 0 75168 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_784
timestamp 1679581782
transform 1 0 75840 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_791
timestamp 1679581782
transform 1 0 76512 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_798
timestamp 1679581782
transform 1 0 77184 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_805
timestamp 1679581782
transform 1 0 77856 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_812
timestamp 1679581782
transform 1 0 78528 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_819
timestamp 1679581782
transform 1 0 79200 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_826
timestamp 1679581782
transform 1 0 79872 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_833
timestamp 1679581782
transform 1 0 80544 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_840
timestamp 1679581782
transform 1 0 81216 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_847
timestamp 1679581782
transform 1 0 81888 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_854
timestamp 1679581782
transform 1 0 82560 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_861
timestamp 1679581782
transform 1 0 83232 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_868
timestamp 1679581782
transform 1 0 83904 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_875
timestamp 1679581782
transform 1 0 84576 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_882
timestamp 1679581782
transform 1 0 85248 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_889
timestamp 1679581782
transform 1 0 85920 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_896
timestamp 1679581782
transform 1 0 86592 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_903
timestamp 1679581782
transform 1 0 87264 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_910
timestamp 1679581782
transform 1 0 87936 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_917
timestamp 1679581782
transform 1 0 88608 0 -1 38556
box -48 -56 720 834
use sg13g2_fill_1  FILLER_49_924
timestamp 1677579658
transform 1 0 89280 0 -1 38556
box -48 -56 144 834
use sg13g2_tielo  heichips25_example_small_25
timestamp 1680000637
transform -1 0 960 0 1 15876
box -48 -56 432 834
use sg13g2_tielo  heichips25_example_small_26
timestamp 1680000637
transform -1 0 960 0 -1 17388
box -48 -56 432 834
use sg13g2_tielo  heichips25_example_small_27
timestamp 1680000637
transform -1 0 960 0 1 17388
box -48 -56 432 834
use sg13g2_tielo  heichips25_example_small_28
timestamp 1680000637
transform -1 0 960 0 -1 18900
box -48 -56 432 834
use sg13g2_tielo  heichips25_example_small_29
timestamp 1680000637
transform -1 0 960 0 1 18900
box -48 -56 432 834
use sg13g2_tielo  heichips25_example_small_30
timestamp 1680000637
transform -1 0 960 0 -1 20412
box -48 -56 432 834
use sg13g2_tielo  heichips25_example_small_31
timestamp 1680000637
transform -1 0 960 0 1 20412
box -48 -56 432 834
use sg13g2_tielo  heichips25_example_small_32
timestamp 1680000637
transform -1 0 960 0 1 21924
box -48 -56 432 834
use sg13g2_tielo  heichips25_example_small_33
timestamp 1680000637
transform -1 0 960 0 -1 9828
box -48 -56 432 834
use sg13g2_tielo  heichips25_example_small_34
timestamp 1680000637
transform -1 0 960 0 1 9828
box -48 -56 432 834
use sg13g2_tielo  heichips25_example_small_35
timestamp 1680000637
transform -1 0 960 0 -1 11340
box -48 -56 432 834
use sg13g2_tielo  heichips25_example_small_36
timestamp 1680000637
transform -1 0 960 0 1 11340
box -48 -56 432 834
use sg13g2_tielo  heichips25_example_small_37
timestamp 1680000637
transform -1 0 960 0 -1 12852
box -48 -56 432 834
use sg13g2_tielo  heichips25_example_small_38
timestamp 1680000637
transform -1 0 960 0 1 12852
box -48 -56 432 834
use sg13g2_tielo  heichips25_example_small_39
timestamp 1680000637
transform -1 0 960 0 1 14364
box -48 -56 432 834
use sg13g2_tielo  heichips25_example_small_40
timestamp 1680000637
transform -1 0 960 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  input1
timestamp 1676381911
transform 1 0 576 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  input2
timestamp 1676381911
transform 1 0 576 0 1 23436
box -48 -56 432 834
use sg13g2_buf_1  input3
timestamp 1676381911
transform 1 0 576 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  input4
timestamp 1676381911
transform 1 0 576 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  input5
timestamp 1676381911
transform 1 0 576 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  input6
timestamp 1676381911
transform 1 0 576 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  input7
timestamp 1676381911
transform 1 0 576 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_1  input8
timestamp 1676381911
transform 1 0 576 0 1 27972
box -48 -56 432 834
use sg13g2_buf_1  input9
timestamp 1676381911
transform 1 0 576 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  input10
timestamp 1676381911
transform 1 0 576 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  input11
timestamp 1676381911
transform 1 0 576 0 1 30996
box -48 -56 432 834
use sg13g2_buf_1  input12
timestamp 1676381911
transform 1 0 576 0 -1 32508
box -48 -56 432 834
use sg13g2_buf_1  input13
timestamp 1676381911
transform 1 0 576 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  input14
timestamp 1676381911
transform 1 0 576 0 -1 34020
box -48 -56 432 834
use sg13g2_buf_1  input15
timestamp 1676381911
transform 1 0 576 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  input16
timestamp 1676381911
transform 1 0 576 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  output17
timestamp 1676381911
transform -1 0 960 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  output18
timestamp 1676381911
transform -1 0 960 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  output19
timestamp 1676381911
transform -1 0 960 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  output20
timestamp 1676381911
transform -1 0 960 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  output21
timestamp 1676381911
transform -1 0 960 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  output22
timestamp 1676381911
transform -1 0 960 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  output23
timestamp 1676381911
transform -1 0 960 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  output24
timestamp 1676381911
transform -1 0 960 0 1 8316
box -48 -56 432 834
<< labels >>
flabel metal6 s 4316 630 4756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 19436 630 19876 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 34556 630 34996 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 49676 630 50116 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 64796 630 65236 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 79916 630 80356 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 3076 712 3516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 18196 712 18636 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 33316 712 33756 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 48436 712 48876 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 63556 712 63996 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 78676 712 79116 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 36668 80 36748 0 FreeSans 320 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 0 35828 80 35908 0 FreeSans 320 0 0 0 ena
port 3 nsew signal input
flabel metal3 s 0 37508 80 37588 0 FreeSans 320 0 0 0 rst_n
port 4 nsew signal input
flabel metal3 s 0 22388 80 22468 0 FreeSans 320 0 0 0 ui_in[0]
port 5 nsew signal input
flabel metal3 s 0 23228 80 23308 0 FreeSans 320 0 0 0 ui_in[1]
port 6 nsew signal input
flabel metal3 s 0 24068 80 24148 0 FreeSans 320 0 0 0 ui_in[2]
port 7 nsew signal input
flabel metal3 s 0 24908 80 24988 0 FreeSans 320 0 0 0 ui_in[3]
port 8 nsew signal input
flabel metal3 s 0 25748 80 25828 0 FreeSans 320 0 0 0 ui_in[4]
port 9 nsew signal input
flabel metal3 s 0 26588 80 26668 0 FreeSans 320 0 0 0 ui_in[5]
port 10 nsew signal input
flabel metal3 s 0 27428 80 27508 0 FreeSans 320 0 0 0 ui_in[6]
port 11 nsew signal input
flabel metal3 s 0 28268 80 28348 0 FreeSans 320 0 0 0 ui_in[7]
port 12 nsew signal input
flabel metal3 s 0 29108 80 29188 0 FreeSans 320 0 0 0 uio_in[0]
port 13 nsew signal input
flabel metal3 s 0 29948 80 30028 0 FreeSans 320 0 0 0 uio_in[1]
port 14 nsew signal input
flabel metal3 s 0 30788 80 30868 0 FreeSans 320 0 0 0 uio_in[2]
port 15 nsew signal input
flabel metal3 s 0 31628 80 31708 0 FreeSans 320 0 0 0 uio_in[3]
port 16 nsew signal input
flabel metal3 s 0 32468 80 32548 0 FreeSans 320 0 0 0 uio_in[4]
port 17 nsew signal input
flabel metal3 s 0 33308 80 33388 0 FreeSans 320 0 0 0 uio_in[5]
port 18 nsew signal input
flabel metal3 s 0 34148 80 34228 0 FreeSans 320 0 0 0 uio_in[6]
port 19 nsew signal input
flabel metal3 s 0 34988 80 35068 0 FreeSans 320 0 0 0 uio_in[7]
port 20 nsew signal input
flabel metal3 s 0 15668 80 15748 0 FreeSans 320 0 0 0 uio_oe[0]
port 21 nsew signal output
flabel metal3 s 0 16508 80 16588 0 FreeSans 320 0 0 0 uio_oe[1]
port 22 nsew signal output
flabel metal3 s 0 17348 80 17428 0 FreeSans 320 0 0 0 uio_oe[2]
port 23 nsew signal output
flabel metal3 s 0 18188 80 18268 0 FreeSans 320 0 0 0 uio_oe[3]
port 24 nsew signal output
flabel metal3 s 0 19028 80 19108 0 FreeSans 320 0 0 0 uio_oe[4]
port 25 nsew signal output
flabel metal3 s 0 19868 80 19948 0 FreeSans 320 0 0 0 uio_oe[5]
port 26 nsew signal output
flabel metal3 s 0 20708 80 20788 0 FreeSans 320 0 0 0 uio_oe[6]
port 27 nsew signal output
flabel metal3 s 0 21548 80 21628 0 FreeSans 320 0 0 0 uio_oe[7]
port 28 nsew signal output
flabel metal3 s 0 8948 80 9028 0 FreeSans 320 0 0 0 uio_out[0]
port 29 nsew signal output
flabel metal3 s 0 9788 80 9868 0 FreeSans 320 0 0 0 uio_out[1]
port 30 nsew signal output
flabel metal3 s 0 10628 80 10708 0 FreeSans 320 0 0 0 uio_out[2]
port 31 nsew signal output
flabel metal3 s 0 11468 80 11548 0 FreeSans 320 0 0 0 uio_out[3]
port 32 nsew signal output
flabel metal3 s 0 12308 80 12388 0 FreeSans 320 0 0 0 uio_out[4]
port 33 nsew signal output
flabel metal3 s 0 13148 80 13228 0 FreeSans 320 0 0 0 uio_out[5]
port 34 nsew signal output
flabel metal3 s 0 13988 80 14068 0 FreeSans 320 0 0 0 uio_out[6]
port 35 nsew signal output
flabel metal3 s 0 14828 80 14908 0 FreeSans 320 0 0 0 uio_out[7]
port 36 nsew signal output
flabel metal3 s 0 2228 80 2308 0 FreeSans 320 0 0 0 uo_out[0]
port 37 nsew signal output
flabel metal3 s 0 3068 80 3148 0 FreeSans 320 0 0 0 uo_out[1]
port 38 nsew signal output
flabel metal3 s 0 3908 80 3988 0 FreeSans 320 0 0 0 uo_out[2]
port 39 nsew signal output
flabel metal3 s 0 4748 80 4828 0 FreeSans 320 0 0 0 uo_out[3]
port 40 nsew signal output
flabel metal3 s 0 5588 80 5668 0 FreeSans 320 0 0 0 uo_out[4]
port 41 nsew signal output
flabel metal3 s 0 6428 80 6508 0 FreeSans 320 0 0 0 uo_out[5]
port 42 nsew signal output
flabel metal3 s 0 7268 80 7348 0 FreeSans 320 0 0 0 uo_out[6]
port 43 nsew signal output
flabel metal3 s 0 8108 80 8188 0 FreeSans 320 0 0 0 uo_out[7]
port 44 nsew signal output
rlabel metal1 44976 38556 44976 38556 0 VGND
rlabel metal1 44976 37800 44976 37800 0 VPWR
rlabel metal2 8544 20706 8544 20706 0 _00_
rlabel metal2 8304 19488 8304 19488 0 _01_
rlabel via2 8352 20244 8352 20244 0 _02_
rlabel metal3 10224 22260 10224 22260 0 _03_
rlabel metal2 12048 23268 12048 23268 0 _04_
rlabel metal2 11328 22302 11328 22302 0 _05_
rlabel metal3 11808 24024 11808 24024 0 _06_
rlabel metal2 11424 26376 11424 26376 0 _07_
rlabel metal2 11136 26754 11136 26754 0 _08_
rlabel metal2 12672 25326 12672 25326 0 _09_
rlabel metal2 12096 25032 12096 25032 0 _10_
rlabel metal3 10416 24780 10416 24780 0 _11_
rlabel metal2 9888 25242 9888 25242 0 _12_
rlabel metal2 4128 23856 4128 23856 0 _13_
rlabel metal2 4320 24318 4320 24318 0 _14_
rlabel metal2 4320 23730 4320 23730 0 _15_
rlabel metal2 5376 25410 5376 25410 0 _16_
rlabel metal2 4176 24024 4176 24024 0 _17_
rlabel metal2 3648 26376 3648 26376 0 _18_
rlabel metal2 5184 26376 5184 26376 0 _19_
rlabel metal3 4848 24612 4848 24612 0 _20_
rlabel metal2 5280 26544 5280 26544 0 _21_
rlabel metal2 3696 25956 3696 25956 0 _22_
rlabel metal3 3600 29820 3600 29820 0 _23_
rlabel metal2 3744 30576 3744 30576 0 _24_
rlabel metal2 3648 30534 3648 30534 0 _25_
rlabel metal2 2784 29778 2784 29778 0 _26_
rlabel metal2 3840 31500 3840 31500 0 _27_
rlabel metal2 4704 32676 4704 32676 0 _28_
rlabel metal3 2352 20748 2352 20748 0 net1
rlabel metal2 864 30156 864 30156 0 net10
rlabel metal2 1056 28308 1056 28308 0 net11
rlabel metal2 576 29442 576 29442 0 net12
rlabel metal2 1824 23814 1824 23814 0 net13
rlabel metal2 624 33096 624 33096 0 net14
rlabel metal2 960 34188 960 34188 0 net15
rlabel metal2 4416 33222 4416 33222 0 net16
rlabel metal2 1056 2688 1056 2688 0 net17
rlabel metal2 816 3360 816 3360 0 net18
rlabel metal2 960 4200 960 4200 0 net19
rlabel metal2 912 23604 912 23604 0 net2
rlabel metal2 912 4872 912 4872 0 net20
rlabel metal3 3648 5712 3648 5712 0 net21
rlabel metal3 1008 7224 1008 7224 0 net22
rlabel metal3 1488 7896 1488 7896 0 net23
rlabel metal2 480 26712 480 26712 0 net24
rlabel metal3 318 15708 318 15708 0 net25
rlabel metal3 366 16548 366 16548 0 net26
rlabel metal3 366 17388 366 17388 0 net27
rlabel metal3 366 18228 366 18228 0 net28
rlabel metal3 366 19068 366 19068 0 net29
rlabel metal2 12384 22764 12384 22764 0 net3
rlabel metal3 366 19908 366 19908 0 net30
rlabel metal3 366 20748 366 20748 0 net31
rlabel metal3 366 21588 366 21588 0 net32
rlabel metal3 366 8988 366 8988 0 net33
rlabel metal3 366 9828 366 9828 0 net34
rlabel metal3 366 10668 366 10668 0 net35
rlabel metal3 366 11508 366 11508 0 net36
rlabel metal3 366 12348 366 12348 0 net37
rlabel metal3 366 13188 366 13188 0 net38
rlabel metal3 366 14028 366 14028 0 net39
rlabel metal3 1008 25536 1008 25536 0 net4
rlabel metal3 366 14868 366 14868 0 net40
rlabel metal3 1392 23772 1392 23772 0 net5
rlabel metal3 2160 26796 2160 26796 0 net6
rlabel metal2 2304 29568 2304 29568 0 net7
rlabel metal2 4320 32802 4320 32802 0 net8
rlabel metal2 3456 20790 3456 20790 0 net9
rlabel metal3 366 22428 366 22428 0 ui_in[0]
rlabel metal3 366 23268 366 23268 0 ui_in[1]
rlabel metal3 366 24108 366 24108 0 ui_in[2]
rlabel metal3 366 24948 366 24948 0 ui_in[3]
rlabel metal3 366 25788 366 25788 0 ui_in[4]
rlabel metal3 366 26628 366 26628 0 ui_in[5]
rlabel metal3 366 27468 366 27468 0 ui_in[6]
rlabel metal3 366 28308 366 28308 0 ui_in[7]
rlabel metal3 366 29148 366 29148 0 uio_in[0]
rlabel metal3 366 29988 366 29988 0 uio_in[1]
rlabel metal3 366 30828 366 30828 0 uio_in[2]
rlabel metal3 366 31668 366 31668 0 uio_in[3]
rlabel metal3 366 32508 366 32508 0 uio_in[4]
rlabel metal3 366 33348 366 33348 0 uio_in[5]
rlabel metal3 366 34188 366 34188 0 uio_in[6]
rlabel metal3 366 35028 366 35028 0 uio_in[7]
rlabel metal3 366 2268 366 2268 0 uo_out[0]
rlabel metal3 366 3108 366 3108 0 uo_out[1]
rlabel metal3 366 3948 366 3948 0 uo_out[2]
rlabel metal3 366 4788 366 4788 0 uo_out[3]
rlabel metal3 366 5628 366 5628 0 uo_out[4]
rlabel metal3 366 6468 366 6468 0 uo_out[5]
rlabel metal3 366 7308 366 7308 0 uo_out[6]
rlabel metal3 366 8148 366 8148 0 uo_out[7]
<< properties >>
string FIXED_BBOX 0 0 90000 40000
<< end >>
