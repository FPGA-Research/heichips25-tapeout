module IHP_SRAM (ADDR_SRAM0,
    ADDR_SRAM1,
    ADDR_SRAM2,
    ADDR_SRAM3,
    ADDR_SRAM4,
    ADDR_SRAM5,
    ADDR_SRAM6,
    ADDR_SRAM7,
    ADDR_SRAM8,
    ADDR_SRAM9,
    BM_SRAM0,
    BM_SRAM1,
    BM_SRAM10,
    BM_SRAM11,
    BM_SRAM12,
    BM_SRAM13,
    BM_SRAM14,
    BM_SRAM15,
    BM_SRAM16,
    BM_SRAM17,
    BM_SRAM18,
    BM_SRAM19,
    BM_SRAM2,
    BM_SRAM20,
    BM_SRAM21,
    BM_SRAM22,
    BM_SRAM23,
    BM_SRAM24,
    BM_SRAM25,
    BM_SRAM26,
    BM_SRAM27,
    BM_SRAM28,
    BM_SRAM29,
    BM_SRAM3,
    BM_SRAM30,
    BM_SRAM31,
    BM_SRAM4,
    BM_SRAM5,
    BM_SRAM6,
    BM_SRAM7,
    BM_SRAM8,
    BM_SRAM9,
    CLK_SRAM,
    CONFIGURED_top,
    DIN_SRAM0,
    DIN_SRAM1,
    DIN_SRAM10,
    DIN_SRAM11,
    DIN_SRAM12,
    DIN_SRAM13,
    DIN_SRAM14,
    DIN_SRAM15,
    DIN_SRAM16,
    DIN_SRAM17,
    DIN_SRAM18,
    DIN_SRAM19,
    DIN_SRAM2,
    DIN_SRAM20,
    DIN_SRAM21,
    DIN_SRAM22,
    DIN_SRAM23,
    DIN_SRAM24,
    DIN_SRAM25,
    DIN_SRAM26,
    DIN_SRAM27,
    DIN_SRAM28,
    DIN_SRAM29,
    DIN_SRAM3,
    DIN_SRAM30,
    DIN_SRAM31,
    DIN_SRAM4,
    DIN_SRAM5,
    DIN_SRAM6,
    DIN_SRAM7,
    DIN_SRAM8,
    DIN_SRAM9,
    DOUT_SRAM0,
    DOUT_SRAM1,
    DOUT_SRAM10,
    DOUT_SRAM11,
    DOUT_SRAM12,
    DOUT_SRAM13,
    DOUT_SRAM14,
    DOUT_SRAM15,
    DOUT_SRAM16,
    DOUT_SRAM17,
    DOUT_SRAM18,
    DOUT_SRAM19,
    DOUT_SRAM2,
    DOUT_SRAM20,
    DOUT_SRAM21,
    DOUT_SRAM22,
    DOUT_SRAM23,
    DOUT_SRAM24,
    DOUT_SRAM25,
    DOUT_SRAM26,
    DOUT_SRAM27,
    DOUT_SRAM28,
    DOUT_SRAM29,
    DOUT_SRAM3,
    DOUT_SRAM30,
    DOUT_SRAM31,
    DOUT_SRAM4,
    DOUT_SRAM5,
    DOUT_SRAM6,
    DOUT_SRAM7,
    DOUT_SRAM8,
    DOUT_SRAM9,
    MEN_SRAM,
    REN_SRAM,
    TIE_HIGH_SRAM,
    TIE_LOW_SRAM,
    Tile_X0Y0_UserCLKo,
    Tile_X0Y1_UserCLK,
    WEN_SRAM,
    Tile_X0Y0_E1END,
    Tile_X0Y0_E2END,
    Tile_X0Y0_E2MID,
    Tile_X0Y0_E6END,
    Tile_X0Y0_EE4END,
    Tile_X0Y0_FrameData,
    Tile_X0Y0_FrameData_O,
    Tile_X0Y0_FrameStrobe_O,
    Tile_X0Y0_N1BEG,
    Tile_X0Y0_N2BEG,
    Tile_X0Y0_N2BEGb,
    Tile_X0Y0_N4BEG,
    Tile_X0Y0_S1END,
    Tile_X0Y0_S2END,
    Tile_X0Y0_S2MID,
    Tile_X0Y0_S4END,
    Tile_X0Y0_W1BEG,
    Tile_X0Y0_W2BEG,
    Tile_X0Y0_W2BEGb,
    Tile_X0Y0_W6BEG,
    Tile_X0Y0_WW4BEG,
    Tile_X0Y1_E1END,
    Tile_X0Y1_E2END,
    Tile_X0Y1_E2MID,
    Tile_X0Y1_E6END,
    Tile_X0Y1_EE4END,
    Tile_X0Y1_FrameData,
    Tile_X0Y1_FrameData_O,
    Tile_X0Y1_FrameStrobe,
    Tile_X0Y1_N1END,
    Tile_X0Y1_N2END,
    Tile_X0Y1_N2MID,
    Tile_X0Y1_N4END,
    Tile_X0Y1_S1BEG,
    Tile_X0Y1_S2BEG,
    Tile_X0Y1_S2BEGb,
    Tile_X0Y1_S4BEG,
    Tile_X0Y1_W1BEG,
    Tile_X0Y1_W2BEG,
    Tile_X0Y1_W2BEGb,
    Tile_X0Y1_W6BEG,
    Tile_X0Y1_WW4BEG);
 output ADDR_SRAM0;
 output ADDR_SRAM1;
 output ADDR_SRAM2;
 output ADDR_SRAM3;
 output ADDR_SRAM4;
 output ADDR_SRAM5;
 output ADDR_SRAM6;
 output ADDR_SRAM7;
 output ADDR_SRAM8;
 output ADDR_SRAM9;
 output BM_SRAM0;
 output BM_SRAM1;
 output BM_SRAM10;
 output BM_SRAM11;
 output BM_SRAM12;
 output BM_SRAM13;
 output BM_SRAM14;
 output BM_SRAM15;
 output BM_SRAM16;
 output BM_SRAM17;
 output BM_SRAM18;
 output BM_SRAM19;
 output BM_SRAM2;
 output BM_SRAM20;
 output BM_SRAM21;
 output BM_SRAM22;
 output BM_SRAM23;
 output BM_SRAM24;
 output BM_SRAM25;
 output BM_SRAM26;
 output BM_SRAM27;
 output BM_SRAM28;
 output BM_SRAM29;
 output BM_SRAM3;
 output BM_SRAM30;
 output BM_SRAM31;
 output BM_SRAM4;
 output BM_SRAM5;
 output BM_SRAM6;
 output BM_SRAM7;
 output BM_SRAM8;
 output BM_SRAM9;
 output CLK_SRAM;
 input CONFIGURED_top;
 output DIN_SRAM0;
 output DIN_SRAM1;
 output DIN_SRAM10;
 output DIN_SRAM11;
 output DIN_SRAM12;
 output DIN_SRAM13;
 output DIN_SRAM14;
 output DIN_SRAM15;
 output DIN_SRAM16;
 output DIN_SRAM17;
 output DIN_SRAM18;
 output DIN_SRAM19;
 output DIN_SRAM2;
 output DIN_SRAM20;
 output DIN_SRAM21;
 output DIN_SRAM22;
 output DIN_SRAM23;
 output DIN_SRAM24;
 output DIN_SRAM25;
 output DIN_SRAM26;
 output DIN_SRAM27;
 output DIN_SRAM28;
 output DIN_SRAM29;
 output DIN_SRAM3;
 output DIN_SRAM30;
 output DIN_SRAM31;
 output DIN_SRAM4;
 output DIN_SRAM5;
 output DIN_SRAM6;
 output DIN_SRAM7;
 output DIN_SRAM8;
 output DIN_SRAM9;
 input DOUT_SRAM0;
 input DOUT_SRAM1;
 input DOUT_SRAM10;
 input DOUT_SRAM11;
 input DOUT_SRAM12;
 input DOUT_SRAM13;
 input DOUT_SRAM14;
 input DOUT_SRAM15;
 input DOUT_SRAM16;
 input DOUT_SRAM17;
 input DOUT_SRAM18;
 input DOUT_SRAM19;
 input DOUT_SRAM2;
 input DOUT_SRAM20;
 input DOUT_SRAM21;
 input DOUT_SRAM22;
 input DOUT_SRAM23;
 input DOUT_SRAM24;
 input DOUT_SRAM25;
 input DOUT_SRAM26;
 input DOUT_SRAM27;
 input DOUT_SRAM28;
 input DOUT_SRAM29;
 input DOUT_SRAM3;
 input DOUT_SRAM30;
 input DOUT_SRAM31;
 input DOUT_SRAM4;
 input DOUT_SRAM5;
 input DOUT_SRAM6;
 input DOUT_SRAM7;
 input DOUT_SRAM8;
 input DOUT_SRAM9;
 output MEN_SRAM;
 output REN_SRAM;
 output TIE_HIGH_SRAM;
 output TIE_LOW_SRAM;
 output Tile_X0Y0_UserCLKo;
 input Tile_X0Y1_UserCLK;
 output WEN_SRAM;
 input [3:0] Tile_X0Y0_E1END;
 input [7:0] Tile_X0Y0_E2END;
 input [7:0] Tile_X0Y0_E2MID;
 input [11:0] Tile_X0Y0_E6END;
 input [15:0] Tile_X0Y0_EE4END;
 input [31:0] Tile_X0Y0_FrameData;
 output [31:0] Tile_X0Y0_FrameData_O;
 output [19:0] Tile_X0Y0_FrameStrobe_O;
 output [3:0] Tile_X0Y0_N1BEG;
 output [7:0] Tile_X0Y0_N2BEG;
 output [7:0] Tile_X0Y0_N2BEGb;
 output [15:0] Tile_X0Y0_N4BEG;
 input [3:0] Tile_X0Y0_S1END;
 input [7:0] Tile_X0Y0_S2END;
 input [7:0] Tile_X0Y0_S2MID;
 input [15:0] Tile_X0Y0_S4END;
 output [3:0] Tile_X0Y0_W1BEG;
 output [7:0] Tile_X0Y0_W2BEG;
 output [7:0] Tile_X0Y0_W2BEGb;
 output [11:0] Tile_X0Y0_W6BEG;
 output [15:0] Tile_X0Y0_WW4BEG;
 input [3:0] Tile_X0Y1_E1END;
 input [7:0] Tile_X0Y1_E2END;
 input [7:0] Tile_X0Y1_E2MID;
 input [11:0] Tile_X0Y1_E6END;
 input [15:0] Tile_X0Y1_EE4END;
 input [31:0] Tile_X0Y1_FrameData;
 output [31:0] Tile_X0Y1_FrameData_O;
 input [19:0] Tile_X0Y1_FrameStrobe;
 input [3:0] Tile_X0Y1_N1END;
 input [7:0] Tile_X0Y1_N2END;
 input [7:0] Tile_X0Y1_N2MID;
 input [15:0] Tile_X0Y1_N4END;
 output [3:0] Tile_X0Y1_S1BEG;
 output [7:0] Tile_X0Y1_S2BEG;
 output [7:0] Tile_X0Y1_S2BEGb;
 output [15:0] Tile_X0Y1_S4BEG;
 output [3:0] Tile_X0Y1_W1BEG;
 output [7:0] Tile_X0Y1_W2BEG;
 output [7:0] Tile_X0Y1_W2BEGb;
 output [11:0] Tile_X0Y1_W6BEG;
 output [15:0] Tile_X0Y1_WW4BEG;

 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit0.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit1.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit10.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit11.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit12.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit13.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit14.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit15.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit16.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit17.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit2.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit3.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit4.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit5.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit6.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit7.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit8.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit9.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit0.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit1.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit10.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit11.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit12.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit13.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit14.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit15.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit16.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit17.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit18.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit19.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit2.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit20.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit21.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit22.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit23.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit24.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit25.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit26.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit27.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit28.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit29.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit3.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit30.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit31.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit4.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit5.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit6.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit7.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit8.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit9.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit0.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit1.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit10.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit11.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit12.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit13.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit14.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit15.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit16.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit17.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit18.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit19.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit2.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit20.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit21.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit22.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit23.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit24.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit25.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit26.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit27.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit28.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit29.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit3.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit30.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit31.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit4.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit5.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit6.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit7.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit8.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit9.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit0.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit1.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit10.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit11.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit12.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit13.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit14.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit15.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit16.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit17.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit18.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit19.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit2.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit20.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit21.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit22.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit23.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit24.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit25.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit26.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit27.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit28.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit29.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit3.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit30.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit31.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit4.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit5.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit6.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit7.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit8.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit9.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit0.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit1.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit10.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit11.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit12.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit13.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit14.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit15.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit16.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit17.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit18.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit19.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit2.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit20.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit21.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit22.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit23.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit24.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit25.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit26.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit27.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit28.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit29.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit3.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit30.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit31.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit4.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit5.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit6.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit7.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit8.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit9.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit0.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit1.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit10.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit11.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit12.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit13.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit14.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit15.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit16.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit17.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit18.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit19.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit2.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit20.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit21.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit22.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit23.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit24.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit25.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit26.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit27.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit28.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit29.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit3.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit30.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit31.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit4.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit5.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit6.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit7.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit8.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit9.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit22.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit23.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit24.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit25.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit26.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit27.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit28.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit29.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit30.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit31.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG4 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG5 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG6 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG7 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG0 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG1 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG2 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG3 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG0 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG1 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG2 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG3 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END0 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END1 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END2 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END3 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG0 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG1 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG2 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG3 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG4 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG5 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG6 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG7 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb0 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb1 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb2 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb3 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb4 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb5 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb6 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb7 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG0 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG1 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG2 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG3 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG0 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG1 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG2 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG3 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG4 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG5 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG6 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG7 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG0 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG1 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG2 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG3 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG0 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG1 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG2 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG3 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG0 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG1 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG2 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG3 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG4 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG5 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG6 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG7 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb0 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb1 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb2 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb3 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb4 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb5 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb6 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb7 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG0 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG1 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG10 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG11 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG2 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG3 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG4 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG5 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG6 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG7 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG8 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG9 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG0 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG1 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG10 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG11 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG12 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG13 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG14 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG15 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG2 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG3 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG4 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG5 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG6 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG7 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG8 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG9 ;
 wire \Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_10.A ;
 wire \Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_11.A ;
 wire \Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_8.A ;
 wire \Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_9.A ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit0.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit1.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit10.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit11.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit12.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit13.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit14.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit15.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit16.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit17.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit2.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit3.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit4.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit5.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit6.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit7.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit8.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit9.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit0.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit1.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit10.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit11.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit12.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit13.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit14.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit15.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit16.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit17.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit18.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit19.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit2.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit20.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit21.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit22.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit23.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit24.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit25.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit26.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit27.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit28.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit29.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit3.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit30.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit31.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit4.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit5.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit6.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit7.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit8.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit9.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit0.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit1.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit10.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit11.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit12.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit13.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit14.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit15.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit16.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit17.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit18.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit19.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit2.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit20.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit21.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit22.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit23.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit24.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit25.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit26.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit27.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit28.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit29.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit3.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit30.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit31.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit4.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit5.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit6.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit7.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit8.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit9.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit0.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit1.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit10.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit11.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit12.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit13.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit14.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit15.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit16.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit17.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit18.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit19.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit2.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit20.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit21.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit22.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit23.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit24.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit25.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit26.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit27.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit28.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit29.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit3.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit30.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit31.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit4.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit5.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit6.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit7.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit8.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit9.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit0.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit1.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit11.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit14.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit17.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit18.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit19.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit2.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit20.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit21.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit22.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit23.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit24.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit25.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit26.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit27.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit28.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit29.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit3.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit30.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit31.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit4.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit5.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit7.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit8.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit0.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit1.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit10.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit12.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit13.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit14.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit15.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit16.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit17.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit18.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit19.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit2.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit20.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit21.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit22.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit23.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit24.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit25.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit26.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit27.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit28.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit29.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit3.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit30.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit31.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit4.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit5.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit6.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit7.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit9.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit10.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit11.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit12.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit13.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit14.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit15.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit16.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit17.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit18.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit19.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit20.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit21.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit22.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit23.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit24.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit25.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit26.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit27.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit28.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit29.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit30.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit31.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG0 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG1 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG2 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG3 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG0 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG1 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG2 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG3 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG4 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG5 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG6 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG7 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG0 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG1 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG2 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG3 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG0 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG1 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG2 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG3 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG0 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG1 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG2 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG3 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG4 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG5 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG6 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG7 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb0 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb1 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb2 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb3 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb4 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb5 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb6 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb7 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG0 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG1 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG10 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG11 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG2 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG3 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG4 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG5 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG6 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG7 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG8 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG9 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG0 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG1 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG10 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG11 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG12 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG13 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG14 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG15 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG2 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG3 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG4 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG5 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG6 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG7 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG8 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG9 ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire clknet_0_Tile_X0Y1_UserCLK;
 wire clknet_1_0__leaf_Tile_X0Y1_UserCLK;
 wire clknet_1_1__leaf_Tile_X0Y1_UserCLK;

 sg13g2_inv_1 _0297_ (.Y(_0000_),
    .A(Tile_X0Y1_E2MID[3]));
 sg13g2_inv_1 _0298_ (.Y(_0001_),
    .A(Tile_X0Y1_E2END[5]));
 sg13g2_inv_1 _0299_ (.Y(_0002_),
    .A(Tile_X0Y0_S2MID[2]));
 sg13g2_inv_1 _0300_ (.Y(_0003_),
    .A(Tile_X0Y0_E6END[1]));
 sg13g2_inv_1 _0301_ (.Y(_0004_),
    .A(Tile_X0Y0_E6END[2]));
 sg13g2_inv_1 _0302_ (.Y(_0005_),
    .A(Tile_X0Y0_E6END[3]));
 sg13g2_inv_1 _0303_ (.Y(_0006_),
    .A(Tile_X0Y0_E6END[0]));
 sg13g2_inv_1 _0304_ (.Y(_0007_),
    .A(Tile_X0Y1_E6END[3]));
 sg13g2_inv_1 _0305_ (.Y(_0008_),
    .A(Tile_X0Y1_E6END[2]));
 sg13g2_inv_1 _0306_ (.Y(_0009_),
    .A(Tile_X0Y1_E6END[1]));
 sg13g2_inv_1 _0307_ (.Y(_0010_),
    .A(Tile_X0Y1_E6END[0]));
 sg13g2_inv_1 _0308_ (.Y(_0011_),
    .A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit15.Q ));
 sg13g2_inv_1 _0309_ (.Y(_0012_),
    .A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit18.Q ));
 sg13g2_inv_1 _0310_ (.Y(_0013_),
    .A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit21.Q ));
 sg13g2_inv_1 _0311_ (.Y(_0014_),
    .A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit24.Q ));
 sg13g2_inv_1 _0312_ (.Y(_0015_),
    .A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit19.Q ));
 sg13g2_inv_1 _0313_ (.Y(_0016_),
    .A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit22.Q ));
 sg13g2_inv_1 _0314_ (.Y(_0017_),
    .A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit25.Q ));
 sg13g2_inv_1 _0315_ (.Y(_0018_),
    .A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit28.Q ));
 sg13g2_inv_1 _0316_ (.Y(_0019_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit2.Q ));
 sg13g2_inv_1 _0317_ (.Y(_0020_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit3.Q ));
 sg13g2_inv_1 _0318_ (.Y(_0021_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit5.Q ));
 sg13g2_inv_1 _0319_ (.Y(_0022_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit6.Q ));
 sg13g2_inv_1 _0320_ (.Y(_0023_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q ));
 sg13g2_inv_1 _0321_ (.Y(_0024_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit9.Q ));
 sg13g2_inv_1 _0322_ (.Y(_0025_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q ));
 sg13g2_inv_1 _0323_ (.Y(_0026_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit12.Q ));
 sg13g2_inv_1 _0324_ (.Y(_0027_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q ));
 sg13g2_inv_1 _0325_ (.Y(_0028_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit7.Q ));
 sg13g2_inv_1 _0326_ (.Y(_0029_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q ));
 sg13g2_inv_1 _0327_ (.Y(_0030_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q ));
 sg13g2_inv_1 _0328_ (.Y(_0031_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q ));
 sg13g2_inv_1 _0329_ (.Y(_0032_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q ));
 sg13g2_inv_1 _0330_ (.Y(_0033_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q ));
 sg13g2_inv_1 _0331_ (.Y(_0034_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q ));
 sg13g2_inv_1 _0332_ (.Y(_0035_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q ));
 sg13g2_inv_1 _0333_ (.Y(_0036_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit31.Q ));
 sg13g2_inv_1 _0334_ (.Y(_0037_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q ));
 sg13g2_inv_1 _0335_ (.Y(_0038_),
    .A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0 ));
 sg13g2_inv_1 _0336_ (.Y(_0039_),
    .A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1 ));
 sg13g2_inv_1 _0337_ (.Y(_0040_),
    .A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2 ));
 sg13g2_inv_1 _0338_ (.Y(_0041_),
    .A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3 ));
 sg13g2_inv_1 _0339_ (.Y(_0042_),
    .A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG4 ));
 sg13g2_mux4_1 _0340_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit2.Q ),
    .A0(Tile_X0Y0_E2MID[7]),
    .A1(Tile_X0Y0_E2END[7]),
    .A2(Tile_X0Y0_E6END[8]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit3.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG0 ));
 sg13g2_mux4_1 _0341_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit8.Q ),
    .A0(Tile_X0Y1_N2MID[0]),
    .A1(Tile_X0Y1_N2END[0]),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG0 ),
    .A3(Tile_X0Y0_S2MID[0]),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit9.Q ),
    .X(_0043_));
 sg13g2_mux4_1 _0342_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit18.Q ),
    .A0(Tile_X0Y1_E2MID[7]),
    .A1(Tile_X0Y1_E2END[7]),
    .A2(Tile_X0Y1_E6END[7]),
    .A3(_0043_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit19.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb0 ));
 sg13g2_mux4_1 _0343_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit9.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb0 ),
    .A1(Tile_X0Y0_S2MID[0]),
    .A2(Tile_X0Y1_N2MID[0]),
    .A3(Tile_X0Y0_S2END[0]),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit8.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0 ));
 sg13g2_o21ai_1 _0344_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .Y(_0044_),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG0 ));
 sg13g2_nor2_1 _0345_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .Y(_0045_));
 sg13g2_a22oi_1 _0346_ (.Y(_0046_),
    .B1(_0045_),
    .B2(Tile_X0Y1_E2END[4]),
    .A2(Tile_X0Y0_S2MID[3]),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q ));
 sg13g2_nand3_1 _0347_ (.B(_0044_),
    .C(_0046_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .Y(_0047_));
 sg13g2_nand2_1 _0348_ (.Y(_0048_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .B(_0002_));
 sg13g2_o21ai_1 _0349_ (.B1(_0048_),
    .Y(_0049_),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .A2(Tile_X0Y1_E2END[3]));
 sg13g2_nand3b_1 _0350_ (.B(Tile_X0Y1_E2END[5]),
    .C(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .Y(_0050_),
    .A_N(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q ));
 sg13g2_o21ai_1 _0351_ (.B1(_0050_),
    .Y(_0051_),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .A2(_0049_));
 sg13g2_o21ai_1 _0352_ (.B1(_0047_),
    .Y(_0052_),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .A2(_0051_));
 sg13g2_mux4_1 _0353_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .A0(Tile_X0Y1_E2MID[3]),
    .A1(Tile_X0Y1_E2MID[6]),
    .A2(Tile_X0Y1_E2END[1]),
    .A3(Tile_X0Y1_E2END[2]),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .X(_0053_));
 sg13g2_mux4_1 _0354_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .A0(Tile_X0Y1_N2MID[6]),
    .A1(Tile_X0Y1_N2END[2]),
    .A2(Tile_X0Y1_N2END[3]),
    .A3(Tile_X0Y1_E2MID[0]),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .X(_0054_));
 sg13g2_mux2_1 _0355_ (.A0(_0054_),
    .A1(_0053_),
    .S(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .X(_0055_));
 sg13g2_o21ai_1 _0356_ (.B1(CONFIGURED_top),
    .Y(_0056_),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit3.Q ),
    .A2(_0055_));
 sg13g2_a21oi_1 _0357_ (.A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit3.Q ),
    .A2(_0052_),
    .Y(MEN_SRAM),
    .B1(_0056_));
 sg13g2_nand2b_1 _0358_ (.Y(_0057_),
    .B(Tile_X0Y0_S1END[1]),
    .A_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_nor3_1 _0359_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit26.Q ),
    .B(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit27.Q ),
    .C(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END1 ),
    .Y(_0058_));
 sg13g2_a221oi_1 _0360_ (.B2(_0057_),
    .C1(_0058_),
    .B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit27.Q ),
    .A1(_0003_),
    .Y(_0059_),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_mux4_1 _0361_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit28.Q ),
    .A0(Tile_X0Y0_E1END[1]),
    .A1(Tile_X0Y0_E6END[9]),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13 ),
    .A3(_0059_),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit29.Q ),
    .X(_0060_));
 sg13g2_nand2b_1 _0362_ (.Y(_0061_),
    .B(_0060_),
    .A_N(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_nor3_1 _0363_ (.A(Tile_X0Y1_N1END[1]),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q ),
    .C(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit27.Q ),
    .Y(_0062_));
 sg13g2_a221oi_1 _0364_ (.B2(_0061_),
    .C1(_0062_),
    .B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit27.Q ),
    .A1(_0009_),
    .Y(_0063_),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_mux4_1 _0365_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit13.Q ),
    .A0(Tile_X0Y1_E1END[1]),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13 ),
    .A2(Tile_X0Y1_E6END[5]),
    .A3(_0063_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit12.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END1 ));
 sg13g2_mux4_1 _0366_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit2.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END1 ),
    .A1(Tile_X0Y1_N4END[5]),
    .A2(Tile_X0Y0_S1END[1]),
    .A3(Tile_X0Y0_S4END[1]),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit3.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13 ));
 sg13g2_mux4_1 _0367_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit24.Q ),
    .A0(Tile_X0Y0_E1END[1]),
    .A1(Tile_X0Y0_E6END[5]),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13 ),
    .A3(_0059_),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit25.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG1 ));
 sg13g2_nand2b_1 _0368_ (.Y(_0064_),
    .B(Tile_X0Y0_S1END[2]),
    .A_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit28.Q ));
 sg13g2_nor3_1 _0369_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit28.Q ),
    .B(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit29.Q ),
    .C(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END2 ),
    .Y(_0065_));
 sg13g2_a221oi_1 _0370_ (.B2(_0064_),
    .C1(_0065_),
    .B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit29.Q ),
    .A1(_0004_),
    .Y(_0066_),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit28.Q ));
 sg13g2_mux4_1 _0371_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit30.Q ),
    .A0(Tile_X0Y0_E1END[2]),
    .A1(Tile_X0Y0_E6END[10]),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14 ),
    .A3(_0066_),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit31.Q ),
    .X(_0067_));
 sg13g2_nor3_1 _0372_ (.A(Tile_X0Y1_N1END[2]),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q ),
    .C(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit29.Q ),
    .Y(_0068_));
 sg13g2_nand2b_1 _0373_ (.Y(_0069_),
    .B(_0067_),
    .A_N(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q ));
 sg13g2_a221oi_1 _0374_ (.B2(_0069_),
    .C1(_0068_),
    .B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit29.Q ),
    .A1(_0008_),
    .Y(_0070_),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q ));
 sg13g2_mux4_1 _0375_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit15.Q ),
    .A0(Tile_X0Y1_E1END[2]),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14 ),
    .A2(Tile_X0Y1_E6END[6]),
    .A3(_0070_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit14.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END2 ));
 sg13g2_mux4_1 _0376_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit4.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END2 ),
    .A1(Tile_X0Y1_N4END[6]),
    .A2(Tile_X0Y0_S1END[2]),
    .A3(Tile_X0Y0_S4END[2]),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit5.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14 ));
 sg13g2_mux4_1 _0377_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit26.Q ),
    .A0(Tile_X0Y0_E1END[2]),
    .A1(Tile_X0Y0_E6END[6]),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14 ),
    .A3(_0066_),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit27.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG2 ));
 sg13g2_nand2b_1 _0378_ (.Y(_0071_),
    .B(Tile_X0Y0_S1END[3]),
    .A_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit30.Q ));
 sg13g2_nor3_1 _0379_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit30.Q ),
    .B(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit31.Q ),
    .C(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END3 ),
    .Y(_0072_));
 sg13g2_a221oi_1 _0380_ (.B2(_0071_),
    .C1(_0072_),
    .B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit31.Q ),
    .A1(_0005_),
    .Y(_0073_),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit30.Q ));
 sg13g2_mux4_1 _0381_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit0.Q ),
    .A0(Tile_X0Y0_E1END[3]),
    .A1(Tile_X0Y0_E6END[11]),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15 ),
    .A3(_0073_),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit1.Q ),
    .X(_0074_));
 sg13g2_nor3_1 _0382_ (.A(Tile_X0Y1_N1END[3]),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q ),
    .C(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit31.Q ),
    .Y(_0075_));
 sg13g2_nand2b_1 _0383_ (.Y(_0076_),
    .B(_0074_),
    .A_N(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q ));
 sg13g2_a221oi_1 _0384_ (.B2(_0076_),
    .C1(_0075_),
    .B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit31.Q ),
    .A1(_0007_),
    .Y(_0077_),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q ));
 sg13g2_mux4_1 _0385_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit17.Q ),
    .A0(Tile_X0Y1_E1END[3]),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15 ),
    .A2(Tile_X0Y1_E6END[7]),
    .A3(_0077_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit16.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END3 ));
 sg13g2_mux4_1 _0386_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit6.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END3 ),
    .A1(Tile_X0Y1_N4END[7]),
    .A2(Tile_X0Y0_S1END[3]),
    .A3(Tile_X0Y0_S4END[3]),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit7.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15 ));
 sg13g2_mux4_1 _0387_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit28.Q ),
    .A0(Tile_X0Y0_E1END[3]),
    .A1(Tile_X0Y0_E6END[7]),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15 ),
    .A3(_0073_),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit29.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG3 ));
 sg13g2_mux4_1 _0388_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit30.Q ),
    .A0(Tile_X0Y0_E2MID[7]),
    .A1(Tile_X0Y0_E2END[7]),
    .A2(Tile_X0Y0_E6END[7]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit31.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG0 ));
 sg13g2_mux4_1 _0389_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit4.Q ),
    .A0(Tile_X0Y0_E2MID[6]),
    .A1(Tile_X0Y0_E2END[6]),
    .A2(Tile_X0Y0_E6END[9]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit5.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG1 ));
 sg13g2_mux4_1 _0390_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit10.Q ),
    .A0(Tile_X0Y1_N2MID[1]),
    .A1(Tile_X0Y1_N2END[1]),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG1 ),
    .A3(Tile_X0Y0_S2MID[1]),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit11.Q ),
    .X(_0078_));
 sg13g2_mux4_1 _0391_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit20.Q ),
    .A0(Tile_X0Y1_E2MID[6]),
    .A1(Tile_X0Y1_E2END[6]),
    .A2(Tile_X0Y1_E6END[6]),
    .A3(_0078_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit21.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb1 ));
 sg13g2_mux4_1 _0392_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit11.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb1 ),
    .A1(Tile_X0Y0_S2MID[1]),
    .A2(Tile_X0Y1_N2MID[1]),
    .A3(Tile_X0Y0_S2END[1]),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit10.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1 ));
 sg13g2_mux4_1 _0393_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit0.Q ),
    .A0(Tile_X0Y0_E2MID[6]),
    .A1(Tile_X0Y0_E2END[6]),
    .A2(Tile_X0Y0_E6END[6]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit1.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG1 ));
 sg13g2_mux4_1 _0394_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit6.Q ),
    .A0(Tile_X0Y0_E2MID[5]),
    .A1(Tile_X0Y0_E2END[5]),
    .A2(Tile_X0Y0_E6END[10]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit7.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG2 ));
 sg13g2_mux4_1 _0395_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit13.Q ),
    .A0(Tile_X0Y1_N2MID[2]),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG2 ),
    .A2(Tile_X0Y1_N2END[2]),
    .A3(Tile_X0Y0_S2MID[2]),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit12.Q ),
    .X(_0079_));
 sg13g2_mux4_1 _0396_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit23.Q ),
    .A0(Tile_X0Y1_E2MID[5]),
    .A1(Tile_X0Y1_E6END[5]),
    .A2(Tile_X0Y1_E2END[5]),
    .A3(_0079_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit22.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb2 ));
 sg13g2_mux4_1 _0397_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit12.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb2 ),
    .A1(Tile_X0Y1_N2MID[2]),
    .A2(Tile_X0Y0_S2MID[2]),
    .A3(Tile_X0Y0_S2END[2]),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit13.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2 ));
 sg13g2_mux4_1 _0398_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit2.Q ),
    .A0(Tile_X0Y0_E2MID[5]),
    .A1(Tile_X0Y0_E2END[5]),
    .A2(Tile_X0Y0_E6END[5]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit3.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG2 ));
 sg13g2_mux4_1 _0399_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit8.Q ),
    .A0(Tile_X0Y0_E2MID[4]),
    .A1(Tile_X0Y0_E2END[4]),
    .A2(Tile_X0Y0_E6END[11]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit9.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG3 ));
 sg13g2_mux4_1 _0400_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit15.Q ),
    .A0(Tile_X0Y1_N2MID[3]),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG3 ),
    .A2(Tile_X0Y1_N2END[3]),
    .A3(Tile_X0Y0_S2MID[3]),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit14.Q ),
    .X(_0080_));
 sg13g2_mux4_1 _0401_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit25.Q ),
    .A0(Tile_X0Y1_E2MID[4]),
    .A1(Tile_X0Y1_E6END[4]),
    .A2(Tile_X0Y1_E2END[4]),
    .A3(_0080_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit24.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb3 ));
 sg13g2_mux4_1 _0402_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit14.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb3 ),
    .A1(Tile_X0Y1_N2MID[3]),
    .A2(Tile_X0Y0_S2MID[3]),
    .A3(Tile_X0Y0_S2END[3]),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit15.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3 ));
 sg13g2_mux4_1 _0403_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit4.Q ),
    .A0(Tile_X0Y0_E2MID[4]),
    .A1(Tile_X0Y0_E2END[4]),
    .A2(Tile_X0Y0_E6END[4]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit5.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG3 ));
 sg13g2_mux4_1 _0404_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit11.Q ),
    .A0(Tile_X0Y0_E1END[0]),
    .A1(Tile_X0Y0_E2END[3]),
    .A2(Tile_X0Y0_E2MID[3]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG4 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit10.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG4 ));
 sg13g2_mux4_1 _0405_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit16.Q ),
    .A0(Tile_X0Y1_N2MID[4]),
    .A1(Tile_X0Y1_N2END[4]),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG4 ),
    .A3(Tile_X0Y0_S2MID[4]),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit17.Q ),
    .X(_0081_));
 sg13g2_mux4_1 _0406_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit26.Q ),
    .A0(Tile_X0Y1_E2MID[3]),
    .A1(Tile_X0Y1_E2END[3]),
    .A2(Tile_X0Y1_E6END[3]),
    .A3(_0081_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit27.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb4 ));
 sg13g2_mux4_1 _0407_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit17.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb4 ),
    .A1(Tile_X0Y0_S2MID[4]),
    .A2(Tile_X0Y1_N2MID[4]),
    .A3(Tile_X0Y0_S2END[4]),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit16.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG4 ));
 sg13g2_mux4_1 _0408_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit6.Q ),
    .A0(Tile_X0Y0_E2MID[3]),
    .A1(Tile_X0Y0_E2END[3]),
    .A2(Tile_X0Y0_E6END[3]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG4 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit7.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG4 ));
 sg13g2_mux4_1 _0409_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit12.Q ),
    .A0(Tile_X0Y0_E1END[1]),
    .A1(Tile_X0Y0_E2MID[2]),
    .A2(Tile_X0Y0_E2END[2]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG5 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit13.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG5 ));
 sg13g2_mux4_1 _0410_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit18.Q ),
    .A0(Tile_X0Y1_N2MID[5]),
    .A1(Tile_X0Y1_N2END[5]),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG5 ),
    .A3(Tile_X0Y0_S2MID[5]),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit19.Q ),
    .X(_0082_));
 sg13g2_mux4_1 _0411_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit29.Q ),
    .A0(Tile_X0Y1_E2MID[2]),
    .A1(Tile_X0Y1_E6END[2]),
    .A2(Tile_X0Y1_E2END[2]),
    .A3(_0082_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit28.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb5 ));
 sg13g2_mux4_1 _0412_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit19.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb5 ),
    .A1(Tile_X0Y0_S2MID[5]),
    .A2(Tile_X0Y1_N2MID[5]),
    .A3(Tile_X0Y0_S2END[5]),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit18.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG5 ));
 sg13g2_mux4_1 _0413_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit8.Q ),
    .A0(Tile_X0Y0_E2MID[2]),
    .A1(Tile_X0Y0_E2END[2]),
    .A2(Tile_X0Y0_E6END[2]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG5 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit9.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG5 ));
 sg13g2_mux4_1 _0414_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit14.Q ),
    .A0(Tile_X0Y0_E1END[2]),
    .A1(Tile_X0Y0_E2MID[1]),
    .A2(Tile_X0Y0_E2END[1]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG6 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit15.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG6 ));
 sg13g2_mux4_1 _0415_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit20.Q ),
    .A0(Tile_X0Y1_N2MID[6]),
    .A1(Tile_X0Y1_N2END[6]),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG6 ),
    .A3(Tile_X0Y0_S2MID[6]),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit21.Q ),
    .X(_0083_));
 sg13g2_mux4_1 _0416_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit31.Q ),
    .A0(Tile_X0Y1_E2MID[1]),
    .A1(Tile_X0Y1_E6END[1]),
    .A2(Tile_X0Y1_E2END[1]),
    .A3(_0083_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit30.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb6 ));
 sg13g2_mux4_1 _0417_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit21.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb6 ),
    .A1(Tile_X0Y0_S2MID[6]),
    .A2(Tile_X0Y1_N2MID[6]),
    .A3(Tile_X0Y0_S2END[6]),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit20.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG6 ));
 sg13g2_mux4_1 _0418_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit10.Q ),
    .A0(Tile_X0Y0_E2MID[1]),
    .A1(Tile_X0Y0_E2END[1]),
    .A2(Tile_X0Y0_E6END[1]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG6 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit11.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG6 ));
 sg13g2_mux4_1 _0419_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit16.Q ),
    .A0(Tile_X0Y0_E1END[3]),
    .A1(Tile_X0Y0_E2MID[0]),
    .A2(Tile_X0Y0_E2END[0]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG7 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit17.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG7 ));
 sg13g2_mux4_1 _0420_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit22.Q ),
    .A0(Tile_X0Y1_N2MID[7]),
    .A1(Tile_X0Y1_N2END[7]),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG7 ),
    .A3(Tile_X0Y0_S2MID[7]),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit23.Q ),
    .X(_0084_));
 sg13g2_mux4_1 _0421_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit0.Q ),
    .A0(Tile_X0Y1_E2MID[0]),
    .A1(Tile_X0Y1_E2END[0]),
    .A2(Tile_X0Y1_E6END[0]),
    .A3(_0084_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit1.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb7 ));
 sg13g2_mux4_1 _0422_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit23.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb7 ),
    .A1(Tile_X0Y0_S2MID[7]),
    .A2(Tile_X0Y1_N2MID[7]),
    .A3(Tile_X0Y0_S2END[7]),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit22.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG7 ));
 sg13g2_mux4_1 _0423_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit12.Q ),
    .A0(Tile_X0Y0_E2MID[0]),
    .A1(Tile_X0Y0_E2END[0]),
    .A2(Tile_X0Y0_E6END[0]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG7 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit13.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG7 ));
 sg13g2_nand2b_1 _0424_ (.Y(_0085_),
    .B(Tile_X0Y0_S1END[0]),
    .A_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_nor3_1 _0425_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit24.Q ),
    .B(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit25.Q ),
    .C(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END0 ),
    .Y(_0086_));
 sg13g2_a221oi_1 _0426_ (.B2(_0085_),
    .C1(_0086_),
    .B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit25.Q ),
    .A1(_0006_),
    .Y(_0087_),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_mux4_1 _0427_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit27.Q ),
    .A0(Tile_X0Y0_E1END[0]),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 ),
    .A2(Tile_X0Y0_E6END[8]),
    .A3(_0087_),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit26.Q ),
    .X(_0088_));
 sg13g2_nor3_1 _0428_ (.A(Tile_X0Y1_N1END[0]),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q ),
    .C(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit25.Q ),
    .Y(_0089_));
 sg13g2_nand2b_1 _0429_ (.Y(_0090_),
    .B(_0088_),
    .A_N(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_a221oi_1 _0430_ (.B2(_0090_),
    .C1(_0089_),
    .B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit25.Q ),
    .A1(_0010_),
    .Y(_0091_),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_mux4_1 _0431_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit11.Q ),
    .A0(Tile_X0Y1_E1END[0]),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12 ),
    .A2(Tile_X0Y1_E6END[4]),
    .A3(_0091_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit10.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END0 ));
 sg13g2_mux4_1 _0432_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit31.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END0 ),
    .A1(DOUT_SRAM18),
    .A2(Tile_X0Y0_S1END[0]),
    .A3(DOUT_SRAM23),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit30.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG0 ));
 sg13g2_mux4_1 _0433_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit1.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END1 ),
    .A1(DOUT_SRAM19),
    .A2(Tile_X0Y0_S1END[1]),
    .A3(DOUT_SRAM22),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit0.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG1 ));
 sg13g2_mux4_1 _0434_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit3.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END2 ),
    .A1(DOUT_SRAM16),
    .A2(Tile_X0Y0_S1END[2]),
    .A3(DOUT_SRAM21),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit2.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG2 ));
 sg13g2_mux4_1 _0435_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit5.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END3 ),
    .A1(DOUT_SRAM17),
    .A2(Tile_X0Y0_S1END[3]),
    .A3(DOUT_SRAM20),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit4.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG3 ));
 sg13g2_mux4_1 _0436_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit6.Q ),
    .A0(DOUT_SRAM16),
    .A1(DOUT_SRAM24),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG7 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit7.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG0 ));
 sg13g2_mux4_1 _0437_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit8.Q ),
    .A0(DOUT_SRAM17),
    .A1(DOUT_SRAM25),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG6 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit9.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG1 ));
 sg13g2_mux4_1 _0438_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit10.Q ),
    .A0(DOUT_SRAM18),
    .A1(DOUT_SRAM26),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG5 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit11.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG2 ));
 sg13g2_mux4_1 _0439_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit12.Q ),
    .A0(DOUT_SRAM19),
    .A1(DOUT_SRAM27),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG4 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit13.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG3 ));
 sg13g2_mux4_1 _0440_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit14.Q ),
    .A0(DOUT_SRAM20),
    .A1(DOUT_SRAM28),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG4 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit15.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG4 ));
 sg13g2_mux4_1 _0441_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit16.Q ),
    .A0(DOUT_SRAM21),
    .A1(DOUT_SRAM29),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG5 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit17.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG5 ));
 sg13g2_mux4_1 _0442_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit18.Q ),
    .A0(DOUT_SRAM22),
    .A1(DOUT_SRAM30),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG6 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit19.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG6 ));
 sg13g2_mux4_1 _0443_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit20.Q ),
    .A0(DOUT_SRAM23),
    .A1(DOUT_SRAM31),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG7 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit21.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG7 ));
 sg13g2_mux4_1 _0444_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit22.Q ),
    .A0(DOUT_SRAM16),
    .A1(DOUT_SRAM24),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG7 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit23.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb0 ));
 sg13g2_mux4_1 _0445_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit24.Q ),
    .A0(DOUT_SRAM17),
    .A1(DOUT_SRAM25),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG6 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit25.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb1 ));
 sg13g2_mux4_1 _0446_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit26.Q ),
    .A0(DOUT_SRAM18),
    .A1(DOUT_SRAM26),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG5 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit27.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb2 ));
 sg13g2_mux4_1 _0447_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit28.Q ),
    .A0(DOUT_SRAM19),
    .A1(DOUT_SRAM27),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG4 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit29.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb3 ));
 sg13g2_mux4_1 _0448_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit30.Q ),
    .A0(DOUT_SRAM20),
    .A1(DOUT_SRAM28),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG4 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit31.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb4 ));
 sg13g2_mux4_1 _0449_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit0.Q ),
    .A0(DOUT_SRAM21),
    .A1(DOUT_SRAM29),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG5 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit1.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb5 ));
 sg13g2_mux4_1 _0450_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit2.Q ),
    .A0(DOUT_SRAM22),
    .A1(DOUT_SRAM30),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG6 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit3.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb6 ));
 sg13g2_mux4_1 _0451_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit4.Q ),
    .A0(DOUT_SRAM23),
    .A1(DOUT_SRAM31),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG7 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit5.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb7 ));
 sg13g2_mux4_1 _0452_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit6.Q ),
    .A0(DOUT_SRAM16),
    .A1(DOUT_SRAM28),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG7 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit7.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG0 ));
 sg13g2_mux4_1 _0453_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit8.Q ),
    .A0(DOUT_SRAM17),
    .A1(DOUT_SRAM29),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG6 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit9.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG1 ));
 sg13g2_mux4_1 _0454_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit10.Q ),
    .A0(DOUT_SRAM18),
    .A1(DOUT_SRAM30),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG5 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit11.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG2 ));
 sg13g2_mux4_1 _0455_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit0.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END0 ),
    .A1(Tile_X0Y1_N4END[4]),
    .A2(Tile_X0Y0_S1END[0]),
    .A3(Tile_X0Y0_S4END[0]),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit1.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 ));
 sg13g2_mux4_1 _0456_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit12.Q ),
    .A0(DOUT_SRAM19),
    .A1(DOUT_SRAM31),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG4 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit13.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG3 ));
 sg13g2_mux4_1 _0457_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit30.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END3 ),
    .A1(Tile_X0Y1_N4END[7]),
    .A2(Tile_X0Y0_S1END[3]),
    .A3(Tile_X0Y0_S4END[3]),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit31.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11 ));
 sg13g2_mux4_1 _0458_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit14.Q ),
    .A0(DOUT_SRAM20),
    .A1(DOUT_SRAM24),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit15.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG4 ));
 sg13g2_mux4_1 _0459_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit28.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END2 ),
    .A1(Tile_X0Y1_N4END[6]),
    .A2(Tile_X0Y0_S1END[2]),
    .A3(Tile_X0Y0_S4END[2]),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit29.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10 ));
 sg13g2_mux4_1 _0460_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit16.Q ),
    .A0(DOUT_SRAM21),
    .A1(DOUT_SRAM24),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit17.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG5 ));
 sg13g2_mux4_1 _0461_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit26.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END1 ),
    .A1(Tile_X0Y1_N4END[5]),
    .A2(Tile_X0Y0_S1END[1]),
    .A3(Tile_X0Y0_S4END[1]),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit27.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9 ));
 sg13g2_mux4_1 _0462_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit18.Q ),
    .A0(DOUT_SRAM22),
    .A1(DOUT_SRAM26),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit19.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG6 ));
 sg13g2_mux4_1 _0463_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit24.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END0 ),
    .A1(Tile_X0Y1_N4END[4]),
    .A2(Tile_X0Y0_S1END[0]),
    .A3(Tile_X0Y0_S4END[0]),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit25.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8 ));
 sg13g2_mux4_1 _0464_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit20.Q ),
    .A0(DOUT_SRAM23),
    .A1(DOUT_SRAM27),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit21.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG7 ));
 sg13g2_mux4_1 _0465_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit22.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END3 ),
    .A1(Tile_X0Y1_N4END[7]),
    .A2(Tile_X0Y0_S1END[3]),
    .A3(Tile_X0Y0_S4END[3]),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit23.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7 ));
 sg13g2_mux4_1 _0466_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit22.Q ),
    .A0(DOUT_SRAM20),
    .A1(DOUT_SRAM24),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG7 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit23.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG8 ));
 sg13g2_mux4_1 _0467_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit20.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END2 ),
    .A1(Tile_X0Y1_N4END[6]),
    .A2(Tile_X0Y0_S1END[2]),
    .A3(Tile_X0Y0_S4END[2]),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit21.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6 ));
 sg13g2_mux4_1 _0468_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit24.Q ),
    .A0(DOUT_SRAM21),
    .A1(DOUT_SRAM25),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG6 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit25.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG9 ));
 sg13g2_mux4_1 _0469_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit18.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END1 ),
    .A1(Tile_X0Y1_N4END[5]),
    .A2(Tile_X0Y0_S1END[1]),
    .A3(Tile_X0Y0_S4END[1]),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit19.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5 ));
 sg13g2_mux4_1 _0470_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit26.Q ),
    .A0(DOUT_SRAM22),
    .A1(DOUT_SRAM26),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG5 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit27.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG10 ));
 sg13g2_mux4_1 _0471_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit16.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END0 ),
    .A1(Tile_X0Y1_N4END[4]),
    .A2(Tile_X0Y0_S1END[0]),
    .A3(Tile_X0Y0_S4END[0]),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit17.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4 ));
 sg13g2_mux4_1 _0472_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit28.Q ),
    .A0(DOUT_SRAM23),
    .A1(DOUT_SRAM27),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG4 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit29.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG11 ));
 sg13g2_mux4_1 _0473_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit14.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END3 ),
    .A1(Tile_X0Y1_N4END[7]),
    .A2(Tile_X0Y0_S1END[3]),
    .A3(Tile_X0Y0_S4END[3]),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit15.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG3 ));
 sg13g2_mux4_1 _0474_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit30.Q ),
    .A0(DOUT_SRAM16),
    .A1(DOUT_SRAM28),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG3 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit31.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG12 ));
 sg13g2_mux4_1 _0475_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit12.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END2 ),
    .A1(Tile_X0Y1_N4END[6]),
    .A2(Tile_X0Y0_S1END[2]),
    .A3(Tile_X0Y0_S4END[2]),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit13.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG2 ));
 sg13g2_mux4_1 _0476_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit0.Q ),
    .A0(DOUT_SRAM17),
    .A1(DOUT_SRAM29),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG2 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit1.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG13 ));
 sg13g2_mux4_1 _0477_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit10.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END1 ),
    .A1(Tile_X0Y1_N4END[5]),
    .A2(Tile_X0Y0_S1END[1]),
    .A3(Tile_X0Y0_S4END[1]),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit11.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG1 ));
 sg13g2_mux4_1 _0478_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit2.Q ),
    .A0(DOUT_SRAM18),
    .A1(DOUT_SRAM30),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG1 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit3.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG14 ));
 sg13g2_mux4_1 _0479_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit8.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END0 ),
    .A1(Tile_X0Y1_N4END[4]),
    .A2(Tile_X0Y0_S1END[0]),
    .A3(Tile_X0Y0_S4END[0]),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit9.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG0 ));
 sg13g2_mux4_1 _0480_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit4.Q ),
    .A0(DOUT_SRAM19),
    .A1(DOUT_SRAM31),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG0 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit5.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG15 ));
 sg13g2_mux4_1 _0481_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit6.Q ),
    .A0(Tile_X0Y1_N4END[4]),
    .A1(Tile_X0Y0_S4END[0]),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit7.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG0 ));
 sg13g2_mux4_1 _0482_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit8.Q ),
    .A0(Tile_X0Y1_N4END[5]),
    .A1(Tile_X0Y0_S4END[1]),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit9.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG1 ));
 sg13g2_mux4_1 _0483_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit10.Q ),
    .A0(Tile_X0Y1_N4END[6]),
    .A1(Tile_X0Y0_S4END[2]),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit11.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG2 ));
 sg13g2_mux4_1 _0484_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit12.Q ),
    .A0(Tile_X0Y1_N4END[7]),
    .A1(Tile_X0Y0_S4END[3]),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit13.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG3 ));
 sg13g2_mux4_1 _0485_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit15.Q ),
    .A0(DOUT_SRAM20),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11 ),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit14.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG4 ));
 sg13g2_mux4_1 _0486_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit17.Q ),
    .A0(DOUT_SRAM21),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10 ),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit16.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG5 ));
 sg13g2_mux4_1 _0487_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit18.Q ),
    .A0(DOUT_SRAM22),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5 ),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit19.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG6 ));
 sg13g2_mux4_1 _0488_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit20.Q ),
    .A0(DOUT_SRAM23),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4 ),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit21.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG7 ));
 sg13g2_mux4_1 _0489_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit23.Q ),
    .A0(DOUT_SRAM16),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7 ),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG3 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG4 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit22.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG8 ));
 sg13g2_mux4_1 _0490_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit25.Q ),
    .A0(DOUT_SRAM17),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6 ),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG2 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG5 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit24.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG9 ));
 sg13g2_mux4_1 _0491_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit27.Q ),
    .A0(DOUT_SRAM18),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5 ),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG1 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG6 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit26.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG10 ));
 sg13g2_mux4_1 _0492_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit29.Q ),
    .A0(DOUT_SRAM19),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4 ),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG0 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG7 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit28.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG11 ));
 sg13g2_mux4_1 _0493_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit30.Q ),
    .A0(Tile_X0Y0_EE4END[0]),
    .A1(Tile_X0Y0_EE4END[8]),
    .A2(Tile_X0Y0_E6END[0]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG0 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit31.Q ),
    .X(DIN_SRAM16));
 sg13g2_mux4_1 _0494_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit0.Q ),
    .A0(Tile_X0Y0_EE4END[1]),
    .A1(Tile_X0Y0_EE4END[9]),
    .A2(Tile_X0Y0_E6END[1]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG1 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit1.Q ),
    .X(DIN_SRAM17));
 sg13g2_mux4_1 _0495_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit2.Q ),
    .A0(Tile_X0Y0_EE4END[2]),
    .A1(Tile_X0Y0_EE4END[10]),
    .A2(Tile_X0Y0_E6END[2]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG2 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit3.Q ),
    .X(DIN_SRAM18));
 sg13g2_mux4_1 _0496_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit4.Q ),
    .A0(Tile_X0Y0_EE4END[3]),
    .A1(Tile_X0Y0_EE4END[11]),
    .A2(Tile_X0Y0_E6END[3]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG3 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit5.Q ),
    .X(DIN_SRAM19));
 sg13g2_mux4_1 _0497_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit6.Q ),
    .A0(Tile_X0Y0_EE4END[4]),
    .A1(Tile_X0Y0_EE4END[12]),
    .A2(Tile_X0Y0_E6END[4]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit7.Q ),
    .X(DIN_SRAM20));
 sg13g2_mux4_1 _0498_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit8.Q ),
    .A0(Tile_X0Y0_EE4END[5]),
    .A1(Tile_X0Y0_EE4END[13]),
    .A2(Tile_X0Y0_E6END[5]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit9.Q ),
    .X(DIN_SRAM21));
 sg13g2_mux4_1 _0499_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit10.Q ),
    .A0(Tile_X0Y0_EE4END[6]),
    .A1(Tile_X0Y0_EE4END[14]),
    .A2(Tile_X0Y0_E6END[6]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit11.Q ),
    .X(DIN_SRAM22));
 sg13g2_mux4_1 _0500_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit12.Q ),
    .A0(Tile_X0Y0_EE4END[7]),
    .A1(Tile_X0Y0_EE4END[15]),
    .A2(Tile_X0Y0_E6END[7]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit13.Q ),
    .X(DIN_SRAM23));
 sg13g2_mux4_1 _0501_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit14.Q ),
    .A0(Tile_X0Y0_EE4END[0]),
    .A1(Tile_X0Y0_EE4END[8]),
    .A2(Tile_X0Y0_E6END[8]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit15.Q ),
    .X(DIN_SRAM24));
 sg13g2_mux4_1 _0502_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit16.Q ),
    .A0(Tile_X0Y0_EE4END[1]),
    .A1(Tile_X0Y0_EE4END[9]),
    .A2(Tile_X0Y0_E6END[9]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit17.Q ),
    .X(DIN_SRAM25));
 sg13g2_mux4_1 _0503_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit18.Q ),
    .A0(Tile_X0Y0_EE4END[2]),
    .A1(Tile_X0Y0_EE4END[10]),
    .A2(Tile_X0Y0_E6END[10]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit19.Q ),
    .X(DIN_SRAM26));
 sg13g2_mux4_1 _0504_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit20.Q ),
    .A0(Tile_X0Y0_EE4END[3]),
    .A1(Tile_X0Y0_EE4END[11]),
    .A2(Tile_X0Y0_E6END[11]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit21.Q ),
    .X(DIN_SRAM27));
 sg13g2_mux4_1 _0505_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit22.Q ),
    .A0(Tile_X0Y0_E1END[0]),
    .A1(Tile_X0Y0_EE4END[4]),
    .A2(Tile_X0Y0_EE4END[12]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit23.Q ),
    .X(DIN_SRAM28));
 sg13g2_mux4_1 _0506_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit24.Q ),
    .A0(Tile_X0Y0_E1END[1]),
    .A1(Tile_X0Y0_EE4END[5]),
    .A2(Tile_X0Y0_EE4END[13]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit25.Q ),
    .X(DIN_SRAM29));
 sg13g2_mux4_1 _0507_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit26.Q ),
    .A0(Tile_X0Y0_E1END[2]),
    .A1(Tile_X0Y0_EE4END[6]),
    .A2(Tile_X0Y0_EE4END[14]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit27.Q ),
    .X(DIN_SRAM30));
 sg13g2_mux4_1 _0508_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit28.Q ),
    .A0(Tile_X0Y0_E1END[3]),
    .A1(Tile_X0Y0_EE4END[7]),
    .A2(Tile_X0Y0_EE4END[15]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit29.Q ),
    .X(DIN_SRAM31));
 sg13g2_mux4_1 _0509_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit30.Q ),
    .A0(Tile_X0Y0_EE4END[0]),
    .A1(Tile_X0Y0_EE4END[8]),
    .A2(Tile_X0Y0_E6END[0]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG0 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit31.Q ),
    .X(BM_SRAM16));
 sg13g2_mux4_1 _0510_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit0.Q ),
    .A0(Tile_X0Y0_EE4END[1]),
    .A1(Tile_X0Y0_EE4END[9]),
    .A2(Tile_X0Y0_E6END[1]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG1 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit1.Q ),
    .X(BM_SRAM17));
 sg13g2_mux4_1 _0511_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit2.Q ),
    .A0(Tile_X0Y0_EE4END[2]),
    .A1(Tile_X0Y0_EE4END[10]),
    .A2(Tile_X0Y0_E6END[2]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG2 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit3.Q ),
    .X(BM_SRAM18));
 sg13g2_mux4_1 _0512_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit4.Q ),
    .A0(Tile_X0Y0_EE4END[3]),
    .A1(Tile_X0Y0_EE4END[11]),
    .A2(Tile_X0Y0_E6END[3]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG3 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit5.Q ),
    .X(BM_SRAM19));
 sg13g2_mux4_1 _0513_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit6.Q ),
    .A0(Tile_X0Y0_EE4END[4]),
    .A1(Tile_X0Y0_EE4END[12]),
    .A2(Tile_X0Y0_E6END[4]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit7.Q ),
    .X(BM_SRAM20));
 sg13g2_mux4_1 _0514_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit8.Q ),
    .A0(Tile_X0Y0_EE4END[5]),
    .A1(Tile_X0Y0_EE4END[13]),
    .A2(Tile_X0Y0_E6END[5]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit9.Q ),
    .X(BM_SRAM21));
 sg13g2_mux4_1 _0515_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit10.Q ),
    .A0(Tile_X0Y0_EE4END[6]),
    .A1(Tile_X0Y0_EE4END[14]),
    .A2(Tile_X0Y0_E6END[6]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit11.Q ),
    .X(BM_SRAM22));
 sg13g2_mux4_1 _0516_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit12.Q ),
    .A0(Tile_X0Y0_EE4END[7]),
    .A1(Tile_X0Y0_EE4END[15]),
    .A2(Tile_X0Y0_E6END[7]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit13.Q ),
    .X(BM_SRAM23));
 sg13g2_mux4_1 _0517_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit14.Q ),
    .A0(Tile_X0Y0_EE4END[0]),
    .A1(Tile_X0Y0_EE4END[8]),
    .A2(Tile_X0Y0_E6END[8]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit15.Q ),
    .X(BM_SRAM24));
 sg13g2_mux4_1 _0518_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit16.Q ),
    .A0(Tile_X0Y0_EE4END[1]),
    .A1(Tile_X0Y0_EE4END[9]),
    .A2(Tile_X0Y0_E6END[9]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit17.Q ),
    .X(BM_SRAM25));
 sg13g2_mux4_1 _0519_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit18.Q ),
    .A0(Tile_X0Y0_EE4END[2]),
    .A1(Tile_X0Y0_EE4END[10]),
    .A2(Tile_X0Y0_E6END[10]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit19.Q ),
    .X(BM_SRAM26));
 sg13g2_mux4_1 _0520_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit20.Q ),
    .A0(Tile_X0Y0_EE4END[3]),
    .A1(Tile_X0Y0_EE4END[11]),
    .A2(Tile_X0Y0_E6END[11]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit21.Q ),
    .X(BM_SRAM27));
 sg13g2_mux4_1 _0521_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit22.Q ),
    .A0(Tile_X0Y0_E1END[0]),
    .A1(Tile_X0Y0_EE4END[4]),
    .A2(Tile_X0Y0_EE4END[12]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit23.Q ),
    .X(BM_SRAM28));
 sg13g2_mux4_1 _0522_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit24.Q ),
    .A0(Tile_X0Y0_E1END[1]),
    .A1(Tile_X0Y0_EE4END[5]),
    .A2(Tile_X0Y0_EE4END[13]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit25.Q ),
    .X(BM_SRAM29));
 sg13g2_mux4_1 _0523_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit26.Q ),
    .A0(Tile_X0Y0_E1END[2]),
    .A1(Tile_X0Y0_EE4END[6]),
    .A2(Tile_X0Y0_EE4END[14]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit27.Q ),
    .X(BM_SRAM30));
 sg13g2_mux4_1 _0524_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit28.Q ),
    .A0(Tile_X0Y0_E1END[3]),
    .A1(Tile_X0Y0_EE4END[7]),
    .A2(Tile_X0Y0_EE4END[15]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit29.Q ),
    .X(BM_SRAM31));
 sg13g2_nor3_1 _0525_ (.A(Tile_X0Y0_E2MID[0]),
    .B(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit30.Q ),
    .C(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit31.Q ),
    .Y(_0092_));
 sg13g2_nand2b_1 _0526_ (.Y(_0093_),
    .B(Tile_X0Y0_E2END[0]),
    .A_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit31.Q ));
 sg13g2_a221oi_1 _0527_ (.B2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit30.Q ),
    .C1(_0092_),
    .B1(_0093_),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit31.Q ),
    .Y(ADDR_SRAM5),
    .A2(_0038_));
 sg13g2_nor3_1 _0528_ (.A(Tile_X0Y0_E2MID[1]),
    .B(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit0.Q ),
    .C(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit1.Q ),
    .Y(_0094_));
 sg13g2_nand2b_1 _0529_ (.Y(_0095_),
    .B(Tile_X0Y0_E2END[1]),
    .A_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit1.Q ));
 sg13g2_a221oi_1 _0530_ (.B2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit0.Q ),
    .C1(_0094_),
    .B1(_0095_),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit1.Q ),
    .Y(ADDR_SRAM6),
    .A2(_0039_));
 sg13g2_nor3_1 _0531_ (.A(Tile_X0Y0_E2MID[2]),
    .B(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit2.Q ),
    .C(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit3.Q ),
    .Y(_0096_));
 sg13g2_nand2b_1 _0532_ (.Y(_0097_),
    .B(Tile_X0Y0_E2END[2]),
    .A_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit3.Q ));
 sg13g2_a221oi_1 _0533_ (.B2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit2.Q ),
    .C1(_0096_),
    .B1(_0097_),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit3.Q ),
    .Y(ADDR_SRAM7),
    .A2(_0040_));
 sg13g2_nor3_1 _0534_ (.A(Tile_X0Y0_E2MID[3]),
    .B(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit4.Q ),
    .C(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit5.Q ),
    .Y(_0098_));
 sg13g2_nand2b_1 _0535_ (.Y(_0099_),
    .B(Tile_X0Y0_E2END[3]),
    .A_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit5.Q ));
 sg13g2_a221oi_1 _0536_ (.B2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit4.Q ),
    .C1(_0098_),
    .B1(_0099_),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit5.Q ),
    .Y(ADDR_SRAM8),
    .A2(_0041_));
 sg13g2_nor3_1 _0537_ (.A(Tile_X0Y0_E2MID[4]),
    .B(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit6.Q ),
    .C(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit7.Q ),
    .Y(_0100_));
 sg13g2_nand2b_1 _0538_ (.Y(_0101_),
    .B(Tile_X0Y0_E2END[4]),
    .A_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit7.Q ));
 sg13g2_a221oi_1 _0539_ (.B2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit6.Q ),
    .C1(_0100_),
    .B1(_0101_),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit7.Q ),
    .Y(ADDR_SRAM9),
    .A2(_0042_));
 sg13g2_mux2_1 _0540_ (.A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4 ),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8 ),
    .S(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit14.Q ),
    .X(_0102_));
 sg13g2_nor2b_1 _0541_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0 ),
    .B_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit14.Q ),
    .Y(_0103_));
 sg13g2_o21ai_1 _0542_ (.B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit15.Q ),
    .Y(_0104_),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit14.Q ),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 ));
 sg13g2_o21ai_1 _0543_ (.B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit16.Q ),
    .Y(_0105_),
    .A1(_0103_),
    .A2(_0104_));
 sg13g2_a21oi_1 _0544_ (.A1(_0011_),
    .A2(_0102_),
    .Y(_0106_),
    .B1(_0105_));
 sg13g2_mux4_1 _0545_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit14.Q ),
    .A0(Tile_X0Y0_E1END[0]),
    .A1(Tile_X0Y0_EE4END[0]),
    .A2(Tile_X0Y0_E6END[8]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG0 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit15.Q ),
    .X(_0107_));
 sg13g2_nor2_1 _0546_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit16.Q ),
    .B(_0107_),
    .Y(_0108_));
 sg13g2_nor2_1 _0547_ (.A(_0106_),
    .B(_0108_),
    .Y(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG0 ));
 sg13g2_mux2_1 _0548_ (.A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5 ),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9 ),
    .S(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit17.Q ),
    .X(_0109_));
 sg13g2_nor2b_1 _0549_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1 ),
    .B_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit17.Q ),
    .Y(_0110_));
 sg13g2_o21ai_1 _0550_ (.B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit18.Q ),
    .Y(_0111_),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit17.Q ),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13 ));
 sg13g2_o21ai_1 _0551_ (.B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit19.Q ),
    .Y(_0112_),
    .A1(_0110_),
    .A2(_0111_));
 sg13g2_a21oi_1 _0552_ (.A1(_0012_),
    .A2(_0109_),
    .Y(_0113_),
    .B1(_0112_));
 sg13g2_mux4_1 _0553_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit18.Q ),
    .A0(Tile_X0Y0_E1END[1]),
    .A1(Tile_X0Y0_E6END[9]),
    .A2(Tile_X0Y0_EE4END[1]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG1 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit17.Q ),
    .X(_0114_));
 sg13g2_nor2_1 _0554_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit19.Q ),
    .B(_0114_),
    .Y(_0115_));
 sg13g2_nor2_1 _0555_ (.A(_0113_),
    .B(_0115_),
    .Y(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG1 ));
 sg13g2_mux2_1 _0556_ (.A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6 ),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10 ),
    .S(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit20.Q ),
    .X(_0116_));
 sg13g2_nor2b_1 _0557_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2 ),
    .B_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit20.Q ),
    .Y(_0117_));
 sg13g2_o21ai_1 _0558_ (.B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit21.Q ),
    .Y(_0118_),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit20.Q ),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14 ));
 sg13g2_o21ai_1 _0559_ (.B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit22.Q ),
    .Y(_0119_),
    .A1(_0117_),
    .A2(_0118_));
 sg13g2_a21oi_1 _0560_ (.A1(_0013_),
    .A2(_0116_),
    .Y(_0120_),
    .B1(_0119_));
 sg13g2_mux4_1 _0561_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit21.Q ),
    .A0(Tile_X0Y0_E1END[2]),
    .A1(Tile_X0Y0_E6END[10]),
    .A2(Tile_X0Y0_EE4END[2]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG2 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit20.Q ),
    .X(_0121_));
 sg13g2_nor2_1 _0562_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit22.Q ),
    .B(_0121_),
    .Y(_0122_));
 sg13g2_nor2_1 _0563_ (.A(_0120_),
    .B(_0122_),
    .Y(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG2 ));
 sg13g2_mux2_1 _0564_ (.A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7 ),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11 ),
    .S(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit23.Q ),
    .X(_0123_));
 sg13g2_nor2b_1 _0565_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3 ),
    .B_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit23.Q ),
    .Y(_0124_));
 sg13g2_o21ai_1 _0566_ (.B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit24.Q ),
    .Y(_0125_),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit23.Q ),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15 ));
 sg13g2_o21ai_1 _0567_ (.B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit25.Q ),
    .Y(_0126_),
    .A1(_0124_),
    .A2(_0125_));
 sg13g2_a21oi_1 _0568_ (.A1(_0014_),
    .A2(_0123_),
    .Y(_0127_),
    .B1(_0126_));
 sg13g2_mux4_1 _0569_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit24.Q ),
    .A0(Tile_X0Y0_E1END[3]),
    .A1(Tile_X0Y0_E6END[11]),
    .A2(Tile_X0Y0_EE4END[3]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG3 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit23.Q ),
    .X(_0128_));
 sg13g2_nor2_1 _0570_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit25.Q ),
    .B(_0128_),
    .Y(_0129_));
 sg13g2_nor2_1 _0571_ (.A(_0127_),
    .B(_0129_),
    .Y(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG3 ));
 sg13g2_mux2_1 _0572_ (.A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4 ),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8 ),
    .S(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit18.Q ),
    .X(_0130_));
 sg13g2_nor2b_1 _0573_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG4 ),
    .B_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit18.Q ),
    .Y(_0131_));
 sg13g2_o21ai_1 _0574_ (.B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit19.Q ),
    .Y(_0132_),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit18.Q ),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 ));
 sg13g2_o21ai_1 _0575_ (.B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit20.Q ),
    .Y(_0133_),
    .A1(_0131_),
    .A2(_0132_));
 sg13g2_a21oi_1 _0576_ (.A1(_0015_),
    .A2(_0130_),
    .Y(_0134_),
    .B1(_0133_));
 sg13g2_mux4_1 _0577_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit18.Q ),
    .A0(Tile_X0Y0_E1END[0]),
    .A1(Tile_X0Y0_EE4END[12]),
    .A2(Tile_X0Y0_E6END[4]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG0 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit19.Q ),
    .X(_0135_));
 sg13g2_nor2_1 _0578_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit20.Q ),
    .B(_0135_),
    .Y(_0136_));
 sg13g2_nor2_1 _0579_ (.A(_0134_),
    .B(_0136_),
    .Y(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG0 ));
 sg13g2_mux2_1 _0580_ (.A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5 ),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9 ),
    .S(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit21.Q ),
    .X(_0137_));
 sg13g2_nor2b_1 _0581_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG5 ),
    .B_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit21.Q ),
    .Y(_0138_));
 sg13g2_o21ai_1 _0582_ (.B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit22.Q ),
    .Y(_0139_),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit21.Q ),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13 ));
 sg13g2_o21ai_1 _0583_ (.B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit23.Q ),
    .Y(_0140_),
    .A1(_0138_),
    .A2(_0139_));
 sg13g2_a21oi_1 _0584_ (.A1(_0016_),
    .A2(_0137_),
    .Y(_0141_),
    .B1(_0140_));
 sg13g2_mux4_1 _0585_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit22.Q ),
    .A0(Tile_X0Y0_E1END[1]),
    .A1(Tile_X0Y0_E6END[5]),
    .A2(Tile_X0Y0_EE4END[13]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG1 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit21.Q ),
    .X(_0142_));
 sg13g2_nor2_1 _0586_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit23.Q ),
    .B(_0142_),
    .Y(_0143_));
 sg13g2_nor2_1 _0587_ (.A(_0141_),
    .B(_0143_),
    .Y(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG1 ));
 sg13g2_mux2_1 _0588_ (.A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6 ),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10 ),
    .S(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit24.Q ),
    .X(_0144_));
 sg13g2_nor2b_1 _0589_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG6 ),
    .B_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit24.Q ),
    .Y(_0145_));
 sg13g2_o21ai_1 _0590_ (.B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit25.Q ),
    .Y(_0146_),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit24.Q ),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14 ));
 sg13g2_o21ai_1 _0591_ (.B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit26.Q ),
    .Y(_0147_),
    .A1(_0145_),
    .A2(_0146_));
 sg13g2_a21oi_1 _0592_ (.A1(_0017_),
    .A2(_0144_),
    .Y(_0148_),
    .B1(_0147_));
 sg13g2_mux4_1 _0593_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit25.Q ),
    .A0(Tile_X0Y0_E1END[2]),
    .A1(Tile_X0Y0_E6END[6]),
    .A2(Tile_X0Y0_EE4END[14]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG2 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit24.Q ),
    .X(_0149_));
 sg13g2_nor2_1 _0594_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit26.Q ),
    .B(_0149_),
    .Y(_0150_));
 sg13g2_nor2_1 _0595_ (.A(_0148_),
    .B(_0150_),
    .Y(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG2 ));
 sg13g2_mux2_1 _0596_ (.A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7 ),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11 ),
    .S(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit27.Q ),
    .X(_0151_));
 sg13g2_nor2b_1 _0597_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG7 ),
    .B_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit27.Q ),
    .Y(_0152_));
 sg13g2_o21ai_1 _0598_ (.B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit28.Q ),
    .Y(_0153_),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit27.Q ),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15 ));
 sg13g2_o21ai_1 _0599_ (.B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit29.Q ),
    .Y(_0154_),
    .A1(_0152_),
    .A2(_0153_));
 sg13g2_a21oi_1 _0600_ (.A1(_0018_),
    .A2(_0151_),
    .Y(_0155_),
    .B1(_0154_));
 sg13g2_mux4_1 _0601_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit28.Q ),
    .A0(Tile_X0Y0_E1END[3]),
    .A1(Tile_X0Y0_E6END[7]),
    .A2(Tile_X0Y0_EE4END[15]),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG3 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit27.Q ),
    .X(_0156_));
 sg13g2_nor2_1 _0602_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit29.Q ),
    .B(_0156_),
    .Y(_0157_));
 sg13g2_nor2_1 _0603_ (.A(_0155_),
    .B(_0157_),
    .Y(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG3 ));
 sg13g2_mux4_1 _0604_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit0.Q ),
    .A0(Tile_X0Y1_N1END[0]),
    .A1(Tile_X0Y1_N4END[0]),
    .A2(_0088_),
    .A3(Tile_X0Y0_S4END[4]),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit1.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12 ));
 sg13g2_mux4_1 _0605_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit2.Q ),
    .A0(Tile_X0Y1_N1END[1]),
    .A1(Tile_X0Y1_N4END[1]),
    .A2(_0060_),
    .A3(Tile_X0Y0_S4END[5]),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit3.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13 ));
 sg13g2_mux4_1 _0606_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit4.Q ),
    .A0(Tile_X0Y1_N1END[2]),
    .A1(Tile_X0Y1_N4END[2]),
    .A2(_0067_),
    .A3(Tile_X0Y0_S4END[6]),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit5.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14 ));
 sg13g2_mux4_1 _0607_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit6.Q ),
    .A0(Tile_X0Y1_N1END[3]),
    .A1(Tile_X0Y1_N4END[3]),
    .A2(_0074_),
    .A3(Tile_X0Y0_S4END[7]),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit7.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15 ));
 sg13g2_mux4_1 _0608_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit23.Q ),
    .A0(Tile_X0Y0_E1END[0]),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 ),
    .A2(Tile_X0Y0_E6END[4]),
    .A3(_0087_),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit22.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG0 ));
 sg13g2_mux4_1 _0609_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit14.Q ),
    .A0(Tile_X0Y1_E1END[0]),
    .A1(Tile_X0Y1_E6END[8]),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12 ),
    .A3(_0091_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit15.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG0 ));
 sg13g2_mux4_1 _0610_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit16.Q ),
    .A0(Tile_X0Y1_E1END[1]),
    .A1(Tile_X0Y1_E6END[9]),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13 ),
    .A3(_0063_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit17.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG1 ));
 sg13g2_mux4_1 _0611_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit18.Q ),
    .A0(Tile_X0Y1_E1END[2]),
    .A1(Tile_X0Y1_E6END[10]),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14 ),
    .A3(_0070_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit19.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG2 ));
 sg13g2_mux4_1 _0612_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit20.Q ),
    .A0(Tile_X0Y1_E1END[3]),
    .A1(Tile_X0Y1_E6END[11]),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15 ),
    .A3(_0077_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit21.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG3 ));
 sg13g2_mux4_1 _0613_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit22.Q ),
    .A0(Tile_X0Y1_E2MID[7]),
    .A1(Tile_X0Y1_E2END[7]),
    .A2(Tile_X0Y1_E6END[8]),
    .A3(_0043_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit23.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG0 ));
 sg13g2_mux4_1 _0614_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit24.Q ),
    .A0(Tile_X0Y1_E2MID[6]),
    .A1(Tile_X0Y1_E2END[6]),
    .A2(Tile_X0Y1_E6END[9]),
    .A3(_0078_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit25.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG1 ));
 sg13g2_mux4_1 _0615_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit27.Q ),
    .A0(Tile_X0Y1_E2MID[5]),
    .A1(Tile_X0Y1_E6END[10]),
    .A2(Tile_X0Y1_E2END[5]),
    .A3(_0079_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit26.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG2 ));
 sg13g2_mux4_1 _0616_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit29.Q ),
    .A0(Tile_X0Y1_E2MID[4]),
    .A1(Tile_X0Y1_E6END[11]),
    .A2(Tile_X0Y1_E2END[4]),
    .A3(_0080_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit28.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG3 ));
 sg13g2_mux4_1 _0617_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit31.Q ),
    .A0(Tile_X0Y1_E1END[0]),
    .A1(Tile_X0Y1_E2END[3]),
    .A2(Tile_X0Y1_E2MID[3]),
    .A3(_0081_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit30.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG4 ));
 sg13g2_mux4_1 _0618_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit0.Q ),
    .A0(Tile_X0Y1_E1END[1]),
    .A1(Tile_X0Y1_E2MID[2]),
    .A2(Tile_X0Y1_E2END[2]),
    .A3(_0082_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit1.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG5 ));
 sg13g2_mux4_1 _0619_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit2.Q ),
    .A0(Tile_X0Y1_E1END[2]),
    .A1(Tile_X0Y1_E2MID[1]),
    .A2(Tile_X0Y1_E2END[1]),
    .A3(_0083_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit3.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG6 ));
 sg13g2_mux4_1 _0620_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit5.Q ),
    .A0(Tile_X0Y1_E1END[3]),
    .A1(Tile_X0Y1_E2END[0]),
    .A2(Tile_X0Y1_E2MID[0]),
    .A3(_0084_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit4.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG7 ));
 sg13g2_mux4_1 _0621_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit19.Q ),
    .A0(Tile_X0Y1_N1END[0]),
    .A1(DOUT_SRAM2),
    .A2(_0088_),
    .A3(DOUT_SRAM7),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit18.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG0 ));
 sg13g2_mux4_1 _0622_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit21.Q ),
    .A0(Tile_X0Y1_N1END[1]),
    .A1(DOUT_SRAM3),
    .A2(_0060_),
    .A3(DOUT_SRAM6),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit20.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG1 ));
 sg13g2_mux4_1 _0623_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit23.Q ),
    .A0(Tile_X0Y1_N1END[2]),
    .A1(DOUT_SRAM0),
    .A2(_0067_),
    .A3(DOUT_SRAM5),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit22.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG2 ));
 sg13g2_mux4_1 _0624_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit25.Q ),
    .A0(Tile_X0Y1_N1END[3]),
    .A1(DOUT_SRAM1),
    .A2(_0074_),
    .A3(DOUT_SRAM4),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit24.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG3 ));
 sg13g2_mux4_1 _0625_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit26.Q ),
    .A0(DOUT_SRAM0),
    .A1(DOUT_SRAM8),
    .A2(_0043_),
    .A3(_0084_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit27.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG0 ));
 sg13g2_mux4_1 _0626_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit28.Q ),
    .A0(DOUT_SRAM1),
    .A1(DOUT_SRAM9),
    .A2(_0078_),
    .A3(_0083_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit29.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG1 ));
 sg13g2_mux4_1 _0627_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit30.Q ),
    .A0(DOUT_SRAM2),
    .A1(DOUT_SRAM10),
    .A2(_0079_),
    .A3(_0082_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit31.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG2 ));
 sg13g2_mux4_1 _0628_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit0.Q ),
    .A0(DOUT_SRAM3),
    .A1(DOUT_SRAM11),
    .A2(_0080_),
    .A3(_0081_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit1.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG3 ));
 sg13g2_mux4_1 _0629_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit2.Q ),
    .A0(DOUT_SRAM4),
    .A1(DOUT_SRAM12),
    .A2(_0080_),
    .A3(_0081_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit3.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG4 ));
 sg13g2_mux4_1 _0630_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit4.Q ),
    .A0(DOUT_SRAM5),
    .A1(DOUT_SRAM13),
    .A2(_0079_),
    .A3(_0082_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit5.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG5 ));
 sg13g2_mux4_1 _0631_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit6.Q ),
    .A0(DOUT_SRAM6),
    .A1(DOUT_SRAM14),
    .A2(_0078_),
    .A3(_0083_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit7.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG6 ));
 sg13g2_mux4_1 _0632_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit8.Q ),
    .A0(DOUT_SRAM7),
    .A1(DOUT_SRAM15),
    .A2(_0043_),
    .A3(_0084_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit9.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG7 ));
 sg13g2_mux4_1 _0633_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit10.Q ),
    .A0(DOUT_SRAM0),
    .A1(DOUT_SRAM8),
    .A2(_0043_),
    .A3(_0084_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit11.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb0 ));
 sg13g2_mux4_1 _0634_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit12.Q ),
    .A0(DOUT_SRAM1),
    .A1(DOUT_SRAM9),
    .A2(_0078_),
    .A3(_0083_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit13.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb1 ));
 sg13g2_mux4_1 _0635_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit14.Q ),
    .A0(DOUT_SRAM2),
    .A1(DOUT_SRAM10),
    .A2(_0079_),
    .A3(_0082_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit15.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb2 ));
 sg13g2_mux4_1 _0636_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit16.Q ),
    .A0(DOUT_SRAM3),
    .A1(DOUT_SRAM11),
    .A2(_0080_),
    .A3(_0081_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit17.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb3 ));
 sg13g2_mux4_1 _0637_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit18.Q ),
    .A0(DOUT_SRAM4),
    .A1(DOUT_SRAM12),
    .A2(_0080_),
    .A3(_0081_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit19.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb4 ));
 sg13g2_mux4_1 _0638_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit20.Q ),
    .A0(DOUT_SRAM5),
    .A1(DOUT_SRAM13),
    .A2(_0079_),
    .A3(_0082_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit21.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb5 ));
 sg13g2_mux4_1 _0639_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit22.Q ),
    .A0(DOUT_SRAM6),
    .A1(DOUT_SRAM14),
    .A2(_0078_),
    .A3(_0083_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit23.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb6 ));
 sg13g2_mux4_1 _0640_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit24.Q ),
    .A0(DOUT_SRAM7),
    .A1(DOUT_SRAM15),
    .A2(_0043_),
    .A3(_0084_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit25.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb7 ));
 sg13g2_mux4_1 _0641_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit26.Q ),
    .A0(DOUT_SRAM0),
    .A1(DOUT_SRAM12),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15 ),
    .A3(_0084_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit27.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG0 ));
 sg13g2_mux4_1 _0642_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit28.Q ),
    .A0(DOUT_SRAM1),
    .A1(DOUT_SRAM13),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14 ),
    .A3(_0083_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit29.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG1 ));
 sg13g2_mux4_1 _0643_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit30.Q ),
    .A0(DOUT_SRAM2),
    .A1(DOUT_SRAM14),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13 ),
    .A3(_0082_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit31.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG2 ));
 sg13g2_mux4_1 _0644_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit0.Q ),
    .A0(DOUT_SRAM3),
    .A1(DOUT_SRAM15),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12 ),
    .A3(_0081_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit1.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG3 ));
 sg13g2_mux4_1 _0645_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit30.Q ),
    .A0(Tile_X0Y1_N1END[3]),
    .A1(Tile_X0Y1_N4END[3]),
    .A2(_0074_),
    .A3(Tile_X0Y0_S4END[7]),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit31.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11 ));
 sg13g2_mux4_1 _0646_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit2.Q ),
    .A0(DOUT_SRAM4),
    .A1(DOUT_SRAM8),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11 ),
    .A3(_0080_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit3.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG4 ));
 sg13g2_mux4_1 _0647_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit28.Q ),
    .A0(Tile_X0Y1_N1END[2]),
    .A1(Tile_X0Y1_N4END[2]),
    .A2(_0067_),
    .A3(Tile_X0Y0_S4END[6]),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit29.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10 ));
 sg13g2_mux4_1 _0648_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit4.Q ),
    .A0(DOUT_SRAM5),
    .A1(DOUT_SRAM9),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10 ),
    .A3(_0079_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit5.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG5 ));
 sg13g2_mux4_1 _0649_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit26.Q ),
    .A0(Tile_X0Y1_N1END[1]),
    .A1(Tile_X0Y1_N4END[1]),
    .A2(_0060_),
    .A3(Tile_X0Y0_S4END[5]),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit27.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9 ));
 sg13g2_mux4_1 _0650_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit6.Q ),
    .A0(DOUT_SRAM6),
    .A1(DOUT_SRAM10),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9 ),
    .A3(_0078_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit7.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG6 ));
 sg13g2_mux4_1 _0651_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit24.Q ),
    .A0(Tile_X0Y1_N1END[0]),
    .A1(Tile_X0Y1_N4END[0]),
    .A2(_0088_),
    .A3(Tile_X0Y0_S4END[4]),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit25.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8 ));
 sg13g2_mux4_1 _0652_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit8.Q ),
    .A0(DOUT_SRAM7),
    .A1(DOUT_SRAM11),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8 ),
    .A3(_0043_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit9.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG7 ));
 sg13g2_mux4_1 _0653_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit22.Q ),
    .A0(Tile_X0Y1_N1END[3]),
    .A1(Tile_X0Y1_N4END[3]),
    .A2(_0074_),
    .A3(Tile_X0Y0_S4END[7]),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit23.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7 ));
 sg13g2_mux4_1 _0654_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit10.Q ),
    .A0(DOUT_SRAM4),
    .A1(DOUT_SRAM8),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7 ),
    .A3(_0084_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit11.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG8 ));
 sg13g2_mux4_1 _0655_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit20.Q ),
    .A0(Tile_X0Y1_N1END[2]),
    .A1(Tile_X0Y1_N4END[2]),
    .A2(_0067_),
    .A3(Tile_X0Y0_S4END[6]),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit21.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6 ));
 sg13g2_mux4_1 _0656_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit12.Q ),
    .A0(DOUT_SRAM5),
    .A1(DOUT_SRAM9),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6 ),
    .A3(_0083_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit13.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG9 ));
 sg13g2_mux4_1 _0657_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit18.Q ),
    .A0(Tile_X0Y1_N1END[1]),
    .A1(Tile_X0Y1_N4END[1]),
    .A2(_0060_),
    .A3(Tile_X0Y0_S4END[5]),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit19.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5 ));
 sg13g2_mux4_1 _0658_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit14.Q ),
    .A0(DOUT_SRAM6),
    .A1(DOUT_SRAM10),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5 ),
    .A3(_0082_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit15.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG10 ));
 sg13g2_mux4_1 _0659_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit16.Q ),
    .A0(Tile_X0Y1_N1END[0]),
    .A1(Tile_X0Y1_N4END[0]),
    .A2(_0088_),
    .A3(Tile_X0Y0_S4END[4]),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit17.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4 ));
 sg13g2_mux4_1 _0660_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit16.Q ),
    .A0(DOUT_SRAM7),
    .A1(DOUT_SRAM11),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4 ),
    .A3(_0081_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit17.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG11 ));
 sg13g2_mux4_1 _0661_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit14.Q ),
    .A0(Tile_X0Y1_N1END[3]),
    .A1(Tile_X0Y1_N4END[3]),
    .A2(_0074_),
    .A3(Tile_X0Y0_S4END[7]),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit15.Q ),
    .X(_0158_));
 sg13g2_mux4_1 _0662_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit18.Q ),
    .A0(DOUT_SRAM0),
    .A1(DOUT_SRAM12),
    .A2(_0158_),
    .A3(_0080_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit19.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG12 ));
 sg13g2_mux4_1 _0663_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit12.Q ),
    .A0(Tile_X0Y1_N1END[2]),
    .A1(Tile_X0Y1_N4END[2]),
    .A2(_0067_),
    .A3(Tile_X0Y0_S4END[6]),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit13.Q ),
    .X(_0159_));
 sg13g2_mux4_1 _0664_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit20.Q ),
    .A0(DOUT_SRAM1),
    .A1(DOUT_SRAM13),
    .A2(_0159_),
    .A3(_0079_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit21.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG13 ));
 sg13g2_mux4_1 _0665_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit10.Q ),
    .A0(Tile_X0Y1_N1END[1]),
    .A1(Tile_X0Y1_N4END[1]),
    .A2(_0060_),
    .A3(Tile_X0Y0_S4END[5]),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit11.Q ),
    .X(_0160_));
 sg13g2_mux4_1 _0666_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit22.Q ),
    .A0(DOUT_SRAM2),
    .A1(DOUT_SRAM14),
    .A2(_0160_),
    .A3(_0078_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit23.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG14 ));
 sg13g2_mux4_1 _0667_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit8.Q ),
    .A0(Tile_X0Y1_N1END[0]),
    .A1(Tile_X0Y1_N4END[0]),
    .A2(_0088_),
    .A3(Tile_X0Y0_S4END[4]),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit9.Q ),
    .X(_0161_));
 sg13g2_mux4_1 _0668_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit24.Q ),
    .A0(DOUT_SRAM3),
    .A1(DOUT_SRAM15),
    .A2(_0161_),
    .A3(_0043_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit25.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG15 ));
 sg13g2_mux4_1 _0669_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit26.Q ),
    .A0(Tile_X0Y1_N4END[0]),
    .A1(Tile_X0Y0_S4END[4]),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11 ),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit27.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG0 ));
 sg13g2_mux4_1 _0670_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit28.Q ),
    .A0(Tile_X0Y1_N4END[1]),
    .A1(Tile_X0Y0_S4END[5]),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10 ),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit29.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG1 ));
 sg13g2_mux4_1 _0671_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit30.Q ),
    .A0(Tile_X0Y1_N4END[2]),
    .A1(Tile_X0Y0_S4END[6]),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9 ),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit31.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG2 ));
 sg13g2_mux4_1 _0672_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit0.Q ),
    .A0(Tile_X0Y1_N4END[3]),
    .A1(Tile_X0Y0_S4END[7]),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8 ),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit1.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG3 ));
 sg13g2_mux4_1 _0673_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit3.Q ),
    .A0(DOUT_SRAM4),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11 ),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7 ),
    .A3(_0043_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit2.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG4 ));
 sg13g2_mux4_1 _0674_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit5.Q ),
    .A0(DOUT_SRAM5),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10 ),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6 ),
    .A3(_0078_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit4.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG5 ));
 sg13g2_mux4_1 _0675_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit6.Q ),
    .A0(DOUT_SRAM6),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5 ),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9 ),
    .A3(_0079_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit7.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG6 ));
 sg13g2_mux4_1 _0676_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit8.Q ),
    .A0(DOUT_SRAM7),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4 ),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8 ),
    .A3(_0080_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit9.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG7 ));
 sg13g2_mux4_1 _0677_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit11.Q ),
    .A0(DOUT_SRAM0),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7 ),
    .A2(_0158_),
    .A3(_0081_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit10.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG8 ));
 sg13g2_mux4_1 _0678_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit13.Q ),
    .A0(DOUT_SRAM1),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6 ),
    .A2(_0159_),
    .A3(_0082_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit12.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG9 ));
 sg13g2_mux4_1 _0679_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit15.Q ),
    .A0(DOUT_SRAM2),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5 ),
    .A2(_0160_),
    .A3(_0083_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit14.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG10 ));
 sg13g2_mux4_1 _0680_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit17.Q ),
    .A0(DOUT_SRAM3),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4 ),
    .A2(_0161_),
    .A3(_0084_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit16.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG11 ));
 sg13g2_nand3b_1 _0681_ (.B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit19.Q ),
    .C(_0043_),
    .Y(_0162_),
    .A_N(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit18.Q ));
 sg13g2_nor2b_1 _0682_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit18.Q ),
    .B_N(Tile_X0Y1_E2MID[0]),
    .Y(_0163_));
 sg13g2_a21oi_1 _0683_ (.A1(Tile_X0Y1_E2END[0]),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit18.Q ),
    .Y(_0164_),
    .B1(_0163_));
 sg13g2_o21ai_1 _0684_ (.B1(_0162_),
    .Y(ADDR_SRAM0),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit19.Q ),
    .A2(_0164_));
 sg13g2_nand3b_1 _0685_ (.B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit21.Q ),
    .C(_0078_),
    .Y(_0165_),
    .A_N(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit20.Q ));
 sg13g2_nor2b_1 _0686_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .B_N(Tile_X0Y1_E2MID[1]),
    .Y(_0166_));
 sg13g2_a21oi_1 _0687_ (.A1(Tile_X0Y1_E2END[1]),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .Y(_0167_),
    .B1(_0166_));
 sg13g2_o21ai_1 _0688_ (.B1(_0165_),
    .Y(ADDR_SRAM1),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit21.Q ),
    .A2(_0167_));
 sg13g2_nand3b_1 _0689_ (.B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit23.Q ),
    .C(_0079_),
    .Y(_0168_),
    .A_N(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit22.Q ));
 sg13g2_nor2b_1 _0690_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit22.Q ),
    .B_N(Tile_X0Y1_E2MID[2]),
    .Y(_0169_));
 sg13g2_a21oi_1 _0691_ (.A1(Tile_X0Y1_E2END[2]),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit22.Q ),
    .Y(_0170_),
    .B1(_0169_));
 sg13g2_o21ai_1 _0692_ (.B1(_0168_),
    .Y(ADDR_SRAM2),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit23.Q ),
    .A2(_0170_));
 sg13g2_nand3b_1 _0693_ (.B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit25.Q ),
    .C(_0080_),
    .Y(_0171_),
    .A_N(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit24.Q ));
 sg13g2_nor2_1 _0694_ (.A(_0000_),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit24.Q ),
    .Y(_0172_));
 sg13g2_a21oi_1 _0695_ (.A1(Tile_X0Y1_E2END[3]),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit24.Q ),
    .Y(_0173_),
    .B1(_0172_));
 sg13g2_o21ai_1 _0696_ (.B1(_0171_),
    .Y(ADDR_SRAM3),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit25.Q ),
    .A2(_0173_));
 sg13g2_nand3b_1 _0697_ (.B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit27.Q ),
    .C(_0081_),
    .Y(_0174_),
    .A_N(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit26.Q ));
 sg13g2_nor2b_1 _0698_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit26.Q ),
    .B_N(Tile_X0Y1_E2MID[4]),
    .Y(_0175_));
 sg13g2_a21oi_1 _0699_ (.A1(Tile_X0Y1_E2END[4]),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit26.Q ),
    .Y(_0176_),
    .B1(_0175_));
 sg13g2_o21ai_1 _0700_ (.B1(_0174_),
    .Y(ADDR_SRAM4),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit27.Q ),
    .A2(_0176_));
 sg13g2_mux4_1 _0701_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit28.Q ),
    .A0(Tile_X0Y1_EE4END[0]),
    .A1(Tile_X0Y1_EE4END[8]),
    .A2(Tile_X0Y1_E6END[0]),
    .A3(_0161_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit29.Q ),
    .X(DIN_SRAM0));
 sg13g2_mux4_1 _0702_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit30.Q ),
    .A0(Tile_X0Y1_EE4END[1]),
    .A1(Tile_X0Y1_EE4END[9]),
    .A2(Tile_X0Y1_E6END[1]),
    .A3(_0160_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit31.Q ),
    .X(DIN_SRAM1));
 sg13g2_mux4_1 _0703_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit0.Q ),
    .A0(Tile_X0Y1_EE4END[2]),
    .A1(Tile_X0Y1_EE4END[10]),
    .A2(Tile_X0Y1_E6END[2]),
    .A3(_0159_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit1.Q ),
    .X(DIN_SRAM2));
 sg13g2_mux4_1 _0704_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit2.Q ),
    .A0(Tile_X0Y1_EE4END[3]),
    .A1(Tile_X0Y1_EE4END[11]),
    .A2(Tile_X0Y1_E6END[3]),
    .A3(_0158_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit3.Q ),
    .X(DIN_SRAM3));
 sg13g2_mux4_1 _0705_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit4.Q ),
    .A0(Tile_X0Y1_EE4END[4]),
    .A1(Tile_X0Y1_EE4END[12]),
    .A2(Tile_X0Y1_E6END[4]),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit5.Q ),
    .X(DIN_SRAM4));
 sg13g2_mux4_1 _0706_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit6.Q ),
    .A0(Tile_X0Y1_EE4END[5]),
    .A1(Tile_X0Y1_EE4END[13]),
    .A2(Tile_X0Y1_E6END[5]),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit7.Q ),
    .X(DIN_SRAM5));
 sg13g2_mux4_1 _0707_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit8.Q ),
    .A0(Tile_X0Y1_EE4END[6]),
    .A1(Tile_X0Y1_EE4END[14]),
    .A2(Tile_X0Y1_E6END[6]),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit9.Q ),
    .X(DIN_SRAM6));
 sg13g2_mux4_1 _0708_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit10.Q ),
    .A0(Tile_X0Y1_EE4END[7]),
    .A1(Tile_X0Y1_EE4END[15]),
    .A2(Tile_X0Y1_E6END[7]),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit11.Q ),
    .X(DIN_SRAM7));
 sg13g2_mux4_1 _0709_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit12.Q ),
    .A0(Tile_X0Y1_EE4END[0]),
    .A1(Tile_X0Y1_EE4END[8]),
    .A2(Tile_X0Y1_E6END[8]),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit13.Q ),
    .X(DIN_SRAM8));
 sg13g2_mux4_1 _0710_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit14.Q ),
    .A0(Tile_X0Y1_EE4END[1]),
    .A1(Tile_X0Y1_EE4END[9]),
    .A2(Tile_X0Y1_E6END[9]),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit15.Q ),
    .X(DIN_SRAM9));
 sg13g2_mux4_1 _0711_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit16.Q ),
    .A0(Tile_X0Y1_EE4END[2]),
    .A1(Tile_X0Y1_EE4END[10]),
    .A2(Tile_X0Y1_E6END[10]),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit17.Q ),
    .X(DIN_SRAM10));
 sg13g2_mux4_1 _0712_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit18.Q ),
    .A0(Tile_X0Y1_EE4END[3]),
    .A1(Tile_X0Y1_EE4END[11]),
    .A2(Tile_X0Y1_E6END[11]),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit19.Q ),
    .X(DIN_SRAM11));
 sg13g2_mux4_1 _0713_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit20.Q ),
    .A0(Tile_X0Y1_E1END[0]),
    .A1(Tile_X0Y1_EE4END[4]),
    .A2(Tile_X0Y1_EE4END[12]),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit21.Q ),
    .X(DIN_SRAM12));
 sg13g2_mux4_1 _0714_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit22.Q ),
    .A0(Tile_X0Y1_E1END[1]),
    .A1(Tile_X0Y1_EE4END[5]),
    .A2(Tile_X0Y1_EE4END[13]),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit23.Q ),
    .X(DIN_SRAM13));
 sg13g2_mux4_1 _0715_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit24.Q ),
    .A0(Tile_X0Y1_E1END[2]),
    .A1(Tile_X0Y1_EE4END[6]),
    .A2(Tile_X0Y1_EE4END[14]),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit25.Q ),
    .X(DIN_SRAM14));
 sg13g2_mux4_1 _0716_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit26.Q ),
    .A0(Tile_X0Y1_E1END[3]),
    .A1(Tile_X0Y1_EE4END[7]),
    .A2(Tile_X0Y1_EE4END[15]),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit27.Q ),
    .X(DIN_SRAM15));
 sg13g2_mux4_1 _0717_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit28.Q ),
    .A0(Tile_X0Y1_EE4END[0]),
    .A1(Tile_X0Y1_EE4END[8]),
    .A2(Tile_X0Y1_E6END[0]),
    .A3(_0161_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit29.Q ),
    .X(BM_SRAM0));
 sg13g2_mux4_1 _0718_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit30.Q ),
    .A0(Tile_X0Y1_EE4END[1]),
    .A1(Tile_X0Y1_EE4END[9]),
    .A2(Tile_X0Y1_E6END[1]),
    .A3(_0160_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit31.Q ),
    .X(BM_SRAM1));
 sg13g2_mux4_1 _0719_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q ),
    .A0(Tile_X0Y1_EE4END[2]),
    .A1(Tile_X0Y1_EE4END[10]),
    .A2(Tile_X0Y1_E6END[2]),
    .A3(_0159_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit1.Q ),
    .X(BM_SRAM2));
 sg13g2_mux4_1 _0720_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit2.Q ),
    .A0(Tile_X0Y1_EE4END[3]),
    .A1(Tile_X0Y1_EE4END[11]),
    .A2(Tile_X0Y1_E6END[3]),
    .A3(_0158_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit3.Q ),
    .X(BM_SRAM3));
 sg13g2_mux4_1 _0721_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q ),
    .A0(Tile_X0Y1_EE4END[4]),
    .A1(Tile_X0Y1_EE4END[12]),
    .A2(Tile_X0Y1_E6END[4]),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit5.Q ),
    .X(BM_SRAM4));
 sg13g2_mux4_1 _0722_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit6.Q ),
    .A0(Tile_X0Y1_EE4END[5]),
    .A1(Tile_X0Y1_EE4END[13]),
    .A2(Tile_X0Y1_E6END[5]),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit7.Q ),
    .X(BM_SRAM5));
 sg13g2_mux4_1 _0723_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit8.Q ),
    .A0(Tile_X0Y1_EE4END[6]),
    .A1(Tile_X0Y1_EE4END[14]),
    .A2(Tile_X0Y1_E6END[6]),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit9.Q ),
    .X(BM_SRAM6));
 sg13g2_mux4_1 _0724_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit10.Q ),
    .A0(Tile_X0Y1_EE4END[7]),
    .A1(Tile_X0Y1_EE4END[15]),
    .A2(Tile_X0Y1_E6END[7]),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit11.Q ),
    .X(BM_SRAM7));
 sg13g2_mux4_1 _0725_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit12.Q ),
    .A0(Tile_X0Y1_EE4END[0]),
    .A1(Tile_X0Y1_EE4END[8]),
    .A2(Tile_X0Y1_E6END[8]),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit13.Q ),
    .X(BM_SRAM8));
 sg13g2_mux4_1 _0726_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit14.Q ),
    .A0(Tile_X0Y1_EE4END[1]),
    .A1(Tile_X0Y1_EE4END[9]),
    .A2(Tile_X0Y1_E6END[9]),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit15.Q ),
    .X(BM_SRAM9));
 sg13g2_mux4_1 _0727_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit16.Q ),
    .A0(Tile_X0Y1_EE4END[2]),
    .A1(Tile_X0Y1_EE4END[10]),
    .A2(Tile_X0Y1_E6END[10]),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit17.Q ),
    .X(BM_SRAM10));
 sg13g2_mux4_1 _0728_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit18.Q ),
    .A0(Tile_X0Y1_EE4END[3]),
    .A1(Tile_X0Y1_EE4END[11]),
    .A2(Tile_X0Y1_E6END[11]),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit19.Q ),
    .X(BM_SRAM11));
 sg13g2_mux4_1 _0729_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit20.Q ),
    .A0(Tile_X0Y1_E1END[0]),
    .A1(Tile_X0Y1_EE4END[4]),
    .A2(Tile_X0Y1_EE4END[12]),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit21.Q ),
    .X(BM_SRAM12));
 sg13g2_mux4_1 _0730_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit22.Q ),
    .A0(Tile_X0Y1_E1END[1]),
    .A1(Tile_X0Y1_EE4END[5]),
    .A2(Tile_X0Y1_EE4END[13]),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit23.Q ),
    .X(BM_SRAM13));
 sg13g2_mux4_1 _0731_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit24.Q ),
    .A0(Tile_X0Y1_E1END[2]),
    .A1(Tile_X0Y1_EE4END[6]),
    .A2(Tile_X0Y1_EE4END[14]),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit25.Q ),
    .X(BM_SRAM14));
 sg13g2_mux4_1 _0732_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit26.Q ),
    .A0(Tile_X0Y1_E1END[3]),
    .A1(Tile_X0Y1_EE4END[7]),
    .A2(Tile_X0Y1_EE4END[15]),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit27.Q ),
    .X(BM_SRAM15));
 sg13g2_o21ai_1 _0733_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit3.Q ),
    .Y(_0177_),
    .A1(Tile_X0Y1_E6END[8]),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit2.Q ));
 sg13g2_inv_1 _0734_ (.Y(_0178_),
    .A(_0177_));
 sg13g2_o21ai_1 _0735_ (.B1(_0178_),
    .Y(_0179_),
    .A1(_0019_),
    .A2(_0161_));
 sg13g2_mux2_1 _0736_ (.A0(Tile_X0Y1_E1END[0]),
    .A1(Tile_X0Y1_EE4END[0]),
    .S(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit2.Q ),
    .X(_0180_));
 sg13g2_a21oi_1 _0737_ (.A1(_0020_),
    .A2(_0180_),
    .Y(_0181_),
    .B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit4.Q ));
 sg13g2_nor2_1 _0738_ (.A(_0019_),
    .B(_0043_),
    .Y(_0182_));
 sg13g2_o21ai_1 _0739_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit3.Q ),
    .Y(_0183_),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit2.Q ),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12 ));
 sg13g2_mux2_1 _0740_ (.A0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4 ),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8 ),
    .S(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit2.Q ),
    .X(_0184_));
 sg13g2_o21ai_1 _0741_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit4.Q ),
    .Y(_0185_),
    .A1(_0182_),
    .A2(_0183_));
 sg13g2_a21oi_1 _0742_ (.A1(_0020_),
    .A2(_0184_),
    .Y(_0186_),
    .B1(_0185_));
 sg13g2_a21oi_1 _0743_ (.A1(_0179_),
    .A2(_0181_),
    .Y(\Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_8.A ),
    .B1(_0186_));
 sg13g2_o21ai_1 _0744_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit6.Q ),
    .Y(_0187_),
    .A1(Tile_X0Y1_E6END[9]),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit5.Q ));
 sg13g2_inv_1 _0745_ (.Y(_0188_),
    .A(_0187_));
 sg13g2_o21ai_1 _0746_ (.B1(_0188_),
    .Y(_0189_),
    .A1(_0021_),
    .A2(_0160_));
 sg13g2_mux2_1 _0747_ (.A0(Tile_X0Y1_E1END[1]),
    .A1(Tile_X0Y1_EE4END[1]),
    .S(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit5.Q ),
    .X(_0190_));
 sg13g2_a21oi_1 _0748_ (.A1(_0022_),
    .A2(_0190_),
    .Y(_0191_),
    .B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit7.Q ));
 sg13g2_nor2_1 _0749_ (.A(_0021_),
    .B(_0078_),
    .Y(_0192_));
 sg13g2_o21ai_1 _0750_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit6.Q ),
    .Y(_0193_),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit5.Q ),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13 ));
 sg13g2_mux2_1 _0751_ (.A0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5 ),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9 ),
    .S(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit5.Q ),
    .X(_0194_));
 sg13g2_o21ai_1 _0752_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit7.Q ),
    .Y(_0195_),
    .A1(_0192_),
    .A2(_0193_));
 sg13g2_a21oi_1 _0753_ (.A1(_0022_),
    .A2(_0194_),
    .Y(_0196_),
    .B1(_0195_));
 sg13g2_a21oi_1 _0754_ (.A1(_0189_),
    .A2(_0191_),
    .Y(\Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_9.A ),
    .B1(_0196_));
 sg13g2_o21ai_1 _0755_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit9.Q ),
    .Y(_0197_),
    .A1(Tile_X0Y1_E6END[10]),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q ));
 sg13g2_inv_1 _0756_ (.Y(_0198_),
    .A(_0197_));
 sg13g2_o21ai_1 _0757_ (.B1(_0198_),
    .Y(_0199_),
    .A1(_0023_),
    .A2(_0159_));
 sg13g2_mux2_1 _0758_ (.A0(Tile_X0Y1_E1END[2]),
    .A1(Tile_X0Y1_EE4END[2]),
    .S(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q ),
    .X(_0200_));
 sg13g2_a21oi_1 _0759_ (.A1(_0024_),
    .A2(_0200_),
    .Y(_0201_),
    .B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit10.Q ));
 sg13g2_nor2_1 _0760_ (.A(_0023_),
    .B(_0079_),
    .Y(_0202_));
 sg13g2_o21ai_1 _0761_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit9.Q ),
    .Y(_0203_),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q ),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14 ));
 sg13g2_mux2_1 _0762_ (.A0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6 ),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10 ),
    .S(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q ),
    .X(_0204_));
 sg13g2_o21ai_1 _0763_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit10.Q ),
    .Y(_0205_),
    .A1(_0202_),
    .A2(_0203_));
 sg13g2_a21oi_1 _0764_ (.A1(_0024_),
    .A2(_0204_),
    .Y(_0206_),
    .B1(_0205_));
 sg13g2_a21oi_1 _0765_ (.A1(_0199_),
    .A2(_0201_),
    .Y(\Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_10.A ),
    .B1(_0206_));
 sg13g2_o21ai_1 _0766_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit12.Q ),
    .Y(_0207_),
    .A1(Tile_X0Y1_E6END[11]),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q ));
 sg13g2_inv_1 _0767_ (.Y(_0208_),
    .A(_0207_));
 sg13g2_o21ai_1 _0768_ (.B1(_0208_),
    .Y(_0209_),
    .A1(_0025_),
    .A2(_0158_));
 sg13g2_mux2_1 _0769_ (.A0(Tile_X0Y1_E1END[3]),
    .A1(Tile_X0Y1_EE4END[3]),
    .S(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q ),
    .X(_0210_));
 sg13g2_a21oi_1 _0770_ (.A1(_0026_),
    .A2(_0210_),
    .Y(_0211_),
    .B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit13.Q ));
 sg13g2_nor2_1 _0771_ (.A(_0025_),
    .B(_0080_),
    .Y(_0212_));
 sg13g2_o21ai_1 _0772_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit12.Q ),
    .Y(_0213_),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q ),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15 ));
 sg13g2_mux2_1 _0773_ (.A0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7 ),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11 ),
    .S(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q ),
    .X(_0214_));
 sg13g2_o21ai_1 _0774_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit13.Q ),
    .Y(_0215_),
    .A1(_0212_),
    .A2(_0213_));
 sg13g2_a21oi_1 _0775_ (.A1(_0026_),
    .A2(_0214_),
    .Y(_0216_),
    .B1(_0215_));
 sg13g2_a21oi_1 _0776_ (.A1(_0209_),
    .A2(_0211_),
    .Y(\Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_11.A ),
    .B1(_0216_));
 sg13g2_o21ai_1 _0777_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit7.Q ),
    .Y(_0217_),
    .A1(Tile_X0Y1_E6END[4]),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q ));
 sg13g2_inv_1 _0778_ (.Y(_0218_),
    .A(_0217_));
 sg13g2_o21ai_1 _0779_ (.B1(_0218_),
    .Y(_0219_),
    .A1(_0027_),
    .A2(_0161_));
 sg13g2_mux2_1 _0780_ (.A0(Tile_X0Y1_E1END[0]),
    .A1(Tile_X0Y1_EE4END[12]),
    .S(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q ),
    .X(_0220_));
 sg13g2_a21oi_1 _0781_ (.A1(_0028_),
    .A2(_0220_),
    .Y(_0221_),
    .B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit8.Q ));
 sg13g2_nor2_1 _0782_ (.A(_0027_),
    .B(_0081_),
    .Y(_0222_));
 sg13g2_o21ai_1 _0783_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit7.Q ),
    .Y(_0223_),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q ),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12 ));
 sg13g2_mux2_1 _0784_ (.A0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4 ),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8 ),
    .S(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q ),
    .X(_0224_));
 sg13g2_o21ai_1 _0785_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit8.Q ),
    .Y(_0225_),
    .A1(_0222_),
    .A2(_0223_));
 sg13g2_a21oi_1 _0786_ (.A1(_0028_),
    .A2(_0224_),
    .Y(_0226_),
    .B1(_0225_));
 sg13g2_a21oi_1 _0787_ (.A1(_0219_),
    .A2(_0221_),
    .Y(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG0 ),
    .B1(_0226_));
 sg13g2_o21ai_1 _0788_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q ),
    .Y(_0227_),
    .A1(Tile_X0Y1_E6END[5]),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q ));
 sg13g2_inv_1 _0789_ (.Y(_0228_),
    .A(_0227_));
 sg13g2_o21ai_1 _0790_ (.B1(_0228_),
    .Y(_0229_),
    .A1(_0029_),
    .A2(_0160_));
 sg13g2_mux2_1 _0791_ (.A0(Tile_X0Y1_E1END[1]),
    .A1(Tile_X0Y1_EE4END[13]),
    .S(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q ),
    .X(_0230_));
 sg13g2_a21oi_1 _0792_ (.A1(_0030_),
    .A2(_0230_),
    .Y(_0231_),
    .B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit11.Q ));
 sg13g2_nor2_1 _0793_ (.A(_0029_),
    .B(_0082_),
    .Y(_0232_));
 sg13g2_o21ai_1 _0794_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q ),
    .Y(_0233_),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q ),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13 ));
 sg13g2_mux2_1 _0795_ (.A0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5 ),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9 ),
    .S(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q ),
    .X(_0234_));
 sg13g2_o21ai_1 _0796_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit11.Q ),
    .Y(_0235_),
    .A1(_0232_),
    .A2(_0233_));
 sg13g2_a21oi_1 _0797_ (.A1(_0030_),
    .A2(_0234_),
    .Y(_0236_),
    .B1(_0235_));
 sg13g2_a21oi_1 _0798_ (.A1(_0229_),
    .A2(_0231_),
    .Y(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG1 ),
    .B1(_0236_));
 sg13g2_o21ai_1 _0799_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q ),
    .Y(_0237_),
    .A1(Tile_X0Y1_E6END[6]),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q ));
 sg13g2_inv_1 _0800_ (.Y(_0238_),
    .A(_0237_));
 sg13g2_o21ai_1 _0801_ (.B1(_0238_),
    .Y(_0239_),
    .A1(_0031_),
    .A2(_0159_));
 sg13g2_mux2_1 _0802_ (.A0(Tile_X0Y1_E1END[2]),
    .A1(Tile_X0Y1_EE4END[14]),
    .S(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q ),
    .X(_0240_));
 sg13g2_a21oi_1 _0803_ (.A1(_0032_),
    .A2(_0240_),
    .Y(_0241_),
    .B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit14.Q ));
 sg13g2_nor2_1 _0804_ (.A(_0031_),
    .B(_0083_),
    .Y(_0242_));
 sg13g2_o21ai_1 _0805_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q ),
    .Y(_0243_),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q ),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14 ));
 sg13g2_mux2_1 _0806_ (.A0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6 ),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10 ),
    .S(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q ),
    .X(_0244_));
 sg13g2_o21ai_1 _0807_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit14.Q ),
    .Y(_0245_),
    .A1(_0242_),
    .A2(_0243_));
 sg13g2_a21oi_1 _0808_ (.A1(_0032_),
    .A2(_0244_),
    .Y(_0246_),
    .B1(_0245_));
 sg13g2_a21oi_1 _0809_ (.A1(_0239_),
    .A2(_0241_),
    .Y(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG2 ),
    .B1(_0246_));
 sg13g2_o21ai_1 _0810_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q ),
    .Y(_0247_),
    .A1(Tile_X0Y1_E6END[7]),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q ));
 sg13g2_inv_1 _0811_ (.Y(_0248_),
    .A(_0247_));
 sg13g2_o21ai_1 _0812_ (.B1(_0248_),
    .Y(_0249_),
    .A1(_0033_),
    .A2(_0158_));
 sg13g2_mux2_1 _0813_ (.A0(Tile_X0Y1_E1END[3]),
    .A1(Tile_X0Y1_EE4END[15]),
    .S(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q ),
    .X(_0250_));
 sg13g2_a21oi_1 _0814_ (.A1(_0034_),
    .A2(_0250_),
    .Y(_0251_),
    .B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit17.Q ));
 sg13g2_nor2_1 _0815_ (.A(_0033_),
    .B(_0084_),
    .Y(_0252_));
 sg13g2_o21ai_1 _0816_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q ),
    .Y(_0253_),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q ),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15 ));
 sg13g2_mux2_1 _0817_ (.A0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7 ),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11 ),
    .S(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q ),
    .X(_0254_));
 sg13g2_o21ai_1 _0818_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit17.Q ),
    .Y(_0255_),
    .A1(_0252_),
    .A2(_0253_));
 sg13g2_a21oi_1 _0819_ (.A1(_0034_),
    .A2(_0254_),
    .Y(_0256_),
    .B1(_0255_));
 sg13g2_a21oi_1 _0820_ (.A1(_0249_),
    .A2(_0251_),
    .Y(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG3 ),
    .B1(_0256_));
 sg13g2_nor2b_1 _0821_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q ),
    .B_N(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .Y(_0257_));
 sg13g2_nand2b_1 _0822_ (.Y(_0258_),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q ),
    .A_N(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q ));
 sg13g2_nand2_1 _0823_ (.Y(_0259_),
    .A(Tile_X0Y1_N2END[2]),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q ));
 sg13g2_or2_1 _0824_ (.X(_0260_),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q ),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q ));
 sg13g2_a21oi_1 _0825_ (.A1(Tile_X0Y1_N2MID[6]),
    .A2(_0035_),
    .Y(_0261_),
    .B1(_0260_));
 sg13g2_nand2_1 _0826_ (.Y(_0262_),
    .A(Tile_X0Y1_E2END[1]),
    .B(_0035_));
 sg13g2_nand2_1 _0827_ (.Y(_0263_),
    .A(Tile_X0Y1_E2END[2]),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q ));
 sg13g2_nand4_1 _0828_ (.B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q ),
    .C(_0262_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .Y(_0264_),
    .D(_0263_));
 sg13g2_a21oi_1 _0829_ (.A1(Tile_X0Y1_E2MID[6]),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .Y(_0265_),
    .B1(_0258_));
 sg13g2_o21ai_1 _0830_ (.B1(_0265_),
    .Y(_0266_),
    .A1(_0000_),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q ));
 sg13g2_and2_1 _0831_ (.A(Tile_X0Y1_E2MID[0]),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .X(_0267_));
 sg13g2_a21oi_1 _0832_ (.A1(Tile_X0Y1_N2END[3]),
    .A2(_0035_),
    .Y(_0268_),
    .B1(_0267_));
 sg13g2_a22oi_1 _0833_ (.Y(_0269_),
    .B1(_0268_),
    .B2(_0257_),
    .A2(_0261_),
    .A1(_0259_));
 sg13g2_nand3_1 _0834_ (.B(_0266_),
    .C(_0269_),
    .A(_0264_),
    .Y(_0270_));
 sg13g2_nand2b_1 _0835_ (.Y(_0271_),
    .B(_0257_),
    .A_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG0 ));
 sg13g2_or3_1 _0836_ (.A(Tile_X0Y1_E2END[4]),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .C(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q ),
    .X(_0272_));
 sg13g2_or2_1 _0837_ (.X(_0273_),
    .B(_0258_),
    .A(Tile_X0Y0_S2MID[3]));
 sg13g2_nand4_1 _0838_ (.B(_0271_),
    .C(_0272_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .Y(_0274_),
    .D(_0273_));
 sg13g2_nand2b_1 _0839_ (.Y(_0275_),
    .B(Tile_X0Y1_E2END[5]),
    .A_N(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q ));
 sg13g2_nor3_1 _0840_ (.A(Tile_X0Y1_E2END[3]),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .C(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q ),
    .Y(_0276_));
 sg13g2_a221oi_1 _0841_ (.B2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .C1(_0276_),
    .B1(_0275_),
    .A1(_0002_),
    .Y(_0277_),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q ));
 sg13g2_a21oi_1 _0842_ (.A1(_0035_),
    .A2(_0277_),
    .Y(_0278_),
    .B1(_0036_));
 sg13g2_a22oi_1 _0843_ (.Y(WEN_SRAM),
    .B1(_0274_),
    .B2(_0278_),
    .A2(_0270_),
    .A1(_0036_));
 sg13g2_mux4_1 _0844_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .A0(Tile_X0Y1_N2END[3]),
    .A1(Tile_X0Y1_E2MID[0]),
    .A2(Tile_X0Y1_E2END[1]),
    .A3(Tile_X0Y1_E2END[2]),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .X(_0279_));
 sg13g2_nand2_1 _0845_ (.Y(_0280_),
    .A(Tile_X0Y1_N2END[2]),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q ));
 sg13g2_nor2b_1 _0846_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .B_N(Tile_X0Y1_N2MID[6]),
    .Y(_0281_));
 sg13g2_nor3_1 _0847_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .C(_0281_),
    .Y(_0282_));
 sg13g2_nand2_1 _0848_ (.Y(_0283_),
    .A(_0037_),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q ));
 sg13g2_nand2b_1 _0849_ (.Y(_0284_),
    .B(Tile_X0Y1_E2MID[3]),
    .A_N(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q ));
 sg13g2_a21oi_1 _0850_ (.A1(Tile_X0Y1_E2MID[6]),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .Y(_0285_),
    .B1(_0283_));
 sg13g2_a22oi_1 _0851_ (.Y(_0286_),
    .B1(_0284_),
    .B2(_0285_),
    .A2(_0282_),
    .A1(_0280_));
 sg13g2_o21ai_1 _0852_ (.B1(_0286_),
    .Y(_0287_),
    .A1(_0037_),
    .A2(_0279_));
 sg13g2_nor3_1 _0853_ (.A(_0037_),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .C(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG0 ),
    .Y(_0288_));
 sg13g2_nor3_1 _0854_ (.A(Tile_X0Y1_E2END[4]),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .C(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .Y(_0289_));
 sg13g2_o21ai_1 _0855_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .Y(_0290_),
    .A1(Tile_X0Y0_S2MID[3]),
    .A2(_0283_));
 sg13g2_nor3_1 _0856_ (.A(_0288_),
    .B(_0289_),
    .C(_0290_),
    .Y(_0291_));
 sg13g2_a21oi_1 _0857_ (.A1(_0001_),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .Y(_0292_),
    .B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q ));
 sg13g2_a21oi_1 _0858_ (.A1(Tile_X0Y0_S2MID[2]),
    .A2(_0037_),
    .Y(_0293_),
    .B1(_0292_));
 sg13g2_nor3_1 _0859_ (.A(Tile_X0Y1_E2END[3]),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .C(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .Y(_0294_));
 sg13g2_nor3_1 _0860_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .B(_0293_),
    .C(_0294_),
    .Y(_0295_));
 sg13g2_o21ai_1 _0861_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit7.Q ),
    .Y(_0296_),
    .A1(_0291_),
    .A2(_0295_));
 sg13g2_o21ai_1 _0862_ (.B1(_0296_),
    .Y(REN_SRAM),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit7.Q ),
    .A2(_0287_));
 sg13g2_dlhq_1 _0863_ (.D(Tile_X0Y0_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit31.Q ));
 sg13g2_dlhq_1 _0864_ (.D(Tile_X0Y0_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit30.Q ));
 sg13g2_dlhq_1 _0865_ (.D(Tile_X0Y0_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit29.Q ));
 sg13g2_dlhq_1 _0866_ (.D(Tile_X0Y0_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit28.Q ));
 sg13g2_dlhq_1 _0867_ (.D(Tile_X0Y0_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit27.Q ));
 sg13g2_dlhq_1 _0868_ (.D(Tile_X0Y0_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_dlhq_1 _0869_ (.D(Tile_X0Y0_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit25.Q ));
 sg13g2_dlhq_1 _0870_ (.D(Tile_X0Y0_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_dlhq_1 _0871_ (.D(Tile_X0Y0_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit23.Q ));
 sg13g2_dlhq_1 _0872_ (.D(Tile_X0Y0_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit22.Q ));
 sg13g2_dlhq_1 _0873_ (.D(Tile_X0Y0_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit21.Q ));
 sg13g2_dlhq_1 _0874_ (.D(Tile_X0Y0_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit20.Q ));
 sg13g2_dlhq_1 _0875_ (.D(Tile_X0Y0_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit19.Q ));
 sg13g2_dlhq_1 _0876_ (.D(Tile_X0Y0_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit18.Q ));
 sg13g2_dlhq_1 _0877_ (.D(Tile_X0Y0_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit17.Q ));
 sg13g2_dlhq_1 _0878_ (.D(Tile_X0Y0_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit16.Q ));
 sg13g2_dlhq_1 _0879_ (.D(Tile_X0Y0_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit15.Q ));
 sg13g2_dlhq_1 _0880_ (.D(Tile_X0Y0_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit14.Q ));
 sg13g2_dlhq_1 _0881_ (.D(Tile_X0Y0_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit13.Q ));
 sg13g2_dlhq_1 _0882_ (.D(Tile_X0Y0_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit12.Q ));
 sg13g2_dlhq_1 _0883_ (.D(Tile_X0Y0_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit11.Q ));
 sg13g2_dlhq_1 _0884_ (.D(Tile_X0Y0_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit10.Q ));
 sg13g2_dlhq_1 _0885_ (.D(Tile_X0Y0_FrameData[9]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit9.Q ));
 sg13g2_dlhq_1 _0886_ (.D(Tile_X0Y0_FrameData[8]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit8.Q ));
 sg13g2_dlhq_1 _0887_ (.D(Tile_X0Y0_FrameData[7]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit7.Q ));
 sg13g2_dlhq_1 _0888_ (.D(Tile_X0Y0_FrameData[6]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit6.Q ));
 sg13g2_dlhq_1 _0889_ (.D(Tile_X0Y0_FrameData[5]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit5.Q ));
 sg13g2_dlhq_1 _0890_ (.D(Tile_X0Y0_FrameData[4]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit4.Q ));
 sg13g2_dlhq_1 _0891_ (.D(Tile_X0Y0_FrameData[3]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit3.Q ));
 sg13g2_dlhq_1 _0892_ (.D(Tile_X0Y0_FrameData[2]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit2.Q ));
 sg13g2_dlhq_1 _0893_ (.D(Tile_X0Y0_FrameData[1]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit1.Q ));
 sg13g2_dlhq_1 _0894_ (.D(Tile_X0Y0_FrameData[0]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit0.Q ));
 sg13g2_dlhq_1 _0895_ (.D(Tile_X0Y0_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit31.Q ));
 sg13g2_dlhq_1 _0896_ (.D(Tile_X0Y0_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit30.Q ));
 sg13g2_dlhq_1 _0897_ (.D(Tile_X0Y0_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit29.Q ));
 sg13g2_dlhq_1 _0898_ (.D(Tile_X0Y0_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit28.Q ));
 sg13g2_dlhq_1 _0899_ (.D(Tile_X0Y0_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit27.Q ));
 sg13g2_dlhq_1 _0900_ (.D(Tile_X0Y0_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit26.Q ));
 sg13g2_dlhq_1 _0901_ (.D(Tile_X0Y0_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit25.Q ));
 sg13g2_dlhq_1 _0902_ (.D(Tile_X0Y0_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit24.Q ));
 sg13g2_dlhq_1 _0903_ (.D(Tile_X0Y0_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit23.Q ));
 sg13g2_dlhq_1 _0904_ (.D(Tile_X0Y0_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit22.Q ));
 sg13g2_dlhq_1 _0905_ (.D(Tile_X0Y0_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit21.Q ));
 sg13g2_dlhq_1 _0906_ (.D(Tile_X0Y0_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit20.Q ));
 sg13g2_dlhq_1 _0907_ (.D(Tile_X0Y0_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit19.Q ));
 sg13g2_dlhq_1 _0908_ (.D(Tile_X0Y0_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit18.Q ));
 sg13g2_dlhq_1 _0909_ (.D(Tile_X0Y0_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit17.Q ));
 sg13g2_dlhq_1 _0910_ (.D(Tile_X0Y0_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit16.Q ));
 sg13g2_dlhq_1 _0911_ (.D(Tile_X0Y0_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit15.Q ));
 sg13g2_dlhq_1 _0912_ (.D(Tile_X0Y0_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit14.Q ));
 sg13g2_dlhq_1 _0913_ (.D(Tile_X0Y0_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit13.Q ));
 sg13g2_dlhq_1 _0914_ (.D(Tile_X0Y0_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit12.Q ));
 sg13g2_dlhq_1 _0915_ (.D(Tile_X0Y0_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit11.Q ));
 sg13g2_dlhq_1 _0916_ (.D(Tile_X0Y0_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit10.Q ));
 sg13g2_dlhq_1 _0917_ (.D(Tile_X0Y0_FrameData[9]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit9.Q ));
 sg13g2_dlhq_1 _0918_ (.D(Tile_X0Y0_FrameData[8]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit8.Q ));
 sg13g2_dlhq_1 _0919_ (.D(Tile_X0Y0_FrameData[7]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit7.Q ));
 sg13g2_dlhq_1 _0920_ (.D(Tile_X0Y0_FrameData[6]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit6.Q ));
 sg13g2_dlhq_1 _0921_ (.D(Tile_X0Y0_FrameData[5]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit5.Q ));
 sg13g2_dlhq_1 _0922_ (.D(Tile_X0Y0_FrameData[4]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit4.Q ));
 sg13g2_dlhq_1 _0923_ (.D(Tile_X0Y0_FrameData[3]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit3.Q ));
 sg13g2_dlhq_1 _0924_ (.D(Tile_X0Y0_FrameData[2]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit2.Q ));
 sg13g2_dlhq_1 _0925_ (.D(Tile_X0Y0_FrameData[1]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit1.Q ));
 sg13g2_dlhq_1 _0926_ (.D(Tile_X0Y0_FrameData[0]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit0.Q ));
 sg13g2_dlhq_1 _0927_ (.D(Tile_X0Y0_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit31.Q ));
 sg13g2_dlhq_1 _0928_ (.D(Tile_X0Y0_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit30.Q ));
 sg13g2_dlhq_1 _0929_ (.D(Tile_X0Y0_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit29.Q ));
 sg13g2_dlhq_1 _0930_ (.D(Tile_X0Y0_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit28.Q ));
 sg13g2_dlhq_1 _0931_ (.D(Tile_X0Y0_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit27.Q ));
 sg13g2_dlhq_1 _0932_ (.D(Tile_X0Y0_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit26.Q ));
 sg13g2_dlhq_1 _0933_ (.D(Tile_X0Y0_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit25.Q ));
 sg13g2_dlhq_1 _0934_ (.D(Tile_X0Y0_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit24.Q ));
 sg13g2_dlhq_1 _0935_ (.D(Tile_X0Y0_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit23.Q ));
 sg13g2_dlhq_1 _0936_ (.D(Tile_X0Y0_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit22.Q ));
 sg13g2_dlhq_1 _0937_ (.D(Tile_X0Y0_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit21.Q ));
 sg13g2_dlhq_1 _0938_ (.D(Tile_X0Y0_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit20.Q ));
 sg13g2_dlhq_1 _0939_ (.D(Tile_X0Y0_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit19.Q ));
 sg13g2_dlhq_1 _0940_ (.D(Tile_X0Y0_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit18.Q ));
 sg13g2_dlhq_1 _0941_ (.D(Tile_X0Y0_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit17.Q ));
 sg13g2_dlhq_1 _0942_ (.D(Tile_X0Y0_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit16.Q ));
 sg13g2_dlhq_1 _0943_ (.D(Tile_X0Y0_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit15.Q ));
 sg13g2_dlhq_1 _0944_ (.D(Tile_X0Y0_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit14.Q ));
 sg13g2_dlhq_1 _0945_ (.D(Tile_X0Y0_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit13.Q ));
 sg13g2_dlhq_1 _0946_ (.D(Tile_X0Y0_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit12.Q ));
 sg13g2_dlhq_1 _0947_ (.D(Tile_X0Y0_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit11.Q ));
 sg13g2_dlhq_1 _0948_ (.D(Tile_X0Y0_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit10.Q ));
 sg13g2_dlhq_1 _0949_ (.D(Tile_X0Y0_FrameData[9]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit9.Q ));
 sg13g2_dlhq_1 _0950_ (.D(Tile_X0Y0_FrameData[8]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit8.Q ));
 sg13g2_dlhq_1 _0951_ (.D(Tile_X0Y0_FrameData[7]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit7.Q ));
 sg13g2_dlhq_1 _0952_ (.D(Tile_X0Y0_FrameData[6]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit6.Q ));
 sg13g2_dlhq_1 _0953_ (.D(Tile_X0Y0_FrameData[5]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit5.Q ));
 sg13g2_dlhq_1 _0954_ (.D(Tile_X0Y0_FrameData[4]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit4.Q ));
 sg13g2_dlhq_1 _0955_ (.D(Tile_X0Y0_FrameData[3]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit3.Q ));
 sg13g2_dlhq_1 _0956_ (.D(Tile_X0Y0_FrameData[2]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit2.Q ));
 sg13g2_dlhq_1 _0957_ (.D(Tile_X0Y0_FrameData[1]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit1.Q ));
 sg13g2_dlhq_1 _0958_ (.D(Tile_X0Y0_FrameData[0]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit0.Q ));
 sg13g2_dlhq_1 _0959_ (.D(Tile_X0Y0_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit31.Q ));
 sg13g2_dlhq_1 _0960_ (.D(Tile_X0Y0_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit30.Q ));
 sg13g2_dlhq_1 _0961_ (.D(Tile_X0Y0_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit29.Q ));
 sg13g2_dlhq_1 _0962_ (.D(Tile_X0Y0_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit28.Q ));
 sg13g2_dlhq_1 _0963_ (.D(Tile_X0Y0_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit27.Q ));
 sg13g2_dlhq_1 _0964_ (.D(Tile_X0Y0_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit26.Q ));
 sg13g2_dlhq_1 _0965_ (.D(Tile_X0Y0_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit25.Q ));
 sg13g2_dlhq_1 _0966_ (.D(Tile_X0Y0_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit24.Q ));
 sg13g2_dlhq_1 _0967_ (.D(Tile_X0Y0_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit23.Q ));
 sg13g2_dlhq_1 _0968_ (.D(Tile_X0Y0_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit22.Q ));
 sg13g2_dlhq_1 _0969_ (.D(Tile_X0Y0_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit21.Q ));
 sg13g2_dlhq_1 _0970_ (.D(Tile_X0Y0_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit20.Q ));
 sg13g2_dlhq_1 _0971_ (.D(Tile_X0Y0_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit19.Q ));
 sg13g2_dlhq_1 _0972_ (.D(Tile_X0Y0_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit18.Q ));
 sg13g2_dlhq_1 _0973_ (.D(Tile_X0Y0_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit17.Q ));
 sg13g2_dlhq_1 _0974_ (.D(Tile_X0Y0_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit16.Q ));
 sg13g2_dlhq_1 _0975_ (.D(Tile_X0Y0_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit15.Q ));
 sg13g2_dlhq_1 _0976_ (.D(Tile_X0Y0_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit14.Q ));
 sg13g2_dlhq_1 _0977_ (.D(Tile_X0Y0_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit13.Q ));
 sg13g2_dlhq_1 _0978_ (.D(Tile_X0Y0_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit12.Q ));
 sg13g2_dlhq_1 _0979_ (.D(Tile_X0Y0_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit11.Q ));
 sg13g2_dlhq_1 _0980_ (.D(Tile_X0Y0_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit10.Q ));
 sg13g2_dlhq_1 _0981_ (.D(Tile_X0Y0_FrameData[9]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit9.Q ));
 sg13g2_dlhq_1 _0982_ (.D(Tile_X0Y0_FrameData[8]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit8.Q ));
 sg13g2_dlhq_1 _0983_ (.D(Tile_X0Y0_FrameData[7]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit7.Q ));
 sg13g2_dlhq_1 _0984_ (.D(Tile_X0Y0_FrameData[6]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit6.Q ));
 sg13g2_dlhq_1 _0985_ (.D(Tile_X0Y0_FrameData[5]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit5.Q ));
 sg13g2_dlhq_1 _0986_ (.D(Tile_X0Y0_FrameData[4]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit4.Q ));
 sg13g2_dlhq_1 _0987_ (.D(Tile_X0Y0_FrameData[3]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit3.Q ));
 sg13g2_dlhq_1 _0988_ (.D(Tile_X0Y0_FrameData[2]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit2.Q ));
 sg13g2_dlhq_1 _0989_ (.D(Tile_X0Y0_FrameData[1]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit1.Q ));
 sg13g2_dlhq_1 _0990_ (.D(Tile_X0Y0_FrameData[0]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit0.Q ));
 sg13g2_dlhq_1 _0991_ (.D(Tile_X0Y0_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit31.Q ));
 sg13g2_dlhq_1 _0992_ (.D(Tile_X0Y0_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit30.Q ));
 sg13g2_dlhq_1 _0993_ (.D(Tile_X0Y0_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit29.Q ));
 sg13g2_dlhq_1 _0994_ (.D(Tile_X0Y0_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit28.Q ));
 sg13g2_dlhq_1 _0995_ (.D(Tile_X0Y0_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit27.Q ));
 sg13g2_dlhq_1 _0996_ (.D(Tile_X0Y0_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit26.Q ));
 sg13g2_dlhq_1 _0997_ (.D(Tile_X0Y0_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit25.Q ));
 sg13g2_dlhq_1 _0998_ (.D(Tile_X0Y0_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit24.Q ));
 sg13g2_dlhq_1 _0999_ (.D(Tile_X0Y0_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit23.Q ));
 sg13g2_dlhq_1 _1000_ (.D(Tile_X0Y0_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit22.Q ));
 sg13g2_dlhq_1 _1001_ (.D(Tile_X0Y0_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit21.Q ));
 sg13g2_dlhq_1 _1002_ (.D(Tile_X0Y0_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit20.Q ));
 sg13g2_dlhq_1 _1003_ (.D(Tile_X0Y0_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit19.Q ));
 sg13g2_dlhq_1 _1004_ (.D(Tile_X0Y0_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit18.Q ));
 sg13g2_dlhq_1 _1005_ (.D(Tile_X0Y0_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit17.Q ));
 sg13g2_dlhq_1 _1006_ (.D(Tile_X0Y0_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit16.Q ));
 sg13g2_dlhq_1 _1007_ (.D(Tile_X0Y0_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit15.Q ));
 sg13g2_dlhq_1 _1008_ (.D(Tile_X0Y0_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit14.Q ));
 sg13g2_dlhq_1 _1009_ (.D(Tile_X0Y0_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit13.Q ));
 sg13g2_dlhq_1 _1010_ (.D(Tile_X0Y0_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit12.Q ));
 sg13g2_dlhq_1 _1011_ (.D(Tile_X0Y0_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit11.Q ));
 sg13g2_dlhq_1 _1012_ (.D(Tile_X0Y0_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit10.Q ));
 sg13g2_dlhq_1 _1013_ (.D(Tile_X0Y0_FrameData[9]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit9.Q ));
 sg13g2_dlhq_1 _1014_ (.D(Tile_X0Y0_FrameData[8]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit8.Q ));
 sg13g2_dlhq_1 _1015_ (.D(Tile_X0Y0_FrameData[7]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit7.Q ));
 sg13g2_dlhq_1 _1016_ (.D(Tile_X0Y0_FrameData[6]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit6.Q ));
 sg13g2_dlhq_1 _1017_ (.D(Tile_X0Y0_FrameData[5]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit5.Q ));
 sg13g2_dlhq_1 _1018_ (.D(Tile_X0Y0_FrameData[4]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit4.Q ));
 sg13g2_dlhq_1 _1019_ (.D(Tile_X0Y0_FrameData[3]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit3.Q ));
 sg13g2_dlhq_1 _1020_ (.D(Tile_X0Y0_FrameData[2]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit2.Q ));
 sg13g2_dlhq_1 _1021_ (.D(Tile_X0Y0_FrameData[1]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit1.Q ));
 sg13g2_dlhq_1 _1022_ (.D(Tile_X0Y0_FrameData[0]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit0.Q ));
 sg13g2_dlhq_1 _1023_ (.D(Tile_X0Y0_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit31.Q ));
 sg13g2_dlhq_1 _1024_ (.D(Tile_X0Y0_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit30.Q ));
 sg13g2_dlhq_1 _1025_ (.D(Tile_X0Y0_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit29.Q ));
 sg13g2_dlhq_1 _1026_ (.D(Tile_X0Y0_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit28.Q ));
 sg13g2_dlhq_1 _1027_ (.D(Tile_X0Y0_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit27.Q ));
 sg13g2_dlhq_1 _1028_ (.D(Tile_X0Y0_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit26.Q ));
 sg13g2_dlhq_1 _1029_ (.D(Tile_X0Y0_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit25.Q ));
 sg13g2_dlhq_1 _1030_ (.D(Tile_X0Y0_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit24.Q ));
 sg13g2_dlhq_1 _1031_ (.D(Tile_X0Y0_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit23.Q ));
 sg13g2_dlhq_1 _1032_ (.D(Tile_X0Y0_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit22.Q ));
 sg13g2_dlhq_1 _1033_ (.D(Tile_X0Y0_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit21.Q ));
 sg13g2_dlhq_1 _1034_ (.D(Tile_X0Y0_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit20.Q ));
 sg13g2_dlhq_1 _1035_ (.D(Tile_X0Y0_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit19.Q ));
 sg13g2_dlhq_1 _1036_ (.D(Tile_X0Y0_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit18.Q ));
 sg13g2_dlhq_1 _1037_ (.D(Tile_X0Y0_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit17.Q ));
 sg13g2_dlhq_1 _1038_ (.D(Tile_X0Y0_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit16.Q ));
 sg13g2_dlhq_1 _1039_ (.D(Tile_X0Y0_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit15.Q ));
 sg13g2_dlhq_1 _1040_ (.D(Tile_X0Y0_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit14.Q ));
 sg13g2_dlhq_1 _1041_ (.D(Tile_X0Y0_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit13.Q ));
 sg13g2_dlhq_1 _1042_ (.D(Tile_X0Y0_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit12.Q ));
 sg13g2_dlhq_1 _1043_ (.D(Tile_X0Y0_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit11.Q ));
 sg13g2_dlhq_1 _1044_ (.D(Tile_X0Y0_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit10.Q ));
 sg13g2_dlhq_1 _1045_ (.D(Tile_X0Y0_FrameData[9]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit9.Q ));
 sg13g2_dlhq_1 _1046_ (.D(Tile_X0Y0_FrameData[8]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit8.Q ));
 sg13g2_dlhq_1 _1047_ (.D(Tile_X0Y0_FrameData[7]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit7.Q ));
 sg13g2_dlhq_1 _1048_ (.D(Tile_X0Y0_FrameData[6]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit6.Q ));
 sg13g2_dlhq_1 _1049_ (.D(Tile_X0Y0_FrameData[5]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit5.Q ));
 sg13g2_dlhq_1 _1050_ (.D(Tile_X0Y0_FrameData[4]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit4.Q ));
 sg13g2_dlhq_1 _1051_ (.D(Tile_X0Y0_FrameData[3]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit3.Q ));
 sg13g2_dlhq_1 _1052_ (.D(Tile_X0Y0_FrameData[2]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit2.Q ));
 sg13g2_dlhq_1 _1053_ (.D(Tile_X0Y0_FrameData[1]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit1.Q ));
 sg13g2_dlhq_1 _1054_ (.D(Tile_X0Y0_FrameData[0]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit0.Q ));
 sg13g2_dlhq_1 _1055_ (.D(Tile_X0Y0_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit31.Q ));
 sg13g2_dlhq_1 _1056_ (.D(Tile_X0Y0_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit30.Q ));
 sg13g2_dlhq_1 _1057_ (.D(Tile_X0Y0_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit29.Q ));
 sg13g2_dlhq_1 _1058_ (.D(Tile_X0Y0_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit28.Q ));
 sg13g2_dlhq_1 _1059_ (.D(Tile_X0Y0_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit27.Q ));
 sg13g2_dlhq_1 _1060_ (.D(Tile_X0Y0_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit26.Q ));
 sg13g2_dlhq_1 _1061_ (.D(Tile_X0Y0_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit25.Q ));
 sg13g2_dlhq_1 _1062_ (.D(Tile_X0Y0_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit24.Q ));
 sg13g2_dlhq_1 _1063_ (.D(Tile_X0Y0_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit23.Q ));
 sg13g2_dlhq_1 _1064_ (.D(Tile_X0Y0_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit22.Q ));
 sg13g2_dlhq_1 _1065_ (.D(Tile_X0Y0_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit21.Q ));
 sg13g2_dlhq_1 _1066_ (.D(Tile_X0Y0_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit20.Q ));
 sg13g2_dlhq_1 _1067_ (.D(Tile_X0Y0_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit19.Q ));
 sg13g2_dlhq_1 _1068_ (.D(Tile_X0Y0_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit18.Q ));
 sg13g2_dlhq_1 _1069_ (.D(Tile_X0Y0_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit17.Q ));
 sg13g2_dlhq_1 _1070_ (.D(Tile_X0Y0_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit16.Q ));
 sg13g2_dlhq_1 _1071_ (.D(Tile_X0Y0_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit15.Q ));
 sg13g2_dlhq_1 _1072_ (.D(Tile_X0Y0_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit14.Q ));
 sg13g2_dlhq_1 _1073_ (.D(Tile_X0Y0_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit13.Q ));
 sg13g2_dlhq_1 _1074_ (.D(Tile_X0Y0_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit12.Q ));
 sg13g2_dlhq_1 _1075_ (.D(Tile_X0Y0_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit11.Q ));
 sg13g2_dlhq_1 _1076_ (.D(Tile_X0Y0_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit10.Q ));
 sg13g2_dlhq_1 _1077_ (.D(Tile_X0Y0_FrameData[9]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit9.Q ));
 sg13g2_dlhq_1 _1078_ (.D(Tile_X0Y0_FrameData[8]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit8.Q ));
 sg13g2_dlhq_1 _1079_ (.D(Tile_X0Y0_FrameData[7]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit7.Q ));
 sg13g2_dlhq_1 _1080_ (.D(Tile_X0Y0_FrameData[6]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit6.Q ));
 sg13g2_dlhq_1 _1081_ (.D(Tile_X0Y0_FrameData[5]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit5.Q ));
 sg13g2_dlhq_1 _1082_ (.D(Tile_X0Y0_FrameData[4]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit4.Q ));
 sg13g2_dlhq_1 _1083_ (.D(Tile_X0Y0_FrameData[3]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit3.Q ));
 sg13g2_dlhq_1 _1084_ (.D(Tile_X0Y0_FrameData[2]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit2.Q ));
 sg13g2_dlhq_1 _1085_ (.D(Tile_X0Y0_FrameData[1]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit1.Q ));
 sg13g2_dlhq_1 _1086_ (.D(Tile_X0Y0_FrameData[0]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit0.Q ));
 sg13g2_dlhq_1 _1087_ (.D(Tile_X0Y0_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit31.Q ));
 sg13g2_dlhq_1 _1088_ (.D(Tile_X0Y0_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit30.Q ));
 sg13g2_dlhq_1 _1089_ (.D(Tile_X0Y0_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit29.Q ));
 sg13g2_dlhq_1 _1090_ (.D(Tile_X0Y0_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit28.Q ));
 sg13g2_dlhq_1 _1091_ (.D(Tile_X0Y0_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit27.Q ));
 sg13g2_dlhq_1 _1092_ (.D(Tile_X0Y0_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit26.Q ));
 sg13g2_dlhq_1 _1093_ (.D(Tile_X0Y0_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit25.Q ));
 sg13g2_dlhq_1 _1094_ (.D(Tile_X0Y0_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit24.Q ));
 sg13g2_dlhq_1 _1095_ (.D(Tile_X0Y0_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit23.Q ));
 sg13g2_dlhq_1 _1096_ (.D(Tile_X0Y0_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit22.Q ));
 sg13g2_dlhq_1 _1097_ (.D(Tile_X0Y0_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit21.Q ));
 sg13g2_dlhq_1 _1098_ (.D(Tile_X0Y0_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit20.Q ));
 sg13g2_dlhq_1 _1099_ (.D(Tile_X0Y0_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit19.Q ));
 sg13g2_dlhq_1 _1100_ (.D(Tile_X0Y0_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit18.Q ));
 sg13g2_dlhq_1 _1101_ (.D(Tile_X0Y0_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit17.Q ));
 sg13g2_dlhq_1 _1102_ (.D(Tile_X0Y0_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit16.Q ));
 sg13g2_dlhq_1 _1103_ (.D(Tile_X0Y0_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit15.Q ));
 sg13g2_dlhq_1 _1104_ (.D(Tile_X0Y0_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit14.Q ));
 sg13g2_dlhq_1 _1105_ (.D(Tile_X0Y0_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit13.Q ));
 sg13g2_dlhq_1 _1106_ (.D(Tile_X0Y0_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit12.Q ));
 sg13g2_dlhq_1 _1107_ (.D(Tile_X0Y0_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit11.Q ));
 sg13g2_dlhq_1 _1108_ (.D(Tile_X0Y0_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit10.Q ));
 sg13g2_dlhq_1 _1109_ (.D(Tile_X0Y0_FrameData[9]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit9.Q ));
 sg13g2_dlhq_1 _1110_ (.D(Tile_X0Y0_FrameData[8]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit8.Q ));
 sg13g2_dlhq_1 _1111_ (.D(Tile_X0Y0_FrameData[7]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit7.Q ));
 sg13g2_dlhq_1 _1112_ (.D(Tile_X0Y0_FrameData[6]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit6.Q ));
 sg13g2_dlhq_1 _1113_ (.D(Tile_X0Y0_FrameData[5]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit5.Q ));
 sg13g2_dlhq_1 _1114_ (.D(Tile_X0Y0_FrameData[4]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit4.Q ));
 sg13g2_dlhq_1 _1115_ (.D(Tile_X0Y0_FrameData[3]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit3.Q ));
 sg13g2_dlhq_1 _1116_ (.D(Tile_X0Y0_FrameData[2]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit2.Q ));
 sg13g2_dlhq_1 _1117_ (.D(Tile_X0Y0_FrameData[1]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit1.Q ));
 sg13g2_dlhq_1 _1118_ (.D(Tile_X0Y0_FrameData[0]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit0.Q ));
 sg13g2_dlhq_1 _1119_ (.D(Tile_X0Y0_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit31.Q ));
 sg13g2_dlhq_1 _1120_ (.D(Tile_X0Y0_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit30.Q ));
 sg13g2_dlhq_1 _1121_ (.D(Tile_X0Y0_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit29.Q ));
 sg13g2_dlhq_1 _1122_ (.D(Tile_X0Y0_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit28.Q ));
 sg13g2_dlhq_1 _1123_ (.D(Tile_X0Y0_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit27.Q ));
 sg13g2_dlhq_1 _1124_ (.D(Tile_X0Y0_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit26.Q ));
 sg13g2_dlhq_1 _1125_ (.D(Tile_X0Y0_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit25.Q ));
 sg13g2_dlhq_1 _1126_ (.D(Tile_X0Y0_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit24.Q ));
 sg13g2_dlhq_1 _1127_ (.D(Tile_X0Y0_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit23.Q ));
 sg13g2_dlhq_1 _1128_ (.D(Tile_X0Y0_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit22.Q ));
 sg13g2_dlhq_1 _1129_ (.D(Tile_X0Y0_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit21.Q ));
 sg13g2_dlhq_1 _1130_ (.D(Tile_X0Y0_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit20.Q ));
 sg13g2_dlhq_1 _1131_ (.D(Tile_X0Y0_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit19.Q ));
 sg13g2_dlhq_1 _1132_ (.D(Tile_X0Y0_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit18.Q ));
 sg13g2_dlhq_1 _1133_ (.D(Tile_X0Y0_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit17.Q ));
 sg13g2_dlhq_1 _1134_ (.D(Tile_X0Y0_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit16.Q ));
 sg13g2_dlhq_1 _1135_ (.D(Tile_X0Y0_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit15.Q ));
 sg13g2_dlhq_1 _1136_ (.D(Tile_X0Y0_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit14.Q ));
 sg13g2_dlhq_1 _1137_ (.D(Tile_X0Y0_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit13.Q ));
 sg13g2_dlhq_1 _1138_ (.D(Tile_X0Y0_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit12.Q ));
 sg13g2_dlhq_1 _1139_ (.D(Tile_X0Y0_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit11.Q ));
 sg13g2_dlhq_1 _1140_ (.D(Tile_X0Y0_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit10.Q ));
 sg13g2_dlhq_1 _1141_ (.D(Tile_X0Y0_FrameData[9]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit9.Q ));
 sg13g2_dlhq_1 _1142_ (.D(Tile_X0Y0_FrameData[8]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit8.Q ));
 sg13g2_dlhq_1 _1143_ (.D(Tile_X0Y0_FrameData[7]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit7.Q ));
 sg13g2_dlhq_1 _1144_ (.D(Tile_X0Y0_FrameData[6]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit6.Q ));
 sg13g2_dlhq_1 _1145_ (.D(Tile_X0Y0_FrameData[5]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit5.Q ));
 sg13g2_dlhq_1 _1146_ (.D(Tile_X0Y0_FrameData[4]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit4.Q ));
 sg13g2_dlhq_1 _1147_ (.D(Tile_X0Y0_FrameData[3]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit3.Q ));
 sg13g2_dlhq_1 _1148_ (.D(Tile_X0Y0_FrameData[2]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit2.Q ));
 sg13g2_dlhq_1 _1149_ (.D(Tile_X0Y0_FrameData[1]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit1.Q ));
 sg13g2_dlhq_1 _1150_ (.D(Tile_X0Y0_FrameData[0]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit0.Q ));
 sg13g2_dlhq_1 _1151_ (.D(Tile_X0Y0_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit31.Q ));
 sg13g2_dlhq_1 _1152_ (.D(Tile_X0Y0_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit30.Q ));
 sg13g2_dlhq_1 _1153_ (.D(Tile_X0Y0_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit29.Q ));
 sg13g2_dlhq_1 _1154_ (.D(Tile_X0Y0_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit28.Q ));
 sg13g2_dlhq_1 _1155_ (.D(Tile_X0Y0_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit27.Q ));
 sg13g2_dlhq_1 _1156_ (.D(Tile_X0Y0_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit26.Q ));
 sg13g2_dlhq_1 _1157_ (.D(Tile_X0Y0_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit25.Q ));
 sg13g2_dlhq_1 _1158_ (.D(Tile_X0Y0_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit24.Q ));
 sg13g2_dlhq_1 _1159_ (.D(Tile_X0Y0_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit23.Q ));
 sg13g2_dlhq_1 _1160_ (.D(Tile_X0Y0_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit22.Q ));
 sg13g2_dlhq_1 _1161_ (.D(Tile_X0Y1_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit31.Q ));
 sg13g2_dlhq_1 _1162_ (.D(Tile_X0Y1_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q ));
 sg13g2_dlhq_1 _1163_ (.D(Tile_X0Y1_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit29.Q ));
 sg13g2_dlhq_1 _1164_ (.D(Tile_X0Y1_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q ));
 sg13g2_dlhq_1 _1165_ (.D(Tile_X0Y1_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit27.Q ));
 sg13g2_dlhq_1 _1166_ (.D(Tile_X0Y1_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_dlhq_1 _1167_ (.D(Tile_X0Y1_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit25.Q ));
 sg13g2_dlhq_1 _1168_ (.D(Tile_X0Y1_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_dlhq_1 _1169_ (.D(Tile_X0Y1_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit23.Q ));
 sg13g2_dlhq_1 _1170_ (.D(Tile_X0Y1_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit22.Q ));
 sg13g2_dlhq_1 _1171_ (.D(Tile_X0Y1_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit21.Q ));
 sg13g2_dlhq_1 _1172_ (.D(Tile_X0Y1_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit20.Q ));
 sg13g2_dlhq_1 _1173_ (.D(Tile_X0Y1_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit19.Q ));
 sg13g2_dlhq_1 _1174_ (.D(Tile_X0Y1_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit18.Q ));
 sg13g2_dlhq_1 _1175_ (.D(Tile_X0Y1_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit17.Q ));
 sg13g2_dlhq_1 _1176_ (.D(Tile_X0Y1_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit16.Q ));
 sg13g2_dlhq_1 _1177_ (.D(Tile_X0Y1_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit15.Q ));
 sg13g2_dlhq_1 _1178_ (.D(Tile_X0Y1_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit14.Q ));
 sg13g2_dlhq_1 _1179_ (.D(Tile_X0Y1_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit13.Q ));
 sg13g2_dlhq_1 _1180_ (.D(Tile_X0Y1_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit12.Q ));
 sg13g2_dlhq_1 _1181_ (.D(Tile_X0Y1_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit11.Q ));
 sg13g2_dlhq_1 _1182_ (.D(Tile_X0Y1_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit10.Q ));
 sg13g2_dlhq_1 _1183_ (.D(Tile_X0Y1_FrameData[9]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit9.Q ));
 sg13g2_dlhq_1 _1184_ (.D(Tile_X0Y1_FrameData[8]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit8.Q ));
 sg13g2_dlhq_1 _1185_ (.D(Tile_X0Y1_FrameData[7]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit7.Q ));
 sg13g2_dlhq_1 _1186_ (.D(Tile_X0Y1_FrameData[6]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit6.Q ));
 sg13g2_dlhq_1 _1187_ (.D(Tile_X0Y1_FrameData[5]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit5.Q ));
 sg13g2_dlhq_1 _1188_ (.D(Tile_X0Y1_FrameData[4]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit4.Q ));
 sg13g2_dlhq_1 _1189_ (.D(Tile_X0Y1_FrameData[3]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit3.Q ));
 sg13g2_dlhq_1 _1190_ (.D(Tile_X0Y1_FrameData[2]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit2.Q ));
 sg13g2_dlhq_1 _1191_ (.D(Tile_X0Y1_FrameData[1]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit1.Q ));
 sg13g2_dlhq_1 _1192_ (.D(Tile_X0Y1_FrameData[0]),
    .GATE(Tile_X0Y1_FrameStrobe[0]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit0.Q ));
 sg13g2_dlhq_1 _1193_ (.D(Tile_X0Y1_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit31.Q ));
 sg13g2_dlhq_1 _1194_ (.D(Tile_X0Y1_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit30.Q ));
 sg13g2_dlhq_1 _1195_ (.D(Tile_X0Y1_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit29.Q ));
 sg13g2_dlhq_1 _1196_ (.D(Tile_X0Y1_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit28.Q ));
 sg13g2_dlhq_1 _1197_ (.D(Tile_X0Y1_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit27.Q ));
 sg13g2_dlhq_1 _1198_ (.D(Tile_X0Y1_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit26.Q ));
 sg13g2_dlhq_1 _1199_ (.D(Tile_X0Y1_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit25.Q ));
 sg13g2_dlhq_1 _1200_ (.D(Tile_X0Y1_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit24.Q ));
 sg13g2_dlhq_1 _1201_ (.D(Tile_X0Y1_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit23.Q ));
 sg13g2_dlhq_1 _1202_ (.D(Tile_X0Y1_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit22.Q ));
 sg13g2_dlhq_1 _1203_ (.D(Tile_X0Y1_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit21.Q ));
 sg13g2_dlhq_1 _1204_ (.D(Tile_X0Y1_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit20.Q ));
 sg13g2_dlhq_1 _1205_ (.D(Tile_X0Y1_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit19.Q ));
 sg13g2_dlhq_1 _1206_ (.D(Tile_X0Y1_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit18.Q ));
 sg13g2_dlhq_1 _1207_ (.D(Tile_X0Y1_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit17.Q ));
 sg13g2_dlhq_1 _1208_ (.D(Tile_X0Y1_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit16.Q ));
 sg13g2_dlhq_1 _1209_ (.D(Tile_X0Y1_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit15.Q ));
 sg13g2_dlhq_1 _1210_ (.D(Tile_X0Y1_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit14.Q ));
 sg13g2_dlhq_1 _1211_ (.D(Tile_X0Y1_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit13.Q ));
 sg13g2_dlhq_1 _1212_ (.D(Tile_X0Y1_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit12.Q ));
 sg13g2_dlhq_1 _1213_ (.D(Tile_X0Y1_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit11.Q ));
 sg13g2_dlhq_1 _1214_ (.D(Tile_X0Y1_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit10.Q ));
 sg13g2_dlhq_1 _1215_ (.D(Tile_X0Y1_FrameData[9]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit9.Q ));
 sg13g2_dlhq_1 _1216_ (.D(Tile_X0Y1_FrameData[8]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit8.Q ));
 sg13g2_dlhq_1 _1217_ (.D(Tile_X0Y1_FrameData[7]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit7.Q ));
 sg13g2_dlhq_1 _1218_ (.D(Tile_X0Y1_FrameData[6]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q ));
 sg13g2_dlhq_1 _1219_ (.D(Tile_X0Y1_FrameData[5]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q ));
 sg13g2_dlhq_1 _1220_ (.D(Tile_X0Y1_FrameData[4]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q ));
 sg13g2_dlhq_1 _1221_ (.D(Tile_X0Y1_FrameData[3]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit3.Q ));
 sg13g2_dlhq_1 _1222_ (.D(Tile_X0Y1_FrameData[2]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q ));
 sg13g2_dlhq_1 _1223_ (.D(Tile_X0Y1_FrameData[1]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q ));
 sg13g2_dlhq_1 _1224_ (.D(Tile_X0Y1_FrameData[0]),
    .GATE(Tile_X0Y1_FrameStrobe[1]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q ));
 sg13g2_dlhq_1 _1225_ (.D(Tile_X0Y1_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit31.Q ));
 sg13g2_dlhq_1 _1226_ (.D(Tile_X0Y1_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q ));
 sg13g2_dlhq_1 _1227_ (.D(Tile_X0Y1_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q ));
 sg13g2_dlhq_1 _1228_ (.D(Tile_X0Y1_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q ));
 sg13g2_dlhq_1 _1229_ (.D(Tile_X0Y1_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit27.Q ));
 sg13g2_dlhq_1 _1230_ (.D(Tile_X0Y1_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit26.Q ));
 sg13g2_dlhq_1 _1231_ (.D(Tile_X0Y1_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit25.Q ));
 sg13g2_dlhq_1 _1232_ (.D(Tile_X0Y1_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit24.Q ));
 sg13g2_dlhq_1 _1233_ (.D(Tile_X0Y1_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit23.Q ));
 sg13g2_dlhq_1 _1234_ (.D(Tile_X0Y1_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit22.Q ));
 sg13g2_dlhq_1 _1235_ (.D(Tile_X0Y1_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit21.Q ));
 sg13g2_dlhq_1 _1236_ (.D(Tile_X0Y1_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit20.Q ));
 sg13g2_dlhq_1 _1237_ (.D(Tile_X0Y1_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit19.Q ));
 sg13g2_dlhq_1 _1238_ (.D(Tile_X0Y1_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit18.Q ));
 sg13g2_dlhq_1 _1239_ (.D(Tile_X0Y1_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit17.Q ));
 sg13g2_dlhq_1 _1240_ (.D(Tile_X0Y1_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit16.Q ));
 sg13g2_dlhq_1 _1241_ (.D(Tile_X0Y1_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit15.Q ));
 sg13g2_dlhq_1 _1242_ (.D(Tile_X0Y1_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit14.Q ));
 sg13g2_dlhq_1 _1243_ (.D(Tile_X0Y1_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit13.Q ));
 sg13g2_dlhq_1 _1244_ (.D(Tile_X0Y1_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit12.Q ));
 sg13g2_dlhq_1 _1245_ (.D(Tile_X0Y1_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit11.Q ));
 sg13g2_dlhq_1 _1246_ (.D(Tile_X0Y1_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit10.Q ));
 sg13g2_dlhq_1 _1247_ (.D(Tile_X0Y1_FrameData[9]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit9.Q ));
 sg13g2_dlhq_1 _1248_ (.D(Tile_X0Y1_FrameData[8]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit8.Q ));
 sg13g2_dlhq_1 _1249_ (.D(Tile_X0Y1_FrameData[7]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit7.Q ));
 sg13g2_dlhq_1 _1250_ (.D(Tile_X0Y1_FrameData[6]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit6.Q ));
 sg13g2_dlhq_1 _1251_ (.D(Tile_X0Y1_FrameData[5]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit5.Q ));
 sg13g2_dlhq_1 _1252_ (.D(Tile_X0Y1_FrameData[4]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q ));
 sg13g2_dlhq_1 _1253_ (.D(Tile_X0Y1_FrameData[3]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit3.Q ));
 sg13g2_dlhq_1 _1254_ (.D(Tile_X0Y1_FrameData[2]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit2.Q ));
 sg13g2_dlhq_1 _1255_ (.D(Tile_X0Y1_FrameData[1]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit1.Q ));
 sg13g2_dlhq_1 _1256_ (.D(Tile_X0Y1_FrameData[0]),
    .GATE(Tile_X0Y1_FrameStrobe[2]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q ));
 sg13g2_dlhq_1 _1257_ (.D(Tile_X0Y1_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit31.Q ));
 sg13g2_dlhq_1 _1258_ (.D(Tile_X0Y1_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit30.Q ));
 sg13g2_dlhq_1 _1259_ (.D(Tile_X0Y1_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit29.Q ));
 sg13g2_dlhq_1 _1260_ (.D(Tile_X0Y1_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit28.Q ));
 sg13g2_dlhq_1 _1261_ (.D(Tile_X0Y1_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit27.Q ));
 sg13g2_dlhq_1 _1262_ (.D(Tile_X0Y1_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit26.Q ));
 sg13g2_dlhq_1 _1263_ (.D(Tile_X0Y1_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit25.Q ));
 sg13g2_dlhq_1 _1264_ (.D(Tile_X0Y1_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit24.Q ));
 sg13g2_dlhq_1 _1265_ (.D(Tile_X0Y1_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit23.Q ));
 sg13g2_dlhq_1 _1266_ (.D(Tile_X0Y1_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit22.Q ));
 sg13g2_dlhq_1 _1267_ (.D(Tile_X0Y1_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit21.Q ));
 sg13g2_dlhq_1 _1268_ (.D(Tile_X0Y1_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit20.Q ));
 sg13g2_dlhq_1 _1269_ (.D(Tile_X0Y1_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit19.Q ));
 sg13g2_dlhq_1 _1270_ (.D(Tile_X0Y1_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit18.Q ));
 sg13g2_dlhq_1 _1271_ (.D(Tile_X0Y1_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit17.Q ));
 sg13g2_dlhq_1 _1272_ (.D(Tile_X0Y1_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit16.Q ));
 sg13g2_dlhq_1 _1273_ (.D(Tile_X0Y1_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit15.Q ));
 sg13g2_dlhq_1 _1274_ (.D(Tile_X0Y1_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit14.Q ));
 sg13g2_dlhq_1 _1275_ (.D(Tile_X0Y1_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit13.Q ));
 sg13g2_dlhq_1 _1276_ (.D(Tile_X0Y1_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit12.Q ));
 sg13g2_dlhq_1 _1277_ (.D(Tile_X0Y1_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit11.Q ));
 sg13g2_dlhq_1 _1278_ (.D(Tile_X0Y1_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit10.Q ));
 sg13g2_dlhq_1 _1279_ (.D(Tile_X0Y1_FrameData[9]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit9.Q ));
 sg13g2_dlhq_1 _1280_ (.D(Tile_X0Y1_FrameData[8]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit8.Q ));
 sg13g2_dlhq_1 _1281_ (.D(Tile_X0Y1_FrameData[7]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit7.Q ));
 sg13g2_dlhq_1 _1282_ (.D(Tile_X0Y1_FrameData[6]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit6.Q ));
 sg13g2_dlhq_1 _1283_ (.D(Tile_X0Y1_FrameData[5]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit5.Q ));
 sg13g2_dlhq_1 _1284_ (.D(Tile_X0Y1_FrameData[4]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit4.Q ));
 sg13g2_dlhq_1 _1285_ (.D(Tile_X0Y1_FrameData[3]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit3.Q ));
 sg13g2_dlhq_1 _1286_ (.D(Tile_X0Y1_FrameData[2]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit2.Q ));
 sg13g2_dlhq_1 _1287_ (.D(Tile_X0Y1_FrameData[1]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit1.Q ));
 sg13g2_dlhq_1 _1288_ (.D(Tile_X0Y1_FrameData[0]),
    .GATE(Tile_X0Y1_FrameStrobe[3]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit0.Q ));
 sg13g2_dlhq_1 _1289_ (.D(Tile_X0Y1_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit31.Q ));
 sg13g2_dlhq_1 _1290_ (.D(Tile_X0Y1_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit30.Q ));
 sg13g2_dlhq_1 _1291_ (.D(Tile_X0Y1_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit29.Q ));
 sg13g2_dlhq_1 _1292_ (.D(Tile_X0Y1_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit28.Q ));
 sg13g2_dlhq_1 _1293_ (.D(Tile_X0Y1_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit27.Q ));
 sg13g2_dlhq_1 _1294_ (.D(Tile_X0Y1_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit26.Q ));
 sg13g2_dlhq_1 _1295_ (.D(Tile_X0Y1_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit25.Q ));
 sg13g2_dlhq_1 _1296_ (.D(Tile_X0Y1_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit24.Q ));
 sg13g2_dlhq_1 _1297_ (.D(Tile_X0Y1_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit23.Q ));
 sg13g2_dlhq_1 _1298_ (.D(Tile_X0Y1_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit22.Q ));
 sg13g2_dlhq_1 _1299_ (.D(Tile_X0Y1_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit21.Q ));
 sg13g2_dlhq_1 _1300_ (.D(Tile_X0Y1_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit20.Q ));
 sg13g2_dlhq_1 _1301_ (.D(Tile_X0Y1_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit19.Q ));
 sg13g2_dlhq_1 _1302_ (.D(Tile_X0Y1_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit18.Q ));
 sg13g2_dlhq_1 _1303_ (.D(Tile_X0Y1_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit17.Q ));
 sg13g2_dlhq_1 _1304_ (.D(Tile_X0Y1_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit16.Q ));
 sg13g2_dlhq_1 _1305_ (.D(Tile_X0Y1_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit15.Q ));
 sg13g2_dlhq_1 _1306_ (.D(Tile_X0Y1_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit14.Q ));
 sg13g2_dlhq_1 _1307_ (.D(Tile_X0Y1_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit13.Q ));
 sg13g2_dlhq_1 _1308_ (.D(Tile_X0Y1_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit12.Q ));
 sg13g2_dlhq_1 _1309_ (.D(Tile_X0Y1_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit11.Q ));
 sg13g2_dlhq_1 _1310_ (.D(Tile_X0Y1_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit10.Q ));
 sg13g2_dlhq_1 _1311_ (.D(Tile_X0Y1_FrameData[9]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit9.Q ));
 sg13g2_dlhq_1 _1312_ (.D(Tile_X0Y1_FrameData[8]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit8.Q ));
 sg13g2_dlhq_1 _1313_ (.D(Tile_X0Y1_FrameData[7]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit7.Q ));
 sg13g2_dlhq_1 _1314_ (.D(Tile_X0Y1_FrameData[6]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit6.Q ));
 sg13g2_dlhq_1 _1315_ (.D(Tile_X0Y1_FrameData[5]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit5.Q ));
 sg13g2_dlhq_1 _1316_ (.D(Tile_X0Y1_FrameData[4]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit4.Q ));
 sg13g2_dlhq_1 _1317_ (.D(Tile_X0Y1_FrameData[3]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit3.Q ));
 sg13g2_dlhq_1 _1318_ (.D(Tile_X0Y1_FrameData[2]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit2.Q ));
 sg13g2_dlhq_1 _1319_ (.D(Tile_X0Y1_FrameData[1]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit1.Q ));
 sg13g2_dlhq_1 _1320_ (.D(Tile_X0Y1_FrameData[0]),
    .GATE(Tile_X0Y1_FrameStrobe[4]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit0.Q ));
 sg13g2_dlhq_1 _1321_ (.D(Tile_X0Y1_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit31.Q ));
 sg13g2_dlhq_1 _1322_ (.D(Tile_X0Y1_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit30.Q ));
 sg13g2_dlhq_1 _1323_ (.D(Tile_X0Y1_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit29.Q ));
 sg13g2_dlhq_1 _1324_ (.D(Tile_X0Y1_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit28.Q ));
 sg13g2_dlhq_1 _1325_ (.D(Tile_X0Y1_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit27.Q ));
 sg13g2_dlhq_1 _1326_ (.D(Tile_X0Y1_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit26.Q ));
 sg13g2_dlhq_1 _1327_ (.D(Tile_X0Y1_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit25.Q ));
 sg13g2_dlhq_1 _1328_ (.D(Tile_X0Y1_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit24.Q ));
 sg13g2_dlhq_1 _1329_ (.D(Tile_X0Y1_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit23.Q ));
 sg13g2_dlhq_1 _1330_ (.D(Tile_X0Y1_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit22.Q ));
 sg13g2_dlhq_1 _1331_ (.D(Tile_X0Y1_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit21.Q ));
 sg13g2_dlhq_1 _1332_ (.D(Tile_X0Y1_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit20.Q ));
 sg13g2_dlhq_1 _1333_ (.D(Tile_X0Y1_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit19.Q ));
 sg13g2_dlhq_1 _1334_ (.D(Tile_X0Y1_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit18.Q ));
 sg13g2_dlhq_1 _1335_ (.D(Tile_X0Y1_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit17.Q ));
 sg13g2_dlhq_1 _1336_ (.D(Tile_X0Y1_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit16.Q ));
 sg13g2_dlhq_1 _1337_ (.D(Tile_X0Y1_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit15.Q ));
 sg13g2_dlhq_1 _1338_ (.D(Tile_X0Y1_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit14.Q ));
 sg13g2_dlhq_1 _1339_ (.D(Tile_X0Y1_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit13.Q ));
 sg13g2_dlhq_1 _1340_ (.D(Tile_X0Y1_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit12.Q ));
 sg13g2_dlhq_1 _1341_ (.D(Tile_X0Y1_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit11.Q ));
 sg13g2_dlhq_1 _1342_ (.D(Tile_X0Y1_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit10.Q ));
 sg13g2_dlhq_1 _1343_ (.D(Tile_X0Y1_FrameData[9]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit9.Q ));
 sg13g2_dlhq_1 _1344_ (.D(Tile_X0Y1_FrameData[8]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit8.Q ));
 sg13g2_dlhq_1 _1345_ (.D(Tile_X0Y1_FrameData[7]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit7.Q ));
 sg13g2_dlhq_1 _1346_ (.D(Tile_X0Y1_FrameData[6]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit6.Q ));
 sg13g2_dlhq_1 _1347_ (.D(Tile_X0Y1_FrameData[5]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit5.Q ));
 sg13g2_dlhq_1 _1348_ (.D(Tile_X0Y1_FrameData[4]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit4.Q ));
 sg13g2_dlhq_1 _1349_ (.D(Tile_X0Y1_FrameData[3]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit3.Q ));
 sg13g2_dlhq_1 _1350_ (.D(Tile_X0Y1_FrameData[2]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit2.Q ));
 sg13g2_dlhq_1 _1351_ (.D(Tile_X0Y1_FrameData[1]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit1.Q ));
 sg13g2_dlhq_1 _1352_ (.D(Tile_X0Y1_FrameData[0]),
    .GATE(Tile_X0Y1_FrameStrobe[5]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit0.Q ));
 sg13g2_dlhq_1 _1353_ (.D(Tile_X0Y1_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit31.Q ));
 sg13g2_dlhq_1 _1354_ (.D(Tile_X0Y1_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit30.Q ));
 sg13g2_dlhq_1 _1355_ (.D(Tile_X0Y1_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit29.Q ));
 sg13g2_dlhq_1 _1356_ (.D(Tile_X0Y1_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit28.Q ));
 sg13g2_dlhq_1 _1357_ (.D(Tile_X0Y1_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit27.Q ));
 sg13g2_dlhq_1 _1358_ (.D(Tile_X0Y1_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit26.Q ));
 sg13g2_dlhq_1 _1359_ (.D(Tile_X0Y1_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit25.Q ));
 sg13g2_dlhq_1 _1360_ (.D(Tile_X0Y1_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit24.Q ));
 sg13g2_dlhq_1 _1361_ (.D(Tile_X0Y1_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit23.Q ));
 sg13g2_dlhq_1 _1362_ (.D(Tile_X0Y1_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit22.Q ));
 sg13g2_dlhq_1 _1363_ (.D(Tile_X0Y1_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit21.Q ));
 sg13g2_dlhq_1 _1364_ (.D(Tile_X0Y1_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit20.Q ));
 sg13g2_dlhq_1 _1365_ (.D(Tile_X0Y1_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit19.Q ));
 sg13g2_dlhq_1 _1366_ (.D(Tile_X0Y1_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit18.Q ));
 sg13g2_dlhq_1 _1367_ (.D(Tile_X0Y1_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit17.Q ));
 sg13g2_dlhq_1 _1368_ (.D(Tile_X0Y1_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit16.Q ));
 sg13g2_dlhq_1 _1369_ (.D(Tile_X0Y1_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit15.Q ));
 sg13g2_dlhq_1 _1370_ (.D(Tile_X0Y1_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit14.Q ));
 sg13g2_dlhq_1 _1371_ (.D(Tile_X0Y1_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit13.Q ));
 sg13g2_dlhq_1 _1372_ (.D(Tile_X0Y1_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit12.Q ));
 sg13g2_dlhq_1 _1373_ (.D(Tile_X0Y1_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit11.Q ));
 sg13g2_dlhq_1 _1374_ (.D(Tile_X0Y1_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit10.Q ));
 sg13g2_dlhq_1 _1375_ (.D(Tile_X0Y1_FrameData[9]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit9.Q ));
 sg13g2_dlhq_1 _1376_ (.D(Tile_X0Y1_FrameData[8]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit8.Q ));
 sg13g2_dlhq_1 _1377_ (.D(Tile_X0Y1_FrameData[7]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit7.Q ));
 sg13g2_dlhq_1 _1378_ (.D(Tile_X0Y1_FrameData[6]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit6.Q ));
 sg13g2_dlhq_1 _1379_ (.D(Tile_X0Y1_FrameData[5]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit5.Q ));
 sg13g2_dlhq_1 _1380_ (.D(Tile_X0Y1_FrameData[4]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit4.Q ));
 sg13g2_dlhq_1 _1381_ (.D(Tile_X0Y1_FrameData[3]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit3.Q ));
 sg13g2_dlhq_1 _1382_ (.D(Tile_X0Y1_FrameData[2]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit2.Q ));
 sg13g2_dlhq_1 _1383_ (.D(Tile_X0Y1_FrameData[1]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit1.Q ));
 sg13g2_dlhq_1 _1384_ (.D(Tile_X0Y1_FrameData[0]),
    .GATE(Tile_X0Y1_FrameStrobe[6]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit0.Q ));
 sg13g2_dlhq_1 _1385_ (.D(Tile_X0Y1_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit31.Q ));
 sg13g2_dlhq_1 _1386_ (.D(Tile_X0Y1_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit30.Q ));
 sg13g2_dlhq_1 _1387_ (.D(Tile_X0Y1_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit29.Q ));
 sg13g2_dlhq_1 _1388_ (.D(Tile_X0Y1_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit28.Q ));
 sg13g2_dlhq_1 _1389_ (.D(Tile_X0Y1_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit27.Q ));
 sg13g2_dlhq_1 _1390_ (.D(Tile_X0Y1_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit26.Q ));
 sg13g2_dlhq_1 _1391_ (.D(Tile_X0Y1_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit25.Q ));
 sg13g2_dlhq_1 _1392_ (.D(Tile_X0Y1_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit24.Q ));
 sg13g2_dlhq_1 _1393_ (.D(Tile_X0Y1_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit23.Q ));
 sg13g2_dlhq_1 _1394_ (.D(Tile_X0Y1_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit22.Q ));
 sg13g2_dlhq_1 _1395_ (.D(Tile_X0Y1_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit21.Q ));
 sg13g2_dlhq_1 _1396_ (.D(Tile_X0Y1_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit20.Q ));
 sg13g2_dlhq_1 _1397_ (.D(Tile_X0Y1_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit19.Q ));
 sg13g2_dlhq_1 _1398_ (.D(Tile_X0Y1_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit18.Q ));
 sg13g2_dlhq_1 _1399_ (.D(Tile_X0Y1_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit17.Q ));
 sg13g2_dlhq_1 _1400_ (.D(Tile_X0Y1_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q ));
 sg13g2_dlhq_1 _1401_ (.D(Tile_X0Y1_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q ));
 sg13g2_dlhq_1 _1402_ (.D(Tile_X0Y1_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit14.Q ));
 sg13g2_dlhq_1 _1403_ (.D(Tile_X0Y1_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q ));
 sg13g2_dlhq_1 _1404_ (.D(Tile_X0Y1_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q ));
 sg13g2_dlhq_1 _1405_ (.D(Tile_X0Y1_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit11.Q ));
 sg13g2_dlhq_1 _1406_ (.D(Tile_X0Y1_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q ));
 sg13g2_dlhq_1 _1407_ (.D(Tile_X0Y1_FrameData[9]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q ));
 sg13g2_dlhq_1 _1408_ (.D(Tile_X0Y1_FrameData[8]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit8.Q ));
 sg13g2_dlhq_1 _1409_ (.D(Tile_X0Y1_FrameData[7]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit7.Q ));
 sg13g2_dlhq_1 _1410_ (.D(Tile_X0Y1_FrameData[6]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q ));
 sg13g2_dlhq_1 _1411_ (.D(Tile_X0Y1_FrameData[5]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit5.Q ));
 sg13g2_dlhq_1 _1412_ (.D(Tile_X0Y1_FrameData[4]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit4.Q ));
 sg13g2_dlhq_1 _1413_ (.D(Tile_X0Y1_FrameData[3]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit3.Q ));
 sg13g2_dlhq_1 _1414_ (.D(Tile_X0Y1_FrameData[2]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit2.Q ));
 sg13g2_dlhq_1 _1415_ (.D(Tile_X0Y1_FrameData[1]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit1.Q ));
 sg13g2_dlhq_1 _1416_ (.D(Tile_X0Y1_FrameData[0]),
    .GATE(Tile_X0Y1_FrameStrobe[7]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit0.Q ));
 sg13g2_dlhq_1 _1417_ (.D(Tile_X0Y1_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit31.Q ));
 sg13g2_dlhq_1 _1418_ (.D(Tile_X0Y1_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit30.Q ));
 sg13g2_dlhq_1 _1419_ (.D(Tile_X0Y1_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit29.Q ));
 sg13g2_dlhq_1 _1420_ (.D(Tile_X0Y1_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit28.Q ));
 sg13g2_dlhq_1 _1421_ (.D(Tile_X0Y1_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit27.Q ));
 sg13g2_dlhq_1 _1422_ (.D(Tile_X0Y1_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit26.Q ));
 sg13g2_dlhq_1 _1423_ (.D(Tile_X0Y1_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit25.Q ));
 sg13g2_dlhq_1 _1424_ (.D(Tile_X0Y1_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit24.Q ));
 sg13g2_dlhq_1 _1425_ (.D(Tile_X0Y1_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit23.Q ));
 sg13g2_dlhq_1 _1426_ (.D(Tile_X0Y1_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit22.Q ));
 sg13g2_dlhq_1 _1427_ (.D(Tile_X0Y1_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit21.Q ));
 sg13g2_dlhq_1 _1428_ (.D(Tile_X0Y1_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit20.Q ));
 sg13g2_dlhq_1 _1429_ (.D(Tile_X0Y1_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit19.Q ));
 sg13g2_dlhq_1 _1430_ (.D(Tile_X0Y1_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit18.Q ));
 sg13g2_dlhq_1 _1431_ (.D(Tile_X0Y1_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit17.Q ));
 sg13g2_dlhq_1 _1432_ (.D(Tile_X0Y1_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit16.Q ));
 sg13g2_dlhq_1 _1433_ (.D(Tile_X0Y1_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit15.Q ));
 sg13g2_dlhq_1 _1434_ (.D(Tile_X0Y1_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit14.Q ));
 sg13g2_dlhq_1 _1435_ (.D(Tile_X0Y1_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit13.Q ));
 sg13g2_dlhq_1 _1436_ (.D(Tile_X0Y1_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit12.Q ));
 sg13g2_dlhq_1 _1437_ (.D(Tile_X0Y1_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q ));
 sg13g2_dlhq_1 _1438_ (.D(Tile_X0Y1_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit10.Q ));
 sg13g2_dlhq_1 _1439_ (.D(Tile_X0Y1_FrameData[9]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit9.Q ));
 sg13g2_dlhq_1 _1440_ (.D(Tile_X0Y1_FrameData[8]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q ));
 sg13g2_dlhq_1 _1441_ (.D(Tile_X0Y1_FrameData[7]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit7.Q ));
 sg13g2_dlhq_1 _1442_ (.D(Tile_X0Y1_FrameData[6]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit6.Q ));
 sg13g2_dlhq_1 _1443_ (.D(Tile_X0Y1_FrameData[5]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit5.Q ));
 sg13g2_dlhq_1 _1444_ (.D(Tile_X0Y1_FrameData[4]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit4.Q ));
 sg13g2_dlhq_1 _1445_ (.D(Tile_X0Y1_FrameData[3]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit3.Q ));
 sg13g2_dlhq_1 _1446_ (.D(Tile_X0Y1_FrameData[2]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit2.Q ));
 sg13g2_dlhq_1 _1447_ (.D(Tile_X0Y1_FrameData[1]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit1.Q ));
 sg13g2_dlhq_1 _1448_ (.D(Tile_X0Y1_FrameData[0]),
    .GATE(Tile_X0Y1_FrameStrobe[8]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit0.Q ));
 sg13g2_dlhq_1 _1449_ (.D(Tile_X0Y1_FrameData[31]),
    .GATE(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit31.Q ));
 sg13g2_dlhq_1 _1450_ (.D(Tile_X0Y1_FrameData[30]),
    .GATE(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit30.Q ));
 sg13g2_dlhq_1 _1451_ (.D(Tile_X0Y1_FrameData[29]),
    .GATE(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit29.Q ));
 sg13g2_dlhq_1 _1452_ (.D(Tile_X0Y1_FrameData[28]),
    .GATE(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit28.Q ));
 sg13g2_dlhq_1 _1453_ (.D(Tile_X0Y1_FrameData[27]),
    .GATE(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit27.Q ));
 sg13g2_dlhq_1 _1454_ (.D(Tile_X0Y1_FrameData[26]),
    .GATE(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit26.Q ));
 sg13g2_dlhq_1 _1455_ (.D(Tile_X0Y1_FrameData[25]),
    .GATE(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit25.Q ));
 sg13g2_dlhq_1 _1456_ (.D(Tile_X0Y1_FrameData[24]),
    .GATE(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit24.Q ));
 sg13g2_dlhq_1 _1457_ (.D(Tile_X0Y1_FrameData[23]),
    .GATE(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit23.Q ));
 sg13g2_dlhq_1 _1458_ (.D(Tile_X0Y1_FrameData[22]),
    .GATE(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit22.Q ));
 sg13g2_dlhq_1 _1459_ (.D(Tile_X0Y1_FrameData[21]),
    .GATE(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit21.Q ));
 sg13g2_dlhq_1 _1460_ (.D(Tile_X0Y1_FrameData[20]),
    .GATE(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit20.Q ));
 sg13g2_dlhq_1 _1461_ (.D(Tile_X0Y1_FrameData[19]),
    .GATE(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit19.Q ));
 sg13g2_dlhq_1 _1462_ (.D(Tile_X0Y1_FrameData[18]),
    .GATE(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit18.Q ));
 sg13g2_dlhq_1 _1463_ (.D(Tile_X0Y1_FrameData[17]),
    .GATE(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit17.Q ));
 sg13g2_dlhq_1 _1464_ (.D(Tile_X0Y1_FrameData[16]),
    .GATE(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit16.Q ));
 sg13g2_dlhq_1 _1465_ (.D(Tile_X0Y1_FrameData[15]),
    .GATE(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit15.Q ));
 sg13g2_dlhq_1 _1466_ (.D(Tile_X0Y1_FrameData[14]),
    .GATE(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit14.Q ));
 sg13g2_dlhq_1 _1467_ (.D(Tile_X0Y1_FrameData[13]),
    .GATE(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit13.Q ));
 sg13g2_dlhq_1 _1468_ (.D(Tile_X0Y1_FrameData[12]),
    .GATE(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit12.Q ));
 sg13g2_dlhq_1 _1469_ (.D(Tile_X0Y1_FrameData[11]),
    .GATE(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit11.Q ));
 sg13g2_dlhq_1 _1470_ (.D(Tile_X0Y1_FrameData[10]),
    .GATE(Tile_X0Y1_FrameStrobe[9]),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit10.Q ));
 sg13g2_tiehi _1471_ (.L_HI(TIE_HIGH_SRAM));
 sg13g2_tielo _1472_ (.L_LO(TIE_LOW_SRAM));
 sg13g2_buf_1 _1473_ (.A(clknet_1_0__leaf_Tile_X0Y1_UserCLK),
    .X(CLK_SRAM));
 sg13g2_buf_1 _1474_ (.A(Tile_X0Y0_FrameData[0]),
    .X(Tile_X0Y0_FrameData_O[0]));
 sg13g2_buf_1 _1475_ (.A(Tile_X0Y0_FrameData[1]),
    .X(Tile_X0Y0_FrameData_O[1]));
 sg13g2_buf_1 _1476_ (.A(Tile_X0Y0_FrameData[2]),
    .X(Tile_X0Y0_FrameData_O[2]));
 sg13g2_buf_1 _1477_ (.A(Tile_X0Y0_FrameData[3]),
    .X(Tile_X0Y0_FrameData_O[3]));
 sg13g2_buf_1 _1478_ (.A(Tile_X0Y0_FrameData[4]),
    .X(Tile_X0Y0_FrameData_O[4]));
 sg13g2_buf_1 _1479_ (.A(Tile_X0Y0_FrameData[5]),
    .X(Tile_X0Y0_FrameData_O[5]));
 sg13g2_buf_1 _1480_ (.A(Tile_X0Y0_FrameData[6]),
    .X(Tile_X0Y0_FrameData_O[6]));
 sg13g2_buf_1 _1481_ (.A(Tile_X0Y0_FrameData[7]),
    .X(Tile_X0Y0_FrameData_O[7]));
 sg13g2_buf_1 _1482_ (.A(Tile_X0Y0_FrameData[8]),
    .X(Tile_X0Y0_FrameData_O[8]));
 sg13g2_buf_1 _1483_ (.A(Tile_X0Y0_FrameData[9]),
    .X(Tile_X0Y0_FrameData_O[9]));
 sg13g2_buf_1 _1484_ (.A(Tile_X0Y0_FrameData[10]),
    .X(Tile_X0Y0_FrameData_O[10]));
 sg13g2_buf_1 _1485_ (.A(Tile_X0Y0_FrameData[11]),
    .X(Tile_X0Y0_FrameData_O[11]));
 sg13g2_buf_1 _1486_ (.A(Tile_X0Y0_FrameData[12]),
    .X(Tile_X0Y0_FrameData_O[12]));
 sg13g2_buf_1 _1487_ (.A(Tile_X0Y0_FrameData[13]),
    .X(Tile_X0Y0_FrameData_O[13]));
 sg13g2_buf_1 _1488_ (.A(Tile_X0Y0_FrameData[14]),
    .X(Tile_X0Y0_FrameData_O[14]));
 sg13g2_buf_1 _1489_ (.A(Tile_X0Y0_FrameData[15]),
    .X(Tile_X0Y0_FrameData_O[15]));
 sg13g2_buf_1 _1490_ (.A(Tile_X0Y0_FrameData[16]),
    .X(Tile_X0Y0_FrameData_O[16]));
 sg13g2_buf_1 _1491_ (.A(Tile_X0Y0_FrameData[17]),
    .X(Tile_X0Y0_FrameData_O[17]));
 sg13g2_buf_1 _1492_ (.A(Tile_X0Y0_FrameData[18]),
    .X(Tile_X0Y0_FrameData_O[18]));
 sg13g2_buf_1 _1493_ (.A(Tile_X0Y0_FrameData[19]),
    .X(Tile_X0Y0_FrameData_O[19]));
 sg13g2_buf_1 _1494_ (.A(Tile_X0Y0_FrameData[20]),
    .X(Tile_X0Y0_FrameData_O[20]));
 sg13g2_buf_1 _1495_ (.A(Tile_X0Y0_FrameData[21]),
    .X(Tile_X0Y0_FrameData_O[21]));
 sg13g2_buf_1 _1496_ (.A(Tile_X0Y0_FrameData[22]),
    .X(Tile_X0Y0_FrameData_O[22]));
 sg13g2_buf_1 _1497_ (.A(Tile_X0Y0_FrameData[23]),
    .X(Tile_X0Y0_FrameData_O[23]));
 sg13g2_buf_1 _1498_ (.A(Tile_X0Y0_FrameData[24]),
    .X(Tile_X0Y0_FrameData_O[24]));
 sg13g2_buf_1 _1499_ (.A(Tile_X0Y0_FrameData[25]),
    .X(Tile_X0Y0_FrameData_O[25]));
 sg13g2_buf_1 _1500_ (.A(Tile_X0Y0_FrameData[26]),
    .X(Tile_X0Y0_FrameData_O[26]));
 sg13g2_buf_1 _1501_ (.A(Tile_X0Y0_FrameData[27]),
    .X(Tile_X0Y0_FrameData_O[27]));
 sg13g2_buf_1 _1502_ (.A(Tile_X0Y0_FrameData[28]),
    .X(Tile_X0Y0_FrameData_O[28]));
 sg13g2_buf_1 _1503_ (.A(Tile_X0Y0_FrameData[29]),
    .X(Tile_X0Y0_FrameData_O[29]));
 sg13g2_buf_1 _1504_ (.A(Tile_X0Y0_FrameData[30]),
    .X(Tile_X0Y0_FrameData_O[30]));
 sg13g2_buf_1 _1505_ (.A(Tile_X0Y0_FrameData[31]),
    .X(Tile_X0Y0_FrameData_O[31]));
 sg13g2_buf_1 _1506_ (.A(Tile_X0Y1_FrameStrobe[0]),
    .X(Tile_X0Y0_FrameStrobe_O[0]));
 sg13g2_buf_1 _1507_ (.A(Tile_X0Y1_FrameStrobe[1]),
    .X(Tile_X0Y0_FrameStrobe_O[1]));
 sg13g2_buf_1 _1508_ (.A(Tile_X0Y1_FrameStrobe[2]),
    .X(Tile_X0Y0_FrameStrobe_O[2]));
 sg13g2_buf_1 _1509_ (.A(Tile_X0Y1_FrameStrobe[3]),
    .X(Tile_X0Y0_FrameStrobe_O[3]));
 sg13g2_buf_1 _1510_ (.A(Tile_X0Y1_FrameStrobe[4]),
    .X(Tile_X0Y0_FrameStrobe_O[4]));
 sg13g2_buf_1 _1511_ (.A(Tile_X0Y1_FrameStrobe[5]),
    .X(Tile_X0Y0_FrameStrobe_O[5]));
 sg13g2_buf_1 _1512_ (.A(Tile_X0Y1_FrameStrobe[6]),
    .X(Tile_X0Y0_FrameStrobe_O[6]));
 sg13g2_buf_1 _1513_ (.A(Tile_X0Y1_FrameStrobe[7]),
    .X(Tile_X0Y0_FrameStrobe_O[7]));
 sg13g2_buf_1 _1514_ (.A(Tile_X0Y1_FrameStrobe[8]),
    .X(Tile_X0Y0_FrameStrobe_O[8]));
 sg13g2_buf_1 _1515_ (.A(Tile_X0Y1_FrameStrobe[9]),
    .X(Tile_X0Y0_FrameStrobe_O[9]));
 sg13g2_buf_1 _1516_ (.A(Tile_X0Y1_FrameStrobe[10]),
    .X(Tile_X0Y0_FrameStrobe_O[10]));
 sg13g2_buf_1 _1517_ (.A(Tile_X0Y1_FrameStrobe[11]),
    .X(Tile_X0Y0_FrameStrobe_O[11]));
 sg13g2_buf_1 _1518_ (.A(Tile_X0Y1_FrameStrobe[12]),
    .X(Tile_X0Y0_FrameStrobe_O[12]));
 sg13g2_buf_1 _1519_ (.A(Tile_X0Y1_FrameStrobe[13]),
    .X(Tile_X0Y0_FrameStrobe_O[13]));
 sg13g2_buf_1 _1520_ (.A(Tile_X0Y1_FrameStrobe[14]),
    .X(Tile_X0Y0_FrameStrobe_O[14]));
 sg13g2_buf_1 _1521_ (.A(Tile_X0Y1_FrameStrobe[15]),
    .X(Tile_X0Y0_FrameStrobe_O[15]));
 sg13g2_buf_1 _1522_ (.A(Tile_X0Y1_FrameStrobe[16]),
    .X(Tile_X0Y0_FrameStrobe_O[16]));
 sg13g2_buf_1 _1523_ (.A(Tile_X0Y1_FrameStrobe[17]),
    .X(Tile_X0Y0_FrameStrobe_O[17]));
 sg13g2_buf_1 _1524_ (.A(Tile_X0Y1_FrameStrobe[18]),
    .X(Tile_X0Y0_FrameStrobe_O[18]));
 sg13g2_buf_1 _1525_ (.A(Tile_X0Y1_FrameStrobe[19]),
    .X(Tile_X0Y0_FrameStrobe_O[19]));
 sg13g2_buf_1 _1526_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG0 ),
    .X(Tile_X0Y0_N1BEG[0]));
 sg13g2_buf_1 _1527_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG1 ),
    .X(Tile_X0Y0_N1BEG[1]));
 sg13g2_buf_1 _1528_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG2 ),
    .X(Tile_X0Y0_N1BEG[2]));
 sg13g2_buf_1 _1529_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG3 ),
    .X(Tile_X0Y0_N1BEG[3]));
 sg13g2_buf_1 _1530_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG0 ),
    .X(Tile_X0Y0_N2BEG[0]));
 sg13g2_buf_1 _1531_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG1 ),
    .X(Tile_X0Y0_N2BEG[1]));
 sg13g2_buf_1 _1532_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG2 ),
    .X(Tile_X0Y0_N2BEG[2]));
 sg13g2_buf_1 _1533_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG3 ),
    .X(Tile_X0Y0_N2BEG[3]));
 sg13g2_buf_1 _1534_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG4 ),
    .X(Tile_X0Y0_N2BEG[4]));
 sg13g2_buf_1 _1535_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG5 ),
    .X(Tile_X0Y0_N2BEG[5]));
 sg13g2_buf_1 _1536_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG6 ),
    .X(Tile_X0Y0_N2BEG[6]));
 sg13g2_buf_1 _1537_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG7 ),
    .X(Tile_X0Y0_N2BEG[7]));
 sg13g2_buf_1 _1538_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb0 ),
    .X(Tile_X0Y0_N2BEGb[0]));
 sg13g2_buf_1 _1539_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb1 ),
    .X(Tile_X0Y0_N2BEGb[1]));
 sg13g2_buf_1 _1540_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb2 ),
    .X(Tile_X0Y0_N2BEGb[2]));
 sg13g2_buf_1 _1541_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb3 ),
    .X(Tile_X0Y0_N2BEGb[3]));
 sg13g2_buf_1 _1542_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb4 ),
    .X(Tile_X0Y0_N2BEGb[4]));
 sg13g2_buf_1 _1543_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb5 ),
    .X(Tile_X0Y0_N2BEGb[5]));
 sg13g2_buf_1 _1544_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb6 ),
    .X(Tile_X0Y0_N2BEGb[6]));
 sg13g2_buf_1 _1545_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb7 ),
    .X(Tile_X0Y0_N2BEGb[7]));
 sg13g2_buf_1 _1546_ (.A(Tile_X0Y1_N4END[8]),
    .X(Tile_X0Y0_N4BEG[0]));
 sg13g2_buf_1 _1547_ (.A(Tile_X0Y1_N4END[9]),
    .X(Tile_X0Y0_N4BEG[1]));
 sg13g2_buf_1 _1548_ (.A(Tile_X0Y1_N4END[10]),
    .X(Tile_X0Y0_N4BEG[2]));
 sg13g2_buf_1 _1549_ (.A(Tile_X0Y1_N4END[11]),
    .X(Tile_X0Y0_N4BEG[3]));
 sg13g2_buf_1 _1550_ (.A(Tile_X0Y1_N4END[12]),
    .X(Tile_X0Y0_N4BEG[4]));
 sg13g2_buf_1 _1551_ (.A(Tile_X0Y1_N4END[13]),
    .X(Tile_X0Y0_N4BEG[5]));
 sg13g2_buf_1 _1552_ (.A(Tile_X0Y1_N4END[14]),
    .X(Tile_X0Y0_N4BEG[6]));
 sg13g2_buf_1 _1553_ (.A(Tile_X0Y1_N4END[15]),
    .X(Tile_X0Y0_N4BEG[7]));
 sg13g2_buf_1 _1554_ (.A(\Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_8.A ),
    .X(Tile_X0Y0_N4BEG[8]));
 sg13g2_buf_1 _1555_ (.A(\Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_9.A ),
    .X(Tile_X0Y0_N4BEG[9]));
 sg13g2_buf_1 _1556_ (.A(\Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_10.A ),
    .X(Tile_X0Y0_N4BEG[10]));
 sg13g2_buf_1 _1557_ (.A(\Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_11.A ),
    .X(Tile_X0Y0_N4BEG[11]));
 sg13g2_buf_1 _1558_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG0 ),
    .X(Tile_X0Y0_N4BEG[12]));
 sg13g2_buf_1 _1559_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG1 ),
    .X(Tile_X0Y0_N4BEG[13]));
 sg13g2_buf_1 _1560_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG2 ),
    .X(Tile_X0Y0_N4BEG[14]));
 sg13g2_buf_1 _1561_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG3 ),
    .X(Tile_X0Y0_N4BEG[15]));
 sg13g2_buf_1 _1562_ (.A(clknet_1_1__leaf_Tile_X0Y1_UserCLK),
    .X(Tile_X0Y0_UserCLKo));
 sg13g2_buf_1 _1563_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG0 ),
    .X(Tile_X0Y0_W1BEG[0]));
 sg13g2_buf_1 _1564_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG1 ),
    .X(Tile_X0Y0_W1BEG[1]));
 sg13g2_buf_1 _1565_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG2 ),
    .X(Tile_X0Y0_W1BEG[2]));
 sg13g2_buf_1 _1566_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG3 ),
    .X(Tile_X0Y0_W1BEG[3]));
 sg13g2_buf_1 _1567_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG0 ),
    .X(Tile_X0Y0_W2BEG[0]));
 sg13g2_buf_1 _1568_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG1 ),
    .X(Tile_X0Y0_W2BEG[1]));
 sg13g2_buf_1 _1569_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG2 ),
    .X(Tile_X0Y0_W2BEG[2]));
 sg13g2_buf_1 _1570_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG3 ),
    .X(Tile_X0Y0_W2BEG[3]));
 sg13g2_buf_1 _1571_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG4 ),
    .X(Tile_X0Y0_W2BEG[4]));
 sg13g2_buf_1 _1572_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG5 ),
    .X(Tile_X0Y0_W2BEG[5]));
 sg13g2_buf_1 _1573_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG6 ),
    .X(Tile_X0Y0_W2BEG[6]));
 sg13g2_buf_1 _1574_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG7 ),
    .X(Tile_X0Y0_W2BEG[7]));
 sg13g2_buf_1 _1575_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb0 ),
    .X(Tile_X0Y0_W2BEGb[0]));
 sg13g2_buf_1 _1576_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb1 ),
    .X(Tile_X0Y0_W2BEGb[1]));
 sg13g2_buf_1 _1577_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb2 ),
    .X(Tile_X0Y0_W2BEGb[2]));
 sg13g2_buf_1 _1578_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb3 ),
    .X(Tile_X0Y0_W2BEGb[3]));
 sg13g2_buf_1 _1579_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb4 ),
    .X(Tile_X0Y0_W2BEGb[4]));
 sg13g2_buf_1 _1580_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb5 ),
    .X(Tile_X0Y0_W2BEGb[5]));
 sg13g2_buf_1 _1581_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb6 ),
    .X(Tile_X0Y0_W2BEGb[6]));
 sg13g2_buf_1 _1582_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb7 ),
    .X(Tile_X0Y0_W2BEGb[7]));
 sg13g2_buf_1 _1583_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG0 ),
    .X(Tile_X0Y0_W6BEG[0]));
 sg13g2_buf_1 _1584_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG1 ),
    .X(Tile_X0Y0_W6BEG[1]));
 sg13g2_buf_1 _1585_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG2 ),
    .X(Tile_X0Y0_W6BEG[2]));
 sg13g2_buf_1 _1586_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG3 ),
    .X(Tile_X0Y0_W6BEG[3]));
 sg13g2_buf_1 _1587_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG4 ),
    .X(Tile_X0Y0_W6BEG[4]));
 sg13g2_buf_1 _1588_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG5 ),
    .X(Tile_X0Y0_W6BEG[5]));
 sg13g2_buf_1 _1589_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG6 ),
    .X(Tile_X0Y0_W6BEG[6]));
 sg13g2_buf_1 _1590_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG7 ),
    .X(Tile_X0Y0_W6BEG[7]));
 sg13g2_buf_1 _1591_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG8 ),
    .X(Tile_X0Y0_W6BEG[8]));
 sg13g2_buf_1 _1592_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG9 ),
    .X(Tile_X0Y0_W6BEG[9]));
 sg13g2_buf_1 _1593_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG10 ),
    .X(Tile_X0Y0_W6BEG[10]));
 sg13g2_buf_1 _1594_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG11 ),
    .X(Tile_X0Y0_W6BEG[11]));
 sg13g2_buf_1 _1595_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG0 ),
    .X(Tile_X0Y0_WW4BEG[0]));
 sg13g2_buf_1 _1596_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG1 ),
    .X(Tile_X0Y0_WW4BEG[1]));
 sg13g2_buf_1 _1597_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG2 ),
    .X(Tile_X0Y0_WW4BEG[2]));
 sg13g2_buf_1 _1598_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG3 ),
    .X(Tile_X0Y0_WW4BEG[3]));
 sg13g2_buf_1 _1599_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG4 ),
    .X(Tile_X0Y0_WW4BEG[4]));
 sg13g2_buf_1 _1600_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG5 ),
    .X(Tile_X0Y0_WW4BEG[5]));
 sg13g2_buf_1 _1601_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG6 ),
    .X(Tile_X0Y0_WW4BEG[6]));
 sg13g2_buf_1 _1602_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG7 ),
    .X(Tile_X0Y0_WW4BEG[7]));
 sg13g2_buf_1 _1603_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG8 ),
    .X(Tile_X0Y0_WW4BEG[8]));
 sg13g2_buf_1 _1604_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG9 ),
    .X(Tile_X0Y0_WW4BEG[9]));
 sg13g2_buf_1 _1605_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG10 ),
    .X(Tile_X0Y0_WW4BEG[10]));
 sg13g2_buf_1 _1606_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG11 ),
    .X(Tile_X0Y0_WW4BEG[11]));
 sg13g2_buf_1 _1607_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG12 ),
    .X(Tile_X0Y0_WW4BEG[12]));
 sg13g2_buf_1 _1608_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG13 ),
    .X(Tile_X0Y0_WW4BEG[13]));
 sg13g2_buf_1 _1609_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG14 ),
    .X(Tile_X0Y0_WW4BEG[14]));
 sg13g2_buf_1 _1610_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG15 ),
    .X(Tile_X0Y0_WW4BEG[15]));
 sg13g2_buf_1 _1611_ (.A(Tile_X0Y1_FrameData[0]),
    .X(Tile_X0Y1_FrameData_O[0]));
 sg13g2_buf_1 _1612_ (.A(Tile_X0Y1_FrameData[1]),
    .X(Tile_X0Y1_FrameData_O[1]));
 sg13g2_buf_1 _1613_ (.A(Tile_X0Y1_FrameData[2]),
    .X(Tile_X0Y1_FrameData_O[2]));
 sg13g2_buf_1 _1614_ (.A(Tile_X0Y1_FrameData[3]),
    .X(Tile_X0Y1_FrameData_O[3]));
 sg13g2_buf_1 _1615_ (.A(Tile_X0Y1_FrameData[4]),
    .X(Tile_X0Y1_FrameData_O[4]));
 sg13g2_buf_1 _1616_ (.A(Tile_X0Y1_FrameData[5]),
    .X(Tile_X0Y1_FrameData_O[5]));
 sg13g2_buf_1 _1617_ (.A(Tile_X0Y1_FrameData[6]),
    .X(Tile_X0Y1_FrameData_O[6]));
 sg13g2_buf_1 _1618_ (.A(Tile_X0Y1_FrameData[7]),
    .X(Tile_X0Y1_FrameData_O[7]));
 sg13g2_buf_1 _1619_ (.A(Tile_X0Y1_FrameData[8]),
    .X(Tile_X0Y1_FrameData_O[8]));
 sg13g2_buf_1 _1620_ (.A(Tile_X0Y1_FrameData[9]),
    .X(Tile_X0Y1_FrameData_O[9]));
 sg13g2_buf_1 _1621_ (.A(Tile_X0Y1_FrameData[10]),
    .X(Tile_X0Y1_FrameData_O[10]));
 sg13g2_buf_1 _1622_ (.A(Tile_X0Y1_FrameData[11]),
    .X(Tile_X0Y1_FrameData_O[11]));
 sg13g2_buf_1 _1623_ (.A(Tile_X0Y1_FrameData[12]),
    .X(Tile_X0Y1_FrameData_O[12]));
 sg13g2_buf_1 _1624_ (.A(Tile_X0Y1_FrameData[13]),
    .X(Tile_X0Y1_FrameData_O[13]));
 sg13g2_buf_1 _1625_ (.A(Tile_X0Y1_FrameData[14]),
    .X(Tile_X0Y1_FrameData_O[14]));
 sg13g2_buf_1 _1626_ (.A(Tile_X0Y1_FrameData[15]),
    .X(Tile_X0Y1_FrameData_O[15]));
 sg13g2_buf_1 _1627_ (.A(Tile_X0Y1_FrameData[16]),
    .X(Tile_X0Y1_FrameData_O[16]));
 sg13g2_buf_1 _1628_ (.A(Tile_X0Y1_FrameData[17]),
    .X(Tile_X0Y1_FrameData_O[17]));
 sg13g2_buf_1 _1629_ (.A(Tile_X0Y1_FrameData[18]),
    .X(Tile_X0Y1_FrameData_O[18]));
 sg13g2_buf_1 _1630_ (.A(Tile_X0Y1_FrameData[19]),
    .X(Tile_X0Y1_FrameData_O[19]));
 sg13g2_buf_1 _1631_ (.A(Tile_X0Y1_FrameData[20]),
    .X(Tile_X0Y1_FrameData_O[20]));
 sg13g2_buf_1 _1632_ (.A(Tile_X0Y1_FrameData[21]),
    .X(Tile_X0Y1_FrameData_O[21]));
 sg13g2_buf_1 _1633_ (.A(Tile_X0Y1_FrameData[22]),
    .X(Tile_X0Y1_FrameData_O[22]));
 sg13g2_buf_1 _1634_ (.A(Tile_X0Y1_FrameData[23]),
    .X(Tile_X0Y1_FrameData_O[23]));
 sg13g2_buf_1 _1635_ (.A(Tile_X0Y1_FrameData[24]),
    .X(Tile_X0Y1_FrameData_O[24]));
 sg13g2_buf_1 _1636_ (.A(Tile_X0Y1_FrameData[25]),
    .X(Tile_X0Y1_FrameData_O[25]));
 sg13g2_buf_1 _1637_ (.A(Tile_X0Y1_FrameData[26]),
    .X(Tile_X0Y1_FrameData_O[26]));
 sg13g2_buf_1 _1638_ (.A(Tile_X0Y1_FrameData[27]),
    .X(Tile_X0Y1_FrameData_O[27]));
 sg13g2_buf_1 _1639_ (.A(Tile_X0Y1_FrameData[28]),
    .X(Tile_X0Y1_FrameData_O[28]));
 sg13g2_buf_1 _1640_ (.A(Tile_X0Y1_FrameData[29]),
    .X(Tile_X0Y1_FrameData_O[29]));
 sg13g2_buf_1 _1641_ (.A(Tile_X0Y1_FrameData[30]),
    .X(Tile_X0Y1_FrameData_O[30]));
 sg13g2_buf_1 _1642_ (.A(Tile_X0Y1_FrameData[31]),
    .X(Tile_X0Y1_FrameData_O[31]));
 sg13g2_buf_1 _1643_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG0 ),
    .X(Tile_X0Y1_S1BEG[0]));
 sg13g2_buf_1 _1644_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG1 ),
    .X(Tile_X0Y1_S1BEG[1]));
 sg13g2_buf_1 _1645_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG2 ),
    .X(Tile_X0Y1_S1BEG[2]));
 sg13g2_buf_1 _1646_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG3 ),
    .X(Tile_X0Y1_S1BEG[3]));
 sg13g2_buf_1 _1647_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG0 ),
    .X(Tile_X0Y1_S2BEG[0]));
 sg13g2_buf_1 _1648_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG1 ),
    .X(Tile_X0Y1_S2BEG[1]));
 sg13g2_buf_1 _1649_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG2 ),
    .X(Tile_X0Y1_S2BEG[2]));
 sg13g2_buf_1 _1650_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG3 ),
    .X(Tile_X0Y1_S2BEG[3]));
 sg13g2_buf_1 _1651_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG4 ),
    .X(Tile_X0Y1_S2BEG[4]));
 sg13g2_buf_1 _1652_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG5 ),
    .X(Tile_X0Y1_S2BEG[5]));
 sg13g2_buf_1 _1653_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG6 ),
    .X(Tile_X0Y1_S2BEG[6]));
 sg13g2_buf_1 _1654_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG7 ),
    .X(Tile_X0Y1_S2BEG[7]));
 sg13g2_buf_1 _1655_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG0 ),
    .X(Tile_X0Y1_S2BEGb[0]));
 sg13g2_buf_1 _1656_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG1 ),
    .X(Tile_X0Y1_S2BEGb[1]));
 sg13g2_buf_1 _1657_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG2 ),
    .X(Tile_X0Y1_S2BEGb[2]));
 sg13g2_buf_1 _1658_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG3 ),
    .X(Tile_X0Y1_S2BEGb[3]));
 sg13g2_buf_1 _1659_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG4 ),
    .X(Tile_X0Y1_S2BEGb[4]));
 sg13g2_buf_1 _1660_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG5 ),
    .X(Tile_X0Y1_S2BEGb[5]));
 sg13g2_buf_1 _1661_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG6 ),
    .X(Tile_X0Y1_S2BEGb[6]));
 sg13g2_buf_1 _1662_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG7 ),
    .X(Tile_X0Y1_S2BEGb[7]));
 sg13g2_buf_1 _1663_ (.A(Tile_X0Y0_S4END[8]),
    .X(Tile_X0Y1_S4BEG[0]));
 sg13g2_buf_1 _1664_ (.A(Tile_X0Y0_S4END[9]),
    .X(Tile_X0Y1_S4BEG[1]));
 sg13g2_buf_1 _1665_ (.A(Tile_X0Y0_S4END[10]),
    .X(Tile_X0Y1_S4BEG[2]));
 sg13g2_buf_1 _1666_ (.A(Tile_X0Y0_S4END[11]),
    .X(Tile_X0Y1_S4BEG[3]));
 sg13g2_buf_1 _1667_ (.A(Tile_X0Y0_S4END[12]),
    .X(Tile_X0Y1_S4BEG[4]));
 sg13g2_buf_1 _1668_ (.A(Tile_X0Y0_S4END[13]),
    .X(Tile_X0Y1_S4BEG[5]));
 sg13g2_buf_1 _1669_ (.A(Tile_X0Y0_S4END[14]),
    .X(Tile_X0Y1_S4BEG[6]));
 sg13g2_buf_1 _1670_ (.A(Tile_X0Y0_S4END[15]),
    .X(Tile_X0Y1_S4BEG[7]));
 sg13g2_buf_1 _1671_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG0 ),
    .X(Tile_X0Y1_S4BEG[8]));
 sg13g2_buf_1 _1672_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG1 ),
    .X(Tile_X0Y1_S4BEG[9]));
 sg13g2_buf_1 _1673_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG2 ),
    .X(Tile_X0Y1_S4BEG[10]));
 sg13g2_buf_1 _1674_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG3 ),
    .X(Tile_X0Y1_S4BEG[11]));
 sg13g2_buf_1 _1675_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG0 ),
    .X(Tile_X0Y1_S4BEG[12]));
 sg13g2_buf_1 _1676_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG1 ),
    .X(Tile_X0Y1_S4BEG[13]));
 sg13g2_buf_1 _1677_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG2 ),
    .X(Tile_X0Y1_S4BEG[14]));
 sg13g2_buf_1 _1678_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG3 ),
    .X(Tile_X0Y1_S4BEG[15]));
 sg13g2_buf_1 _1679_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG0 ),
    .X(Tile_X0Y1_W1BEG[0]));
 sg13g2_buf_1 _1680_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG1 ),
    .X(Tile_X0Y1_W1BEG[1]));
 sg13g2_buf_1 _1681_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG2 ),
    .X(Tile_X0Y1_W1BEG[2]));
 sg13g2_buf_1 _1682_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG3 ),
    .X(Tile_X0Y1_W1BEG[3]));
 sg13g2_buf_1 _1683_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG0 ),
    .X(Tile_X0Y1_W2BEG[0]));
 sg13g2_buf_1 _1684_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG1 ),
    .X(Tile_X0Y1_W2BEG[1]));
 sg13g2_buf_1 _1685_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG2 ),
    .X(Tile_X0Y1_W2BEG[2]));
 sg13g2_buf_1 _1686_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG3 ),
    .X(Tile_X0Y1_W2BEG[3]));
 sg13g2_buf_1 _1687_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG4 ),
    .X(Tile_X0Y1_W2BEG[4]));
 sg13g2_buf_1 _1688_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG5 ),
    .X(Tile_X0Y1_W2BEG[5]));
 sg13g2_buf_1 _1689_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG6 ),
    .X(Tile_X0Y1_W2BEG[6]));
 sg13g2_buf_1 _1690_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG7 ),
    .X(Tile_X0Y1_W2BEG[7]));
 sg13g2_buf_1 _1691_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb0 ),
    .X(Tile_X0Y1_W2BEGb[0]));
 sg13g2_buf_1 _1692_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb1 ),
    .X(Tile_X0Y1_W2BEGb[1]));
 sg13g2_buf_1 _1693_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb2 ),
    .X(Tile_X0Y1_W2BEGb[2]));
 sg13g2_buf_1 _1694_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb3 ),
    .X(Tile_X0Y1_W2BEGb[3]));
 sg13g2_buf_1 _1695_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb4 ),
    .X(Tile_X0Y1_W2BEGb[4]));
 sg13g2_buf_1 _1696_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb5 ),
    .X(Tile_X0Y1_W2BEGb[5]));
 sg13g2_buf_1 _1697_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb6 ),
    .X(Tile_X0Y1_W2BEGb[6]));
 sg13g2_buf_1 _1698_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb7 ),
    .X(Tile_X0Y1_W2BEGb[7]));
 sg13g2_buf_1 _1699_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG0 ),
    .X(Tile_X0Y1_W6BEG[0]));
 sg13g2_buf_1 _1700_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG1 ),
    .X(Tile_X0Y1_W6BEG[1]));
 sg13g2_buf_1 _1701_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG2 ),
    .X(Tile_X0Y1_W6BEG[2]));
 sg13g2_buf_1 _1702_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG3 ),
    .X(Tile_X0Y1_W6BEG[3]));
 sg13g2_buf_1 _1703_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG4 ),
    .X(Tile_X0Y1_W6BEG[4]));
 sg13g2_buf_1 _1704_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG5 ),
    .X(Tile_X0Y1_W6BEG[5]));
 sg13g2_buf_1 _1705_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG6 ),
    .X(Tile_X0Y1_W6BEG[6]));
 sg13g2_buf_1 _1706_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG7 ),
    .X(Tile_X0Y1_W6BEG[7]));
 sg13g2_buf_1 _1707_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG8 ),
    .X(Tile_X0Y1_W6BEG[8]));
 sg13g2_buf_1 _1708_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG9 ),
    .X(Tile_X0Y1_W6BEG[9]));
 sg13g2_buf_1 _1709_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG10 ),
    .X(Tile_X0Y1_W6BEG[10]));
 sg13g2_buf_1 _1710_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG11 ),
    .X(Tile_X0Y1_W6BEG[11]));
 sg13g2_buf_1 _1711_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG0 ),
    .X(Tile_X0Y1_WW4BEG[0]));
 sg13g2_buf_1 _1712_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG1 ),
    .X(Tile_X0Y1_WW4BEG[1]));
 sg13g2_buf_1 _1713_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG2 ),
    .X(Tile_X0Y1_WW4BEG[2]));
 sg13g2_buf_1 _1714_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG3 ),
    .X(Tile_X0Y1_WW4BEG[3]));
 sg13g2_buf_1 _1715_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG4 ),
    .X(Tile_X0Y1_WW4BEG[4]));
 sg13g2_buf_1 _1716_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG5 ),
    .X(Tile_X0Y1_WW4BEG[5]));
 sg13g2_buf_1 _1717_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG6 ),
    .X(Tile_X0Y1_WW4BEG[6]));
 sg13g2_buf_1 _1718_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG7 ),
    .X(Tile_X0Y1_WW4BEG[7]));
 sg13g2_buf_1 _1719_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG8 ),
    .X(Tile_X0Y1_WW4BEG[8]));
 sg13g2_buf_1 _1720_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG9 ),
    .X(Tile_X0Y1_WW4BEG[9]));
 sg13g2_buf_1 _1721_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG10 ),
    .X(Tile_X0Y1_WW4BEG[10]));
 sg13g2_buf_1 _1722_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG11 ),
    .X(Tile_X0Y1_WW4BEG[11]));
 sg13g2_buf_1 _1723_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG12 ),
    .X(Tile_X0Y1_WW4BEG[12]));
 sg13g2_buf_1 _1724_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG13 ),
    .X(Tile_X0Y1_WW4BEG[13]));
 sg13g2_buf_1 _1725_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG14 ),
    .X(Tile_X0Y1_WW4BEG[14]));
 sg13g2_buf_1 _1726_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG15 ),
    .X(Tile_X0Y1_WW4BEG[15]));
 sg13g2_buf_8 clkbuf_0_Tile_X0Y1_UserCLK (.A(Tile_X0Y1_UserCLK),
    .X(clknet_0_Tile_X0Y1_UserCLK));
 sg13g2_buf_8 clkbuf_1_0__f_Tile_X0Y1_UserCLK (.A(clknet_0_Tile_X0Y1_UserCLK),
    .X(clknet_1_0__leaf_Tile_X0Y1_UserCLK));
 sg13g2_buf_8 clkbuf_1_1__f_Tile_X0Y1_UserCLK (.A(clknet_0_Tile_X0Y1_UserCLK),
    .X(clknet_1_1__leaf_Tile_X0Y1_UserCLK));
 sg13g2_antennanp ANTENNA_1 (.A(\Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_9.A ));
 sg13g2_antennanp ANTENNA_2 (.A(Tile_X0Y0_S2MID[3]));
 sg13g2_antennanp ANTENNA_3 (.A(Tile_X0Y0_S2MID[3]));
 sg13g2_antennanp ANTENNA_4 (.A(Tile_X0Y0_S2MID[3]));
 sg13g2_antennanp ANTENNA_5 (.A(Tile_X0Y0_S2MID[3]));
 sg13g2_antennanp ANTENNA_6 (.A(Tile_X0Y0_S2MID[3]));
 sg13g2_antennanp ANTENNA_7 (.A(Tile_X0Y0_S2MID[3]));
 sg13g2_antennanp ANTENNA_8 (.A(Tile_X0Y0_S2MID[4]));
 sg13g2_antennanp ANTENNA_9 (.A(Tile_X0Y0_S2MID[4]));
 sg13g2_antennanp ANTENNA_10 (.A(Tile_X0Y0_S2MID[4]));
 sg13g2_antennanp ANTENNA_11 (.A(Tile_X0Y0_S2MID[4]));
 sg13g2_antennanp ANTENNA_12 (.A(Tile_X0Y0_S2MID[5]));
 sg13g2_antennanp ANTENNA_13 (.A(Tile_X0Y0_S2MID[5]));
 sg13g2_antennanp ANTENNA_14 (.A(Tile_X0Y0_S2MID[5]));
 sg13g2_antennanp ANTENNA_15 (.A(Tile_X0Y1_FrameStrobe[10]));
 sg13g2_antennanp ANTENNA_16 (.A(Tile_X0Y1_FrameStrobe[11]));
 sg13g2_antennanp ANTENNA_17 (.A(Tile_X0Y1_FrameStrobe[12]));
 sg13g2_antennanp ANTENNA_18 (.A(Tile_X0Y1_FrameStrobe[13]));
 sg13g2_antennanp ANTENNA_19 (.A(Tile_X0Y1_FrameStrobe[14]));
 sg13g2_antennanp ANTENNA_20 (.A(Tile_X0Y1_FrameStrobe[16]));
 sg13g2_antennanp ANTENNA_21 (.A(Tile_X0Y1_FrameStrobe[16]));
 sg13g2_antennanp ANTENNA_22 (.A(Tile_X0Y1_FrameStrobe[16]));
 sg13g2_antennanp ANTENNA_23 (.A(Tile_X0Y1_FrameStrobe[17]));
 sg13g2_antennanp ANTENNA_24 (.A(Tile_X0Y1_FrameStrobe[18]));
 sg13g2_antennanp ANTENNA_25 (.A(Tile_X0Y1_FrameStrobe[18]));
 sg13g2_antennanp ANTENNA_26 (.A(Tile_X0Y1_FrameStrobe[18]));
 sg13g2_antennanp ANTENNA_27 (.A(Tile_X0Y1_FrameStrobe[19]));
 sg13g2_antennanp ANTENNA_28 (.A(Tile_X0Y1_N2MID[0]));
 sg13g2_antennanp ANTENNA_29 (.A(Tile_X0Y1_N2MID[0]));
 sg13g2_antennanp ANTENNA_30 (.A(Tile_X0Y1_N2MID[0]));
 sg13g2_antennanp ANTENNA_31 (.A(Tile_X0Y1_N2MID[3]));
 sg13g2_antennanp ANTENNA_32 (.A(Tile_X0Y1_N2MID[3]));
 sg13g2_antennanp ANTENNA_33 (.A(Tile_X0Y1_N2MID[4]));
 sg13g2_antennanp ANTENNA_34 (.A(Tile_X0Y1_N2MID[4]));
 sg13g2_antennanp ANTENNA_35 (.A(Tile_X0Y1_N2MID[5]));
 sg13g2_antennanp ANTENNA_36 (.A(Tile_X0Y1_N2MID[5]));
 sg13g2_antennanp ANTENNA_37 (.A(Tile_X0Y1_N2MID[7]));
 sg13g2_antennanp ANTENNA_38 (.A(Tile_X0Y1_N2MID[7]));
 sg13g2_antennanp ANTENNA_39 (.A(Tile_X0Y1_N2MID[7]));
 sg13g2_antennanp ANTENNA_40 (.A(Tile_X0Y1_N2MID[7]));
 sg13g2_antennanp ANTENNA_41 (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG0 ));
 sg13g2_antennanp ANTENNA_42 (.A(Tile_X0Y0_S2MID[6]));
 sg13g2_antennanp ANTENNA_43 (.A(Tile_X0Y0_S2MID[6]));
 sg13g2_antennanp ANTENNA_44 (.A(Tile_X0Y0_S2MID[6]));
 sg13g2_antennanp ANTENNA_45 (.A(Tile_X0Y0_S2MID[6]));
 sg13g2_antennanp ANTENNA_46 (.A(Tile_X0Y1_FrameStrobe[15]));
 sg13g2_fill_1 FILLER_0_0 ();
 sg13g2_fill_2 FILLER_0_22 ();
 sg13g2_fill_1 FILLER_0_41 ();
 sg13g2_fill_2 FILLER_0_172 ();
 sg13g2_fill_1 FILLER_0_174 ();
 sg13g2_decap_4 FILLER_0_196 ();
 sg13g2_fill_1 FILLER_1_158 ();
 sg13g2_fill_2 FILLER_1_176 ();
 sg13g2_fill_1 FILLER_1_178 ();
 sg13g2_fill_2 FILLER_2_0 ();
 sg13g2_fill_2 FILLER_2_19 ();
 sg13g2_fill_2 FILLER_2_141 ();
 sg13g2_fill_1 FILLER_2_143 ();
 sg13g2_fill_1 FILLER_2_182 ();
 sg13g2_fill_1 FILLER_3_28 ();
 sg13g2_fill_1 FILLER_3_67 ();
 sg13g2_fill_2 FILLER_3_134 ();
 sg13g2_fill_1 FILLER_3_136 ();
 sg13g2_fill_2 FILLER_3_170 ();
 sg13g2_fill_1 FILLER_3_172 ();
 sg13g2_decap_4 FILLER_3_194 ();
 sg13g2_fill_2 FILLER_3_198 ();
 sg13g2_fill_2 FILLER_4_37 ();
 sg13g2_fill_1 FILLER_4_110 ();
 sg13g2_fill_2 FILLER_4_128 ();
 sg13g2_decap_8 FILLER_4_164 ();
 sg13g2_fill_1 FILLER_4_171 ();
 sg13g2_decap_8 FILLER_4_193 ();
 sg13g2_fill_1 FILLER_5_117 ();
 sg13g2_fill_1 FILLER_5_135 ();
 sg13g2_decap_8 FILLER_5_170 ();
 sg13g2_fill_1 FILLER_5_177 ();
 sg13g2_fill_1 FILLER_5_199 ();
 sg13g2_fill_2 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_2 ();
 sg13g2_fill_1 FILLER_6_11 ();
 sg13g2_fill_2 FILLER_6_78 ();
 sg13g2_decap_8 FILLER_6_153 ();
 sg13g2_fill_1 FILLER_6_160 ();
 sg13g2_fill_1 FILLER_6_199 ();
 sg13g2_fill_1 FILLER_7_17 ();
 sg13g2_fill_2 FILLER_7_47 ();
 sg13g2_fill_1 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_fill_2 FILLER_7_140 ();
 sg13g2_decap_4 FILLER_7_176 ();
 sg13g2_fill_2 FILLER_7_197 ();
 sg13g2_fill_1 FILLER_7_199 ();
 sg13g2_fill_2 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_2 ();
 sg13g2_fill_2 FILLER_8_91 ();
 sg13g2_fill_1 FILLER_8_93 ();
 sg13g2_decap_8 FILLER_8_111 ();
 sg13g2_fill_2 FILLER_8_118 ();
 sg13g2_fill_1 FILLER_8_120 ();
 sg13g2_fill_1 FILLER_8_159 ();
 sg13g2_decap_4 FILLER_8_177 ();
 sg13g2_fill_2 FILLER_8_198 ();
 sg13g2_fill_2 FILLER_9_25 ();
 sg13g2_decap_4 FILLER_9_111 ();
 sg13g2_fill_2 FILLER_9_115 ();
 sg13g2_decap_4 FILLER_9_168 ();
 sg13g2_fill_1 FILLER_9_172 ();
 sg13g2_decap_4 FILLER_9_194 ();
 sg13g2_fill_2 FILLER_9_198 ();
 sg13g2_fill_2 FILLER_10_34 ();
 sg13g2_fill_2 FILLER_10_61 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_4 FILLER_10_136 ();
 sg13g2_fill_2 FILLER_10_140 ();
 sg13g2_fill_2 FILLER_10_180 ();
 sg13g2_fill_1 FILLER_10_199 ();
 sg13g2_fill_2 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_43 ();
 sg13g2_fill_1 FILLER_11_45 ();
 sg13g2_decap_8 FILLER_11_80 ();
 sg13g2_fill_2 FILLER_11_87 ();
 sg13g2_fill_1 FILLER_11_89 ();
 sg13g2_decap_4 FILLER_11_132 ();
 sg13g2_fill_1 FILLER_11_136 ();
 sg13g2_decap_4 FILLER_11_154 ();
 sg13g2_fill_1 FILLER_11_158 ();
 sg13g2_fill_2 FILLER_11_197 ();
 sg13g2_fill_1 FILLER_11_199 ();
 sg13g2_fill_2 FILLER_12_21 ();
 sg13g2_fill_1 FILLER_12_23 ();
 sg13g2_fill_1 FILLER_12_45 ();
 sg13g2_decap_8 FILLER_12_67 ();
 sg13g2_decap_4 FILLER_12_74 ();
 sg13g2_decap_8 FILLER_12_95 ();
 sg13g2_fill_2 FILLER_12_102 ();
 sg13g2_fill_1 FILLER_12_104 ();
 sg13g2_fill_1 FILLER_12_122 ();
 sg13g2_fill_1 FILLER_12_140 ();
 sg13g2_fill_1 FILLER_12_175 ();
 sg13g2_fill_2 FILLER_12_197 ();
 sg13g2_fill_1 FILLER_12_199 ();
 sg13g2_fill_2 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_2 ();
 sg13g2_fill_2 FILLER_13_11 ();
 sg13g2_fill_1 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_64 ();
 sg13g2_decap_4 FILLER_13_71 ();
 sg13g2_fill_1 FILLER_13_75 ();
 sg13g2_fill_2 FILLER_13_114 ();
 sg13g2_fill_1 FILLER_13_116 ();
 sg13g2_decap_8 FILLER_13_142 ();
 sg13g2_fill_1 FILLER_13_149 ();
 sg13g2_decap_8 FILLER_13_171 ();
 sg13g2_decap_4 FILLER_13_178 ();
 sg13g2_fill_1 FILLER_13_199 ();
 sg13g2_fill_1 FILLER_14_29 ();
 sg13g2_decap_8 FILLER_14_68 ();
 sg13g2_fill_1 FILLER_14_96 ();
 sg13g2_fill_1 FILLER_14_118 ();
 sg13g2_fill_2 FILLER_14_136 ();
 sg13g2_decap_8 FILLER_14_159 ();
 sg13g2_fill_1 FILLER_14_166 ();
 sg13g2_decap_8 FILLER_14_184 ();
 sg13g2_decap_8 FILLER_14_191 ();
 sg13g2_fill_2 FILLER_14_198 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_2 ();
 sg13g2_fill_1 FILLER_15_15 ();
 sg13g2_fill_2 FILLER_15_33 ();
 sg13g2_fill_1 FILLER_15_35 ();
 sg13g2_decap_4 FILLER_15_53 ();
 sg13g2_fill_1 FILLER_15_57 ();
 sg13g2_decap_4 FILLER_15_75 ();
 sg13g2_fill_2 FILLER_15_100 ();
 sg13g2_fill_1 FILLER_15_102 ();
 sg13g2_decap_8 FILLER_15_124 ();
 sg13g2_fill_2 FILLER_15_131 ();
 sg13g2_fill_2 FILLER_15_137 ();
 sg13g2_fill_1 FILLER_15_156 ();
 sg13g2_fill_2 FILLER_15_174 ();
 sg13g2_fill_1 FILLER_15_176 ();
 sg13g2_fill_2 FILLER_15_198 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_fill_1 FILLER_16_42 ();
 sg13g2_fill_1 FILLER_16_64 ();
 sg13g2_decap_4 FILLER_16_82 ();
 sg13g2_decap_4 FILLER_16_120 ();
 sg13g2_decap_8 FILLER_16_141 ();
 sg13g2_decap_4 FILLER_16_148 ();
 sg13g2_fill_1 FILLER_16_152 ();
 sg13g2_decap_4 FILLER_16_178 ();
 sg13g2_fill_1 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_17_38 ();
 sg13g2_decap_4 FILLER_17_45 ();
 sg13g2_fill_2 FILLER_17_49 ();
 sg13g2_decap_4 FILLER_17_72 ();
 sg13g2_decap_4 FILLER_17_97 ();
 sg13g2_fill_2 FILLER_17_101 ();
 sg13g2_decap_8 FILLER_17_162 ();
 sg13g2_decap_8 FILLER_17_169 ();
 sg13g2_fill_2 FILLER_17_176 ();
 sg13g2_fill_1 FILLER_17_199 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_2 ();
 sg13g2_fill_1 FILLER_18_7 ();
 sg13g2_fill_2 FILLER_18_29 ();
 sg13g2_fill_2 FILLER_18_48 ();
 sg13g2_decap_8 FILLER_18_67 ();
 sg13g2_fill_1 FILLER_18_74 ();
 sg13g2_decap_4 FILLER_18_92 ();
 sg13g2_fill_1 FILLER_18_96 ();
 sg13g2_decap_8 FILLER_18_114 ();
 sg13g2_fill_2 FILLER_18_121 ();
 sg13g2_fill_1 FILLER_18_123 ();
 sg13g2_fill_2 FILLER_18_141 ();
 sg13g2_fill_1 FILLER_18_143 ();
 sg13g2_fill_1 FILLER_18_169 ();
 sg13g2_decap_4 FILLER_18_195 ();
 sg13g2_fill_1 FILLER_18_199 ();
 sg13g2_decap_4 FILLER_19_21 ();
 sg13g2_fill_1 FILLER_19_25 ();
 sg13g2_fill_2 FILLER_19_77 ();
 sg13g2_decap_4 FILLER_19_96 ();
 sg13g2_fill_2 FILLER_19_100 ();
 sg13g2_fill_2 FILLER_19_174 ();
 sg13g2_fill_2 FILLER_19_198 ();
 sg13g2_decap_8 FILLER_20_4 ();
 sg13g2_fill_2 FILLER_20_11 ();
 sg13g2_fill_1 FILLER_20_13 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_fill_2 FILLER_20_42 ();
 sg13g2_fill_1 FILLER_20_44 ();
 sg13g2_decap_4 FILLER_20_66 ();
 sg13g2_fill_2 FILLER_20_70 ();
 sg13g2_decap_4 FILLER_20_114 ();
 sg13g2_fill_1 FILLER_20_118 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_fill_1 FILLER_20_147 ();
 sg13g2_fill_2 FILLER_20_198 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_7 ();
 sg13g2_fill_1 FILLER_21_9 ();
 sg13g2_decap_8 FILLER_21_31 ();
 sg13g2_fill_2 FILLER_21_38 ();
 sg13g2_fill_1 FILLER_21_40 ();
 sg13g2_decap_4 FILLER_21_79 ();
 sg13g2_decap_4 FILLER_21_100 ();
 sg13g2_fill_1 FILLER_21_104 ();
 sg13g2_decap_4 FILLER_21_122 ();
 sg13g2_decap_8 FILLER_21_143 ();
 sg13g2_fill_1 FILLER_21_150 ();
 sg13g2_decap_8 FILLER_22_17 ();
 sg13g2_decap_8 FILLER_22_24 ();
 sg13g2_fill_2 FILLER_22_31 ();
 sg13g2_decap_8 FILLER_22_50 ();
 sg13g2_decap_4 FILLER_22_57 ();
 sg13g2_decap_8 FILLER_22_99 ();
 sg13g2_decap_8 FILLER_22_106 ();
 sg13g2_decap_8 FILLER_22_113 ();
 sg13g2_decap_8 FILLER_22_120 ();
 sg13g2_decap_4 FILLER_22_144 ();
 sg13g2_decap_4 FILLER_22_165 ();
 sg13g2_fill_2 FILLER_22_169 ();
 sg13g2_fill_1 FILLER_22_199 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_4 FILLER_23_7 ();
 sg13g2_fill_2 FILLER_23_11 ();
 sg13g2_decap_8 FILLER_23_34 ();
 sg13g2_decap_4 FILLER_23_41 ();
 sg13g2_decap_8 FILLER_23_66 ();
 sg13g2_decap_8 FILLER_23_73 ();
 sg13g2_fill_2 FILLER_23_80 ();
 sg13g2_fill_2 FILLER_23_99 ();
 sg13g2_fill_1 FILLER_23_101 ();
 sg13g2_decap_4 FILLER_23_140 ();
 sg13g2_decap_4 FILLER_23_174 ();
 sg13g2_fill_1 FILLER_23_178 ();
 sg13g2_decap_4 FILLER_24_38 ();
 sg13g2_fill_1 FILLER_24_42 ();
 sg13g2_fill_2 FILLER_24_98 ();
 sg13g2_fill_2 FILLER_24_138 ();
 sg13g2_fill_2 FILLER_24_198 ();
 sg13g2_decap_8 FILLER_25_17 ();
 sg13g2_fill_2 FILLER_25_24 ();
 sg13g2_fill_1 FILLER_25_77 ();
 sg13g2_decap_4 FILLER_25_95 ();
 sg13g2_fill_1 FILLER_25_99 ();
 sg13g2_decap_4 FILLER_25_117 ();
 sg13g2_decap_4 FILLER_25_138 ();
 sg13g2_fill_2 FILLER_25_177 ();
 sg13g2_decap_8 FILLER_26_17 ();
 sg13g2_decap_4 FILLER_26_24 ();
 sg13g2_fill_1 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_67 ();
 sg13g2_fill_1 FILLER_26_74 ();
 sg13g2_decap_8 FILLER_26_117 ();
 sg13g2_decap_4 FILLER_26_124 ();
 sg13g2_fill_2 FILLER_26_128 ();
 sg13g2_fill_2 FILLER_26_152 ();
 sg13g2_decap_8 FILLER_26_167 ();
 sg13g2_decap_4 FILLER_26_174 ();
 sg13g2_fill_2 FILLER_26_178 ();
 sg13g2_fill_2 FILLER_26_197 ();
 sg13g2_fill_1 FILLER_26_199 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_11 ();
 sg13g2_fill_2 FILLER_27_34 ();
 sg13g2_fill_1 FILLER_27_36 ();
 sg13g2_decap_8 FILLER_27_54 ();
 sg13g2_decap_8 FILLER_27_61 ();
 sg13g2_fill_1 FILLER_27_68 ();
 sg13g2_decap_8 FILLER_27_103 ();
 sg13g2_decap_4 FILLER_27_110 ();
 sg13g2_fill_1 FILLER_27_114 ();
 sg13g2_decap_4 FILLER_27_157 ();
 sg13g2_fill_1 FILLER_27_199 ();
 sg13g2_fill_2 FILLER_28_34 ();
 sg13g2_decap_8 FILLER_28_57 ();
 sg13g2_fill_2 FILLER_28_64 ();
 sg13g2_fill_1 FILLER_28_66 ();
 sg13g2_decap_8 FILLER_28_88 ();
 sg13g2_fill_2 FILLER_28_95 ();
 sg13g2_fill_2 FILLER_28_135 ();
 sg13g2_decap_8 FILLER_29_17 ();
 sg13g2_fill_2 FILLER_29_24 ();
 sg13g2_decap_4 FILLER_29_70 ();
 sg13g2_fill_1 FILLER_29_74 ();
 sg13g2_fill_1 FILLER_29_109 ();
 sg13g2_decap_8 FILLER_29_115 ();
 sg13g2_fill_2 FILLER_29_139 ();
 sg13g2_decap_4 FILLER_29_177 ();
 sg13g2_fill_1 FILLER_29_181 ();
 sg13g2_fill_1 FILLER_29_199 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_7 ();
 sg13g2_fill_1 FILLER_30_9 ();
 sg13g2_fill_1 FILLER_30_72 ();
 sg13g2_fill_2 FILLER_30_94 ();
 sg13g2_fill_2 FILLER_30_164 ();
 sg13g2_decap_4 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_30 ();
 sg13g2_fill_2 FILLER_31_49 ();
 sg13g2_fill_2 FILLER_31_89 ();
 sg13g2_fill_2 FILLER_31_137 ();
 sg13g2_fill_1 FILLER_31_139 ();
 sg13g2_decap_4 FILLER_32_95 ();
 sg13g2_fill_1 FILLER_32_99 ();
 sg13g2_decap_8 FILLER_32_138 ();
 sg13g2_fill_2 FILLER_32_159 ();
 sg13g2_decap_4 FILLER_32_195 ();
 sg13g2_fill_1 FILLER_32_199 ();
 sg13g2_fill_2 FILLER_33_17 ();
 sg13g2_decap_4 FILLER_33_60 ();
 sg13g2_decap_8 FILLER_33_115 ();
 sg13g2_decap_8 FILLER_33_122 ();
 sg13g2_fill_2 FILLER_33_197 ();
 sg13g2_fill_1 FILLER_33_199 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_4 FILLER_34_7 ();
 sg13g2_fill_1 FILLER_34_54 ();
 sg13g2_decap_4 FILLER_34_70 ();
 sg13g2_fill_2 FILLER_34_74 ();
 sg13g2_decap_4 FILLER_34_120 ();
 sg13g2_fill_2 FILLER_34_124 ();
 sg13g2_fill_1 FILLER_34_148 ();
 sg13g2_decap_8 FILLER_34_187 ();
 sg13g2_decap_4 FILLER_34_194 ();
 sg13g2_fill_2 FILLER_34_198 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_fill_2 FILLER_35_14 ();
 sg13g2_fill_1 FILLER_35_37 ();
 sg13g2_fill_1 FILLER_35_64 ();
 sg13g2_decap_4 FILLER_35_103 ();
 sg13g2_fill_2 FILLER_35_123 ();
 sg13g2_fill_2 FILLER_35_135 ();
 sg13g2_decap_4 FILLER_35_179 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_fill_1 FILLER_36_14 ();
 sg13g2_decap_4 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_73 ();
 sg13g2_decap_4 FILLER_36_80 ();
 sg13g2_fill_1 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_102 ();
 sg13g2_decap_8 FILLER_36_109 ();
 sg13g2_decap_4 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_4 ();
 sg13g2_decap_8 FILLER_37_22 ();
 sg13g2_fill_2 FILLER_37_29 ();
 sg13g2_fill_1 FILLER_37_31 ();
 sg13g2_fill_1 FILLER_37_49 ();
 sg13g2_fill_1 FILLER_37_104 ();
 sg13g2_fill_2 FILLER_37_151 ();
 sg13g2_fill_1 FILLER_37_153 ();
 sg13g2_fill_2 FILLER_37_171 ();
 sg13g2_decap_4 FILLER_37_194 ();
 sg13g2_fill_2 FILLER_37_198 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_4 FILLER_38_7 ();
 sg13g2_fill_2 FILLER_38_49 ();
 sg13g2_fill_1 FILLER_38_51 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_fill_2 FILLER_38_64 ();
 sg13g2_decap_8 FILLER_38_83 ();
 sg13g2_decap_8 FILLER_38_90 ();
 sg13g2_decap_8 FILLER_38_97 ();
 sg13g2_fill_1 FILLER_38_104 ();
 sg13g2_fill_1 FILLER_38_125 ();
 sg13g2_fill_1 FILLER_38_136 ();
 sg13g2_decap_8 FILLER_38_192 ();
 sg13g2_fill_1 FILLER_38_199 ();
 sg13g2_decap_8 FILLER_39_17 ();
 sg13g2_fill_2 FILLER_39_24 ();
 sg13g2_fill_1 FILLER_39_26 ();
 sg13g2_fill_2 FILLER_39_47 ();
 sg13g2_fill_1 FILLER_39_49 ();
 sg13g2_decap_4 FILLER_39_67 ();
 sg13g2_fill_2 FILLER_39_71 ();
 sg13g2_fill_2 FILLER_39_180 ();
 sg13g2_fill_1 FILLER_39_182 ();
 sg13g2_decap_4 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_107 ();
 sg13g2_decap_4 FILLER_40_114 ();
 sg13g2_fill_1 FILLER_40_118 ();
 sg13g2_fill_1 FILLER_40_139 ();
 sg13g2_fill_1 FILLER_40_199 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_fill_2 FILLER_41_42 ();
 sg13g2_fill_2 FILLER_41_64 ();
 sg13g2_fill_1 FILLER_41_66 ();
 sg13g2_decap_4 FILLER_41_95 ();
 sg13g2_decap_8 FILLER_41_137 ();
 sg13g2_decap_8 FILLER_41_161 ();
 sg13g2_fill_2 FILLER_41_168 ();
 sg13g2_fill_1 FILLER_41_170 ();
 sg13g2_decap_8 FILLER_41_192 ();
 sg13g2_fill_1 FILLER_41_199 ();
 sg13g2_decap_8 FILLER_42_17 ();
 sg13g2_decap_8 FILLER_42_24 ();
 sg13g2_fill_1 FILLER_42_67 ();
 sg13g2_decap_8 FILLER_42_119 ();
 sg13g2_decap_8 FILLER_42_126 ();
 sg13g2_decap_8 FILLER_42_133 ();
 sg13g2_decap_8 FILLER_42_161 ();
 sg13g2_decap_4 FILLER_42_168 ();
 sg13g2_fill_2 FILLER_42_172 ();
 sg13g2_decap_8 FILLER_42_191 ();
 sg13g2_fill_2 FILLER_42_198 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_fill_2 FILLER_43_7 ();
 sg13g2_fill_1 FILLER_43_9 ();
 sg13g2_fill_1 FILLER_43_31 ();
 sg13g2_fill_1 FILLER_43_72 ();
 sg13g2_fill_1 FILLER_43_121 ();
 sg13g2_fill_2 FILLER_43_177 ();
 sg13g2_decap_4 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_4 ();
 sg13g2_decap_4 FILLER_44_23 ();
 sg13g2_fill_2 FILLER_44_27 ();
 sg13g2_fill_1 FILLER_44_46 ();
 sg13g2_fill_1 FILLER_44_65 ();
 sg13g2_decap_8 FILLER_44_104 ();
 sg13g2_decap_4 FILLER_44_111 ();
 sg13g2_fill_1 FILLER_44_115 ();
 sg13g2_decap_4 FILLER_44_167 ();
 sg13g2_fill_1 FILLER_44_171 ();
 sg13g2_decap_8 FILLER_44_193 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_65 ();
 sg13g2_decap_8 FILLER_45_72 ();
 sg13g2_decap_8 FILLER_45_79 ();
 sg13g2_fill_2 FILLER_45_86 ();
 sg13g2_decap_8 FILLER_45_105 ();
 sg13g2_fill_2 FILLER_45_112 ();
 sg13g2_decap_8 FILLER_45_135 ();
 sg13g2_decap_8 FILLER_45_142 ();
 sg13g2_fill_1 FILLER_45_149 ();
 sg13g2_decap_8 FILLER_45_184 ();
 sg13g2_decap_8 FILLER_45_191 ();
 sg13g2_fill_2 FILLER_45_198 ();
 sg13g2_decap_8 FILLER_46_17 ();
 sg13g2_decap_4 FILLER_46_24 ();
 sg13g2_fill_1 FILLER_46_28 ();
 sg13g2_fill_1 FILLER_46_46 ();
 sg13g2_decap_4 FILLER_46_123 ();
 sg13g2_fill_2 FILLER_46_161 ();
 sg13g2_fill_2 FILLER_46_197 ();
 sg13g2_fill_1 FILLER_46_199 ();
 sg13g2_fill_2 FILLER_47_70 ();
 sg13g2_fill_1 FILLER_47_72 ();
 sg13g2_decap_4 FILLER_47_94 ();
 sg13g2_fill_2 FILLER_47_98 ();
 sg13g2_fill_2 FILLER_47_117 ();
 sg13g2_decap_8 FILLER_47_140 ();
 sg13g2_fill_2 FILLER_47_147 ();
 sg13g2_decap_8 FILLER_47_170 ();
 sg13g2_fill_2 FILLER_47_198 ();
 sg13g2_decap_4 FILLER_48_38 ();
 sg13g2_fill_2 FILLER_48_42 ();
 sg13g2_decap_4 FILLER_48_91 ();
 sg13g2_fill_2 FILLER_48_95 ();
 sg13g2_fill_1 FILLER_48_135 ();
 sg13g2_decap_8 FILLER_48_170 ();
 sg13g2_fill_2 FILLER_48_177 ();
 sg13g2_fill_1 FILLER_48_179 ();
 sg13g2_fill_2 FILLER_48_197 ();
 sg13g2_fill_1 FILLER_48_199 ();
 sg13g2_fill_1 FILLER_49_17 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_62 ();
 sg13g2_decap_8 FILLER_49_69 ();
 sg13g2_decap_8 FILLER_49_76 ();
 sg13g2_fill_1 FILLER_49_83 ();
 sg13g2_fill_2 FILLER_49_101 ();
 sg13g2_decap_8 FILLER_49_108 ();
 sg13g2_decap_4 FILLER_49_115 ();
 sg13g2_decap_8 FILLER_49_136 ();
 sg13g2_decap_4 FILLER_49_143 ();
 sg13g2_fill_1 FILLER_49_147 ();
 sg13g2_fill_2 FILLER_49_186 ();
 sg13g2_fill_1 FILLER_49_188 ();
 sg13g2_fill_2 FILLER_49_197 ();
 sg13g2_fill_1 FILLER_49_199 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_fill_1 FILLER_50_14 ();
 sg13g2_fill_2 FILLER_50_39 ();
 sg13g2_decap_4 FILLER_50_83 ();
 sg13g2_decap_8 FILLER_50_141 ();
 sg13g2_decap_8 FILLER_50_148 ();
 sg13g2_fill_2 FILLER_50_155 ();
 sg13g2_decap_4 FILLER_50_174 ();
 sg13g2_fill_1 FILLER_50_199 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_4 FILLER_51_7 ();
 sg13g2_fill_2 FILLER_51_11 ();
 sg13g2_fill_1 FILLER_51_83 ();
 sg13g2_fill_1 FILLER_51_94 ();
 sg13g2_decap_4 FILLER_51_100 ();
 sg13g2_fill_1 FILLER_51_104 ();
 sg13g2_fill_1 FILLER_51_150 ();
 sg13g2_decap_8 FILLER_51_168 ();
 sg13g2_decap_4 FILLER_51_196 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_fill_1 FILLER_52_7 ();
 sg13g2_fill_2 FILLER_52_44 ();
 sg13g2_fill_1 FILLER_52_46 ();
 sg13g2_fill_2 FILLER_52_67 ();
 sg13g2_fill_1 FILLER_52_79 ();
 sg13g2_decap_4 FILLER_52_102 ();
 sg13g2_fill_1 FILLER_52_106 ();
 sg13g2_fill_2 FILLER_52_124 ();
 sg13g2_fill_2 FILLER_52_131 ();
 sg13g2_decap_4 FILLER_52_171 ();
 sg13g2_fill_2 FILLER_52_175 ();
 sg13g2_fill_1 FILLER_52_199 ();
 sg13g2_fill_2 FILLER_53_66 ();
 sg13g2_decap_8 FILLER_53_106 ();
 sg13g2_decap_8 FILLER_53_113 ();
 sg13g2_decap_4 FILLER_53_120 ();
 sg13g2_fill_1 FILLER_53_124 ();
 sg13g2_fill_1 FILLER_53_134 ();
 sg13g2_fill_1 FILLER_53_152 ();
 sg13g2_fill_2 FILLER_54_40 ();
 sg13g2_fill_1 FILLER_54_82 ();
 sg13g2_fill_2 FILLER_54_147 ();
 sg13g2_fill_1 FILLER_54_149 ();
 sg13g2_fill_1 FILLER_54_199 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_fill_2 FILLER_55_14 ();
 sg13g2_fill_2 FILLER_55_40 ();
 sg13g2_fill_1 FILLER_55_59 ();
 sg13g2_decap_4 FILLER_55_103 ();
 sg13g2_fill_2 FILLER_55_141 ();
 sg13g2_decap_8 FILLER_55_147 ();
 sg13g2_fill_1 FILLER_55_154 ();
 sg13g2_fill_1 FILLER_55_159 ();
 sg13g2_fill_2 FILLER_55_164 ();
 sg13g2_fill_2 FILLER_55_170 ();
 sg13g2_fill_2 FILLER_55_180 ();
 sg13g2_fill_1 FILLER_55_182 ();
 sg13g2_fill_2 FILLER_55_187 ();
 sg13g2_fill_2 FILLER_55_197 ();
 sg13g2_fill_1 FILLER_55_199 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_fill_2 FILLER_56_7 ();
 sg13g2_fill_1 FILLER_56_9 ();
 sg13g2_decap_8 FILLER_56_32 ();
 sg13g2_decap_8 FILLER_56_39 ();
 sg13g2_decap_8 FILLER_56_46 ();
 sg13g2_fill_1 FILLER_56_53 ();
 sg13g2_decap_8 FILLER_56_76 ();
 sg13g2_fill_1 FILLER_56_83 ();
 sg13g2_decap_8 FILLER_56_87 ();
 sg13g2_decap_8 FILLER_56_94 ();
 sg13g2_decap_8 FILLER_56_101 ();
 sg13g2_fill_1 FILLER_56_108 ();
 sg13g2_decap_8 FILLER_56_113 ();
 sg13g2_decap_4 FILLER_56_120 ();
 sg13g2_fill_2 FILLER_56_128 ();
 sg13g2_fill_1 FILLER_56_130 ();
 sg13g2_decap_8 FILLER_56_148 ();
 sg13g2_decap_8 FILLER_56_155 ();
 sg13g2_decap_8 FILLER_56_162 ();
 sg13g2_fill_1 FILLER_56_169 ();
 sg13g2_fill_2 FILLER_56_178 ();
 sg13g2_fill_1 FILLER_56_180 ();
 sg13g2_fill_2 FILLER_56_197 ();
 sg13g2_fill_1 FILLER_56_199 ();
 sg13g2_decap_4 FILLER_57_0 ();
 sg13g2_fill_1 FILLER_57_25 ();
 sg13g2_decap_8 FILLER_57_47 ();
 sg13g2_fill_1 FILLER_57_71 ();
 sg13g2_decap_4 FILLER_57_89 ();
 sg13g2_fill_1 FILLER_57_93 ();
 sg13g2_decap_8 FILLER_57_132 ();
 sg13g2_decap_4 FILLER_57_139 ();
 sg13g2_decap_4 FILLER_57_168 ();
 sg13g2_fill_1 FILLER_57_180 ();
 sg13g2_fill_2 FILLER_57_198 ();
 sg13g2_decap_4 FILLER_58_46 ();
 sg13g2_fill_1 FILLER_58_50 ();
 sg13g2_fill_2 FILLER_58_89 ();
 sg13g2_fill_1 FILLER_58_91 ();
 sg13g2_fill_1 FILLER_58_113 ();
 sg13g2_decap_8 FILLER_58_131 ();
 sg13g2_decap_8 FILLER_58_138 ();
 sg13g2_fill_2 FILLER_58_145 ();
 sg13g2_decap_8 FILLER_58_168 ();
 sg13g2_fill_1 FILLER_58_175 ();
 sg13g2_fill_2 FILLER_58_197 ();
 sg13g2_fill_1 FILLER_58_199 ();
 sg13g2_fill_2 FILLER_59_0 ();
 sg13g2_fill_1 FILLER_59_2 ();
 sg13g2_decap_8 FILLER_59_19 ();
 sg13g2_decap_8 FILLER_59_26 ();
 sg13g2_decap_8 FILLER_59_50 ();
 sg13g2_decap_8 FILLER_59_57 ();
 sg13g2_decap_8 FILLER_59_64 ();
 sg13g2_decap_8 FILLER_59_71 ();
 sg13g2_decap_8 FILLER_59_112 ();
 sg13g2_decap_8 FILLER_59_119 ();
 sg13g2_decap_4 FILLER_59_126 ();
 sg13g2_decap_4 FILLER_59_147 ();
 sg13g2_fill_1 FILLER_59_151 ();
 sg13g2_fill_2 FILLER_59_186 ();
 sg13g2_fill_1 FILLER_59_188 ();
 sg13g2_fill_2 FILLER_59_197 ();
 sg13g2_fill_1 FILLER_59_199 ();
 sg13g2_decap_4 FILLER_60_25 ();
 sg13g2_fill_1 FILLER_60_29 ();
 sg13g2_decap_8 FILLER_60_47 ();
 sg13g2_decap_8 FILLER_60_92 ();
 sg13g2_fill_2 FILLER_60_99 ();
 sg13g2_decap_8 FILLER_60_139 ();
 sg13g2_decap_4 FILLER_60_146 ();
 sg13g2_fill_1 FILLER_60_150 ();
 sg13g2_decap_8 FILLER_60_168 ();
 sg13g2_fill_2 FILLER_60_175 ();
 sg13g2_fill_1 FILLER_60_177 ();
 sg13g2_fill_1 FILLER_60_199 ();
 sg13g2_fill_2 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_2 ();
 sg13g2_fill_2 FILLER_61_24 ();
 sg13g2_decap_4 FILLER_61_47 ();
 sg13g2_decap_4 FILLER_61_72 ();
 sg13g2_fill_1 FILLER_61_93 ();
 sg13g2_decap_8 FILLER_61_115 ();
 sg13g2_decap_8 FILLER_61_139 ();
 sg13g2_fill_1 FILLER_61_146 ();
 sg13g2_decap_8 FILLER_61_168 ();
 sg13g2_fill_2 FILLER_61_175 ();
 sg13g2_fill_2 FILLER_61_198 ();
 sg13g2_fill_2 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_2 ();
 sg13g2_fill_1 FILLER_62_36 ();
 sg13g2_decap_4 FILLER_62_71 ();
 sg13g2_fill_2 FILLER_62_75 ();
 sg13g2_decap_4 FILLER_62_98 ();
 sg13g2_decap_8 FILLER_62_191 ();
 sg13g2_fill_2 FILLER_62_198 ();
 sg13g2_fill_2 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_2 ();
 sg13g2_fill_2 FILLER_63_11 ();
 sg13g2_fill_1 FILLER_63_13 ();
 sg13g2_fill_1 FILLER_63_69 ();
 sg13g2_fill_1 FILLER_63_97 ();
 sg13g2_decap_8 FILLER_63_115 ();
 sg13g2_fill_2 FILLER_63_122 ();
 sg13g2_decap_8 FILLER_63_141 ();
 sg13g2_decap_4 FILLER_63_169 ();
 sg13g2_fill_1 FILLER_63_173 ();
 sg13g2_decap_4 FILLER_63_195 ();
 sg13g2_fill_1 FILLER_63_199 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_fill_1 FILLER_64_14 ();
 sg13g2_decap_4 FILLER_64_53 ();
 sg13g2_decap_8 FILLER_64_159 ();
 sg13g2_decap_8 FILLER_64_166 ();
 sg13g2_fill_1 FILLER_64_173 ();
 sg13g2_decap_4 FILLER_64_195 ();
 sg13g2_fill_1 FILLER_64_199 ();
 sg13g2_fill_2 FILLER_65_0 ();
 sg13g2_fill_1 FILLER_65_2 ();
 sg13g2_fill_2 FILLER_65_66 ();
 sg13g2_fill_2 FILLER_65_98 ();
 sg13g2_fill_2 FILLER_65_197 ();
 sg13g2_fill_1 FILLER_65_199 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_4 FILLER_66_49 ();
 sg13g2_fill_2 FILLER_66_53 ();
 sg13g2_decap_4 FILLER_66_72 ();
 sg13g2_fill_2 FILLER_66_93 ();
 sg13g2_decap_8 FILLER_66_112 ();
 sg13g2_fill_1 FILLER_66_119 ();
 sg13g2_fill_1 FILLER_66_137 ();
 sg13g2_decap_4 FILLER_66_153 ();
 sg13g2_decap_4 FILLER_66_174 ();
 sg13g2_fill_1 FILLER_66_199 ();
 sg13g2_fill_2 FILLER_67_0 ();
 sg13g2_fill_1 FILLER_67_2 ();
 sg13g2_decap_4 FILLER_67_79 ();
 sg13g2_fill_1 FILLER_67_83 ();
 sg13g2_fill_1 FILLER_67_89 ();
 sg13g2_decap_4 FILLER_67_111 ();
 sg13g2_fill_2 FILLER_67_132 ();
 sg13g2_fill_2 FILLER_67_164 ();
 sg13g2_fill_1 FILLER_67_166 ();
 sg13g2_fill_1 FILLER_67_188 ();
 sg13g2_fill_2 FILLER_67_197 ();
 sg13g2_fill_1 FILLER_67_199 ();
 sg13g2_fill_2 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_2 ();
 sg13g2_decap_8 FILLER_68_41 ();
 sg13g2_decap_8 FILLER_68_48 ();
 sg13g2_fill_1 FILLER_68_55 ();
 sg13g2_decap_8 FILLER_68_94 ();
 sg13g2_decap_8 FILLER_68_101 ();
 sg13g2_decap_8 FILLER_68_108 ();
 sg13g2_decap_8 FILLER_68_115 ();
 sg13g2_fill_2 FILLER_68_139 ();
 sg13g2_fill_2 FILLER_68_197 ();
 sg13g2_fill_1 FILLER_68_199 ();
 sg13g2_fill_1 FILLER_69_0 ();
 sg13g2_fill_2 FILLER_69_26 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_fill_2 FILLER_69_70 ();
 sg13g2_fill_1 FILLER_69_72 ();
 sg13g2_fill_1 FILLER_69_128 ();
 sg13g2_decap_8 FILLER_69_170 ();
 sg13g2_fill_1 FILLER_69_177 ();
 sg13g2_fill_1 FILLER_69_199 ();
 sg13g2_fill_2 FILLER_70_0 ();
 sg13g2_fill_1 FILLER_70_2 ();
 sg13g2_fill_2 FILLER_70_11 ();
 sg13g2_fill_1 FILLER_70_13 ();
 sg13g2_fill_2 FILLER_70_31 ();
 sg13g2_fill_2 FILLER_70_50 ();
 sg13g2_fill_1 FILLER_70_52 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_decap_4 FILLER_70_98 ();
 sg13g2_fill_2 FILLER_70_102 ();
 sg13g2_decap_8 FILLER_70_159 ();
 sg13g2_decap_4 FILLER_70_166 ();
 sg13g2_fill_1 FILLER_70_170 ();
 sg13g2_fill_2 FILLER_71_0 ();
 sg13g2_fill_1 FILLER_71_2 ();
 sg13g2_fill_2 FILLER_71_11 ();
 sg13g2_decap_8 FILLER_71_34 ();
 sg13g2_decap_8 FILLER_71_41 ();
 sg13g2_fill_1 FILLER_71_48 ();
 sg13g2_decap_4 FILLER_71_70 ();
 sg13g2_fill_1 FILLER_71_74 ();
 sg13g2_fill_1 FILLER_71_109 ();
 sg13g2_decap_4 FILLER_71_131 ();
 sg13g2_fill_1 FILLER_71_135 ();
 sg13g2_decap_4 FILLER_71_167 ();
 sg13g2_fill_1 FILLER_71_171 ();
 sg13g2_fill_2 FILLER_71_197 ();
 sg13g2_fill_1 FILLER_71_199 ();
 sg13g2_decap_8 FILLER_72_25 ();
 sg13g2_decap_4 FILLER_72_32 ();
 sg13g2_fill_2 FILLER_72_53 ();
 sg13g2_decap_8 FILLER_72_93 ();
 sg13g2_decap_4 FILLER_72_100 ();
 sg13g2_fill_2 FILLER_72_104 ();
 sg13g2_decap_8 FILLER_72_131 ();
 sg13g2_decap_8 FILLER_72_138 ();
 sg13g2_decap_8 FILLER_72_145 ();
 sg13g2_fill_2 FILLER_72_186 ();
 sg13g2_fill_1 FILLER_72_188 ();
 sg13g2_fill_2 FILLER_72_197 ();
 sg13g2_fill_1 FILLER_72_199 ();
 sg13g2_fill_2 FILLER_73_21 ();
 sg13g2_fill_1 FILLER_73_23 ();
 sg13g2_decap_4 FILLER_73_45 ();
 sg13g2_fill_1 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_67 ();
 sg13g2_fill_2 FILLER_73_74 ();
 sg13g2_fill_2 FILLER_73_114 ();
 sg13g2_decap_8 FILLER_73_133 ();
 sg13g2_decap_4 FILLER_73_140 ();
 sg13g2_fill_1 FILLER_73_144 ();
 sg13g2_fill_1 FILLER_73_175 ();
 sg13g2_fill_2 FILLER_73_197 ();
 sg13g2_fill_1 FILLER_73_199 ();
 sg13g2_fill_2 FILLER_74_0 ();
 sg13g2_fill_1 FILLER_74_2 ();
 sg13g2_fill_1 FILLER_74_11 ();
 sg13g2_fill_1 FILLER_74_50 ();
 sg13g2_fill_2 FILLER_74_148 ();
 sg13g2_fill_2 FILLER_74_197 ();
 sg13g2_fill_1 FILLER_74_199 ();
 sg13g2_fill_1 FILLER_75_0 ();
 sg13g2_fill_1 FILLER_75_22 ();
 sg13g2_decap_8 FILLER_75_44 ();
 sg13g2_fill_1 FILLER_75_51 ();
 sg13g2_fill_2 FILLER_75_90 ();
 sg13g2_fill_1 FILLER_75_92 ();
 sg13g2_fill_1 FILLER_75_110 ();
 sg13g2_decap_4 FILLER_75_128 ();
 sg13g2_fill_2 FILLER_75_132 ();
 sg13g2_fill_2 FILLER_75_198 ();
 sg13g2_fill_2 FILLER_76_0 ();
 sg13g2_fill_1 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_109 ();
 sg13g2_decap_4 FILLER_76_116 ();
 sg13g2_decap_4 FILLER_76_124 ();
 sg13g2_fill_2 FILLER_76_128 ();
 sg13g2_fill_2 FILLER_76_164 ();
 sg13g2_fill_1 FILLER_76_166 ();
 sg13g2_fill_1 FILLER_77_17 ();
 sg13g2_decap_8 FILLER_77_43 ();
 sg13g2_fill_2 FILLER_77_50 ();
 sg13g2_fill_1 FILLER_77_73 ();
 sg13g2_decap_4 FILLER_77_112 ();
 sg13g2_fill_2 FILLER_77_116 ();
 sg13g2_decap_4 FILLER_77_160 ();
 sg13g2_fill_2 FILLER_77_197 ();
 sg13g2_fill_1 FILLER_77_199 ();
 sg13g2_fill_2 FILLER_78_0 ();
 sg13g2_fill_1 FILLER_78_2 ();
 sg13g2_decap_8 FILLER_78_41 ();
 sg13g2_decap_8 FILLER_78_48 ();
 sg13g2_decap_8 FILLER_78_76 ();
 sg13g2_decap_8 FILLER_78_83 ();
 sg13g2_decap_4 FILLER_78_90 ();
 sg13g2_fill_2 FILLER_78_94 ();
 sg13g2_fill_2 FILLER_78_117 ();
 sg13g2_fill_2 FILLER_78_157 ();
 sg13g2_fill_1 FILLER_78_159 ();
 sg13g2_fill_2 FILLER_78_197 ();
 sg13g2_fill_1 FILLER_78_199 ();
 sg13g2_fill_2 FILLER_79_0 ();
 sg13g2_fill_1 FILLER_79_2 ();
 sg13g2_fill_1 FILLER_79_58 ();
 sg13g2_fill_2 FILLER_79_76 ();
 sg13g2_fill_1 FILLER_79_78 ();
 sg13g2_decap_4 FILLER_79_117 ();
 sg13g2_decap_4 FILLER_79_151 ();
 sg13g2_fill_2 FILLER_79_155 ();
 sg13g2_fill_2 FILLER_79_174 ();
 sg13g2_fill_2 FILLER_79_193 ();
 sg13g2_fill_1 FILLER_79_195 ();
 sg13g2_fill_1 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_39 ();
 sg13g2_decap_8 FILLER_80_46 ();
 sg13g2_fill_2 FILLER_80_53 ();
 sg13g2_decap_8 FILLER_80_72 ();
 sg13g2_fill_1 FILLER_80_79 ();
 sg13g2_decap_4 FILLER_80_97 ();
 sg13g2_fill_1 FILLER_80_101 ();
 sg13g2_decap_4 FILLER_80_119 ();
 sg13g2_fill_2 FILLER_80_123 ();
 sg13g2_decap_8 FILLER_80_146 ();
 sg13g2_fill_2 FILLER_80_174 ();
 sg13g2_fill_2 FILLER_80_197 ();
 sg13g2_fill_1 FILLER_80_199 ();
 sg13g2_fill_1 FILLER_81_0 ();
 sg13g2_fill_2 FILLER_81_18 ();
 sg13g2_fill_1 FILLER_81_20 ();
 sg13g2_decap_8 FILLER_81_42 ();
 sg13g2_decap_4 FILLER_81_49 ();
 sg13g2_fill_2 FILLER_81_53 ();
 sg13g2_decap_8 FILLER_81_93 ();
 sg13g2_fill_2 FILLER_81_100 ();
 sg13g2_fill_1 FILLER_81_102 ();
 sg13g2_fill_2 FILLER_81_120 ();
 sg13g2_fill_1 FILLER_81_122 ();
 sg13g2_decap_8 FILLER_81_127 ();
 sg13g2_fill_2 FILLER_81_134 ();
 sg13g2_decap_4 FILLER_81_157 ();
 sg13g2_decap_8 FILLER_81_165 ();
 sg13g2_fill_1 FILLER_81_172 ();
 sg13g2_fill_2 FILLER_81_198 ();
 sg13g2_fill_2 FILLER_82_0 ();
 sg13g2_fill_1 FILLER_82_2 ();
 sg13g2_fill_1 FILLER_82_70 ();
 sg13g2_decap_8 FILLER_82_130 ();
 sg13g2_decap_4 FILLER_82_137 ();
 sg13g2_fill_1 FILLER_82_141 ();
 sg13g2_decap_8 FILLER_82_159 ();
 sg13g2_decap_8 FILLER_82_166 ();
 sg13g2_fill_2 FILLER_82_198 ();
 sg13g2_fill_2 FILLER_83_0 ();
 sg13g2_decap_8 FILLER_83_19 ();
 sg13g2_fill_1 FILLER_83_26 ();
 sg13g2_decap_4 FILLER_83_44 ();
 sg13g2_fill_2 FILLER_83_48 ();
 sg13g2_decap_4 FILLER_83_67 ();
 sg13g2_fill_2 FILLER_83_71 ();
 sg13g2_fill_2 FILLER_83_112 ();
 sg13g2_fill_1 FILLER_83_114 ();
 sg13g2_decap_4 FILLER_83_153 ();
 sg13g2_fill_2 FILLER_83_191 ();
 sg13g2_fill_2 FILLER_83_197 ();
 sg13g2_fill_1 FILLER_83_199 ();
 sg13g2_decap_8 FILLER_84_0 ();
 sg13g2_fill_1 FILLER_84_7 ();
 sg13g2_fill_2 FILLER_84_67 ();
 sg13g2_fill_1 FILLER_84_97 ();
 sg13g2_decap_4 FILLER_84_115 ();
 sg13g2_fill_2 FILLER_84_136 ();
 sg13g2_decap_8 FILLER_84_155 ();
 sg13g2_decap_8 FILLER_84_162 ();
 sg13g2_decap_4 FILLER_84_190 ();
 sg13g2_fill_2 FILLER_84_198 ();
 sg13g2_decap_8 FILLER_85_0 ();
 sg13g2_decap_8 FILLER_85_7 ();
 sg13g2_fill_2 FILLER_85_14 ();
 sg13g2_decap_8 FILLER_85_37 ();
 sg13g2_fill_2 FILLER_85_44 ();
 sg13g2_decap_8 FILLER_85_123 ();
 sg13g2_decap_4 FILLER_85_130 ();
 sg13g2_fill_1 FILLER_85_134 ();
 sg13g2_fill_2 FILLER_85_156 ();
 sg13g2_fill_1 FILLER_85_158 ();
 sg13g2_decap_4 FILLER_85_163 ();
 sg13g2_fill_1 FILLER_85_167 ();
 sg13g2_decap_8 FILLER_85_189 ();
 sg13g2_decap_4 FILLER_85_196 ();
 sg13g2_fill_2 FILLER_86_0 ();
 sg13g2_fill_2 FILLER_86_19 ();
 sg13g2_fill_1 FILLER_86_21 ();
 sg13g2_fill_1 FILLER_86_39 ();
 sg13g2_decap_8 FILLER_86_70 ();
 sg13g2_fill_1 FILLER_86_77 ();
 sg13g2_decap_8 FILLER_86_86 ();
 sg13g2_decap_8 FILLER_86_93 ();
 sg13g2_decap_4 FILLER_86_100 ();
 sg13g2_decap_4 FILLER_86_155 ();
 sg13g2_fill_2 FILLER_86_159 ();
 sg13g2_decap_4 FILLER_86_195 ();
 sg13g2_fill_1 FILLER_86_199 ();
 sg13g2_decap_8 FILLER_87_0 ();
 sg13g2_decap_4 FILLER_87_7 ();
 sg13g2_fill_1 FILLER_87_11 ();
 sg13g2_decap_8 FILLER_87_33 ();
 sg13g2_fill_1 FILLER_87_40 ();
 sg13g2_fill_1 FILLER_87_58 ();
 sg13g2_decap_8 FILLER_87_127 ();
 sg13g2_fill_2 FILLER_87_134 ();
 sg13g2_fill_2 FILLER_87_157 ();
 sg13g2_fill_1 FILLER_87_159 ();
 sg13g2_decap_4 FILLER_87_194 ();
 sg13g2_fill_2 FILLER_87_198 ();
 sg13g2_decap_4 FILLER_88_0 ();
 sg13g2_fill_2 FILLER_88_4 ();
 sg13g2_decap_8 FILLER_88_23 ();
 sg13g2_decap_4 FILLER_88_30 ();
 sg13g2_fill_1 FILLER_88_34 ();
 sg13g2_decap_8 FILLER_88_56 ();
 sg13g2_fill_1 FILLER_88_63 ();
 sg13g2_decap_4 FILLER_88_100 ();
 sg13g2_fill_2 FILLER_88_104 ();
 sg13g2_decap_8 FILLER_88_144 ();
 sg13g2_fill_2 FILLER_88_151 ();
 sg13g2_fill_2 FILLER_88_170 ();
 sg13g2_fill_1 FILLER_88_172 ();
 sg13g2_decap_4 FILLER_88_194 ();
 sg13g2_fill_2 FILLER_88_198 ();
 sg13g2_decap_4 FILLER_89_0 ();
 sg13g2_decap_8 FILLER_89_25 ();
 sg13g2_decap_4 FILLER_89_32 ();
 sg13g2_fill_1 FILLER_89_36 ();
 sg13g2_fill_1 FILLER_89_54 ();
 sg13g2_decap_4 FILLER_89_110 ();
 sg13g2_fill_2 FILLER_89_114 ();
 sg13g2_fill_2 FILLER_89_150 ();
 sg13g2_fill_1 FILLER_89_152 ();
 sg13g2_decap_8 FILLER_89_170 ();
 sg13g2_fill_2 FILLER_89_177 ();
 sg13g2_decap_4 FILLER_89_196 ();
 sg13g2_fill_1 FILLER_90_51 ();
 sg13g2_decap_4 FILLER_90_69 ();
 sg13g2_fill_2 FILLER_90_73 ();
 sg13g2_fill_2 FILLER_90_84 ();
 sg13g2_fill_1 FILLER_90_86 ();
 sg13g2_decap_4 FILLER_90_121 ();
 sg13g2_decap_8 FILLER_90_163 ();
 sg13g2_decap_8 FILLER_90_170 ();
 sg13g2_fill_2 FILLER_90_198 ();
 sg13g2_decap_4 FILLER_91_17 ();
 sg13g2_fill_1 FILLER_91_21 ();
 sg13g2_decap_8 FILLER_91_43 ();
 sg13g2_fill_1 FILLER_91_50 ();
 sg13g2_decap_4 FILLER_91_72 ();
 sg13g2_fill_2 FILLER_91_76 ();
 sg13g2_decap_8 FILLER_91_95 ();
 sg13g2_fill_2 FILLER_91_123 ();
 sg13g2_decap_8 FILLER_91_163 ();
 sg13g2_decap_4 FILLER_91_170 ();
 sg13g2_fill_2 FILLER_91_174 ();
 sg13g2_fill_2 FILLER_91_197 ();
 sg13g2_fill_1 FILLER_91_199 ();
 sg13g2_fill_2 FILLER_92_17 ();
 sg13g2_fill_1 FILLER_92_19 ();
 sg13g2_fill_2 FILLER_92_54 ();
 sg13g2_fill_1 FILLER_92_94 ();
 sg13g2_decap_4 FILLER_92_106 ();
 sg13g2_fill_2 FILLER_92_110 ();
 sg13g2_decap_8 FILLER_92_148 ();
 sg13g2_fill_1 FILLER_92_155 ();
 sg13g2_decap_8 FILLER_92_173 ();
 sg13g2_fill_2 FILLER_92_197 ();
 sg13g2_fill_1 FILLER_92_199 ();
 sg13g2_fill_2 FILLER_93_0 ();
 sg13g2_decap_8 FILLER_93_23 ();
 sg13g2_fill_1 FILLER_93_30 ();
 sg13g2_fill_2 FILLER_93_112 ();
 sg13g2_decap_4 FILLER_93_173 ();
 sg13g2_fill_1 FILLER_93_177 ();
 sg13g2_decap_4 FILLER_93_195 ();
 sg13g2_fill_1 FILLER_93_199 ();
 sg13g2_decap_4 FILLER_94_0 ();
 sg13g2_fill_1 FILLER_94_4 ();
 sg13g2_decap_8 FILLER_94_22 ();
 sg13g2_fill_2 FILLER_94_29 ();
 sg13g2_fill_1 FILLER_94_31 ();
 sg13g2_fill_2 FILLER_94_66 ();
 sg13g2_fill_1 FILLER_94_107 ();
 sg13g2_decap_8 FILLER_94_171 ();
 sg13g2_fill_1 FILLER_94_178 ();
 sg13g2_decap_8 FILLER_95_17 ();
 sg13g2_fill_1 FILLER_95_24 ();
 sg13g2_decap_4 FILLER_95_46 ();
 sg13g2_fill_2 FILLER_95_72 ();
 sg13g2_decap_8 FILLER_95_99 ();
 sg13g2_fill_2 FILLER_95_106 ();
 sg13g2_fill_1 FILLER_95_108 ();
 sg13g2_fill_2 FILLER_95_131 ();
 sg13g2_decap_8 FILLER_95_171 ();
 sg13g2_fill_1 FILLER_95_178 ();
 sg13g2_decap_4 FILLER_95_196 ();
 sg13g2_fill_2 FILLER_96_0 ();
 sg13g2_fill_1 FILLER_96_2 ();
 sg13g2_fill_1 FILLER_96_74 ();
 sg13g2_fill_2 FILLER_96_134 ();
 sg13g2_fill_1 FILLER_96_153 ();
 sg13g2_decap_4 FILLER_96_157 ();
 sg13g2_fill_2 FILLER_96_161 ();
 sg13g2_fill_2 FILLER_96_197 ();
 sg13g2_fill_1 FILLER_96_199 ();
 sg13g2_decap_8 FILLER_97_0 ();
 sg13g2_decap_4 FILLER_97_24 ();
 sg13g2_fill_1 FILLER_97_28 ();
 sg13g2_fill_2 FILLER_97_46 ();
 sg13g2_fill_1 FILLER_97_48 ();
 sg13g2_decap_8 FILLER_97_70 ();
 sg13g2_decap_8 FILLER_97_77 ();
 sg13g2_decap_4 FILLER_97_84 ();
 sg13g2_fill_2 FILLER_97_114 ();
 sg13g2_fill_1 FILLER_97_116 ();
 sg13g2_fill_2 FILLER_97_147 ();
 sg13g2_fill_2 FILLER_98_0 ();
 sg13g2_decap_4 FILLER_98_6 ();
 sg13g2_fill_1 FILLER_98_127 ();
 sg13g2_fill_1 FILLER_98_145 ();
 sg13g2_fill_1 FILLER_98_159 ();
 sg13g2_decap_8 FILLER_98_181 ();
 sg13g2_decap_8 FILLER_98_188 ();
 sg13g2_fill_1 FILLER_98_195 ();
 sg13g2_fill_1 FILLER_98_199 ();
 sg13g2_fill_1 FILLER_99_38 ();
 sg13g2_decap_8 FILLER_99_74 ();
 sg13g2_decap_8 FILLER_99_81 ();
 sg13g2_decap_4 FILLER_99_88 ();
 sg13g2_fill_1 FILLER_99_92 ();
 sg13g2_decap_4 FILLER_99_110 ();
 sg13g2_fill_2 FILLER_99_131 ();
 sg13g2_fill_1 FILLER_99_155 ();
 sg13g2_fill_2 FILLER_99_190 ();
 sg13g2_fill_1 FILLER_99_195 ();
 sg13g2_fill_1 FILLER_100_0 ();
 sg13g2_fill_1 FILLER_100_39 ();
 sg13g2_decap_8 FILLER_100_95 ();
 sg13g2_fill_1 FILLER_100_102 ();
 sg13g2_decap_8 FILLER_100_120 ();
 sg13g2_decap_8 FILLER_100_127 ();
 sg13g2_decap_4 FILLER_100_134 ();
 sg13g2_fill_1 FILLER_100_138 ();
 sg13g2_fill_1 FILLER_100_173 ();
 sg13g2_fill_1 FILLER_100_199 ();
 sg13g2_fill_1 FILLER_101_17 ();
 sg13g2_decap_8 FILLER_101_43 ();
 sg13g2_fill_2 FILLER_101_79 ();
 sg13g2_decap_8 FILLER_101_119 ();
 sg13g2_fill_1 FILLER_101_126 ();
 sg13g2_fill_1 FILLER_101_148 ();
 sg13g2_fill_2 FILLER_101_198 ();
 sg13g2_fill_2 FILLER_102_73 ();
 sg13g2_decap_4 FILLER_102_92 ();
 sg13g2_decap_8 FILLER_102_117 ();
 sg13g2_fill_1 FILLER_102_124 ();
 sg13g2_fill_1 FILLER_102_199 ();
 sg13g2_fill_1 FILLER_103_38 ();
 sg13g2_fill_2 FILLER_103_56 ();
 sg13g2_fill_1 FILLER_103_58 ();
 sg13g2_fill_1 FILLER_103_67 ();
 sg13g2_fill_2 FILLER_103_77 ();
 sg13g2_fill_1 FILLER_103_96 ();
 sg13g2_fill_1 FILLER_103_152 ();
 sg13g2_fill_1 FILLER_103_199 ();
 sg13g2_fill_1 FILLER_104_0 ();
 sg13g2_fill_1 FILLER_104_26 ();
 sg13g2_fill_2 FILLER_104_67 ();
 sg13g2_decap_8 FILLER_104_120 ();
 sg13g2_fill_2 FILLER_104_127 ();
 sg13g2_fill_1 FILLER_104_129 ();
 sg13g2_fill_2 FILLER_104_198 ();
 sg13g2_fill_1 FILLER_105_21 ();
 sg13g2_fill_1 FILLER_105_25 ();
 sg13g2_fill_2 FILLER_105_54 ();
 sg13g2_fill_2 FILLER_105_85 ();
 sg13g2_fill_1 FILLER_105_87 ();
 sg13g2_fill_1 FILLER_105_109 ();
 sg13g2_fill_1 FILLER_105_151 ();
 sg13g2_fill_1 FILLER_105_178 ();
 sg13g2_fill_1 FILLER_105_199 ();
 sg13g2_fill_2 FILLER_106_17 ();
 sg13g2_fill_2 FILLER_106_101 ();
 sg13g2_fill_1 FILLER_106_103 ();
 sg13g2_fill_1 FILLER_106_179 ();
 sg13g2_fill_2 FILLER_107_21 ();
 sg13g2_fill_1 FILLER_107_136 ();
 sg13g2_fill_1 FILLER_107_161 ();
 sg13g2_fill_2 FILLER_107_179 ();
 sg13g2_fill_2 FILLER_107_198 ();
 sg13g2_fill_1 FILLER_108_0 ();
 sg13g2_fill_1 FILLER_108_18 ();
 sg13g2_fill_1 FILLER_108_43 ();
 sg13g2_fill_1 FILLER_108_77 ();
 sg13g2_fill_2 FILLER_108_112 ();
 sg13g2_fill_2 FILLER_108_125 ();
 sg13g2_fill_1 FILLER_109_0 ();
 sg13g2_fill_2 FILLER_109_59 ();
 sg13g2_fill_2 FILLER_109_112 ();
 sg13g2_fill_1 FILLER_109_158 ();
 sg13g2_fill_2 FILLER_109_184 ();
 sg13g2_fill_1 FILLER_109_199 ();
 sg13g2_fill_1 FILLER_110_0 ();
 sg13g2_fill_1 FILLER_110_60 ();
 sg13g2_fill_2 FILLER_110_65 ();
 sg13g2_fill_2 FILLER_110_113 ();
endmodule
