VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO eFPGA
  CLASS BLOCK ;
  FOREIGN eFPGA ;
  ORIGIN 0.000 0.000 ;
  SIZE 1076.160 BY 1832.520 ;
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1778.500 0.880 1778.900 ;
    END
  END FrameData[0]
  PIN FrameData[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1265.260 0.860 1265.660 ;
    END
  END FrameData[100]
  PIN FrameData[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1267.780 0.880 1268.180 ;
    END
  END FrameData[101]
  PIN FrameData[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1270.300 0.880 1270.700 ;
    END
  END FrameData[102]
  PIN FrameData[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1272.820 0.880 1273.220 ;
    END
  END FrameData[103]
  PIN FrameData[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1275.340 0.880 1275.740 ;
    END
  END FrameData[104]
  PIN FrameData[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1277.860 0.880 1278.260 ;
    END
  END FrameData[105]
  PIN FrameData[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1280.380 0.880 1280.780 ;
    END
  END FrameData[106]
  PIN FrameData[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1282.900 0.880 1283.300 ;
    END
  END FrameData[107]
  PIN FrameData[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1285.420 0.880 1285.820 ;
    END
  END FrameData[108]
  PIN FrameData[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1287.940 0.880 1288.340 ;
    END
  END FrameData[109]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1795.300 0.880 1795.700 ;
    END
  END FrameData[10]
  PIN FrameData[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1290.460 0.880 1290.860 ;
    END
  END FrameData[110]
  PIN FrameData[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1292.980 0.880 1293.380 ;
    END
  END FrameData[111]
  PIN FrameData[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1295.500 0.880 1295.900 ;
    END
  END FrameData[112]
  PIN FrameData[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1298.020 0.880 1298.420 ;
    END
  END FrameData[113]
  PIN FrameData[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1300.540 0.880 1300.940 ;
    END
  END FrameData[114]
  PIN FrameData[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1303.060 0.880 1303.460 ;
    END
  END FrameData[115]
  PIN FrameData[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1305.580 0.880 1305.980 ;
    END
  END FrameData[116]
  PIN FrameData[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1308.100 0.880 1308.500 ;
    END
  END FrameData[117]
  PIN FrameData[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1310.620 0.880 1311.020 ;
    END
  END FrameData[118]
  PIN FrameData[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1313.140 0.880 1313.540 ;
    END
  END FrameData[119]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1796.980 0.880 1797.380 ;
    END
  END FrameData[11]
  PIN FrameData[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1315.660 0.880 1316.060 ;
    END
  END FrameData[120]
  PIN FrameData[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1318.180 0.880 1318.580 ;
    END
  END FrameData[121]
  PIN FrameData[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1320.700 0.880 1321.100 ;
    END
  END FrameData[122]
  PIN FrameData[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1323.220 0.880 1323.620 ;
    END
  END FrameData[123]
  PIN FrameData[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1325.740 0.880 1326.140 ;
    END
  END FrameData[124]
  PIN FrameData[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1328.260 0.880 1328.660 ;
    END
  END FrameData[125]
  PIN FrameData[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1330.780 0.880 1331.180 ;
    END
  END FrameData[126]
  PIN FrameData[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1333.300 0.880 1333.700 ;
    END
  END FrameData[127]
  PIN FrameData[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1040.140 0.880 1040.540 ;
    END
  END FrameData[128]
  PIN FrameData[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1042.660 0.880 1043.060 ;
    END
  END FrameData[129]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1798.660 0.880 1799.060 ;
    END
  END FrameData[12]
  PIN FrameData[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1045.180 0.880 1045.580 ;
    END
  END FrameData[130]
  PIN FrameData[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1047.700 0.880 1048.100 ;
    END
  END FrameData[131]
  PIN FrameData[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1050.220 0.860 1050.620 ;
    END
  END FrameData[132]
  PIN FrameData[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1052.740 0.880 1053.140 ;
    END
  END FrameData[133]
  PIN FrameData[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1055.260 0.880 1055.660 ;
    END
  END FrameData[134]
  PIN FrameData[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1057.780 0.880 1058.180 ;
    END
  END FrameData[135]
  PIN FrameData[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1060.300 0.880 1060.700 ;
    END
  END FrameData[136]
  PIN FrameData[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1062.820 0.880 1063.220 ;
    END
  END FrameData[137]
  PIN FrameData[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1065.340 0.880 1065.740 ;
    END
  END FrameData[138]
  PIN FrameData[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1067.860 0.880 1068.260 ;
    END
  END FrameData[139]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1800.340 0.880 1800.740 ;
    END
  END FrameData[13]
  PIN FrameData[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1070.380 0.880 1070.780 ;
    END
  END FrameData[140]
  PIN FrameData[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1072.900 0.880 1073.300 ;
    END
  END FrameData[141]
  PIN FrameData[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1075.420 0.880 1075.820 ;
    END
  END FrameData[142]
  PIN FrameData[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1077.940 0.880 1078.340 ;
    END
  END FrameData[143]
  PIN FrameData[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1080.460 0.880 1080.860 ;
    END
  END FrameData[144]
  PIN FrameData[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1082.980 0.880 1083.380 ;
    END
  END FrameData[145]
  PIN FrameData[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1085.500 0.880 1085.900 ;
    END
  END FrameData[146]
  PIN FrameData[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1088.020 0.880 1088.420 ;
    END
  END FrameData[147]
  PIN FrameData[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1090.540 0.880 1090.940 ;
    END
  END FrameData[148]
  PIN FrameData[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1093.060 0.880 1093.460 ;
    END
  END FrameData[149]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1802.020 0.880 1802.420 ;
    END
  END FrameData[14]
  PIN FrameData[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1095.580 0.880 1095.980 ;
    END
  END FrameData[150]
  PIN FrameData[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1098.100 0.880 1098.500 ;
    END
  END FrameData[151]
  PIN FrameData[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1100.620 0.880 1101.020 ;
    END
  END FrameData[152]
  PIN FrameData[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1103.140 0.880 1103.540 ;
    END
  END FrameData[153]
  PIN FrameData[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1105.660 0.880 1106.060 ;
    END
  END FrameData[154]
  PIN FrameData[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1108.180 0.880 1108.580 ;
    END
  END FrameData[155]
  PIN FrameData[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1110.700 0.880 1111.100 ;
    END
  END FrameData[156]
  PIN FrameData[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1113.220 0.880 1113.620 ;
    END
  END FrameData[157]
  PIN FrameData[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1115.740 0.880 1116.140 ;
    END
  END FrameData[158]
  PIN FrameData[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1118.260 0.880 1118.660 ;
    END
  END FrameData[159]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1803.700 0.880 1804.100 ;
    END
  END FrameData[15]
  PIN FrameData[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 825.100 0.880 825.500 ;
    END
  END FrameData[160]
  PIN FrameData[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 827.620 0.880 828.020 ;
    END
  END FrameData[161]
  PIN FrameData[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 830.140 0.880 830.540 ;
    END
  END FrameData[162]
  PIN FrameData[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 832.660 0.880 833.060 ;
    END
  END FrameData[163]
  PIN FrameData[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 835.180 0.860 835.580 ;
    END
  END FrameData[164]
  PIN FrameData[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 837.700 0.880 838.100 ;
    END
  END FrameData[165]
  PIN FrameData[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 840.220 0.880 840.620 ;
    END
  END FrameData[166]
  PIN FrameData[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 842.740 0.880 843.140 ;
    END
  END FrameData[167]
  PIN FrameData[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 845.260 0.880 845.660 ;
    END
  END FrameData[168]
  PIN FrameData[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 847.780 0.880 848.180 ;
    END
  END FrameData[169]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1805.380 0.880 1805.780 ;
    END
  END FrameData[16]
  PIN FrameData[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 850.300 0.880 850.700 ;
    END
  END FrameData[170]
  PIN FrameData[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 852.820 0.880 853.220 ;
    END
  END FrameData[171]
  PIN FrameData[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 855.340 0.880 855.740 ;
    END
  END FrameData[172]
  PIN FrameData[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 857.860 0.880 858.260 ;
    END
  END FrameData[173]
  PIN FrameData[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 860.380 0.880 860.780 ;
    END
  END FrameData[174]
  PIN FrameData[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 862.900 0.880 863.300 ;
    END
  END FrameData[175]
  PIN FrameData[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 865.420 0.880 865.820 ;
    END
  END FrameData[176]
  PIN FrameData[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 867.940 0.880 868.340 ;
    END
  END FrameData[177]
  PIN FrameData[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 870.460 0.880 870.860 ;
    END
  END FrameData[178]
  PIN FrameData[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 872.980 0.880 873.380 ;
    END
  END FrameData[179]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1807.060 0.880 1807.460 ;
    END
  END FrameData[17]
  PIN FrameData[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 875.500 0.880 875.900 ;
    END
  END FrameData[180]
  PIN FrameData[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 878.020 0.880 878.420 ;
    END
  END FrameData[181]
  PIN FrameData[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 880.540 0.880 880.940 ;
    END
  END FrameData[182]
  PIN FrameData[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 883.060 0.880 883.460 ;
    END
  END FrameData[183]
  PIN FrameData[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 885.580 0.880 885.980 ;
    END
  END FrameData[184]
  PIN FrameData[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 888.100 0.880 888.500 ;
    END
  END FrameData[185]
  PIN FrameData[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 890.620 0.880 891.020 ;
    END
  END FrameData[186]
  PIN FrameData[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 893.140 0.880 893.540 ;
    END
  END FrameData[187]
  PIN FrameData[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 895.660 0.880 896.060 ;
    END
  END FrameData[188]
  PIN FrameData[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 898.180 0.880 898.580 ;
    END
  END FrameData[189]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1808.740 0.880 1809.140 ;
    END
  END FrameData[18]
  PIN FrameData[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 900.700 0.880 901.100 ;
    END
  END FrameData[190]
  PIN FrameData[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 903.220 0.880 903.620 ;
    END
  END FrameData[191]
  PIN FrameData[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 610.060 0.880 610.460 ;
    END
  END FrameData[192]
  PIN FrameData[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 612.580 0.880 612.980 ;
    END
  END FrameData[193]
  PIN FrameData[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 615.100 0.880 615.500 ;
    END
  END FrameData[194]
  PIN FrameData[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 617.620 0.880 618.020 ;
    END
  END FrameData[195]
  PIN FrameData[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 620.140 0.860 620.540 ;
    END
  END FrameData[196]
  PIN FrameData[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 622.660 0.880 623.060 ;
    END
  END FrameData[197]
  PIN FrameData[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 625.180 0.880 625.580 ;
    END
  END FrameData[198]
  PIN FrameData[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 627.700 0.880 628.100 ;
    END
  END FrameData[199]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1810.420 0.880 1810.820 ;
    END
  END FrameData[19]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1780.180 0.880 1780.580 ;
    END
  END FrameData[1]
  PIN FrameData[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 630.220 0.880 630.620 ;
    END
  END FrameData[200]
  PIN FrameData[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 632.740 0.880 633.140 ;
    END
  END FrameData[201]
  PIN FrameData[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 635.260 0.880 635.660 ;
    END
  END FrameData[202]
  PIN FrameData[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 637.780 0.880 638.180 ;
    END
  END FrameData[203]
  PIN FrameData[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 640.300 0.880 640.700 ;
    END
  END FrameData[204]
  PIN FrameData[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 642.820 0.880 643.220 ;
    END
  END FrameData[205]
  PIN FrameData[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 645.340 0.880 645.740 ;
    END
  END FrameData[206]
  PIN FrameData[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 647.860 0.880 648.260 ;
    END
  END FrameData[207]
  PIN FrameData[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 650.380 0.880 650.780 ;
    END
  END FrameData[208]
  PIN FrameData[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 652.900 0.880 653.300 ;
    END
  END FrameData[209]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1812.100 0.880 1812.500 ;
    END
  END FrameData[20]
  PIN FrameData[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 655.420 0.880 655.820 ;
    END
  END FrameData[210]
  PIN FrameData[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 657.940 0.880 658.340 ;
    END
  END FrameData[211]
  PIN FrameData[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 660.460 0.880 660.860 ;
    END
  END FrameData[212]
  PIN FrameData[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 662.980 0.880 663.380 ;
    END
  END FrameData[213]
  PIN FrameData[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 665.500 0.880 665.900 ;
    END
  END FrameData[214]
  PIN FrameData[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 668.020 0.880 668.420 ;
    END
  END FrameData[215]
  PIN FrameData[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 670.540 0.880 670.940 ;
    END
  END FrameData[216]
  PIN FrameData[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 673.060 0.880 673.460 ;
    END
  END FrameData[217]
  PIN FrameData[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 675.580 0.880 675.980 ;
    END
  END FrameData[218]
  PIN FrameData[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 678.100 0.880 678.500 ;
    END
  END FrameData[219]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1813.780 0.880 1814.180 ;
    END
  END FrameData[21]
  PIN FrameData[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 680.620 0.880 681.020 ;
    END
  END FrameData[220]
  PIN FrameData[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 683.140 0.880 683.540 ;
    END
  END FrameData[221]
  PIN FrameData[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 685.660 0.880 686.060 ;
    END
  END FrameData[222]
  PIN FrameData[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 688.180 0.880 688.580 ;
    END
  END FrameData[223]
  PIN FrameData[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 395.020 0.880 395.420 ;
    END
  END FrameData[224]
  PIN FrameData[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 397.540 0.880 397.940 ;
    END
  END FrameData[225]
  PIN FrameData[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 400.060 0.880 400.460 ;
    END
  END FrameData[226]
  PIN FrameData[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 402.580 0.880 402.980 ;
    END
  END FrameData[227]
  PIN FrameData[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 405.100 0.860 405.500 ;
    END
  END FrameData[228]
  PIN FrameData[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 407.620 0.880 408.020 ;
    END
  END FrameData[229]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1815.460 0.880 1815.860 ;
    END
  END FrameData[22]
  PIN FrameData[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 410.140 0.880 410.540 ;
    END
  END FrameData[230]
  PIN FrameData[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 412.660 0.880 413.060 ;
    END
  END FrameData[231]
  PIN FrameData[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 415.180 0.880 415.580 ;
    END
  END FrameData[232]
  PIN FrameData[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 417.700 0.880 418.100 ;
    END
  END FrameData[233]
  PIN FrameData[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 420.220 0.880 420.620 ;
    END
  END FrameData[234]
  PIN FrameData[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 422.740 0.880 423.140 ;
    END
  END FrameData[235]
  PIN FrameData[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 425.260 0.880 425.660 ;
    END
  END FrameData[236]
  PIN FrameData[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 427.780 0.880 428.180 ;
    END
  END FrameData[237]
  PIN FrameData[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 430.300 0.880 430.700 ;
    END
  END FrameData[238]
  PIN FrameData[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 432.820 0.880 433.220 ;
    END
  END FrameData[239]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1817.140 0.880 1817.540 ;
    END
  END FrameData[23]
  PIN FrameData[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 435.340 0.880 435.740 ;
    END
  END FrameData[240]
  PIN FrameData[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 437.860 0.880 438.260 ;
    END
  END FrameData[241]
  PIN FrameData[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 440.380 0.880 440.780 ;
    END
  END FrameData[242]
  PIN FrameData[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 442.900 0.880 443.300 ;
    END
  END FrameData[243]
  PIN FrameData[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 445.420 0.880 445.820 ;
    END
  END FrameData[244]
  PIN FrameData[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 447.940 0.880 448.340 ;
    END
  END FrameData[245]
  PIN FrameData[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 450.460 0.880 450.860 ;
    END
  END FrameData[246]
  PIN FrameData[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 452.980 0.880 453.380 ;
    END
  END FrameData[247]
  PIN FrameData[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 455.500 0.880 455.900 ;
    END
  END FrameData[248]
  PIN FrameData[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 458.020 0.880 458.420 ;
    END
  END FrameData[249]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1818.820 0.880 1819.220 ;
    END
  END FrameData[24]
  PIN FrameData[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 460.540 0.880 460.940 ;
    END
  END FrameData[250]
  PIN FrameData[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 463.060 0.880 463.460 ;
    END
  END FrameData[251]
  PIN FrameData[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 465.580 0.880 465.980 ;
    END
  END FrameData[252]
  PIN FrameData[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 468.100 0.880 468.500 ;
    END
  END FrameData[253]
  PIN FrameData[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 470.620 0.880 471.020 ;
    END
  END FrameData[254]
  PIN FrameData[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 473.140 0.880 473.540 ;
    END
  END FrameData[255]
  PIN FrameData[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 179.980 0.880 180.380 ;
    END
  END FrameData[256]
  PIN FrameData[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 182.500 0.880 182.900 ;
    END
  END FrameData[257]
  PIN FrameData[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 185.020 0.880 185.420 ;
    END
  END FrameData[258]
  PIN FrameData[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 187.540 0.880 187.940 ;
    END
  END FrameData[259]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1820.500 0.880 1820.900 ;
    END
  END FrameData[25]
  PIN FrameData[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 190.060 0.860 190.460 ;
    END
  END FrameData[260]
  PIN FrameData[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 192.580 0.880 192.980 ;
    END
  END FrameData[261]
  PIN FrameData[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 195.100 0.880 195.500 ;
    END
  END FrameData[262]
  PIN FrameData[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 197.620 0.880 198.020 ;
    END
  END FrameData[263]
  PIN FrameData[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 200.140 0.880 200.540 ;
    END
  END FrameData[264]
  PIN FrameData[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 202.660 0.880 203.060 ;
    END
  END FrameData[265]
  PIN FrameData[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 205.180 0.880 205.580 ;
    END
  END FrameData[266]
  PIN FrameData[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 207.700 0.880 208.100 ;
    END
  END FrameData[267]
  PIN FrameData[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 210.220 0.880 210.620 ;
    END
  END FrameData[268]
  PIN FrameData[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 212.740 0.880 213.140 ;
    END
  END FrameData[269]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1822.180 0.880 1822.580 ;
    END
  END FrameData[26]
  PIN FrameData[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 215.260 0.880 215.660 ;
    END
  END FrameData[270]
  PIN FrameData[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 217.780 0.880 218.180 ;
    END
  END FrameData[271]
  PIN FrameData[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 220.300 0.880 220.700 ;
    END
  END FrameData[272]
  PIN FrameData[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 222.820 0.880 223.220 ;
    END
  END FrameData[273]
  PIN FrameData[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 225.340 0.880 225.740 ;
    END
  END FrameData[274]
  PIN FrameData[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 227.860 0.880 228.260 ;
    END
  END FrameData[275]
  PIN FrameData[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 230.380 0.880 230.780 ;
    END
  END FrameData[276]
  PIN FrameData[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 232.900 0.880 233.300 ;
    END
  END FrameData[277]
  PIN FrameData[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 235.420 0.880 235.820 ;
    END
  END FrameData[278]
  PIN FrameData[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 237.940 0.880 238.340 ;
    END
  END FrameData[279]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1823.860 0.880 1824.260 ;
    END
  END FrameData[27]
  PIN FrameData[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 240.460 0.880 240.860 ;
    END
  END FrameData[280]
  PIN FrameData[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 242.980 0.880 243.380 ;
    END
  END FrameData[281]
  PIN FrameData[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 245.500 0.880 245.900 ;
    END
  END FrameData[282]
  PIN FrameData[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 248.020 0.880 248.420 ;
    END
  END FrameData[283]
  PIN FrameData[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 250.540 0.880 250.940 ;
    END
  END FrameData[284]
  PIN FrameData[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 253.060 0.880 253.460 ;
    END
  END FrameData[285]
  PIN FrameData[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 255.580 0.880 255.980 ;
    END
  END FrameData[286]
  PIN FrameData[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 258.100 0.880 258.500 ;
    END
  END FrameData[287]
  PIN FrameData[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 4.420 0.880 4.820 ;
    END
  END FrameData[288]
  PIN FrameData[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 6.100 0.880 6.500 ;
    END
  END FrameData[289]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1825.540 0.880 1825.940 ;
    END
  END FrameData[28]
  PIN FrameData[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 7.780 0.880 8.180 ;
    END
  END FrameData[290]
  PIN FrameData[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 9.460 0.880 9.860 ;
    END
  END FrameData[291]
  PIN FrameData[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 11.140 0.880 11.540 ;
    END
  END FrameData[292]
  PIN FrameData[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 12.820 0.880 13.220 ;
    END
  END FrameData[293]
  PIN FrameData[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 14.500 0.880 14.900 ;
    END
  END FrameData[294]
  PIN FrameData[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 16.180 0.880 16.580 ;
    END
  END FrameData[295]
  PIN FrameData[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 17.860 0.880 18.260 ;
    END
  END FrameData[296]
  PIN FrameData[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 19.540 0.880 19.940 ;
    END
  END FrameData[297]
  PIN FrameData[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 21.220 0.880 21.620 ;
    END
  END FrameData[298]
  PIN FrameData[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 22.900 0.880 23.300 ;
    END
  END FrameData[299]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1827.220 0.880 1827.620 ;
    END
  END FrameData[29]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1781.860 0.880 1782.260 ;
    END
  END FrameData[2]
  PIN FrameData[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 24.580 0.880 24.980 ;
    END
  END FrameData[300]
  PIN FrameData[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 26.260 0.880 26.660 ;
    END
  END FrameData[301]
  PIN FrameData[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 27.940 0.880 28.340 ;
    END
  END FrameData[302]
  PIN FrameData[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 29.620 0.880 30.020 ;
    END
  END FrameData[303]
  PIN FrameData[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 31.300 0.880 31.700 ;
    END
  END FrameData[304]
  PIN FrameData[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 32.980 0.880 33.380 ;
    END
  END FrameData[305]
  PIN FrameData[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 34.660 0.880 35.060 ;
    END
  END FrameData[306]
  PIN FrameData[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 36.340 0.880 36.740 ;
    END
  END FrameData[307]
  PIN FrameData[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 38.020 0.880 38.420 ;
    END
  END FrameData[308]
  PIN FrameData[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 39.700 0.880 40.100 ;
    END
  END FrameData[309]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1828.900 0.880 1829.300 ;
    END
  END FrameData[30]
  PIN FrameData[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 41.380 0.880 41.780 ;
    END
  END FrameData[310]
  PIN FrameData[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 43.060 0.880 43.460 ;
    END
  END FrameData[311]
  PIN FrameData[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 44.740 0.880 45.140 ;
    END
  END FrameData[312]
  PIN FrameData[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 46.420 0.880 46.820 ;
    END
  END FrameData[313]
  PIN FrameData[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 48.100 0.880 48.500 ;
    END
  END FrameData[314]
  PIN FrameData[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 49.780 0.880 50.180 ;
    END
  END FrameData[315]
  PIN FrameData[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 51.460 0.880 51.860 ;
    END
  END FrameData[316]
  PIN FrameData[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 53.140 0.880 53.540 ;
    END
  END FrameData[317]
  PIN FrameData[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 54.820 0.880 55.220 ;
    END
  END FrameData[318]
  PIN FrameData[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 56.500 0.880 56.900 ;
    END
  END FrameData[319]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1830.580 0.880 1830.980 ;
    END
  END FrameData[31]
  PIN FrameData[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1685.260 0.880 1685.660 ;
    END
  END FrameData[32]
  PIN FrameData[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1687.780 0.880 1688.180 ;
    END
  END FrameData[33]
  PIN FrameData[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1690.300 0.880 1690.700 ;
    END
  END FrameData[34]
  PIN FrameData[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1692.820 0.880 1693.220 ;
    END
  END FrameData[35]
  PIN FrameData[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1695.340 0.860 1695.740 ;
    END
  END FrameData[36]
  PIN FrameData[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1697.860 0.880 1698.260 ;
    END
  END FrameData[37]
  PIN FrameData[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1700.380 0.880 1700.780 ;
    END
  END FrameData[38]
  PIN FrameData[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1702.900 0.880 1703.300 ;
    END
  END FrameData[39]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1783.540 0.880 1783.940 ;
    END
  END FrameData[3]
  PIN FrameData[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1705.420 0.880 1705.820 ;
    END
  END FrameData[40]
  PIN FrameData[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1707.940 0.880 1708.340 ;
    END
  END FrameData[41]
  PIN FrameData[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1710.460 0.880 1710.860 ;
    END
  END FrameData[42]
  PIN FrameData[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1712.980 0.880 1713.380 ;
    END
  END FrameData[43]
  PIN FrameData[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1715.500 0.880 1715.900 ;
    END
  END FrameData[44]
  PIN FrameData[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1718.020 0.880 1718.420 ;
    END
  END FrameData[45]
  PIN FrameData[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1720.540 0.880 1720.940 ;
    END
  END FrameData[46]
  PIN FrameData[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1723.060 0.880 1723.460 ;
    END
  END FrameData[47]
  PIN FrameData[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1725.580 0.880 1725.980 ;
    END
  END FrameData[48]
  PIN FrameData[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1728.100 0.880 1728.500 ;
    END
  END FrameData[49]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1785.220 0.880 1785.620 ;
    END
  END FrameData[4]
  PIN FrameData[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1730.620 0.880 1731.020 ;
    END
  END FrameData[50]
  PIN FrameData[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1733.140 0.880 1733.540 ;
    END
  END FrameData[51]
  PIN FrameData[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1735.660 0.880 1736.060 ;
    END
  END FrameData[52]
  PIN FrameData[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1738.180 0.880 1738.580 ;
    END
  END FrameData[53]
  PIN FrameData[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1740.700 0.880 1741.100 ;
    END
  END FrameData[54]
  PIN FrameData[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1743.220 0.880 1743.620 ;
    END
  END FrameData[55]
  PIN FrameData[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1745.740 0.880 1746.140 ;
    END
  END FrameData[56]
  PIN FrameData[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1748.260 0.880 1748.660 ;
    END
  END FrameData[57]
  PIN FrameData[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1750.780 0.880 1751.180 ;
    END
  END FrameData[58]
  PIN FrameData[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1753.300 0.880 1753.700 ;
    END
  END FrameData[59]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1786.900 0.880 1787.300 ;
    END
  END FrameData[5]
  PIN FrameData[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1755.820 0.880 1756.220 ;
    END
  END FrameData[60]
  PIN FrameData[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1758.340 0.880 1758.740 ;
    END
  END FrameData[61]
  PIN FrameData[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1760.860 0.880 1761.260 ;
    END
  END FrameData[62]
  PIN FrameData[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1763.380 0.880 1763.780 ;
    END
  END FrameData[63]
  PIN FrameData[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1470.220 0.880 1470.620 ;
    END
  END FrameData[64]
  PIN FrameData[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1472.740 0.880 1473.140 ;
    END
  END FrameData[65]
  PIN FrameData[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1475.260 0.880 1475.660 ;
    END
  END FrameData[66]
  PIN FrameData[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1477.780 0.880 1478.180 ;
    END
  END FrameData[67]
  PIN FrameData[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1480.300 0.860 1480.700 ;
    END
  END FrameData[68]
  PIN FrameData[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1482.820 0.880 1483.220 ;
    END
  END FrameData[69]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1788.580 0.880 1788.980 ;
    END
  END FrameData[6]
  PIN FrameData[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1485.340 0.880 1485.740 ;
    END
  END FrameData[70]
  PIN FrameData[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1487.860 0.880 1488.260 ;
    END
  END FrameData[71]
  PIN FrameData[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1490.380 0.880 1490.780 ;
    END
  END FrameData[72]
  PIN FrameData[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1492.900 0.880 1493.300 ;
    END
  END FrameData[73]
  PIN FrameData[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1495.420 0.880 1495.820 ;
    END
  END FrameData[74]
  PIN FrameData[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1497.940 0.880 1498.340 ;
    END
  END FrameData[75]
  PIN FrameData[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1500.460 0.880 1500.860 ;
    END
  END FrameData[76]
  PIN FrameData[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1502.980 0.880 1503.380 ;
    END
  END FrameData[77]
  PIN FrameData[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1505.500 0.880 1505.900 ;
    END
  END FrameData[78]
  PIN FrameData[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1508.020 0.880 1508.420 ;
    END
  END FrameData[79]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1790.260 0.880 1790.660 ;
    END
  END FrameData[7]
  PIN FrameData[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1510.540 0.880 1510.940 ;
    END
  END FrameData[80]
  PIN FrameData[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1513.060 0.880 1513.460 ;
    END
  END FrameData[81]
  PIN FrameData[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1515.580 0.880 1515.980 ;
    END
  END FrameData[82]
  PIN FrameData[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1518.100 0.880 1518.500 ;
    END
  END FrameData[83]
  PIN FrameData[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1520.620 0.880 1521.020 ;
    END
  END FrameData[84]
  PIN FrameData[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1523.140 0.880 1523.540 ;
    END
  END FrameData[85]
  PIN FrameData[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1525.660 0.880 1526.060 ;
    END
  END FrameData[86]
  PIN FrameData[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1528.180 0.880 1528.580 ;
    END
  END FrameData[87]
  PIN FrameData[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1530.700 0.880 1531.100 ;
    END
  END FrameData[88]
  PIN FrameData[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1533.220 0.880 1533.620 ;
    END
  END FrameData[89]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1791.940 0.880 1792.340 ;
    END
  END FrameData[8]
  PIN FrameData[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1535.740 0.880 1536.140 ;
    END
  END FrameData[90]
  PIN FrameData[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1538.260 0.880 1538.660 ;
    END
  END FrameData[91]
  PIN FrameData[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1540.780 0.880 1541.180 ;
    END
  END FrameData[92]
  PIN FrameData[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1543.300 0.880 1543.700 ;
    END
  END FrameData[93]
  PIN FrameData[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1545.820 0.880 1546.220 ;
    END
  END FrameData[94]
  PIN FrameData[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1548.340 0.880 1548.740 ;
    END
  END FrameData[95]
  PIN FrameData[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1255.180 0.880 1255.580 ;
    END
  END FrameData[96]
  PIN FrameData[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1257.700 0.880 1258.100 ;
    END
  END FrameData[97]
  PIN FrameData[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1260.220 0.880 1260.620 ;
    END
  END FrameData[98]
  PIN FrameData[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1262.740 0.880 1263.140 ;
    END
  END FrameData[99]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1793.620 0.880 1794.020 ;
    END
  END FrameData[9]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 10.360 0.000 10.760 0.480 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 978.040 0.000 978.440 0.480 ;
    END
  END FrameStrobe[100]
  PIN FrameStrobe[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 982.840 0.000 983.240 0.480 ;
    END
  END FrameStrobe[101]
  PIN FrameStrobe[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 987.640 0.000 988.040 0.480 ;
    END
  END FrameStrobe[102]
  PIN FrameStrobe[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 992.440 0.000 992.840 0.480 ;
    END
  END FrameStrobe[103]
  PIN FrameStrobe[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 997.240 0.000 997.640 0.480 ;
    END
  END FrameStrobe[104]
  PIN FrameStrobe[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 1002.040 0.000 1002.440 0.480 ;
    END
  END FrameStrobe[105]
  PIN FrameStrobe[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 1006.840 0.000 1007.240 0.480 ;
    END
  END FrameStrobe[106]
  PIN FrameStrobe[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 1011.640 0.000 1012.040 0.480 ;
    END
  END FrameStrobe[107]
  PIN FrameStrobe[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 1016.440 0.000 1016.840 0.480 ;
    END
  END FrameStrobe[108]
  PIN FrameStrobe[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 1021.240 0.000 1021.640 0.480 ;
    END
  END FrameStrobe[109]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 58.360 0.000 58.760 0.480 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 1026.040 0.000 1026.440 0.480 ;
    END
  END FrameStrobe[110]
  PIN FrameStrobe[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 1030.840 0.000 1031.240 0.480 ;
    END
  END FrameStrobe[111]
  PIN FrameStrobe[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 1035.640 0.000 1036.040 0.480 ;
    END
  END FrameStrobe[112]
  PIN FrameStrobe[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 1040.440 0.000 1040.840 0.480 ;
    END
  END FrameStrobe[113]
  PIN FrameStrobe[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 1045.240 0.000 1045.640 0.480 ;
    END
  END FrameStrobe[114]
  PIN FrameStrobe[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 1050.040 0.000 1050.440 0.480 ;
    END
  END FrameStrobe[115]
  PIN FrameStrobe[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 1054.840 0.000 1055.240 0.480 ;
    END
  END FrameStrobe[116]
  PIN FrameStrobe[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 1059.640 0.000 1060.040 0.480 ;
    END
  END FrameStrobe[117]
  PIN FrameStrobe[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 1064.440 0.000 1064.840 0.480 ;
    END
  END FrameStrobe[118]
  PIN FrameStrobe[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 1069.240 0.000 1069.640 0.480 ;
    END
  END FrameStrobe[119]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 63.160 0.000 63.560 0.480 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 67.960 0.000 68.360 0.480 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 72.760 0.000 73.160 0.480 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 77.560 0.000 77.960 0.480 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 82.360 0.000 82.760 0.480 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 87.160 0.000 87.560 0.480 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 91.960 0.000 92.360 0.480 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 96.760 0.000 97.160 0.480 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 101.560 0.000 101.960 0.480 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 15.160 0.000 15.560 0.480 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.753500 ;
    PORT
      LAYER Metal2 ;
        RECT 197.560 0.000 197.960 0.480 ;
    END
  END FrameStrobe[20]
  PIN FrameStrobe[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.753500 ;
    PORT
      LAYER Metal2 ;
        RECT 203.320 0.000 203.720 0.480 ;
    END
  END FrameStrobe[21]
  PIN FrameStrobe[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.753500 ;
    PORT
      LAYER Metal2 ;
        RECT 209.080 0.000 209.480 0.480 ;
    END
  END FrameStrobe[22]
  PIN FrameStrobe[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.753500 ;
    PORT
      LAYER Metal2 ;
        RECT 214.840 0.000 215.240 0.480 ;
    END
  END FrameStrobe[23]
  PIN FrameStrobe[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.002300 ;
    PORT
      LAYER Metal2 ;
        RECT 220.600 0.000 221.000 0.480 ;
    END
  END FrameStrobe[24]
  PIN FrameStrobe[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 226.360 0.000 226.760 0.480 ;
    END
  END FrameStrobe[25]
  PIN FrameStrobe[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 232.120 0.000 232.520 0.480 ;
    END
  END FrameStrobe[26]
  PIN FrameStrobe[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 237.880 0.000 238.280 0.480 ;
    END
  END FrameStrobe[27]
  PIN FrameStrobe[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 243.640 0.000 244.040 0.480 ;
    END
  END FrameStrobe[28]
  PIN FrameStrobe[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 249.400 0.000 249.800 0.480 ;
    END
  END FrameStrobe[29]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 19.960 0.000 20.360 0.480 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 255.160 0.000 255.560 0.480 ;
    END
  END FrameStrobe[30]
  PIN FrameStrobe[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 260.920 0.000 261.320 0.480 ;
    END
  END FrameStrobe[31]
  PIN FrameStrobe[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 266.680 0.000 267.080 0.480 ;
    END
  END FrameStrobe[32]
  PIN FrameStrobe[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 272.440 0.000 272.840 0.480 ;
    END
  END FrameStrobe[33]
  PIN FrameStrobe[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 278.200 0.000 278.600 0.480 ;
    END
  END FrameStrobe[34]
  PIN FrameStrobe[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 283.960 0.000 284.360 0.480 ;
    END
  END FrameStrobe[35]
  PIN FrameStrobe[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 289.720 0.000 290.120 0.480 ;
    END
  END FrameStrobe[36]
  PIN FrameStrobe[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 295.480 0.000 295.880 0.480 ;
    END
  END FrameStrobe[37]
  PIN FrameStrobe[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 301.240 0.000 301.640 0.480 ;
    END
  END FrameStrobe[38]
  PIN FrameStrobe[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 307.000 0.000 307.400 0.480 ;
    END
  END FrameStrobe[39]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 24.760 0.000 25.160 0.480 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.753500 ;
    PORT
      LAYER Metal2 ;
        RECT 412.600 0.000 413.000 0.480 ;
    END
  END FrameStrobe[40]
  PIN FrameStrobe[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.753500 ;
    PORT
      LAYER Metal2 ;
        RECT 418.360 0.000 418.760 0.480 ;
    END
  END FrameStrobe[41]
  PIN FrameStrobe[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.753500 ;
    PORT
      LAYER Metal2 ;
        RECT 424.120 0.000 424.520 0.480 ;
    END
  END FrameStrobe[42]
  PIN FrameStrobe[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.753500 ;
    PORT
      LAYER Metal2 ;
        RECT 429.880 0.000 430.280 0.480 ;
    END
  END FrameStrobe[43]
  PIN FrameStrobe[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.002300 ;
    PORT
      LAYER Metal2 ;
        RECT 435.640 0.000 436.040 0.480 ;
    END
  END FrameStrobe[44]
  PIN FrameStrobe[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 441.400 0.000 441.800 0.480 ;
    END
  END FrameStrobe[45]
  PIN FrameStrobe[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 447.160 0.000 447.560 0.480 ;
    END
  END FrameStrobe[46]
  PIN FrameStrobe[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 452.920 0.000 453.320 0.480 ;
    END
  END FrameStrobe[47]
  PIN FrameStrobe[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 458.680 0.000 459.080 0.480 ;
    END
  END FrameStrobe[48]
  PIN FrameStrobe[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 464.440 0.000 464.840 0.480 ;
    END
  END FrameStrobe[49]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 29.560 0.000 29.960 0.480 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 470.200 0.000 470.600 0.480 ;
    END
  END FrameStrobe[50]
  PIN FrameStrobe[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 475.960 0.000 476.360 0.480 ;
    END
  END FrameStrobe[51]
  PIN FrameStrobe[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 481.720 0.000 482.120 0.480 ;
    END
  END FrameStrobe[52]
  PIN FrameStrobe[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 487.480 0.000 487.880 0.480 ;
    END
  END FrameStrobe[53]
  PIN FrameStrobe[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 493.240 0.000 493.640 0.480 ;
    END
  END FrameStrobe[54]
  PIN FrameStrobe[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 499.000 0.000 499.400 0.480 ;
    END
  END FrameStrobe[55]
  PIN FrameStrobe[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 504.760 0.000 505.160 0.480 ;
    END
  END FrameStrobe[56]
  PIN FrameStrobe[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 510.520 0.000 510.920 0.480 ;
    END
  END FrameStrobe[57]
  PIN FrameStrobe[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 516.280 0.000 516.680 0.480 ;
    END
  END FrameStrobe[58]
  PIN FrameStrobe[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 522.040 0.000 522.440 0.480 ;
    END
  END FrameStrobe[59]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 34.360 0.000 34.760 0.480 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.753500 ;
    PORT
      LAYER Metal2 ;
        RECT 627.640 0.000 628.040 0.480 ;
    END
  END FrameStrobe[60]
  PIN FrameStrobe[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.753500 ;
    PORT
      LAYER Metal2 ;
        RECT 633.400 0.000 633.800 0.480 ;
    END
  END FrameStrobe[61]
  PIN FrameStrobe[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.753500 ;
    PORT
      LAYER Metal2 ;
        RECT 639.160 0.000 639.560 0.480 ;
    END
  END FrameStrobe[62]
  PIN FrameStrobe[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.753500 ;
    PORT
      LAYER Metal2 ;
        RECT 644.920 0.000 645.320 0.480 ;
    END
  END FrameStrobe[63]
  PIN FrameStrobe[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.002300 ;
    PORT
      LAYER Metal2 ;
        RECT 650.680 0.000 651.080 0.480 ;
    END
  END FrameStrobe[64]
  PIN FrameStrobe[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 656.440 0.000 656.840 0.480 ;
    END
  END FrameStrobe[65]
  PIN FrameStrobe[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 662.200 0.000 662.600 0.480 ;
    END
  END FrameStrobe[66]
  PIN FrameStrobe[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 667.960 0.000 668.360 0.480 ;
    END
  END FrameStrobe[67]
  PIN FrameStrobe[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 673.720 0.000 674.120 0.480 ;
    END
  END FrameStrobe[68]
  PIN FrameStrobe[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 679.480 0.000 679.880 0.480 ;
    END
  END FrameStrobe[69]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 39.160 0.000 39.560 0.480 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 685.240 0.000 685.640 0.480 ;
    END
  END FrameStrobe[70]
  PIN FrameStrobe[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 691.000 0.000 691.400 0.480 ;
    END
  END FrameStrobe[71]
  PIN FrameStrobe[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 696.760 0.000 697.160 0.480 ;
    END
  END FrameStrobe[72]
  PIN FrameStrobe[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 702.520 0.000 702.920 0.480 ;
    END
  END FrameStrobe[73]
  PIN FrameStrobe[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 708.280 0.000 708.680 0.480 ;
    END
  END FrameStrobe[74]
  PIN FrameStrobe[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 714.040 0.000 714.440 0.480 ;
    END
  END FrameStrobe[75]
  PIN FrameStrobe[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 719.800 0.000 720.200 0.480 ;
    END
  END FrameStrobe[76]
  PIN FrameStrobe[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 725.560 0.000 725.960 0.480 ;
    END
  END FrameStrobe[77]
  PIN FrameStrobe[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 731.320 0.000 731.720 0.480 ;
    END
  END FrameStrobe[78]
  PIN FrameStrobe[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 737.080 0.000 737.480 0.480 ;
    END
  END FrameStrobe[79]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 43.960 0.000 44.360 0.480 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.753500 ;
    PORT
      LAYER Metal2 ;
        RECT 842.680 0.000 843.080 0.480 ;
    END
  END FrameStrobe[80]
  PIN FrameStrobe[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.753500 ;
    PORT
      LAYER Metal2 ;
        RECT 848.440 0.000 848.840 0.480 ;
    END
  END FrameStrobe[81]
  PIN FrameStrobe[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.753500 ;
    PORT
      LAYER Metal2 ;
        RECT 854.200 0.000 854.600 0.480 ;
    END
  END FrameStrobe[82]
  PIN FrameStrobe[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.753500 ;
    PORT
      LAYER Metal2 ;
        RECT 859.960 0.000 860.360 0.480 ;
    END
  END FrameStrobe[83]
  PIN FrameStrobe[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.002300 ;
    PORT
      LAYER Metal2 ;
        RECT 865.720 0.000 866.120 0.480 ;
    END
  END FrameStrobe[84]
  PIN FrameStrobe[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 871.480 0.000 871.880 0.480 ;
    END
  END FrameStrobe[85]
  PIN FrameStrobe[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 877.240 0.000 877.640 0.480 ;
    END
  END FrameStrobe[86]
  PIN FrameStrobe[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 883.000 0.000 883.400 0.480 ;
    END
  END FrameStrobe[87]
  PIN FrameStrobe[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 888.760 0.000 889.160 0.480 ;
    END
  END FrameStrobe[88]
  PIN FrameStrobe[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 894.520 0.000 894.920 0.480 ;
    END
  END FrameStrobe[89]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 48.760 0.000 49.160 0.480 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 900.280 0.000 900.680 0.480 ;
    END
  END FrameStrobe[90]
  PIN FrameStrobe[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 906.040 0.000 906.440 0.480 ;
    END
  END FrameStrobe[91]
  PIN FrameStrobe[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 911.800 0.000 912.200 0.480 ;
    END
  END FrameStrobe[92]
  PIN FrameStrobe[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 917.560 0.000 917.960 0.480 ;
    END
  END FrameStrobe[93]
  PIN FrameStrobe[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 923.320 0.000 923.720 0.480 ;
    END
  END FrameStrobe[94]
  PIN FrameStrobe[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 929.080 0.000 929.480 0.480 ;
    END
  END FrameStrobe[95]
  PIN FrameStrobe[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 934.840 0.000 935.240 0.480 ;
    END
  END FrameStrobe[96]
  PIN FrameStrobe[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 940.600 0.000 941.000 0.480 ;
    END
  END FrameStrobe[97]
  PIN FrameStrobe[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 946.360 0.000 946.760 0.480 ;
    END
  END FrameStrobe[98]
  PIN FrameStrobe[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 952.120 0.000 952.520 0.480 ;
    END
  END FrameStrobe[99]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 53.560 0.000 53.960 0.480 ;
    END
  END FrameStrobe[9]
  PIN Tile_X0Y1_CLK_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1680.220 0.880 1680.620 ;
    END
  END Tile_X0Y1_CLK_TT_PROJECT
  PIN Tile_X0Y1_ENA_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1677.700 0.880 1678.100 ;
    END
  END Tile_X0Y1_ENA_TT_PROJECT
  PIN Tile_X0Y1_RST_N_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.615900 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1682.740 0.860 1683.140 ;
    END
  END Tile_X0Y1_RST_N_TT_PROJECT
  PIN Tile_X0Y1_UIO_IN_TT_PROJECT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1657.540 0.880 1657.940 ;
    END
  END Tile_X0Y1_UIO_IN_TT_PROJECT0
  PIN Tile_X0Y1_UIO_IN_TT_PROJECT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1660.060 0.880 1660.460 ;
    END
  END Tile_X0Y1_UIO_IN_TT_PROJECT1
  PIN Tile_X0Y1_UIO_IN_TT_PROJECT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1662.580 0.880 1662.980 ;
    END
  END Tile_X0Y1_UIO_IN_TT_PROJECT2
  PIN Tile_X0Y1_UIO_IN_TT_PROJECT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1665.100 0.880 1665.500 ;
    END
  END Tile_X0Y1_UIO_IN_TT_PROJECT3
  PIN Tile_X0Y1_UIO_IN_TT_PROJECT4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1667.620 0.880 1668.020 ;
    END
  END Tile_X0Y1_UIO_IN_TT_PROJECT4
  PIN Tile_X0Y1_UIO_IN_TT_PROJECT5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1670.140 0.880 1670.540 ;
    END
  END Tile_X0Y1_UIO_IN_TT_PROJECT5
  PIN Tile_X0Y1_UIO_IN_TT_PROJECT6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1672.660 0.880 1673.060 ;
    END
  END Tile_X0Y1_UIO_IN_TT_PROJECT6
  PIN Tile_X0Y1_UIO_IN_TT_PROJECT7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1675.180 0.880 1675.580 ;
    END
  END Tile_X0Y1_UIO_IN_TT_PROJECT7
  PIN Tile_X0Y1_UIO_OE_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1617.220 0.880 1617.620 ;
    END
  END Tile_X0Y1_UIO_OE_TT_PROJECT0
  PIN Tile_X0Y1_UIO_OE_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1619.740 0.880 1620.140 ;
    END
  END Tile_X0Y1_UIO_OE_TT_PROJECT1
  PIN Tile_X0Y1_UIO_OE_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1622.260 0.880 1622.660 ;
    END
  END Tile_X0Y1_UIO_OE_TT_PROJECT2
  PIN Tile_X0Y1_UIO_OE_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1624.780 0.880 1625.180 ;
    END
  END Tile_X0Y1_UIO_OE_TT_PROJECT3
  PIN Tile_X0Y1_UIO_OE_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1627.300 0.880 1627.700 ;
    END
  END Tile_X0Y1_UIO_OE_TT_PROJECT4
  PIN Tile_X0Y1_UIO_OE_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1629.820 0.880 1630.220 ;
    END
  END Tile_X0Y1_UIO_OE_TT_PROJECT5
  PIN Tile_X0Y1_UIO_OE_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1632.340 0.880 1632.740 ;
    END
  END Tile_X0Y1_UIO_OE_TT_PROJECT6
  PIN Tile_X0Y1_UIO_OE_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1634.860 0.880 1635.260 ;
    END
  END Tile_X0Y1_UIO_OE_TT_PROJECT7
  PIN Tile_X0Y1_UIO_OUT_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1597.060 0.880 1597.460 ;
    END
  END Tile_X0Y1_UIO_OUT_TT_PROJECT0
  PIN Tile_X0Y1_UIO_OUT_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1599.580 0.880 1599.980 ;
    END
  END Tile_X0Y1_UIO_OUT_TT_PROJECT1
  PIN Tile_X0Y1_UIO_OUT_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1602.100 0.880 1602.500 ;
    END
  END Tile_X0Y1_UIO_OUT_TT_PROJECT2
  PIN Tile_X0Y1_UIO_OUT_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1604.620 0.880 1605.020 ;
    END
  END Tile_X0Y1_UIO_OUT_TT_PROJECT3
  PIN Tile_X0Y1_UIO_OUT_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1607.140 0.880 1607.540 ;
    END
  END Tile_X0Y1_UIO_OUT_TT_PROJECT4
  PIN Tile_X0Y1_UIO_OUT_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1609.660 0.880 1610.060 ;
    END
  END Tile_X0Y1_UIO_OUT_TT_PROJECT5
  PIN Tile_X0Y1_UIO_OUT_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1612.180 0.880 1612.580 ;
    END
  END Tile_X0Y1_UIO_OUT_TT_PROJECT6
  PIN Tile_X0Y1_UIO_OUT_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1614.700 0.880 1615.100 ;
    END
  END Tile_X0Y1_UIO_OUT_TT_PROJECT7
  PIN Tile_X0Y1_UI_IN_TT_PROJECT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1637.380 0.880 1637.780 ;
    END
  END Tile_X0Y1_UI_IN_TT_PROJECT0
  PIN Tile_X0Y1_UI_IN_TT_PROJECT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1639.900 0.880 1640.300 ;
    END
  END Tile_X0Y1_UI_IN_TT_PROJECT1
  PIN Tile_X0Y1_UI_IN_TT_PROJECT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1642.420 0.880 1642.820 ;
    END
  END Tile_X0Y1_UI_IN_TT_PROJECT2
  PIN Tile_X0Y1_UI_IN_TT_PROJECT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1644.940 0.880 1645.340 ;
    END
  END Tile_X0Y1_UI_IN_TT_PROJECT3
  PIN Tile_X0Y1_UI_IN_TT_PROJECT4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1647.460 0.880 1647.860 ;
    END
  END Tile_X0Y1_UI_IN_TT_PROJECT4
  PIN Tile_X0Y1_UI_IN_TT_PROJECT5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1649.980 0.880 1650.380 ;
    END
  END Tile_X0Y1_UI_IN_TT_PROJECT5
  PIN Tile_X0Y1_UI_IN_TT_PROJECT6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1652.500 0.860 1652.900 ;
    END
  END Tile_X0Y1_UI_IN_TT_PROJECT6
  PIN Tile_X0Y1_UI_IN_TT_PROJECT7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1655.020 0.880 1655.420 ;
    END
  END Tile_X0Y1_UI_IN_TT_PROJECT7
  PIN Tile_X0Y1_UO_OUT_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1576.900 0.880 1577.300 ;
    END
  END Tile_X0Y1_UO_OUT_TT_PROJECT0
  PIN Tile_X0Y1_UO_OUT_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1579.420 0.880 1579.820 ;
    END
  END Tile_X0Y1_UO_OUT_TT_PROJECT1
  PIN Tile_X0Y1_UO_OUT_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1581.940 0.880 1582.340 ;
    END
  END Tile_X0Y1_UO_OUT_TT_PROJECT2
  PIN Tile_X0Y1_UO_OUT_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1584.460 0.880 1584.860 ;
    END
  END Tile_X0Y1_UO_OUT_TT_PROJECT3
  PIN Tile_X0Y1_UO_OUT_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1586.980 0.880 1587.380 ;
    END
  END Tile_X0Y1_UO_OUT_TT_PROJECT4
  PIN Tile_X0Y1_UO_OUT_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1589.500 0.880 1589.900 ;
    END
  END Tile_X0Y1_UO_OUT_TT_PROJECT5
  PIN Tile_X0Y1_UO_OUT_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1592.020 0.880 1592.420 ;
    END
  END Tile_X0Y1_UO_OUT_TT_PROJECT6
  PIN Tile_X0Y1_UO_OUT_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1594.540 0.880 1594.940 ;
    END
  END Tile_X0Y1_UO_OUT_TT_PROJECT7
  PIN Tile_X0Y2_CLK_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1465.180 0.880 1465.580 ;
    END
  END Tile_X0Y2_CLK_TT_PROJECT
  PIN Tile_X0Y2_ENA_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1462.660 0.880 1463.060 ;
    END
  END Tile_X0Y2_ENA_TT_PROJECT
  PIN Tile_X0Y2_RST_N_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.615900 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1467.700 0.860 1468.100 ;
    END
  END Tile_X0Y2_RST_N_TT_PROJECT
  PIN Tile_X0Y2_UIO_IN_TT_PROJECT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1442.500 0.880 1442.900 ;
    END
  END Tile_X0Y2_UIO_IN_TT_PROJECT0
  PIN Tile_X0Y2_UIO_IN_TT_PROJECT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1445.020 0.880 1445.420 ;
    END
  END Tile_X0Y2_UIO_IN_TT_PROJECT1
  PIN Tile_X0Y2_UIO_IN_TT_PROJECT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1447.540 0.880 1447.940 ;
    END
  END Tile_X0Y2_UIO_IN_TT_PROJECT2
  PIN Tile_X0Y2_UIO_IN_TT_PROJECT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1450.060 0.880 1450.460 ;
    END
  END Tile_X0Y2_UIO_IN_TT_PROJECT3
  PIN Tile_X0Y2_UIO_IN_TT_PROJECT4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1452.580 0.880 1452.980 ;
    END
  END Tile_X0Y2_UIO_IN_TT_PROJECT4
  PIN Tile_X0Y2_UIO_IN_TT_PROJECT5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1455.100 0.880 1455.500 ;
    END
  END Tile_X0Y2_UIO_IN_TT_PROJECT5
  PIN Tile_X0Y2_UIO_IN_TT_PROJECT6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1457.620 0.880 1458.020 ;
    END
  END Tile_X0Y2_UIO_IN_TT_PROJECT6
  PIN Tile_X0Y2_UIO_IN_TT_PROJECT7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1460.140 0.880 1460.540 ;
    END
  END Tile_X0Y2_UIO_IN_TT_PROJECT7
  PIN Tile_X0Y2_UIO_OE_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1402.180 0.880 1402.580 ;
    END
  END Tile_X0Y2_UIO_OE_TT_PROJECT0
  PIN Tile_X0Y2_UIO_OE_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1404.700 0.880 1405.100 ;
    END
  END Tile_X0Y2_UIO_OE_TT_PROJECT1
  PIN Tile_X0Y2_UIO_OE_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1407.220 0.880 1407.620 ;
    END
  END Tile_X0Y2_UIO_OE_TT_PROJECT2
  PIN Tile_X0Y2_UIO_OE_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1409.740 0.880 1410.140 ;
    END
  END Tile_X0Y2_UIO_OE_TT_PROJECT3
  PIN Tile_X0Y2_UIO_OE_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1412.260 0.880 1412.660 ;
    END
  END Tile_X0Y2_UIO_OE_TT_PROJECT4
  PIN Tile_X0Y2_UIO_OE_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1414.780 0.880 1415.180 ;
    END
  END Tile_X0Y2_UIO_OE_TT_PROJECT5
  PIN Tile_X0Y2_UIO_OE_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1417.300 0.880 1417.700 ;
    END
  END Tile_X0Y2_UIO_OE_TT_PROJECT6
  PIN Tile_X0Y2_UIO_OE_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1419.820 0.880 1420.220 ;
    END
  END Tile_X0Y2_UIO_OE_TT_PROJECT7
  PIN Tile_X0Y2_UIO_OUT_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1382.020 0.880 1382.420 ;
    END
  END Tile_X0Y2_UIO_OUT_TT_PROJECT0
  PIN Tile_X0Y2_UIO_OUT_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1384.540 0.880 1384.940 ;
    END
  END Tile_X0Y2_UIO_OUT_TT_PROJECT1
  PIN Tile_X0Y2_UIO_OUT_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1387.060 0.880 1387.460 ;
    END
  END Tile_X0Y2_UIO_OUT_TT_PROJECT2
  PIN Tile_X0Y2_UIO_OUT_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1389.580 0.880 1389.980 ;
    END
  END Tile_X0Y2_UIO_OUT_TT_PROJECT3
  PIN Tile_X0Y2_UIO_OUT_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1392.100 0.880 1392.500 ;
    END
  END Tile_X0Y2_UIO_OUT_TT_PROJECT4
  PIN Tile_X0Y2_UIO_OUT_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1394.620 0.880 1395.020 ;
    END
  END Tile_X0Y2_UIO_OUT_TT_PROJECT5
  PIN Tile_X0Y2_UIO_OUT_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1397.140 0.880 1397.540 ;
    END
  END Tile_X0Y2_UIO_OUT_TT_PROJECT6
  PIN Tile_X0Y2_UIO_OUT_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1399.660 0.880 1400.060 ;
    END
  END Tile_X0Y2_UIO_OUT_TT_PROJECT7
  PIN Tile_X0Y2_UI_IN_TT_PROJECT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1422.340 0.880 1422.740 ;
    END
  END Tile_X0Y2_UI_IN_TT_PROJECT0
  PIN Tile_X0Y2_UI_IN_TT_PROJECT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1424.860 0.880 1425.260 ;
    END
  END Tile_X0Y2_UI_IN_TT_PROJECT1
  PIN Tile_X0Y2_UI_IN_TT_PROJECT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1427.380 0.880 1427.780 ;
    END
  END Tile_X0Y2_UI_IN_TT_PROJECT2
  PIN Tile_X0Y2_UI_IN_TT_PROJECT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1429.900 0.880 1430.300 ;
    END
  END Tile_X0Y2_UI_IN_TT_PROJECT3
  PIN Tile_X0Y2_UI_IN_TT_PROJECT4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1432.420 0.880 1432.820 ;
    END
  END Tile_X0Y2_UI_IN_TT_PROJECT4
  PIN Tile_X0Y2_UI_IN_TT_PROJECT5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1434.940 0.880 1435.340 ;
    END
  END Tile_X0Y2_UI_IN_TT_PROJECT5
  PIN Tile_X0Y2_UI_IN_TT_PROJECT6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1437.460 0.860 1437.860 ;
    END
  END Tile_X0Y2_UI_IN_TT_PROJECT6
  PIN Tile_X0Y2_UI_IN_TT_PROJECT7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1439.980 0.880 1440.380 ;
    END
  END Tile_X0Y2_UI_IN_TT_PROJECT7
  PIN Tile_X0Y2_UO_OUT_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1361.860 0.880 1362.260 ;
    END
  END Tile_X0Y2_UO_OUT_TT_PROJECT0
  PIN Tile_X0Y2_UO_OUT_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1364.380 0.880 1364.780 ;
    END
  END Tile_X0Y2_UO_OUT_TT_PROJECT1
  PIN Tile_X0Y2_UO_OUT_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1366.900 0.880 1367.300 ;
    END
  END Tile_X0Y2_UO_OUT_TT_PROJECT2
  PIN Tile_X0Y2_UO_OUT_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1369.420 0.880 1369.820 ;
    END
  END Tile_X0Y2_UO_OUT_TT_PROJECT3
  PIN Tile_X0Y2_UO_OUT_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1371.940 0.880 1372.340 ;
    END
  END Tile_X0Y2_UO_OUT_TT_PROJECT4
  PIN Tile_X0Y2_UO_OUT_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1374.460 0.880 1374.860 ;
    END
  END Tile_X0Y2_UO_OUT_TT_PROJECT5
  PIN Tile_X0Y2_UO_OUT_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1376.980 0.880 1377.380 ;
    END
  END Tile_X0Y2_UO_OUT_TT_PROJECT6
  PIN Tile_X0Y2_UO_OUT_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1379.500 0.880 1379.900 ;
    END
  END Tile_X0Y2_UO_OUT_TT_PROJECT7
  PIN Tile_X0Y3_CLK_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1250.140 0.880 1250.540 ;
    END
  END Tile_X0Y3_CLK_TT_PROJECT
  PIN Tile_X0Y3_ENA_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1247.620 0.880 1248.020 ;
    END
  END Tile_X0Y3_ENA_TT_PROJECT
  PIN Tile_X0Y3_RST_N_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.615900 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1252.660 0.860 1253.060 ;
    END
  END Tile_X0Y3_RST_N_TT_PROJECT
  PIN Tile_X0Y3_UIO_IN_TT_PROJECT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1227.460 0.880 1227.860 ;
    END
  END Tile_X0Y3_UIO_IN_TT_PROJECT0
  PIN Tile_X0Y3_UIO_IN_TT_PROJECT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1229.980 0.880 1230.380 ;
    END
  END Tile_X0Y3_UIO_IN_TT_PROJECT1
  PIN Tile_X0Y3_UIO_IN_TT_PROJECT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1232.500 0.880 1232.900 ;
    END
  END Tile_X0Y3_UIO_IN_TT_PROJECT2
  PIN Tile_X0Y3_UIO_IN_TT_PROJECT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1235.020 0.880 1235.420 ;
    END
  END Tile_X0Y3_UIO_IN_TT_PROJECT3
  PIN Tile_X0Y3_UIO_IN_TT_PROJECT4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1237.540 0.880 1237.940 ;
    END
  END Tile_X0Y3_UIO_IN_TT_PROJECT4
  PIN Tile_X0Y3_UIO_IN_TT_PROJECT5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1240.060 0.880 1240.460 ;
    END
  END Tile_X0Y3_UIO_IN_TT_PROJECT5
  PIN Tile_X0Y3_UIO_IN_TT_PROJECT6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1242.580 0.880 1242.980 ;
    END
  END Tile_X0Y3_UIO_IN_TT_PROJECT6
  PIN Tile_X0Y3_UIO_IN_TT_PROJECT7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1245.100 0.880 1245.500 ;
    END
  END Tile_X0Y3_UIO_IN_TT_PROJECT7
  PIN Tile_X0Y3_UIO_OE_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1187.140 0.880 1187.540 ;
    END
  END Tile_X0Y3_UIO_OE_TT_PROJECT0
  PIN Tile_X0Y3_UIO_OE_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1189.660 0.880 1190.060 ;
    END
  END Tile_X0Y3_UIO_OE_TT_PROJECT1
  PIN Tile_X0Y3_UIO_OE_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1192.180 0.880 1192.580 ;
    END
  END Tile_X0Y3_UIO_OE_TT_PROJECT2
  PIN Tile_X0Y3_UIO_OE_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1194.700 0.880 1195.100 ;
    END
  END Tile_X0Y3_UIO_OE_TT_PROJECT3
  PIN Tile_X0Y3_UIO_OE_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1197.220 0.880 1197.620 ;
    END
  END Tile_X0Y3_UIO_OE_TT_PROJECT4
  PIN Tile_X0Y3_UIO_OE_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1199.740 0.880 1200.140 ;
    END
  END Tile_X0Y3_UIO_OE_TT_PROJECT5
  PIN Tile_X0Y3_UIO_OE_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1202.260 0.880 1202.660 ;
    END
  END Tile_X0Y3_UIO_OE_TT_PROJECT6
  PIN Tile_X0Y3_UIO_OE_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1204.780 0.880 1205.180 ;
    END
  END Tile_X0Y3_UIO_OE_TT_PROJECT7
  PIN Tile_X0Y3_UIO_OUT_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1166.980 0.880 1167.380 ;
    END
  END Tile_X0Y3_UIO_OUT_TT_PROJECT0
  PIN Tile_X0Y3_UIO_OUT_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1169.500 0.880 1169.900 ;
    END
  END Tile_X0Y3_UIO_OUT_TT_PROJECT1
  PIN Tile_X0Y3_UIO_OUT_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1172.020 0.880 1172.420 ;
    END
  END Tile_X0Y3_UIO_OUT_TT_PROJECT2
  PIN Tile_X0Y3_UIO_OUT_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1174.540 0.880 1174.940 ;
    END
  END Tile_X0Y3_UIO_OUT_TT_PROJECT3
  PIN Tile_X0Y3_UIO_OUT_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1177.060 0.880 1177.460 ;
    END
  END Tile_X0Y3_UIO_OUT_TT_PROJECT4
  PIN Tile_X0Y3_UIO_OUT_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1179.580 0.880 1179.980 ;
    END
  END Tile_X0Y3_UIO_OUT_TT_PROJECT5
  PIN Tile_X0Y3_UIO_OUT_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1182.100 0.880 1182.500 ;
    END
  END Tile_X0Y3_UIO_OUT_TT_PROJECT6
  PIN Tile_X0Y3_UIO_OUT_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1184.620 0.880 1185.020 ;
    END
  END Tile_X0Y3_UIO_OUT_TT_PROJECT7
  PIN Tile_X0Y3_UI_IN_TT_PROJECT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1207.300 0.880 1207.700 ;
    END
  END Tile_X0Y3_UI_IN_TT_PROJECT0
  PIN Tile_X0Y3_UI_IN_TT_PROJECT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1209.820 0.880 1210.220 ;
    END
  END Tile_X0Y3_UI_IN_TT_PROJECT1
  PIN Tile_X0Y3_UI_IN_TT_PROJECT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1212.340 0.880 1212.740 ;
    END
  END Tile_X0Y3_UI_IN_TT_PROJECT2
  PIN Tile_X0Y3_UI_IN_TT_PROJECT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1214.860 0.880 1215.260 ;
    END
  END Tile_X0Y3_UI_IN_TT_PROJECT3
  PIN Tile_X0Y3_UI_IN_TT_PROJECT4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1217.380 0.880 1217.780 ;
    END
  END Tile_X0Y3_UI_IN_TT_PROJECT4
  PIN Tile_X0Y3_UI_IN_TT_PROJECT5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1219.900 0.880 1220.300 ;
    END
  END Tile_X0Y3_UI_IN_TT_PROJECT5
  PIN Tile_X0Y3_UI_IN_TT_PROJECT6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1222.420 0.860 1222.820 ;
    END
  END Tile_X0Y3_UI_IN_TT_PROJECT6
  PIN Tile_X0Y3_UI_IN_TT_PROJECT7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1224.940 0.880 1225.340 ;
    END
  END Tile_X0Y3_UI_IN_TT_PROJECT7
  PIN Tile_X0Y3_UO_OUT_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1146.820 0.880 1147.220 ;
    END
  END Tile_X0Y3_UO_OUT_TT_PROJECT0
  PIN Tile_X0Y3_UO_OUT_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1149.340 0.880 1149.740 ;
    END
  END Tile_X0Y3_UO_OUT_TT_PROJECT1
  PIN Tile_X0Y3_UO_OUT_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1151.860 0.880 1152.260 ;
    END
  END Tile_X0Y3_UO_OUT_TT_PROJECT2
  PIN Tile_X0Y3_UO_OUT_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1154.380 0.880 1154.780 ;
    END
  END Tile_X0Y3_UO_OUT_TT_PROJECT3
  PIN Tile_X0Y3_UO_OUT_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1156.900 0.880 1157.300 ;
    END
  END Tile_X0Y3_UO_OUT_TT_PROJECT4
  PIN Tile_X0Y3_UO_OUT_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1159.420 0.880 1159.820 ;
    END
  END Tile_X0Y3_UO_OUT_TT_PROJECT5
  PIN Tile_X0Y3_UO_OUT_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1161.940 0.880 1162.340 ;
    END
  END Tile_X0Y3_UO_OUT_TT_PROJECT6
  PIN Tile_X0Y3_UO_OUT_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1164.460 0.880 1164.860 ;
    END
  END Tile_X0Y3_UO_OUT_TT_PROJECT7
  PIN Tile_X0Y4_CLK_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1035.100 0.880 1035.500 ;
    END
  END Tile_X0Y4_CLK_TT_PROJECT
  PIN Tile_X0Y4_ENA_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1032.580 0.880 1032.980 ;
    END
  END Tile_X0Y4_ENA_TT_PROJECT
  PIN Tile_X0Y4_RST_N_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.615900 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1037.620 0.860 1038.020 ;
    END
  END Tile_X0Y4_RST_N_TT_PROJECT
  PIN Tile_X0Y4_UIO_IN_TT_PROJECT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1012.420 0.880 1012.820 ;
    END
  END Tile_X0Y4_UIO_IN_TT_PROJECT0
  PIN Tile_X0Y4_UIO_IN_TT_PROJECT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1014.940 0.880 1015.340 ;
    END
  END Tile_X0Y4_UIO_IN_TT_PROJECT1
  PIN Tile_X0Y4_UIO_IN_TT_PROJECT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1017.460 0.880 1017.860 ;
    END
  END Tile_X0Y4_UIO_IN_TT_PROJECT2
  PIN Tile_X0Y4_UIO_IN_TT_PROJECT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1019.980 0.880 1020.380 ;
    END
  END Tile_X0Y4_UIO_IN_TT_PROJECT3
  PIN Tile_X0Y4_UIO_IN_TT_PROJECT4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1022.500 0.880 1022.900 ;
    END
  END Tile_X0Y4_UIO_IN_TT_PROJECT4
  PIN Tile_X0Y4_UIO_IN_TT_PROJECT5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1025.020 0.880 1025.420 ;
    END
  END Tile_X0Y4_UIO_IN_TT_PROJECT5
  PIN Tile_X0Y4_UIO_IN_TT_PROJECT6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1027.540 0.880 1027.940 ;
    END
  END Tile_X0Y4_UIO_IN_TT_PROJECT6
  PIN Tile_X0Y4_UIO_IN_TT_PROJECT7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1030.060 0.880 1030.460 ;
    END
  END Tile_X0Y4_UIO_IN_TT_PROJECT7
  PIN Tile_X0Y4_UIO_OE_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 972.100 0.880 972.500 ;
    END
  END Tile_X0Y4_UIO_OE_TT_PROJECT0
  PIN Tile_X0Y4_UIO_OE_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 974.620 0.880 975.020 ;
    END
  END Tile_X0Y4_UIO_OE_TT_PROJECT1
  PIN Tile_X0Y4_UIO_OE_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 977.140 0.880 977.540 ;
    END
  END Tile_X0Y4_UIO_OE_TT_PROJECT2
  PIN Tile_X0Y4_UIO_OE_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 979.660 0.880 980.060 ;
    END
  END Tile_X0Y4_UIO_OE_TT_PROJECT3
  PIN Tile_X0Y4_UIO_OE_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 982.180 0.880 982.580 ;
    END
  END Tile_X0Y4_UIO_OE_TT_PROJECT4
  PIN Tile_X0Y4_UIO_OE_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 984.700 0.880 985.100 ;
    END
  END Tile_X0Y4_UIO_OE_TT_PROJECT5
  PIN Tile_X0Y4_UIO_OE_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 987.220 0.880 987.620 ;
    END
  END Tile_X0Y4_UIO_OE_TT_PROJECT6
  PIN Tile_X0Y4_UIO_OE_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 989.740 0.880 990.140 ;
    END
  END Tile_X0Y4_UIO_OE_TT_PROJECT7
  PIN Tile_X0Y4_UIO_OUT_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 951.940 0.880 952.340 ;
    END
  END Tile_X0Y4_UIO_OUT_TT_PROJECT0
  PIN Tile_X0Y4_UIO_OUT_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 954.460 0.880 954.860 ;
    END
  END Tile_X0Y4_UIO_OUT_TT_PROJECT1
  PIN Tile_X0Y4_UIO_OUT_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 956.980 0.880 957.380 ;
    END
  END Tile_X0Y4_UIO_OUT_TT_PROJECT2
  PIN Tile_X0Y4_UIO_OUT_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 959.500 0.880 959.900 ;
    END
  END Tile_X0Y4_UIO_OUT_TT_PROJECT3
  PIN Tile_X0Y4_UIO_OUT_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 962.020 0.880 962.420 ;
    END
  END Tile_X0Y4_UIO_OUT_TT_PROJECT4
  PIN Tile_X0Y4_UIO_OUT_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 964.540 0.880 964.940 ;
    END
  END Tile_X0Y4_UIO_OUT_TT_PROJECT5
  PIN Tile_X0Y4_UIO_OUT_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 967.060 0.880 967.460 ;
    END
  END Tile_X0Y4_UIO_OUT_TT_PROJECT6
  PIN Tile_X0Y4_UIO_OUT_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 969.580 0.880 969.980 ;
    END
  END Tile_X0Y4_UIO_OUT_TT_PROJECT7
  PIN Tile_X0Y4_UI_IN_TT_PROJECT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 992.260 0.880 992.660 ;
    END
  END Tile_X0Y4_UI_IN_TT_PROJECT0
  PIN Tile_X0Y4_UI_IN_TT_PROJECT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 994.780 0.880 995.180 ;
    END
  END Tile_X0Y4_UI_IN_TT_PROJECT1
  PIN Tile_X0Y4_UI_IN_TT_PROJECT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 997.300 0.880 997.700 ;
    END
  END Tile_X0Y4_UI_IN_TT_PROJECT2
  PIN Tile_X0Y4_UI_IN_TT_PROJECT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 999.820 0.880 1000.220 ;
    END
  END Tile_X0Y4_UI_IN_TT_PROJECT3
  PIN Tile_X0Y4_UI_IN_TT_PROJECT4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1002.340 0.880 1002.740 ;
    END
  END Tile_X0Y4_UI_IN_TT_PROJECT4
  PIN Tile_X0Y4_UI_IN_TT_PROJECT5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1004.860 0.880 1005.260 ;
    END
  END Tile_X0Y4_UI_IN_TT_PROJECT5
  PIN Tile_X0Y4_UI_IN_TT_PROJECT6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1007.380 0.860 1007.780 ;
    END
  END Tile_X0Y4_UI_IN_TT_PROJECT6
  PIN Tile_X0Y4_UI_IN_TT_PROJECT7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1009.900 0.880 1010.300 ;
    END
  END Tile_X0Y4_UI_IN_TT_PROJECT7
  PIN Tile_X0Y4_UO_OUT_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 931.780 0.880 932.180 ;
    END
  END Tile_X0Y4_UO_OUT_TT_PROJECT0
  PIN Tile_X0Y4_UO_OUT_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 934.300 0.880 934.700 ;
    END
  END Tile_X0Y4_UO_OUT_TT_PROJECT1
  PIN Tile_X0Y4_UO_OUT_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 936.820 0.880 937.220 ;
    END
  END Tile_X0Y4_UO_OUT_TT_PROJECT2
  PIN Tile_X0Y4_UO_OUT_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 939.340 0.880 939.740 ;
    END
  END Tile_X0Y4_UO_OUT_TT_PROJECT3
  PIN Tile_X0Y4_UO_OUT_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 941.860 0.880 942.260 ;
    END
  END Tile_X0Y4_UO_OUT_TT_PROJECT4
  PIN Tile_X0Y4_UO_OUT_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 944.380 0.880 944.780 ;
    END
  END Tile_X0Y4_UO_OUT_TT_PROJECT5
  PIN Tile_X0Y4_UO_OUT_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 946.900 0.880 947.300 ;
    END
  END Tile_X0Y4_UO_OUT_TT_PROJECT6
  PIN Tile_X0Y4_UO_OUT_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 949.420 0.880 949.820 ;
    END
  END Tile_X0Y4_UO_OUT_TT_PROJECT7
  PIN Tile_X0Y5_CLK_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 820.060 0.880 820.460 ;
    END
  END Tile_X0Y5_CLK_TT_PROJECT
  PIN Tile_X0Y5_ENA_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 817.540 0.880 817.940 ;
    END
  END Tile_X0Y5_ENA_TT_PROJECT
  PIN Tile_X0Y5_RST_N_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.615900 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 822.580 0.860 822.980 ;
    END
  END Tile_X0Y5_RST_N_TT_PROJECT
  PIN Tile_X0Y5_UIO_IN_TT_PROJECT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 797.380 0.880 797.780 ;
    END
  END Tile_X0Y5_UIO_IN_TT_PROJECT0
  PIN Tile_X0Y5_UIO_IN_TT_PROJECT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 799.900 0.880 800.300 ;
    END
  END Tile_X0Y5_UIO_IN_TT_PROJECT1
  PIN Tile_X0Y5_UIO_IN_TT_PROJECT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 802.420 0.880 802.820 ;
    END
  END Tile_X0Y5_UIO_IN_TT_PROJECT2
  PIN Tile_X0Y5_UIO_IN_TT_PROJECT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 804.940 0.880 805.340 ;
    END
  END Tile_X0Y5_UIO_IN_TT_PROJECT3
  PIN Tile_X0Y5_UIO_IN_TT_PROJECT4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 807.460 0.880 807.860 ;
    END
  END Tile_X0Y5_UIO_IN_TT_PROJECT4
  PIN Tile_X0Y5_UIO_IN_TT_PROJECT5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 809.980 0.880 810.380 ;
    END
  END Tile_X0Y5_UIO_IN_TT_PROJECT5
  PIN Tile_X0Y5_UIO_IN_TT_PROJECT6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 812.500 0.880 812.900 ;
    END
  END Tile_X0Y5_UIO_IN_TT_PROJECT6
  PIN Tile_X0Y5_UIO_IN_TT_PROJECT7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 815.020 0.880 815.420 ;
    END
  END Tile_X0Y5_UIO_IN_TT_PROJECT7
  PIN Tile_X0Y5_UIO_OE_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 757.060 0.880 757.460 ;
    END
  END Tile_X0Y5_UIO_OE_TT_PROJECT0
  PIN Tile_X0Y5_UIO_OE_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 759.580 0.880 759.980 ;
    END
  END Tile_X0Y5_UIO_OE_TT_PROJECT1
  PIN Tile_X0Y5_UIO_OE_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 762.100 0.880 762.500 ;
    END
  END Tile_X0Y5_UIO_OE_TT_PROJECT2
  PIN Tile_X0Y5_UIO_OE_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 764.620 0.880 765.020 ;
    END
  END Tile_X0Y5_UIO_OE_TT_PROJECT3
  PIN Tile_X0Y5_UIO_OE_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 767.140 0.880 767.540 ;
    END
  END Tile_X0Y5_UIO_OE_TT_PROJECT4
  PIN Tile_X0Y5_UIO_OE_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 769.660 0.880 770.060 ;
    END
  END Tile_X0Y5_UIO_OE_TT_PROJECT5
  PIN Tile_X0Y5_UIO_OE_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 772.180 0.880 772.580 ;
    END
  END Tile_X0Y5_UIO_OE_TT_PROJECT6
  PIN Tile_X0Y5_UIO_OE_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 774.700 0.880 775.100 ;
    END
  END Tile_X0Y5_UIO_OE_TT_PROJECT7
  PIN Tile_X0Y5_UIO_OUT_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 736.900 0.880 737.300 ;
    END
  END Tile_X0Y5_UIO_OUT_TT_PROJECT0
  PIN Tile_X0Y5_UIO_OUT_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 739.420 0.880 739.820 ;
    END
  END Tile_X0Y5_UIO_OUT_TT_PROJECT1
  PIN Tile_X0Y5_UIO_OUT_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 741.940 0.880 742.340 ;
    END
  END Tile_X0Y5_UIO_OUT_TT_PROJECT2
  PIN Tile_X0Y5_UIO_OUT_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 744.460 0.880 744.860 ;
    END
  END Tile_X0Y5_UIO_OUT_TT_PROJECT3
  PIN Tile_X0Y5_UIO_OUT_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 746.980 0.880 747.380 ;
    END
  END Tile_X0Y5_UIO_OUT_TT_PROJECT4
  PIN Tile_X0Y5_UIO_OUT_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 749.500 0.880 749.900 ;
    END
  END Tile_X0Y5_UIO_OUT_TT_PROJECT5
  PIN Tile_X0Y5_UIO_OUT_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 752.020 0.880 752.420 ;
    END
  END Tile_X0Y5_UIO_OUT_TT_PROJECT6
  PIN Tile_X0Y5_UIO_OUT_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 754.540 0.880 754.940 ;
    END
  END Tile_X0Y5_UIO_OUT_TT_PROJECT7
  PIN Tile_X0Y5_UI_IN_TT_PROJECT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 777.220 0.880 777.620 ;
    END
  END Tile_X0Y5_UI_IN_TT_PROJECT0
  PIN Tile_X0Y5_UI_IN_TT_PROJECT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 779.740 0.880 780.140 ;
    END
  END Tile_X0Y5_UI_IN_TT_PROJECT1
  PIN Tile_X0Y5_UI_IN_TT_PROJECT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 782.260 0.880 782.660 ;
    END
  END Tile_X0Y5_UI_IN_TT_PROJECT2
  PIN Tile_X0Y5_UI_IN_TT_PROJECT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 784.780 0.880 785.180 ;
    END
  END Tile_X0Y5_UI_IN_TT_PROJECT3
  PIN Tile_X0Y5_UI_IN_TT_PROJECT4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 787.300 0.880 787.700 ;
    END
  END Tile_X0Y5_UI_IN_TT_PROJECT4
  PIN Tile_X0Y5_UI_IN_TT_PROJECT5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 789.820 0.880 790.220 ;
    END
  END Tile_X0Y5_UI_IN_TT_PROJECT5
  PIN Tile_X0Y5_UI_IN_TT_PROJECT6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 792.340 0.860 792.740 ;
    END
  END Tile_X0Y5_UI_IN_TT_PROJECT6
  PIN Tile_X0Y5_UI_IN_TT_PROJECT7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 794.860 0.880 795.260 ;
    END
  END Tile_X0Y5_UI_IN_TT_PROJECT7
  PIN Tile_X0Y5_UO_OUT_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 716.740 0.880 717.140 ;
    END
  END Tile_X0Y5_UO_OUT_TT_PROJECT0
  PIN Tile_X0Y5_UO_OUT_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 719.260 0.880 719.660 ;
    END
  END Tile_X0Y5_UO_OUT_TT_PROJECT1
  PIN Tile_X0Y5_UO_OUT_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 721.780 0.880 722.180 ;
    END
  END Tile_X0Y5_UO_OUT_TT_PROJECT2
  PIN Tile_X0Y5_UO_OUT_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 724.300 0.880 724.700 ;
    END
  END Tile_X0Y5_UO_OUT_TT_PROJECT3
  PIN Tile_X0Y5_UO_OUT_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 726.820 0.880 727.220 ;
    END
  END Tile_X0Y5_UO_OUT_TT_PROJECT4
  PIN Tile_X0Y5_UO_OUT_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 729.340 0.880 729.740 ;
    END
  END Tile_X0Y5_UO_OUT_TT_PROJECT5
  PIN Tile_X0Y5_UO_OUT_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 731.860 0.880 732.260 ;
    END
  END Tile_X0Y5_UO_OUT_TT_PROJECT6
  PIN Tile_X0Y5_UO_OUT_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 734.380 0.880 734.780 ;
    END
  END Tile_X0Y5_UO_OUT_TT_PROJECT7
  PIN Tile_X0Y6_CLK_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 605.020 0.880 605.420 ;
    END
  END Tile_X0Y6_CLK_TT_PROJECT
  PIN Tile_X0Y6_ENA_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 602.500 0.880 602.900 ;
    END
  END Tile_X0Y6_ENA_TT_PROJECT
  PIN Tile_X0Y6_RST_N_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.615900 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 607.540 0.860 607.940 ;
    END
  END Tile_X0Y6_RST_N_TT_PROJECT
  PIN Tile_X0Y6_UIO_IN_TT_PROJECT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 582.340 0.880 582.740 ;
    END
  END Tile_X0Y6_UIO_IN_TT_PROJECT0
  PIN Tile_X0Y6_UIO_IN_TT_PROJECT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 584.860 0.880 585.260 ;
    END
  END Tile_X0Y6_UIO_IN_TT_PROJECT1
  PIN Tile_X0Y6_UIO_IN_TT_PROJECT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 587.380 0.880 587.780 ;
    END
  END Tile_X0Y6_UIO_IN_TT_PROJECT2
  PIN Tile_X0Y6_UIO_IN_TT_PROJECT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 589.900 0.880 590.300 ;
    END
  END Tile_X0Y6_UIO_IN_TT_PROJECT3
  PIN Tile_X0Y6_UIO_IN_TT_PROJECT4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 592.420 0.880 592.820 ;
    END
  END Tile_X0Y6_UIO_IN_TT_PROJECT4
  PIN Tile_X0Y6_UIO_IN_TT_PROJECT5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 594.940 0.880 595.340 ;
    END
  END Tile_X0Y6_UIO_IN_TT_PROJECT5
  PIN Tile_X0Y6_UIO_IN_TT_PROJECT6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 597.460 0.880 597.860 ;
    END
  END Tile_X0Y6_UIO_IN_TT_PROJECT6
  PIN Tile_X0Y6_UIO_IN_TT_PROJECT7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 599.980 0.880 600.380 ;
    END
  END Tile_X0Y6_UIO_IN_TT_PROJECT7
  PIN Tile_X0Y6_UIO_OE_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 542.020 0.880 542.420 ;
    END
  END Tile_X0Y6_UIO_OE_TT_PROJECT0
  PIN Tile_X0Y6_UIO_OE_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 544.540 0.880 544.940 ;
    END
  END Tile_X0Y6_UIO_OE_TT_PROJECT1
  PIN Tile_X0Y6_UIO_OE_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 547.060 0.880 547.460 ;
    END
  END Tile_X0Y6_UIO_OE_TT_PROJECT2
  PIN Tile_X0Y6_UIO_OE_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 549.580 0.880 549.980 ;
    END
  END Tile_X0Y6_UIO_OE_TT_PROJECT3
  PIN Tile_X0Y6_UIO_OE_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 552.100 0.880 552.500 ;
    END
  END Tile_X0Y6_UIO_OE_TT_PROJECT4
  PIN Tile_X0Y6_UIO_OE_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 554.620 0.880 555.020 ;
    END
  END Tile_X0Y6_UIO_OE_TT_PROJECT5
  PIN Tile_X0Y6_UIO_OE_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 557.140 0.880 557.540 ;
    END
  END Tile_X0Y6_UIO_OE_TT_PROJECT6
  PIN Tile_X0Y6_UIO_OE_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 559.660 0.880 560.060 ;
    END
  END Tile_X0Y6_UIO_OE_TT_PROJECT7
  PIN Tile_X0Y6_UIO_OUT_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 521.860 0.880 522.260 ;
    END
  END Tile_X0Y6_UIO_OUT_TT_PROJECT0
  PIN Tile_X0Y6_UIO_OUT_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 524.380 0.880 524.780 ;
    END
  END Tile_X0Y6_UIO_OUT_TT_PROJECT1
  PIN Tile_X0Y6_UIO_OUT_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 526.900 0.880 527.300 ;
    END
  END Tile_X0Y6_UIO_OUT_TT_PROJECT2
  PIN Tile_X0Y6_UIO_OUT_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 529.420 0.880 529.820 ;
    END
  END Tile_X0Y6_UIO_OUT_TT_PROJECT3
  PIN Tile_X0Y6_UIO_OUT_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 531.940 0.880 532.340 ;
    END
  END Tile_X0Y6_UIO_OUT_TT_PROJECT4
  PIN Tile_X0Y6_UIO_OUT_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 534.460 0.880 534.860 ;
    END
  END Tile_X0Y6_UIO_OUT_TT_PROJECT5
  PIN Tile_X0Y6_UIO_OUT_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 536.980 0.880 537.380 ;
    END
  END Tile_X0Y6_UIO_OUT_TT_PROJECT6
  PIN Tile_X0Y6_UIO_OUT_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 539.500 0.880 539.900 ;
    END
  END Tile_X0Y6_UIO_OUT_TT_PROJECT7
  PIN Tile_X0Y6_UI_IN_TT_PROJECT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 562.180 0.880 562.580 ;
    END
  END Tile_X0Y6_UI_IN_TT_PROJECT0
  PIN Tile_X0Y6_UI_IN_TT_PROJECT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 564.700 0.880 565.100 ;
    END
  END Tile_X0Y6_UI_IN_TT_PROJECT1
  PIN Tile_X0Y6_UI_IN_TT_PROJECT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 567.220 0.880 567.620 ;
    END
  END Tile_X0Y6_UI_IN_TT_PROJECT2
  PIN Tile_X0Y6_UI_IN_TT_PROJECT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 569.740 0.880 570.140 ;
    END
  END Tile_X0Y6_UI_IN_TT_PROJECT3
  PIN Tile_X0Y6_UI_IN_TT_PROJECT4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 572.260 0.880 572.660 ;
    END
  END Tile_X0Y6_UI_IN_TT_PROJECT4
  PIN Tile_X0Y6_UI_IN_TT_PROJECT5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 574.780 0.880 575.180 ;
    END
  END Tile_X0Y6_UI_IN_TT_PROJECT5
  PIN Tile_X0Y6_UI_IN_TT_PROJECT6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 577.300 0.860 577.700 ;
    END
  END Tile_X0Y6_UI_IN_TT_PROJECT6
  PIN Tile_X0Y6_UI_IN_TT_PROJECT7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 579.820 0.880 580.220 ;
    END
  END Tile_X0Y6_UI_IN_TT_PROJECT7
  PIN Tile_X0Y6_UO_OUT_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 501.700 0.880 502.100 ;
    END
  END Tile_X0Y6_UO_OUT_TT_PROJECT0
  PIN Tile_X0Y6_UO_OUT_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 504.220 0.880 504.620 ;
    END
  END Tile_X0Y6_UO_OUT_TT_PROJECT1
  PIN Tile_X0Y6_UO_OUT_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 506.740 0.880 507.140 ;
    END
  END Tile_X0Y6_UO_OUT_TT_PROJECT2
  PIN Tile_X0Y6_UO_OUT_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 509.260 0.880 509.660 ;
    END
  END Tile_X0Y6_UO_OUT_TT_PROJECT3
  PIN Tile_X0Y6_UO_OUT_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 511.780 0.880 512.180 ;
    END
  END Tile_X0Y6_UO_OUT_TT_PROJECT4
  PIN Tile_X0Y6_UO_OUT_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 514.300 0.880 514.700 ;
    END
  END Tile_X0Y6_UO_OUT_TT_PROJECT5
  PIN Tile_X0Y6_UO_OUT_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 516.820 0.880 517.220 ;
    END
  END Tile_X0Y6_UO_OUT_TT_PROJECT6
  PIN Tile_X0Y6_UO_OUT_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 519.340 0.880 519.740 ;
    END
  END Tile_X0Y6_UO_OUT_TT_PROJECT7
  PIN Tile_X0Y7_CLK_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 389.980 0.880 390.380 ;
    END
  END Tile_X0Y7_CLK_TT_PROJECT
  PIN Tile_X0Y7_ENA_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 387.460 0.880 387.860 ;
    END
  END Tile_X0Y7_ENA_TT_PROJECT
  PIN Tile_X0Y7_RST_N_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.615900 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 392.500 0.860 392.900 ;
    END
  END Tile_X0Y7_RST_N_TT_PROJECT
  PIN Tile_X0Y7_UIO_IN_TT_PROJECT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 367.300 0.880 367.700 ;
    END
  END Tile_X0Y7_UIO_IN_TT_PROJECT0
  PIN Tile_X0Y7_UIO_IN_TT_PROJECT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 369.820 0.880 370.220 ;
    END
  END Tile_X0Y7_UIO_IN_TT_PROJECT1
  PIN Tile_X0Y7_UIO_IN_TT_PROJECT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 372.340 0.880 372.740 ;
    END
  END Tile_X0Y7_UIO_IN_TT_PROJECT2
  PIN Tile_X0Y7_UIO_IN_TT_PROJECT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 374.860 0.880 375.260 ;
    END
  END Tile_X0Y7_UIO_IN_TT_PROJECT3
  PIN Tile_X0Y7_UIO_IN_TT_PROJECT4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 377.380 0.880 377.780 ;
    END
  END Tile_X0Y7_UIO_IN_TT_PROJECT4
  PIN Tile_X0Y7_UIO_IN_TT_PROJECT5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 379.900 0.880 380.300 ;
    END
  END Tile_X0Y7_UIO_IN_TT_PROJECT5
  PIN Tile_X0Y7_UIO_IN_TT_PROJECT6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 382.420 0.880 382.820 ;
    END
  END Tile_X0Y7_UIO_IN_TT_PROJECT6
  PIN Tile_X0Y7_UIO_IN_TT_PROJECT7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 384.940 0.880 385.340 ;
    END
  END Tile_X0Y7_UIO_IN_TT_PROJECT7
  PIN Tile_X0Y7_UIO_OE_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 326.980 0.880 327.380 ;
    END
  END Tile_X0Y7_UIO_OE_TT_PROJECT0
  PIN Tile_X0Y7_UIO_OE_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 329.500 0.880 329.900 ;
    END
  END Tile_X0Y7_UIO_OE_TT_PROJECT1
  PIN Tile_X0Y7_UIO_OE_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 332.020 0.880 332.420 ;
    END
  END Tile_X0Y7_UIO_OE_TT_PROJECT2
  PIN Tile_X0Y7_UIO_OE_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 334.540 0.880 334.940 ;
    END
  END Tile_X0Y7_UIO_OE_TT_PROJECT3
  PIN Tile_X0Y7_UIO_OE_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 337.060 0.880 337.460 ;
    END
  END Tile_X0Y7_UIO_OE_TT_PROJECT4
  PIN Tile_X0Y7_UIO_OE_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 339.580 0.880 339.980 ;
    END
  END Tile_X0Y7_UIO_OE_TT_PROJECT5
  PIN Tile_X0Y7_UIO_OE_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 342.100 0.880 342.500 ;
    END
  END Tile_X0Y7_UIO_OE_TT_PROJECT6
  PIN Tile_X0Y7_UIO_OE_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 344.620 0.880 345.020 ;
    END
  END Tile_X0Y7_UIO_OE_TT_PROJECT7
  PIN Tile_X0Y7_UIO_OUT_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 306.820 0.880 307.220 ;
    END
  END Tile_X0Y7_UIO_OUT_TT_PROJECT0
  PIN Tile_X0Y7_UIO_OUT_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 309.340 0.880 309.740 ;
    END
  END Tile_X0Y7_UIO_OUT_TT_PROJECT1
  PIN Tile_X0Y7_UIO_OUT_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 311.860 0.880 312.260 ;
    END
  END Tile_X0Y7_UIO_OUT_TT_PROJECT2
  PIN Tile_X0Y7_UIO_OUT_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 314.380 0.880 314.780 ;
    END
  END Tile_X0Y7_UIO_OUT_TT_PROJECT3
  PIN Tile_X0Y7_UIO_OUT_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 316.900 0.880 317.300 ;
    END
  END Tile_X0Y7_UIO_OUT_TT_PROJECT4
  PIN Tile_X0Y7_UIO_OUT_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 319.420 0.880 319.820 ;
    END
  END Tile_X0Y7_UIO_OUT_TT_PROJECT5
  PIN Tile_X0Y7_UIO_OUT_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 321.940 0.880 322.340 ;
    END
  END Tile_X0Y7_UIO_OUT_TT_PROJECT6
  PIN Tile_X0Y7_UIO_OUT_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 324.460 0.880 324.860 ;
    END
  END Tile_X0Y7_UIO_OUT_TT_PROJECT7
  PIN Tile_X0Y7_UI_IN_TT_PROJECT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 347.140 0.880 347.540 ;
    END
  END Tile_X0Y7_UI_IN_TT_PROJECT0
  PIN Tile_X0Y7_UI_IN_TT_PROJECT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 349.660 0.880 350.060 ;
    END
  END Tile_X0Y7_UI_IN_TT_PROJECT1
  PIN Tile_X0Y7_UI_IN_TT_PROJECT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 352.180 0.880 352.580 ;
    END
  END Tile_X0Y7_UI_IN_TT_PROJECT2
  PIN Tile_X0Y7_UI_IN_TT_PROJECT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 354.700 0.880 355.100 ;
    END
  END Tile_X0Y7_UI_IN_TT_PROJECT3
  PIN Tile_X0Y7_UI_IN_TT_PROJECT4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 357.220 0.880 357.620 ;
    END
  END Tile_X0Y7_UI_IN_TT_PROJECT4
  PIN Tile_X0Y7_UI_IN_TT_PROJECT5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 359.740 0.880 360.140 ;
    END
  END Tile_X0Y7_UI_IN_TT_PROJECT5
  PIN Tile_X0Y7_UI_IN_TT_PROJECT6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 362.260 0.860 362.660 ;
    END
  END Tile_X0Y7_UI_IN_TT_PROJECT6
  PIN Tile_X0Y7_UI_IN_TT_PROJECT7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 364.780 0.880 365.180 ;
    END
  END Tile_X0Y7_UI_IN_TT_PROJECT7
  PIN Tile_X0Y7_UO_OUT_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 286.660 0.880 287.060 ;
    END
  END Tile_X0Y7_UO_OUT_TT_PROJECT0
  PIN Tile_X0Y7_UO_OUT_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 289.180 0.880 289.580 ;
    END
  END Tile_X0Y7_UO_OUT_TT_PROJECT1
  PIN Tile_X0Y7_UO_OUT_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 291.700 0.880 292.100 ;
    END
  END Tile_X0Y7_UO_OUT_TT_PROJECT2
  PIN Tile_X0Y7_UO_OUT_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 294.220 0.880 294.620 ;
    END
  END Tile_X0Y7_UO_OUT_TT_PROJECT3
  PIN Tile_X0Y7_UO_OUT_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 296.740 0.880 297.140 ;
    END
  END Tile_X0Y7_UO_OUT_TT_PROJECT4
  PIN Tile_X0Y7_UO_OUT_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 299.260 0.880 299.660 ;
    END
  END Tile_X0Y7_UO_OUT_TT_PROJECT5
  PIN Tile_X0Y7_UO_OUT_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 301.780 0.880 302.180 ;
    END
  END Tile_X0Y7_UO_OUT_TT_PROJECT6
  PIN Tile_X0Y7_UO_OUT_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 304.300 0.880 304.700 ;
    END
  END Tile_X0Y7_UO_OUT_TT_PROJECT7
  PIN Tile_X0Y8_CLK_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 174.940 0.880 175.340 ;
    END
  END Tile_X0Y8_CLK_TT_PROJECT
  PIN Tile_X0Y8_ENA_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 172.420 0.880 172.820 ;
    END
  END Tile_X0Y8_ENA_TT_PROJECT
  PIN Tile_X0Y8_RST_N_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.615900 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 177.460 0.860 177.860 ;
    END
  END Tile_X0Y8_RST_N_TT_PROJECT
  PIN Tile_X0Y8_UIO_IN_TT_PROJECT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 152.260 0.880 152.660 ;
    END
  END Tile_X0Y8_UIO_IN_TT_PROJECT0
  PIN Tile_X0Y8_UIO_IN_TT_PROJECT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 154.780 0.880 155.180 ;
    END
  END Tile_X0Y8_UIO_IN_TT_PROJECT1
  PIN Tile_X0Y8_UIO_IN_TT_PROJECT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 157.300 0.880 157.700 ;
    END
  END Tile_X0Y8_UIO_IN_TT_PROJECT2
  PIN Tile_X0Y8_UIO_IN_TT_PROJECT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 159.820 0.880 160.220 ;
    END
  END Tile_X0Y8_UIO_IN_TT_PROJECT3
  PIN Tile_X0Y8_UIO_IN_TT_PROJECT4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 162.340 0.880 162.740 ;
    END
  END Tile_X0Y8_UIO_IN_TT_PROJECT4
  PIN Tile_X0Y8_UIO_IN_TT_PROJECT5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 164.860 0.880 165.260 ;
    END
  END Tile_X0Y8_UIO_IN_TT_PROJECT5
  PIN Tile_X0Y8_UIO_IN_TT_PROJECT6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 167.380 0.880 167.780 ;
    END
  END Tile_X0Y8_UIO_IN_TT_PROJECT6
  PIN Tile_X0Y8_UIO_IN_TT_PROJECT7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 169.900 0.880 170.300 ;
    END
  END Tile_X0Y8_UIO_IN_TT_PROJECT7
  PIN Tile_X0Y8_UIO_OE_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 111.940 0.880 112.340 ;
    END
  END Tile_X0Y8_UIO_OE_TT_PROJECT0
  PIN Tile_X0Y8_UIO_OE_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 114.460 0.880 114.860 ;
    END
  END Tile_X0Y8_UIO_OE_TT_PROJECT1
  PIN Tile_X0Y8_UIO_OE_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 116.980 0.880 117.380 ;
    END
  END Tile_X0Y8_UIO_OE_TT_PROJECT2
  PIN Tile_X0Y8_UIO_OE_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 119.500 0.880 119.900 ;
    END
  END Tile_X0Y8_UIO_OE_TT_PROJECT3
  PIN Tile_X0Y8_UIO_OE_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 122.020 0.880 122.420 ;
    END
  END Tile_X0Y8_UIO_OE_TT_PROJECT4
  PIN Tile_X0Y8_UIO_OE_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 124.540 0.880 124.940 ;
    END
  END Tile_X0Y8_UIO_OE_TT_PROJECT5
  PIN Tile_X0Y8_UIO_OE_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 127.060 0.880 127.460 ;
    END
  END Tile_X0Y8_UIO_OE_TT_PROJECT6
  PIN Tile_X0Y8_UIO_OE_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 129.580 0.880 129.980 ;
    END
  END Tile_X0Y8_UIO_OE_TT_PROJECT7
  PIN Tile_X0Y8_UIO_OUT_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 91.780 0.880 92.180 ;
    END
  END Tile_X0Y8_UIO_OUT_TT_PROJECT0
  PIN Tile_X0Y8_UIO_OUT_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 94.300 0.880 94.700 ;
    END
  END Tile_X0Y8_UIO_OUT_TT_PROJECT1
  PIN Tile_X0Y8_UIO_OUT_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 96.820 0.880 97.220 ;
    END
  END Tile_X0Y8_UIO_OUT_TT_PROJECT2
  PIN Tile_X0Y8_UIO_OUT_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 99.340 0.880 99.740 ;
    END
  END Tile_X0Y8_UIO_OUT_TT_PROJECT3
  PIN Tile_X0Y8_UIO_OUT_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 101.860 0.880 102.260 ;
    END
  END Tile_X0Y8_UIO_OUT_TT_PROJECT4
  PIN Tile_X0Y8_UIO_OUT_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 104.380 0.880 104.780 ;
    END
  END Tile_X0Y8_UIO_OUT_TT_PROJECT5
  PIN Tile_X0Y8_UIO_OUT_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 106.900 0.880 107.300 ;
    END
  END Tile_X0Y8_UIO_OUT_TT_PROJECT6
  PIN Tile_X0Y8_UIO_OUT_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 109.420 0.880 109.820 ;
    END
  END Tile_X0Y8_UIO_OUT_TT_PROJECT7
  PIN Tile_X0Y8_UI_IN_TT_PROJECT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 132.100 0.880 132.500 ;
    END
  END Tile_X0Y8_UI_IN_TT_PROJECT0
  PIN Tile_X0Y8_UI_IN_TT_PROJECT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 134.620 0.880 135.020 ;
    END
  END Tile_X0Y8_UI_IN_TT_PROJECT1
  PIN Tile_X0Y8_UI_IN_TT_PROJECT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 137.140 0.880 137.540 ;
    END
  END Tile_X0Y8_UI_IN_TT_PROJECT2
  PIN Tile_X0Y8_UI_IN_TT_PROJECT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 139.660 0.880 140.060 ;
    END
  END Tile_X0Y8_UI_IN_TT_PROJECT3
  PIN Tile_X0Y8_UI_IN_TT_PROJECT4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 142.180 0.880 142.580 ;
    END
  END Tile_X0Y8_UI_IN_TT_PROJECT4
  PIN Tile_X0Y8_UI_IN_TT_PROJECT5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 144.700 0.880 145.100 ;
    END
  END Tile_X0Y8_UI_IN_TT_PROJECT5
  PIN Tile_X0Y8_UI_IN_TT_PROJECT6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 147.220 0.860 147.620 ;
    END
  END Tile_X0Y8_UI_IN_TT_PROJECT6
  PIN Tile_X0Y8_UI_IN_TT_PROJECT7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 149.740 0.880 150.140 ;
    END
  END Tile_X0Y8_UI_IN_TT_PROJECT7
  PIN Tile_X0Y8_UO_OUT_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 71.620 0.880 72.020 ;
    END
  END Tile_X0Y8_UO_OUT_TT_PROJECT0
  PIN Tile_X0Y8_UO_OUT_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 74.140 0.880 74.540 ;
    END
  END Tile_X0Y8_UO_OUT_TT_PROJECT1
  PIN Tile_X0Y8_UO_OUT_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 76.660 0.880 77.060 ;
    END
  END Tile_X0Y8_UO_OUT_TT_PROJECT2
  PIN Tile_X0Y8_UO_OUT_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 79.180 0.880 79.580 ;
    END
  END Tile_X0Y8_UO_OUT_TT_PROJECT3
  PIN Tile_X0Y8_UO_OUT_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 81.700 0.880 82.100 ;
    END
  END Tile_X0Y8_UO_OUT_TT_PROJECT4
  PIN Tile_X0Y8_UO_OUT_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 84.220 0.880 84.620 ;
    END
  END Tile_X0Y8_UO_OUT_TT_PROJECT5
  PIN Tile_X0Y8_UO_OUT_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 86.740 0.880 87.140 ;
    END
  END Tile_X0Y8_UO_OUT_TT_PROJECT6
  PIN Tile_X0Y8_UO_OUT_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 89.260 0.880 89.660 ;
    END
  END Tile_X0Y8_UO_OUT_TT_PROJECT7
  PIN Tile_X1Y0_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 128.440 1831.640 128.840 1832.520 ;
    END
  END Tile_X1Y0_A_I_top
  PIN Tile_X1Y0_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 122.680 1831.640 123.080 1832.520 ;
    END
  END Tile_X1Y0_A_O_top
  PIN Tile_X1Y0_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 134.200 1831.640 134.600 1832.520 ;
    END
  END Tile_X1Y0_A_T_top
  PIN Tile_X1Y0_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 145.720 1831.640 146.120 1832.520 ;
    END
  END Tile_X1Y0_B_I_top
  PIN Tile_X1Y0_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 139.960 1831.640 140.360 1832.520 ;
    END
  END Tile_X1Y0_B_O_top
  PIN Tile_X1Y0_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 151.480 1831.640 151.880 1832.520 ;
    END
  END Tile_X1Y0_B_T_top
  PIN Tile_X1Y0_C_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.615900 ;
    PORT
      LAYER Metal2 ;
        RECT 163.000 1831.640 163.400 1832.520 ;
    END
  END Tile_X1Y0_C_I_top
  PIN Tile_X1Y0_C_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 157.240 1831.640 157.640 1832.520 ;
    END
  END Tile_X1Y0_C_O_top
  PIN Tile_X1Y0_C_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 168.760 1831.640 169.160 1832.520 ;
    END
  END Tile_X1Y0_C_T_top
  PIN Tile_X1Y0_D_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 180.280 1831.640 180.680 1832.520 ;
    END
  END Tile_X1Y0_D_I_top
  PIN Tile_X1Y0_D_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 174.520 1831.640 174.920 1832.520 ;
    END
  END Tile_X1Y0_D_O_top
  PIN Tile_X1Y0_D_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 186.040 1831.640 186.440 1832.520 ;
    END
  END Tile_X1Y0_D_T_top
  PIN Tile_X1Y9_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 128.440 0.000 128.840 0.480 ;
    END
  END Tile_X1Y9_A_I_top
  PIN Tile_X1Y9_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 122.680 0.000 123.080 0.480 ;
    END
  END Tile_X1Y9_A_O_top
  PIN Tile_X1Y9_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 134.200 0.000 134.600 0.480 ;
    END
  END Tile_X1Y9_A_T_top
  PIN Tile_X1Y9_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 145.720 0.000 146.120 0.480 ;
    END
  END Tile_X1Y9_B_I_top
  PIN Tile_X1Y9_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 139.960 0.000 140.360 0.480 ;
    END
  END Tile_X1Y9_B_O_top
  PIN Tile_X1Y9_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 151.480 0.000 151.880 0.480 ;
    END
  END Tile_X1Y9_B_T_top
  PIN Tile_X1Y9_C_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.615900 ;
    PORT
      LAYER Metal2 ;
        RECT 163.000 0.000 163.400 0.480 ;
    END
  END Tile_X1Y9_C_I_top
  PIN Tile_X1Y9_C_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 157.240 0.000 157.640 0.480 ;
    END
  END Tile_X1Y9_C_O_top
  PIN Tile_X1Y9_C_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 168.760 0.000 169.160 0.480 ;
    END
  END Tile_X1Y9_C_T_top
  PIN Tile_X1Y9_D_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 180.280 0.000 180.680 0.480 ;
    END
  END Tile_X1Y9_D_I_top
  PIN Tile_X1Y9_D_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 174.520 0.000 174.920 0.480 ;
    END
  END Tile_X1Y9_D_O_top
  PIN Tile_X1Y9_D_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 186.040 0.000 186.440 0.480 ;
    END
  END Tile_X1Y9_D_T_top
  PIN Tile_X2Y0_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 343.480 1831.640 343.880 1832.520 ;
    END
  END Tile_X2Y0_A_I_top
  PIN Tile_X2Y0_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 337.720 1831.640 338.120 1832.520 ;
    END
  END Tile_X2Y0_A_O_top
  PIN Tile_X2Y0_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 349.240 1831.640 349.640 1832.520 ;
    END
  END Tile_X2Y0_A_T_top
  PIN Tile_X2Y0_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 360.760 1831.640 361.160 1832.520 ;
    END
  END Tile_X2Y0_B_I_top
  PIN Tile_X2Y0_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 355.000 1831.640 355.400 1832.520 ;
    END
  END Tile_X2Y0_B_O_top
  PIN Tile_X2Y0_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 366.520 1831.640 366.920 1832.520 ;
    END
  END Tile_X2Y0_B_T_top
  PIN Tile_X2Y0_C_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.615900 ;
    PORT
      LAYER Metal2 ;
        RECT 378.040 1831.640 378.440 1832.520 ;
    END
  END Tile_X2Y0_C_I_top
  PIN Tile_X2Y0_C_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 372.280 1831.640 372.680 1832.520 ;
    END
  END Tile_X2Y0_C_O_top
  PIN Tile_X2Y0_C_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 383.800 1831.640 384.200 1832.520 ;
    END
  END Tile_X2Y0_C_T_top
  PIN Tile_X2Y0_D_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 395.320 1831.640 395.720 1832.520 ;
    END
  END Tile_X2Y0_D_I_top
  PIN Tile_X2Y0_D_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 389.560 1831.640 389.960 1832.520 ;
    END
  END Tile_X2Y0_D_O_top
  PIN Tile_X2Y0_D_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 401.080 1831.640 401.480 1832.520 ;
    END
  END Tile_X2Y0_D_T_top
  PIN Tile_X2Y9_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 343.480 0.000 343.880 0.480 ;
    END
  END Tile_X2Y9_A_I_top
  PIN Tile_X2Y9_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 337.720 0.000 338.120 0.480 ;
    END
  END Tile_X2Y9_A_O_top
  PIN Tile_X2Y9_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 349.240 0.000 349.640 0.480 ;
    END
  END Tile_X2Y9_A_T_top
  PIN Tile_X2Y9_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 360.760 0.000 361.160 0.480 ;
    END
  END Tile_X2Y9_B_I_top
  PIN Tile_X2Y9_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 355.000 0.000 355.400 0.480 ;
    END
  END Tile_X2Y9_B_O_top
  PIN Tile_X2Y9_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 366.520 0.000 366.920 0.480 ;
    END
  END Tile_X2Y9_B_T_top
  PIN Tile_X2Y9_C_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.615900 ;
    PORT
      LAYER Metal2 ;
        RECT 378.040 0.000 378.440 0.480 ;
    END
  END Tile_X2Y9_C_I_top
  PIN Tile_X2Y9_C_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 372.280 0.000 372.680 0.480 ;
    END
  END Tile_X2Y9_C_O_top
  PIN Tile_X2Y9_C_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 383.800 0.000 384.200 0.480 ;
    END
  END Tile_X2Y9_C_T_top
  PIN Tile_X2Y9_D_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 395.320 0.000 395.720 0.480 ;
    END
  END Tile_X2Y9_D_I_top
  PIN Tile_X2Y9_D_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 389.560 0.000 389.960 0.480 ;
    END
  END Tile_X2Y9_D_O_top
  PIN Tile_X2Y9_D_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 401.080 0.000 401.480 0.480 ;
    END
  END Tile_X2Y9_D_T_top
  PIN Tile_X3Y0_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 558.520 1831.640 558.920 1832.520 ;
    END
  END Tile_X3Y0_A_I_top
  PIN Tile_X3Y0_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 552.760 1831.640 553.160 1832.520 ;
    END
  END Tile_X3Y0_A_O_top
  PIN Tile_X3Y0_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 564.280 1831.640 564.680 1832.520 ;
    END
  END Tile_X3Y0_A_T_top
  PIN Tile_X3Y0_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 575.800 1831.640 576.200 1832.520 ;
    END
  END Tile_X3Y0_B_I_top
  PIN Tile_X3Y0_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 570.040 1831.640 570.440 1832.520 ;
    END
  END Tile_X3Y0_B_O_top
  PIN Tile_X3Y0_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 581.560 1831.640 581.960 1832.520 ;
    END
  END Tile_X3Y0_B_T_top
  PIN Tile_X3Y0_C_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.615900 ;
    PORT
      LAYER Metal2 ;
        RECT 593.080 1831.640 593.480 1832.520 ;
    END
  END Tile_X3Y0_C_I_top
  PIN Tile_X3Y0_C_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 587.320 1831.640 587.720 1832.520 ;
    END
  END Tile_X3Y0_C_O_top
  PIN Tile_X3Y0_C_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 598.840 1831.640 599.240 1832.520 ;
    END
  END Tile_X3Y0_C_T_top
  PIN Tile_X3Y0_D_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 610.360 1831.640 610.760 1832.520 ;
    END
  END Tile_X3Y0_D_I_top
  PIN Tile_X3Y0_D_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 604.600 1831.640 605.000 1832.520 ;
    END
  END Tile_X3Y0_D_O_top
  PIN Tile_X3Y0_D_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 616.120 1831.640 616.520 1832.520 ;
    END
  END Tile_X3Y0_D_T_top
  PIN Tile_X3Y9_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 558.520 0.000 558.920 0.480 ;
    END
  END Tile_X3Y9_A_I_top
  PIN Tile_X3Y9_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 552.760 0.000 553.160 0.480 ;
    END
  END Tile_X3Y9_A_O_top
  PIN Tile_X3Y9_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 564.280 0.000 564.680 0.480 ;
    END
  END Tile_X3Y9_A_T_top
  PIN Tile_X3Y9_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 575.800 0.000 576.200 0.480 ;
    END
  END Tile_X3Y9_B_I_top
  PIN Tile_X3Y9_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 570.040 0.000 570.440 0.480 ;
    END
  END Tile_X3Y9_B_O_top
  PIN Tile_X3Y9_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 581.560 0.000 581.960 0.480 ;
    END
  END Tile_X3Y9_B_T_top
  PIN Tile_X3Y9_C_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.615900 ;
    PORT
      LAYER Metal2 ;
        RECT 593.080 0.000 593.480 0.480 ;
    END
  END Tile_X3Y9_C_I_top
  PIN Tile_X3Y9_C_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 587.320 0.000 587.720 0.480 ;
    END
  END Tile_X3Y9_C_O_top
  PIN Tile_X3Y9_C_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 598.840 0.000 599.240 0.480 ;
    END
  END Tile_X3Y9_C_T_top
  PIN Tile_X3Y9_D_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 610.360 0.000 610.760 0.480 ;
    END
  END Tile_X3Y9_D_I_top
  PIN Tile_X3Y9_D_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 604.600 0.000 605.000 0.480 ;
    END
  END Tile_X3Y9_D_O_top
  PIN Tile_X3Y9_D_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 616.120 0.000 616.520 0.480 ;
    END
  END Tile_X3Y9_D_T_top
  PIN Tile_X4Y0_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 773.560 1831.640 773.960 1832.520 ;
    END
  END Tile_X4Y0_A_I_top
  PIN Tile_X4Y0_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 767.800 1831.640 768.200 1832.520 ;
    END
  END Tile_X4Y0_A_O_top
  PIN Tile_X4Y0_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 779.320 1831.640 779.720 1832.520 ;
    END
  END Tile_X4Y0_A_T_top
  PIN Tile_X4Y0_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 790.840 1831.640 791.240 1832.520 ;
    END
  END Tile_X4Y0_B_I_top
  PIN Tile_X4Y0_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 785.080 1831.640 785.480 1832.520 ;
    END
  END Tile_X4Y0_B_O_top
  PIN Tile_X4Y0_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 796.600 1831.640 797.000 1832.520 ;
    END
  END Tile_X4Y0_B_T_top
  PIN Tile_X4Y0_C_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.615900 ;
    PORT
      LAYER Metal2 ;
        RECT 808.120 1831.640 808.520 1832.520 ;
    END
  END Tile_X4Y0_C_I_top
  PIN Tile_X4Y0_C_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 802.360 1831.640 802.760 1832.520 ;
    END
  END Tile_X4Y0_C_O_top
  PIN Tile_X4Y0_C_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 813.880 1831.640 814.280 1832.520 ;
    END
  END Tile_X4Y0_C_T_top
  PIN Tile_X4Y0_D_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 825.400 1831.640 825.800 1832.520 ;
    END
  END Tile_X4Y0_D_I_top
  PIN Tile_X4Y0_D_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 819.640 1831.640 820.040 1832.520 ;
    END
  END Tile_X4Y0_D_O_top
  PIN Tile_X4Y0_D_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 831.160 1831.640 831.560 1832.520 ;
    END
  END Tile_X4Y0_D_T_top
  PIN Tile_X4Y9_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 773.560 0.000 773.960 0.480 ;
    END
  END Tile_X4Y9_A_I_top
  PIN Tile_X4Y9_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 767.800 0.000 768.200 0.480 ;
    END
  END Tile_X4Y9_A_O_top
  PIN Tile_X4Y9_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 779.320 0.000 779.720 0.480 ;
    END
  END Tile_X4Y9_A_T_top
  PIN Tile_X4Y9_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 790.840 0.000 791.240 0.480 ;
    END
  END Tile_X4Y9_B_I_top
  PIN Tile_X4Y9_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 785.080 0.000 785.480 0.480 ;
    END
  END Tile_X4Y9_B_O_top
  PIN Tile_X4Y9_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 796.600 0.000 797.000 0.480 ;
    END
  END Tile_X4Y9_B_T_top
  PIN Tile_X4Y9_C_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.615900 ;
    PORT
      LAYER Metal2 ;
        RECT 808.120 0.000 808.520 0.480 ;
    END
  END Tile_X4Y9_C_I_top
  PIN Tile_X4Y9_C_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 802.360 0.000 802.760 0.480 ;
    END
  END Tile_X4Y9_C_O_top
  PIN Tile_X4Y9_C_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 813.880 0.000 814.280 0.480 ;
    END
  END Tile_X4Y9_C_T_top
  PIN Tile_X4Y9_D_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 825.400 0.000 825.800 0.480 ;
    END
  END Tile_X4Y9_D_I_top
  PIN Tile_X4Y9_D_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 819.640 0.000 820.040 0.480 ;
    END
  END Tile_X4Y9_D_O_top
  PIN Tile_X4Y9_D_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 831.160 0.000 831.560 0.480 ;
    END
  END Tile_X4Y9_D_T_top
  PIN Tile_X5Y2_ADDR_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1470.220 1076.160 1470.620 ;
    END
  END Tile_X5Y2_ADDR_SRAM0
  PIN Tile_X5Y2_ADDR_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1471.900 1076.160 1472.300 ;
    END
  END Tile_X5Y2_ADDR_SRAM1
  PIN Tile_X5Y2_ADDR_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1473.580 1076.160 1473.980 ;
    END
  END Tile_X5Y2_ADDR_SRAM2
  PIN Tile_X5Y2_ADDR_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1475.260 1076.160 1475.660 ;
    END
  END Tile_X5Y2_ADDR_SRAM3
  PIN Tile_X5Y2_ADDR_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1476.940 1076.160 1477.340 ;
    END
  END Tile_X5Y2_ADDR_SRAM4
  PIN Tile_X5Y2_ADDR_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.135600 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1478.620 1076.160 1479.020 ;
    END
  END Tile_X5Y2_ADDR_SRAM5
  PIN Tile_X5Y2_ADDR_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.135600 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1480.300 1076.160 1480.700 ;
    END
  END Tile_X5Y2_ADDR_SRAM6
  PIN Tile_X5Y2_ADDR_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.135600 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1481.980 1076.160 1482.380 ;
    END
  END Tile_X5Y2_ADDR_SRAM7
  PIN Tile_X5Y2_ADDR_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.135600 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1483.660 1076.160 1484.060 ;
    END
  END Tile_X5Y2_ADDR_SRAM8
  PIN Tile_X5Y2_ADDR_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.135600 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1485.340 1076.160 1485.740 ;
    END
  END Tile_X5Y2_ADDR_SRAM9
  PIN Tile_X5Y2_BM_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1540.780 1076.160 1541.180 ;
    END
  END Tile_X5Y2_BM_SRAM0
  PIN Tile_X5Y2_BM_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1542.460 1076.160 1542.860 ;
    END
  END Tile_X5Y2_BM_SRAM1
  PIN Tile_X5Y2_BM_SRAM10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1557.580 1076.160 1557.980 ;
    END
  END Tile_X5Y2_BM_SRAM10
  PIN Tile_X5Y2_BM_SRAM11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1559.260 1076.160 1559.660 ;
    END
  END Tile_X5Y2_BM_SRAM11
  PIN Tile_X5Y2_BM_SRAM12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1560.940 1076.160 1561.340 ;
    END
  END Tile_X5Y2_BM_SRAM12
  PIN Tile_X5Y2_BM_SRAM13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1562.620 1076.160 1563.020 ;
    END
  END Tile_X5Y2_BM_SRAM13
  PIN Tile_X5Y2_BM_SRAM14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1564.300 1076.160 1564.700 ;
    END
  END Tile_X5Y2_BM_SRAM14
  PIN Tile_X5Y2_BM_SRAM15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1565.980 1076.160 1566.380 ;
    END
  END Tile_X5Y2_BM_SRAM15
  PIN Tile_X5Y2_BM_SRAM16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1567.660 1076.160 1568.060 ;
    END
  END Tile_X5Y2_BM_SRAM16
  PIN Tile_X5Y2_BM_SRAM17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1569.340 1076.160 1569.740 ;
    END
  END Tile_X5Y2_BM_SRAM17
  PIN Tile_X5Y2_BM_SRAM18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1571.020 1076.160 1571.420 ;
    END
  END Tile_X5Y2_BM_SRAM18
  PIN Tile_X5Y2_BM_SRAM19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1572.700 1076.160 1573.100 ;
    END
  END Tile_X5Y2_BM_SRAM19
  PIN Tile_X5Y2_BM_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1544.140 1076.160 1544.540 ;
    END
  END Tile_X5Y2_BM_SRAM2
  PIN Tile_X5Y2_BM_SRAM20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1574.380 1076.160 1574.780 ;
    END
  END Tile_X5Y2_BM_SRAM20
  PIN Tile_X5Y2_BM_SRAM21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1576.060 1076.160 1576.460 ;
    END
  END Tile_X5Y2_BM_SRAM21
  PIN Tile_X5Y2_BM_SRAM22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1577.740 1076.160 1578.140 ;
    END
  END Tile_X5Y2_BM_SRAM22
  PIN Tile_X5Y2_BM_SRAM23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1579.420 1076.160 1579.820 ;
    END
  END Tile_X5Y2_BM_SRAM23
  PIN Tile_X5Y2_BM_SRAM24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1581.100 1076.160 1581.500 ;
    END
  END Tile_X5Y2_BM_SRAM24
  PIN Tile_X5Y2_BM_SRAM25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1582.780 1076.160 1583.180 ;
    END
  END Tile_X5Y2_BM_SRAM25
  PIN Tile_X5Y2_BM_SRAM26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1584.460 1076.160 1584.860 ;
    END
  END Tile_X5Y2_BM_SRAM26
  PIN Tile_X5Y2_BM_SRAM27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1586.140 1076.160 1586.540 ;
    END
  END Tile_X5Y2_BM_SRAM27
  PIN Tile_X5Y2_BM_SRAM28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1587.820 1076.160 1588.220 ;
    END
  END Tile_X5Y2_BM_SRAM28
  PIN Tile_X5Y2_BM_SRAM29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1589.500 1076.160 1589.900 ;
    END
  END Tile_X5Y2_BM_SRAM29
  PIN Tile_X5Y2_BM_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1545.820 1076.160 1546.220 ;
    END
  END Tile_X5Y2_BM_SRAM3
  PIN Tile_X5Y2_BM_SRAM30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1591.180 1076.160 1591.580 ;
    END
  END Tile_X5Y2_BM_SRAM30
  PIN Tile_X5Y2_BM_SRAM31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1592.860 1076.160 1593.260 ;
    END
  END Tile_X5Y2_BM_SRAM31
  PIN Tile_X5Y2_BM_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1547.500 1076.160 1547.900 ;
    END
  END Tile_X5Y2_BM_SRAM4
  PIN Tile_X5Y2_BM_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1549.180 1076.160 1549.580 ;
    END
  END Tile_X5Y2_BM_SRAM5
  PIN Tile_X5Y2_BM_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1550.860 1076.160 1551.260 ;
    END
  END Tile_X5Y2_BM_SRAM6
  PIN Tile_X5Y2_BM_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1552.540 1076.160 1552.940 ;
    END
  END Tile_X5Y2_BM_SRAM7
  PIN Tile_X5Y2_BM_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1554.220 1076.160 1554.620 ;
    END
  END Tile_X5Y2_BM_SRAM8
  PIN Tile_X5Y2_BM_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1555.900 1076.160 1556.300 ;
    END
  END Tile_X5Y2_BM_SRAM9
  PIN Tile_X5Y2_CLK_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1599.580 1076.160 1599.980 ;
    END
  END Tile_X5Y2_CLK_SRAM
  PIN Tile_X5Y2_CONFIGURED_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.300 1468.540 1076.160 1468.940 ;
    END
  END Tile_X5Y2_CONFIGURED_top
  PIN Tile_X5Y2_DIN_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1487.020 1076.160 1487.420 ;
    END
  END Tile_X5Y2_DIN_SRAM0
  PIN Tile_X5Y2_DIN_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1488.700 1076.160 1489.100 ;
    END
  END Tile_X5Y2_DIN_SRAM1
  PIN Tile_X5Y2_DIN_SRAM10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1503.820 1076.160 1504.220 ;
    END
  END Tile_X5Y2_DIN_SRAM10
  PIN Tile_X5Y2_DIN_SRAM11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1505.500 1076.160 1505.900 ;
    END
  END Tile_X5Y2_DIN_SRAM11
  PIN Tile_X5Y2_DIN_SRAM12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1507.180 1076.160 1507.580 ;
    END
  END Tile_X5Y2_DIN_SRAM12
  PIN Tile_X5Y2_DIN_SRAM13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1508.860 1076.160 1509.260 ;
    END
  END Tile_X5Y2_DIN_SRAM13
  PIN Tile_X5Y2_DIN_SRAM14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1510.540 1076.160 1510.940 ;
    END
  END Tile_X5Y2_DIN_SRAM14
  PIN Tile_X5Y2_DIN_SRAM15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1512.220 1076.160 1512.620 ;
    END
  END Tile_X5Y2_DIN_SRAM15
  PIN Tile_X5Y2_DIN_SRAM16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1513.900 1076.160 1514.300 ;
    END
  END Tile_X5Y2_DIN_SRAM16
  PIN Tile_X5Y2_DIN_SRAM17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1515.580 1076.160 1515.980 ;
    END
  END Tile_X5Y2_DIN_SRAM17
  PIN Tile_X5Y2_DIN_SRAM18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1517.260 1076.160 1517.660 ;
    END
  END Tile_X5Y2_DIN_SRAM18
  PIN Tile_X5Y2_DIN_SRAM19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1518.940 1076.160 1519.340 ;
    END
  END Tile_X5Y2_DIN_SRAM19
  PIN Tile_X5Y2_DIN_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1490.380 1076.160 1490.780 ;
    END
  END Tile_X5Y2_DIN_SRAM2
  PIN Tile_X5Y2_DIN_SRAM20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1520.620 1076.160 1521.020 ;
    END
  END Tile_X5Y2_DIN_SRAM20
  PIN Tile_X5Y2_DIN_SRAM21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1522.300 1076.160 1522.700 ;
    END
  END Tile_X5Y2_DIN_SRAM21
  PIN Tile_X5Y2_DIN_SRAM22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1523.980 1076.160 1524.380 ;
    END
  END Tile_X5Y2_DIN_SRAM22
  PIN Tile_X5Y2_DIN_SRAM23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1525.660 1076.160 1526.060 ;
    END
  END Tile_X5Y2_DIN_SRAM23
  PIN Tile_X5Y2_DIN_SRAM24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1527.340 1076.160 1527.740 ;
    END
  END Tile_X5Y2_DIN_SRAM24
  PIN Tile_X5Y2_DIN_SRAM25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1529.020 1076.160 1529.420 ;
    END
  END Tile_X5Y2_DIN_SRAM25
  PIN Tile_X5Y2_DIN_SRAM26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1530.700 1076.160 1531.100 ;
    END
  END Tile_X5Y2_DIN_SRAM26
  PIN Tile_X5Y2_DIN_SRAM27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1532.380 1076.160 1532.780 ;
    END
  END Tile_X5Y2_DIN_SRAM27
  PIN Tile_X5Y2_DIN_SRAM28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1534.060 1076.160 1534.460 ;
    END
  END Tile_X5Y2_DIN_SRAM28
  PIN Tile_X5Y2_DIN_SRAM29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1535.740 1076.160 1536.140 ;
    END
  END Tile_X5Y2_DIN_SRAM29
  PIN Tile_X5Y2_DIN_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1492.060 1076.160 1492.460 ;
    END
  END Tile_X5Y2_DIN_SRAM3
  PIN Tile_X5Y2_DIN_SRAM30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1537.420 1076.160 1537.820 ;
    END
  END Tile_X5Y2_DIN_SRAM30
  PIN Tile_X5Y2_DIN_SRAM31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1539.100 1076.160 1539.500 ;
    END
  END Tile_X5Y2_DIN_SRAM31
  PIN Tile_X5Y2_DIN_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1493.740 1076.160 1494.140 ;
    END
  END Tile_X5Y2_DIN_SRAM4
  PIN Tile_X5Y2_DIN_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1495.420 1076.160 1495.820 ;
    END
  END Tile_X5Y2_DIN_SRAM5
  PIN Tile_X5Y2_DIN_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1497.100 1076.160 1497.500 ;
    END
  END Tile_X5Y2_DIN_SRAM6
  PIN Tile_X5Y2_DIN_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1498.780 1076.160 1499.180 ;
    END
  END Tile_X5Y2_DIN_SRAM7
  PIN Tile_X5Y2_DIN_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1500.460 1076.160 1500.860 ;
    END
  END Tile_X5Y2_DIN_SRAM8
  PIN Tile_X5Y2_DIN_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1502.140 1076.160 1502.540 ;
    END
  END Tile_X5Y2_DIN_SRAM9
  PIN Tile_X5Y2_DOUT_SRAM0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.279200 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1414.780 1076.160 1415.180 ;
    END
  END Tile_X5Y2_DOUT_SRAM0
  PIN Tile_X5Y2_DOUT_SRAM1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.279200 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1416.460 1076.160 1416.860 ;
    END
  END Tile_X5Y2_DOUT_SRAM1
  PIN Tile_X5Y2_DOUT_SRAM10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1431.580 1076.160 1431.980 ;
    END
  END Tile_X5Y2_DOUT_SRAM10
  PIN Tile_X5Y2_DOUT_SRAM11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.300 1433.260 1076.160 1433.660 ;
    END
  END Tile_X5Y2_DOUT_SRAM11
  PIN Tile_X5Y2_DOUT_SRAM12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1434.940 1076.160 1435.340 ;
    END
  END Tile_X5Y2_DOUT_SRAM12
  PIN Tile_X5Y2_DOUT_SRAM13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1436.620 1076.160 1437.020 ;
    END
  END Tile_X5Y2_DOUT_SRAM13
  PIN Tile_X5Y2_DOUT_SRAM14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1438.300 1076.160 1438.700 ;
    END
  END Tile_X5Y2_DOUT_SRAM14
  PIN Tile_X5Y2_DOUT_SRAM15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1439.980 1076.160 1440.380 ;
    END
  END Tile_X5Y2_DOUT_SRAM15
  PIN Tile_X5Y2_DOUT_SRAM16
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.279200 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1441.660 1076.160 1442.060 ;
    END
  END Tile_X5Y2_DOUT_SRAM16
  PIN Tile_X5Y2_DOUT_SRAM17
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.279200 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1443.340 1076.160 1443.740 ;
    END
  END Tile_X5Y2_DOUT_SRAM17
  PIN Tile_X5Y2_DOUT_SRAM18
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.279200 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1445.020 1076.160 1445.420 ;
    END
  END Tile_X5Y2_DOUT_SRAM18
  PIN Tile_X5Y2_DOUT_SRAM19
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.279200 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1446.700 1076.160 1447.100 ;
    END
  END Tile_X5Y2_DOUT_SRAM19
  PIN Tile_X5Y2_DOUT_SRAM2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.279200 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1418.140 1076.160 1418.540 ;
    END
  END Tile_X5Y2_DOUT_SRAM2
  PIN Tile_X5Y2_DOUT_SRAM20
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.279200 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1448.380 1076.160 1448.780 ;
    END
  END Tile_X5Y2_DOUT_SRAM20
  PIN Tile_X5Y2_DOUT_SRAM21
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.279200 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1450.060 1076.160 1450.460 ;
    END
  END Tile_X5Y2_DOUT_SRAM21
  PIN Tile_X5Y2_DOUT_SRAM22
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.279200 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1451.740 1076.160 1452.140 ;
    END
  END Tile_X5Y2_DOUT_SRAM22
  PIN Tile_X5Y2_DOUT_SRAM23
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.279200 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1453.420 1076.160 1453.820 ;
    END
  END Tile_X5Y2_DOUT_SRAM23
  PIN Tile_X5Y2_DOUT_SRAM24
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.066000 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1455.100 1076.160 1455.500 ;
    END
  END Tile_X5Y2_DOUT_SRAM24
  PIN Tile_X5Y2_DOUT_SRAM25
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.639600 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1456.780 1076.160 1457.180 ;
    END
  END Tile_X5Y2_DOUT_SRAM25
  PIN Tile_X5Y2_DOUT_SRAM26
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1458.460 1076.160 1458.860 ;
    END
  END Tile_X5Y2_DOUT_SRAM26
  PIN Tile_X5Y2_DOUT_SRAM27
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1460.140 1076.160 1460.540 ;
    END
  END Tile_X5Y2_DOUT_SRAM27
  PIN Tile_X5Y2_DOUT_SRAM28
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1461.820 1076.160 1462.220 ;
    END
  END Tile_X5Y2_DOUT_SRAM28
  PIN Tile_X5Y2_DOUT_SRAM29
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1463.500 1076.160 1463.900 ;
    END
  END Tile_X5Y2_DOUT_SRAM29
  PIN Tile_X5Y2_DOUT_SRAM3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.279200 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1419.820 1076.160 1420.220 ;
    END
  END Tile_X5Y2_DOUT_SRAM3
  PIN Tile_X5Y2_DOUT_SRAM30
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1465.180 1076.160 1465.580 ;
    END
  END Tile_X5Y2_DOUT_SRAM30
  PIN Tile_X5Y2_DOUT_SRAM31
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1466.860 1076.160 1467.260 ;
    END
  END Tile_X5Y2_DOUT_SRAM31
  PIN Tile_X5Y2_DOUT_SRAM4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.279200 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1421.500 1076.160 1421.900 ;
    END
  END Tile_X5Y2_DOUT_SRAM4
  PIN Tile_X5Y2_DOUT_SRAM5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.279200 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1423.180 1076.160 1423.580 ;
    END
  END Tile_X5Y2_DOUT_SRAM5
  PIN Tile_X5Y2_DOUT_SRAM6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.279200 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1424.860 1076.160 1425.260 ;
    END
  END Tile_X5Y2_DOUT_SRAM6
  PIN Tile_X5Y2_DOUT_SRAM7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.279200 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1426.540 1076.160 1426.940 ;
    END
  END Tile_X5Y2_DOUT_SRAM7
  PIN Tile_X5Y2_DOUT_SRAM8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1428.220 1076.160 1428.620 ;
    END
  END Tile_X5Y2_DOUT_SRAM8
  PIN Tile_X5Y2_DOUT_SRAM9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1429.900 1076.160 1430.300 ;
    END
  END Tile_X5Y2_DOUT_SRAM9
  PIN Tile_X5Y2_MEN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.662000 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1596.220 1076.160 1596.620 ;
    END
  END Tile_X5Y2_MEN_SRAM
  PIN Tile_X5Y2_REN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1597.900 1076.160 1598.300 ;
    END
  END Tile_X5Y2_REN_SRAM
  PIN Tile_X5Y2_TIE_HIGH_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1601.260 1076.160 1601.660 ;
    END
  END Tile_X5Y2_TIE_HIGH_SRAM
  PIN Tile_X5Y2_TIE_LOW_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1602.940 1076.160 1603.340 ;
    END
  END Tile_X5Y2_TIE_LOW_SRAM
  PIN Tile_X5Y2_WEN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.958400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.300 1594.540 1076.160 1594.940 ;
    END
  END Tile_X5Y2_WEN_SRAM
  PIN Tile_X5Y3_CLK_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1250.140 1076.160 1250.540 ;
    END
  END Tile_X5Y3_CLK_TT_PROJECT
  PIN Tile_X5Y3_ENA_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1247.620 1076.160 1248.020 ;
    END
  END Tile_X5Y3_ENA_TT_PROJECT
  PIN Tile_X5Y3_RST_N_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.615900 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.300 1252.660 1076.160 1253.060 ;
    END
  END Tile_X5Y3_RST_N_TT_PROJECT
  PIN Tile_X5Y3_UIO_IN_TT_PROJECT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1227.460 1076.160 1227.860 ;
    END
  END Tile_X5Y3_UIO_IN_TT_PROJECT0
  PIN Tile_X5Y3_UIO_IN_TT_PROJECT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1229.980 1076.160 1230.380 ;
    END
  END Tile_X5Y3_UIO_IN_TT_PROJECT1
  PIN Tile_X5Y3_UIO_IN_TT_PROJECT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1232.500 1076.160 1232.900 ;
    END
  END Tile_X5Y3_UIO_IN_TT_PROJECT2
  PIN Tile_X5Y3_UIO_IN_TT_PROJECT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1235.020 1076.160 1235.420 ;
    END
  END Tile_X5Y3_UIO_IN_TT_PROJECT3
  PIN Tile_X5Y3_UIO_IN_TT_PROJECT4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1237.540 1076.160 1237.940 ;
    END
  END Tile_X5Y3_UIO_IN_TT_PROJECT4
  PIN Tile_X5Y3_UIO_IN_TT_PROJECT5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1240.060 1076.160 1240.460 ;
    END
  END Tile_X5Y3_UIO_IN_TT_PROJECT5
  PIN Tile_X5Y3_UIO_IN_TT_PROJECT6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1242.580 1076.160 1242.980 ;
    END
  END Tile_X5Y3_UIO_IN_TT_PROJECT6
  PIN Tile_X5Y3_UIO_IN_TT_PROJECT7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1245.100 1076.160 1245.500 ;
    END
  END Tile_X5Y3_UIO_IN_TT_PROJECT7
  PIN Tile_X5Y3_UIO_OE_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1187.140 1076.160 1187.540 ;
    END
  END Tile_X5Y3_UIO_OE_TT_PROJECT0
  PIN Tile_X5Y3_UIO_OE_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1189.660 1076.160 1190.060 ;
    END
  END Tile_X5Y3_UIO_OE_TT_PROJECT1
  PIN Tile_X5Y3_UIO_OE_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1192.180 1076.160 1192.580 ;
    END
  END Tile_X5Y3_UIO_OE_TT_PROJECT2
  PIN Tile_X5Y3_UIO_OE_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1194.700 1076.160 1195.100 ;
    END
  END Tile_X5Y3_UIO_OE_TT_PROJECT3
  PIN Tile_X5Y3_UIO_OE_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1197.220 1076.160 1197.620 ;
    END
  END Tile_X5Y3_UIO_OE_TT_PROJECT4
  PIN Tile_X5Y3_UIO_OE_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1199.740 1076.160 1200.140 ;
    END
  END Tile_X5Y3_UIO_OE_TT_PROJECT5
  PIN Tile_X5Y3_UIO_OE_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1202.260 1076.160 1202.660 ;
    END
  END Tile_X5Y3_UIO_OE_TT_PROJECT6
  PIN Tile_X5Y3_UIO_OE_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1204.780 1076.160 1205.180 ;
    END
  END Tile_X5Y3_UIO_OE_TT_PROJECT7
  PIN Tile_X5Y3_UIO_OUT_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1166.980 1076.160 1167.380 ;
    END
  END Tile_X5Y3_UIO_OUT_TT_PROJECT0
  PIN Tile_X5Y3_UIO_OUT_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1169.500 1076.160 1169.900 ;
    END
  END Tile_X5Y3_UIO_OUT_TT_PROJECT1
  PIN Tile_X5Y3_UIO_OUT_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1172.020 1076.160 1172.420 ;
    END
  END Tile_X5Y3_UIO_OUT_TT_PROJECT2
  PIN Tile_X5Y3_UIO_OUT_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1174.540 1076.160 1174.940 ;
    END
  END Tile_X5Y3_UIO_OUT_TT_PROJECT3
  PIN Tile_X5Y3_UIO_OUT_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1177.060 1076.160 1177.460 ;
    END
  END Tile_X5Y3_UIO_OUT_TT_PROJECT4
  PIN Tile_X5Y3_UIO_OUT_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1179.580 1076.160 1179.980 ;
    END
  END Tile_X5Y3_UIO_OUT_TT_PROJECT5
  PIN Tile_X5Y3_UIO_OUT_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1182.100 1076.160 1182.500 ;
    END
  END Tile_X5Y3_UIO_OUT_TT_PROJECT6
  PIN Tile_X5Y3_UIO_OUT_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1184.620 1076.160 1185.020 ;
    END
  END Tile_X5Y3_UIO_OUT_TT_PROJECT7
  PIN Tile_X5Y3_UI_IN_TT_PROJECT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1207.300 1076.160 1207.700 ;
    END
  END Tile_X5Y3_UI_IN_TT_PROJECT0
  PIN Tile_X5Y3_UI_IN_TT_PROJECT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1209.820 1076.160 1210.220 ;
    END
  END Tile_X5Y3_UI_IN_TT_PROJECT1
  PIN Tile_X5Y3_UI_IN_TT_PROJECT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1212.340 1076.160 1212.740 ;
    END
  END Tile_X5Y3_UI_IN_TT_PROJECT2
  PIN Tile_X5Y3_UI_IN_TT_PROJECT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1214.860 1076.160 1215.260 ;
    END
  END Tile_X5Y3_UI_IN_TT_PROJECT3
  PIN Tile_X5Y3_UI_IN_TT_PROJECT4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1217.380 1076.160 1217.780 ;
    END
  END Tile_X5Y3_UI_IN_TT_PROJECT4
  PIN Tile_X5Y3_UI_IN_TT_PROJECT5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1219.900 1076.160 1220.300 ;
    END
  END Tile_X5Y3_UI_IN_TT_PROJECT5
  PIN Tile_X5Y3_UI_IN_TT_PROJECT6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1222.420 1076.160 1222.820 ;
    END
  END Tile_X5Y3_UI_IN_TT_PROJECT6
  PIN Tile_X5Y3_UI_IN_TT_PROJECT7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1224.940 1076.160 1225.340 ;
    END
  END Tile_X5Y3_UI_IN_TT_PROJECT7
  PIN Tile_X5Y3_UO_OUT_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1146.820 1076.160 1147.220 ;
    END
  END Tile_X5Y3_UO_OUT_TT_PROJECT0
  PIN Tile_X5Y3_UO_OUT_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1149.340 1076.160 1149.740 ;
    END
  END Tile_X5Y3_UO_OUT_TT_PROJECT1
  PIN Tile_X5Y3_UO_OUT_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1151.860 1076.160 1152.260 ;
    END
  END Tile_X5Y3_UO_OUT_TT_PROJECT2
  PIN Tile_X5Y3_UO_OUT_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1154.380 1076.160 1154.780 ;
    END
  END Tile_X5Y3_UO_OUT_TT_PROJECT3
  PIN Tile_X5Y3_UO_OUT_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.300 1156.900 1076.160 1157.300 ;
    END
  END Tile_X5Y3_UO_OUT_TT_PROJECT4
  PIN Tile_X5Y3_UO_OUT_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1159.420 1076.160 1159.820 ;
    END
  END Tile_X5Y3_UO_OUT_TT_PROJECT5
  PIN Tile_X5Y3_UO_OUT_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1161.940 1076.160 1162.340 ;
    END
  END Tile_X5Y3_UO_OUT_TT_PROJECT6
  PIN Tile_X5Y3_UO_OUT_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1164.460 1076.160 1164.860 ;
    END
  END Tile_X5Y3_UO_OUT_TT_PROJECT7
  PIN Tile_X5Y4_CLK_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1035.100 1076.160 1035.500 ;
    END
  END Tile_X5Y4_CLK_TT_PROJECT
  PIN Tile_X5Y4_ENA_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1032.580 1076.160 1032.980 ;
    END
  END Tile_X5Y4_ENA_TT_PROJECT
  PIN Tile_X5Y4_RST_N_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.615900 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.300 1037.620 1076.160 1038.020 ;
    END
  END Tile_X5Y4_RST_N_TT_PROJECT
  PIN Tile_X5Y4_UIO_IN_TT_PROJECT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1012.420 1076.160 1012.820 ;
    END
  END Tile_X5Y4_UIO_IN_TT_PROJECT0
  PIN Tile_X5Y4_UIO_IN_TT_PROJECT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1014.940 1076.160 1015.340 ;
    END
  END Tile_X5Y4_UIO_IN_TT_PROJECT1
  PIN Tile_X5Y4_UIO_IN_TT_PROJECT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1017.460 1076.160 1017.860 ;
    END
  END Tile_X5Y4_UIO_IN_TT_PROJECT2
  PIN Tile_X5Y4_UIO_IN_TT_PROJECT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1019.980 1076.160 1020.380 ;
    END
  END Tile_X5Y4_UIO_IN_TT_PROJECT3
  PIN Tile_X5Y4_UIO_IN_TT_PROJECT4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1022.500 1076.160 1022.900 ;
    END
  END Tile_X5Y4_UIO_IN_TT_PROJECT4
  PIN Tile_X5Y4_UIO_IN_TT_PROJECT5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1025.020 1076.160 1025.420 ;
    END
  END Tile_X5Y4_UIO_IN_TT_PROJECT5
  PIN Tile_X5Y4_UIO_IN_TT_PROJECT6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1027.540 1076.160 1027.940 ;
    END
  END Tile_X5Y4_UIO_IN_TT_PROJECT6
  PIN Tile_X5Y4_UIO_IN_TT_PROJECT7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1030.060 1076.160 1030.460 ;
    END
  END Tile_X5Y4_UIO_IN_TT_PROJECT7
  PIN Tile_X5Y4_UIO_OE_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 972.100 1076.160 972.500 ;
    END
  END Tile_X5Y4_UIO_OE_TT_PROJECT0
  PIN Tile_X5Y4_UIO_OE_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 974.620 1076.160 975.020 ;
    END
  END Tile_X5Y4_UIO_OE_TT_PROJECT1
  PIN Tile_X5Y4_UIO_OE_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 977.140 1076.160 977.540 ;
    END
  END Tile_X5Y4_UIO_OE_TT_PROJECT2
  PIN Tile_X5Y4_UIO_OE_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 979.660 1076.160 980.060 ;
    END
  END Tile_X5Y4_UIO_OE_TT_PROJECT3
  PIN Tile_X5Y4_UIO_OE_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 982.180 1076.160 982.580 ;
    END
  END Tile_X5Y4_UIO_OE_TT_PROJECT4
  PIN Tile_X5Y4_UIO_OE_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 984.700 1076.160 985.100 ;
    END
  END Tile_X5Y4_UIO_OE_TT_PROJECT5
  PIN Tile_X5Y4_UIO_OE_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 987.220 1076.160 987.620 ;
    END
  END Tile_X5Y4_UIO_OE_TT_PROJECT6
  PIN Tile_X5Y4_UIO_OE_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 989.740 1076.160 990.140 ;
    END
  END Tile_X5Y4_UIO_OE_TT_PROJECT7
  PIN Tile_X5Y4_UIO_OUT_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 951.940 1076.160 952.340 ;
    END
  END Tile_X5Y4_UIO_OUT_TT_PROJECT0
  PIN Tile_X5Y4_UIO_OUT_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 954.460 1076.160 954.860 ;
    END
  END Tile_X5Y4_UIO_OUT_TT_PROJECT1
  PIN Tile_X5Y4_UIO_OUT_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 956.980 1076.160 957.380 ;
    END
  END Tile_X5Y4_UIO_OUT_TT_PROJECT2
  PIN Tile_X5Y4_UIO_OUT_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 959.500 1076.160 959.900 ;
    END
  END Tile_X5Y4_UIO_OUT_TT_PROJECT3
  PIN Tile_X5Y4_UIO_OUT_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 962.020 1076.160 962.420 ;
    END
  END Tile_X5Y4_UIO_OUT_TT_PROJECT4
  PIN Tile_X5Y4_UIO_OUT_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 964.540 1076.160 964.940 ;
    END
  END Tile_X5Y4_UIO_OUT_TT_PROJECT5
  PIN Tile_X5Y4_UIO_OUT_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 967.060 1076.160 967.460 ;
    END
  END Tile_X5Y4_UIO_OUT_TT_PROJECT6
  PIN Tile_X5Y4_UIO_OUT_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 969.580 1076.160 969.980 ;
    END
  END Tile_X5Y4_UIO_OUT_TT_PROJECT7
  PIN Tile_X5Y4_UI_IN_TT_PROJECT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 992.260 1076.160 992.660 ;
    END
  END Tile_X5Y4_UI_IN_TT_PROJECT0
  PIN Tile_X5Y4_UI_IN_TT_PROJECT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 994.780 1076.160 995.180 ;
    END
  END Tile_X5Y4_UI_IN_TT_PROJECT1
  PIN Tile_X5Y4_UI_IN_TT_PROJECT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 997.300 1076.160 997.700 ;
    END
  END Tile_X5Y4_UI_IN_TT_PROJECT2
  PIN Tile_X5Y4_UI_IN_TT_PROJECT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 999.820 1076.160 1000.220 ;
    END
  END Tile_X5Y4_UI_IN_TT_PROJECT3
  PIN Tile_X5Y4_UI_IN_TT_PROJECT4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1002.340 1076.160 1002.740 ;
    END
  END Tile_X5Y4_UI_IN_TT_PROJECT4
  PIN Tile_X5Y4_UI_IN_TT_PROJECT5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1004.860 1076.160 1005.260 ;
    END
  END Tile_X5Y4_UI_IN_TT_PROJECT5
  PIN Tile_X5Y4_UI_IN_TT_PROJECT6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1007.380 1076.160 1007.780 ;
    END
  END Tile_X5Y4_UI_IN_TT_PROJECT6
  PIN Tile_X5Y4_UI_IN_TT_PROJECT7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 1009.900 1076.160 1010.300 ;
    END
  END Tile_X5Y4_UI_IN_TT_PROJECT7
  PIN Tile_X5Y4_UO_OUT_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 931.780 1076.160 932.180 ;
    END
  END Tile_X5Y4_UO_OUT_TT_PROJECT0
  PIN Tile_X5Y4_UO_OUT_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 934.300 1076.160 934.700 ;
    END
  END Tile_X5Y4_UO_OUT_TT_PROJECT1
  PIN Tile_X5Y4_UO_OUT_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 936.820 1076.160 937.220 ;
    END
  END Tile_X5Y4_UO_OUT_TT_PROJECT2
  PIN Tile_X5Y4_UO_OUT_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 939.340 1076.160 939.740 ;
    END
  END Tile_X5Y4_UO_OUT_TT_PROJECT3
  PIN Tile_X5Y4_UO_OUT_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.300 941.860 1076.160 942.260 ;
    END
  END Tile_X5Y4_UO_OUT_TT_PROJECT4
  PIN Tile_X5Y4_UO_OUT_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 944.380 1076.160 944.780 ;
    END
  END Tile_X5Y4_UO_OUT_TT_PROJECT5
  PIN Tile_X5Y4_UO_OUT_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 946.900 1076.160 947.300 ;
    END
  END Tile_X5Y4_UO_OUT_TT_PROJECT6
  PIN Tile_X5Y4_UO_OUT_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 949.420 1076.160 949.820 ;
    END
  END Tile_X5Y4_UO_OUT_TT_PROJECT7
  PIN Tile_X5Y5_CLK_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 820.060 1076.160 820.460 ;
    END
  END Tile_X5Y5_CLK_TT_PROJECT
  PIN Tile_X5Y5_ENA_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 817.540 1076.160 817.940 ;
    END
  END Tile_X5Y5_ENA_TT_PROJECT
  PIN Tile_X5Y5_RST_N_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.615900 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.300 822.580 1076.160 822.980 ;
    END
  END Tile_X5Y5_RST_N_TT_PROJECT
  PIN Tile_X5Y5_UIO_IN_TT_PROJECT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 797.380 1076.160 797.780 ;
    END
  END Tile_X5Y5_UIO_IN_TT_PROJECT0
  PIN Tile_X5Y5_UIO_IN_TT_PROJECT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 799.900 1076.160 800.300 ;
    END
  END Tile_X5Y5_UIO_IN_TT_PROJECT1
  PIN Tile_X5Y5_UIO_IN_TT_PROJECT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 802.420 1076.160 802.820 ;
    END
  END Tile_X5Y5_UIO_IN_TT_PROJECT2
  PIN Tile_X5Y5_UIO_IN_TT_PROJECT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 804.940 1076.160 805.340 ;
    END
  END Tile_X5Y5_UIO_IN_TT_PROJECT3
  PIN Tile_X5Y5_UIO_IN_TT_PROJECT4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 807.460 1076.160 807.860 ;
    END
  END Tile_X5Y5_UIO_IN_TT_PROJECT4
  PIN Tile_X5Y5_UIO_IN_TT_PROJECT5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 809.980 1076.160 810.380 ;
    END
  END Tile_X5Y5_UIO_IN_TT_PROJECT5
  PIN Tile_X5Y5_UIO_IN_TT_PROJECT6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 812.500 1076.160 812.900 ;
    END
  END Tile_X5Y5_UIO_IN_TT_PROJECT6
  PIN Tile_X5Y5_UIO_IN_TT_PROJECT7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 815.020 1076.160 815.420 ;
    END
  END Tile_X5Y5_UIO_IN_TT_PROJECT7
  PIN Tile_X5Y5_UIO_OE_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 757.060 1076.160 757.460 ;
    END
  END Tile_X5Y5_UIO_OE_TT_PROJECT0
  PIN Tile_X5Y5_UIO_OE_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 759.580 1076.160 759.980 ;
    END
  END Tile_X5Y5_UIO_OE_TT_PROJECT1
  PIN Tile_X5Y5_UIO_OE_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 762.100 1076.160 762.500 ;
    END
  END Tile_X5Y5_UIO_OE_TT_PROJECT2
  PIN Tile_X5Y5_UIO_OE_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 764.620 1076.160 765.020 ;
    END
  END Tile_X5Y5_UIO_OE_TT_PROJECT3
  PIN Tile_X5Y5_UIO_OE_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 767.140 1076.160 767.540 ;
    END
  END Tile_X5Y5_UIO_OE_TT_PROJECT4
  PIN Tile_X5Y5_UIO_OE_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 769.660 1076.160 770.060 ;
    END
  END Tile_X5Y5_UIO_OE_TT_PROJECT5
  PIN Tile_X5Y5_UIO_OE_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 772.180 1076.160 772.580 ;
    END
  END Tile_X5Y5_UIO_OE_TT_PROJECT6
  PIN Tile_X5Y5_UIO_OE_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 774.700 1076.160 775.100 ;
    END
  END Tile_X5Y5_UIO_OE_TT_PROJECT7
  PIN Tile_X5Y5_UIO_OUT_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 736.900 1076.160 737.300 ;
    END
  END Tile_X5Y5_UIO_OUT_TT_PROJECT0
  PIN Tile_X5Y5_UIO_OUT_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 739.420 1076.160 739.820 ;
    END
  END Tile_X5Y5_UIO_OUT_TT_PROJECT1
  PIN Tile_X5Y5_UIO_OUT_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 741.940 1076.160 742.340 ;
    END
  END Tile_X5Y5_UIO_OUT_TT_PROJECT2
  PIN Tile_X5Y5_UIO_OUT_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 744.460 1076.160 744.860 ;
    END
  END Tile_X5Y5_UIO_OUT_TT_PROJECT3
  PIN Tile_X5Y5_UIO_OUT_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 746.980 1076.160 747.380 ;
    END
  END Tile_X5Y5_UIO_OUT_TT_PROJECT4
  PIN Tile_X5Y5_UIO_OUT_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 749.500 1076.160 749.900 ;
    END
  END Tile_X5Y5_UIO_OUT_TT_PROJECT5
  PIN Tile_X5Y5_UIO_OUT_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 752.020 1076.160 752.420 ;
    END
  END Tile_X5Y5_UIO_OUT_TT_PROJECT6
  PIN Tile_X5Y5_UIO_OUT_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 754.540 1076.160 754.940 ;
    END
  END Tile_X5Y5_UIO_OUT_TT_PROJECT7
  PIN Tile_X5Y5_UI_IN_TT_PROJECT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 777.220 1076.160 777.620 ;
    END
  END Tile_X5Y5_UI_IN_TT_PROJECT0
  PIN Tile_X5Y5_UI_IN_TT_PROJECT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 779.740 1076.160 780.140 ;
    END
  END Tile_X5Y5_UI_IN_TT_PROJECT1
  PIN Tile_X5Y5_UI_IN_TT_PROJECT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 782.260 1076.160 782.660 ;
    END
  END Tile_X5Y5_UI_IN_TT_PROJECT2
  PIN Tile_X5Y5_UI_IN_TT_PROJECT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 784.780 1076.160 785.180 ;
    END
  END Tile_X5Y5_UI_IN_TT_PROJECT3
  PIN Tile_X5Y5_UI_IN_TT_PROJECT4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 787.300 1076.160 787.700 ;
    END
  END Tile_X5Y5_UI_IN_TT_PROJECT4
  PIN Tile_X5Y5_UI_IN_TT_PROJECT5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 789.820 1076.160 790.220 ;
    END
  END Tile_X5Y5_UI_IN_TT_PROJECT5
  PIN Tile_X5Y5_UI_IN_TT_PROJECT6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 792.340 1076.160 792.740 ;
    END
  END Tile_X5Y5_UI_IN_TT_PROJECT6
  PIN Tile_X5Y5_UI_IN_TT_PROJECT7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 794.860 1076.160 795.260 ;
    END
  END Tile_X5Y5_UI_IN_TT_PROJECT7
  PIN Tile_X5Y5_UO_OUT_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 716.740 1076.160 717.140 ;
    END
  END Tile_X5Y5_UO_OUT_TT_PROJECT0
  PIN Tile_X5Y5_UO_OUT_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 719.260 1076.160 719.660 ;
    END
  END Tile_X5Y5_UO_OUT_TT_PROJECT1
  PIN Tile_X5Y5_UO_OUT_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 721.780 1076.160 722.180 ;
    END
  END Tile_X5Y5_UO_OUT_TT_PROJECT2
  PIN Tile_X5Y5_UO_OUT_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 724.300 1076.160 724.700 ;
    END
  END Tile_X5Y5_UO_OUT_TT_PROJECT3
  PIN Tile_X5Y5_UO_OUT_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.300 726.820 1076.160 727.220 ;
    END
  END Tile_X5Y5_UO_OUT_TT_PROJECT4
  PIN Tile_X5Y5_UO_OUT_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 729.340 1076.160 729.740 ;
    END
  END Tile_X5Y5_UO_OUT_TT_PROJECT5
  PIN Tile_X5Y5_UO_OUT_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 731.860 1076.160 732.260 ;
    END
  END Tile_X5Y5_UO_OUT_TT_PROJECT6
  PIN Tile_X5Y5_UO_OUT_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 734.380 1076.160 734.780 ;
    END
  END Tile_X5Y5_UO_OUT_TT_PROJECT7
  PIN Tile_X5Y6_CLK_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 605.020 1076.160 605.420 ;
    END
  END Tile_X5Y6_CLK_TT_PROJECT
  PIN Tile_X5Y6_ENA_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 602.500 1076.160 602.900 ;
    END
  END Tile_X5Y6_ENA_TT_PROJECT
  PIN Tile_X5Y6_RST_N_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.615900 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.300 607.540 1076.160 607.940 ;
    END
  END Tile_X5Y6_RST_N_TT_PROJECT
  PIN Tile_X5Y6_UIO_IN_TT_PROJECT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 582.340 1076.160 582.740 ;
    END
  END Tile_X5Y6_UIO_IN_TT_PROJECT0
  PIN Tile_X5Y6_UIO_IN_TT_PROJECT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 584.860 1076.160 585.260 ;
    END
  END Tile_X5Y6_UIO_IN_TT_PROJECT1
  PIN Tile_X5Y6_UIO_IN_TT_PROJECT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 587.380 1076.160 587.780 ;
    END
  END Tile_X5Y6_UIO_IN_TT_PROJECT2
  PIN Tile_X5Y6_UIO_IN_TT_PROJECT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 589.900 1076.160 590.300 ;
    END
  END Tile_X5Y6_UIO_IN_TT_PROJECT3
  PIN Tile_X5Y6_UIO_IN_TT_PROJECT4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 592.420 1076.160 592.820 ;
    END
  END Tile_X5Y6_UIO_IN_TT_PROJECT4
  PIN Tile_X5Y6_UIO_IN_TT_PROJECT5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 594.940 1076.160 595.340 ;
    END
  END Tile_X5Y6_UIO_IN_TT_PROJECT5
  PIN Tile_X5Y6_UIO_IN_TT_PROJECT6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 597.460 1076.160 597.860 ;
    END
  END Tile_X5Y6_UIO_IN_TT_PROJECT6
  PIN Tile_X5Y6_UIO_IN_TT_PROJECT7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 599.980 1076.160 600.380 ;
    END
  END Tile_X5Y6_UIO_IN_TT_PROJECT7
  PIN Tile_X5Y6_UIO_OE_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 542.020 1076.160 542.420 ;
    END
  END Tile_X5Y6_UIO_OE_TT_PROJECT0
  PIN Tile_X5Y6_UIO_OE_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 544.540 1076.160 544.940 ;
    END
  END Tile_X5Y6_UIO_OE_TT_PROJECT1
  PIN Tile_X5Y6_UIO_OE_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 547.060 1076.160 547.460 ;
    END
  END Tile_X5Y6_UIO_OE_TT_PROJECT2
  PIN Tile_X5Y6_UIO_OE_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 549.580 1076.160 549.980 ;
    END
  END Tile_X5Y6_UIO_OE_TT_PROJECT3
  PIN Tile_X5Y6_UIO_OE_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 552.100 1076.160 552.500 ;
    END
  END Tile_X5Y6_UIO_OE_TT_PROJECT4
  PIN Tile_X5Y6_UIO_OE_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 554.620 1076.160 555.020 ;
    END
  END Tile_X5Y6_UIO_OE_TT_PROJECT5
  PIN Tile_X5Y6_UIO_OE_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 557.140 1076.160 557.540 ;
    END
  END Tile_X5Y6_UIO_OE_TT_PROJECT6
  PIN Tile_X5Y6_UIO_OE_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 559.660 1076.160 560.060 ;
    END
  END Tile_X5Y6_UIO_OE_TT_PROJECT7
  PIN Tile_X5Y6_UIO_OUT_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 521.860 1076.160 522.260 ;
    END
  END Tile_X5Y6_UIO_OUT_TT_PROJECT0
  PIN Tile_X5Y6_UIO_OUT_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 524.380 1076.160 524.780 ;
    END
  END Tile_X5Y6_UIO_OUT_TT_PROJECT1
  PIN Tile_X5Y6_UIO_OUT_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 526.900 1076.160 527.300 ;
    END
  END Tile_X5Y6_UIO_OUT_TT_PROJECT2
  PIN Tile_X5Y6_UIO_OUT_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 529.420 1076.160 529.820 ;
    END
  END Tile_X5Y6_UIO_OUT_TT_PROJECT3
  PIN Tile_X5Y6_UIO_OUT_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 531.940 1076.160 532.340 ;
    END
  END Tile_X5Y6_UIO_OUT_TT_PROJECT4
  PIN Tile_X5Y6_UIO_OUT_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 534.460 1076.160 534.860 ;
    END
  END Tile_X5Y6_UIO_OUT_TT_PROJECT5
  PIN Tile_X5Y6_UIO_OUT_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 536.980 1076.160 537.380 ;
    END
  END Tile_X5Y6_UIO_OUT_TT_PROJECT6
  PIN Tile_X5Y6_UIO_OUT_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 539.500 1076.160 539.900 ;
    END
  END Tile_X5Y6_UIO_OUT_TT_PROJECT7
  PIN Tile_X5Y6_UI_IN_TT_PROJECT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 562.180 1076.160 562.580 ;
    END
  END Tile_X5Y6_UI_IN_TT_PROJECT0
  PIN Tile_X5Y6_UI_IN_TT_PROJECT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 564.700 1076.160 565.100 ;
    END
  END Tile_X5Y6_UI_IN_TT_PROJECT1
  PIN Tile_X5Y6_UI_IN_TT_PROJECT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 567.220 1076.160 567.620 ;
    END
  END Tile_X5Y6_UI_IN_TT_PROJECT2
  PIN Tile_X5Y6_UI_IN_TT_PROJECT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 569.740 1076.160 570.140 ;
    END
  END Tile_X5Y6_UI_IN_TT_PROJECT3
  PIN Tile_X5Y6_UI_IN_TT_PROJECT4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 572.260 1076.160 572.660 ;
    END
  END Tile_X5Y6_UI_IN_TT_PROJECT4
  PIN Tile_X5Y6_UI_IN_TT_PROJECT5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 574.780 1076.160 575.180 ;
    END
  END Tile_X5Y6_UI_IN_TT_PROJECT5
  PIN Tile_X5Y6_UI_IN_TT_PROJECT6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 577.300 1076.160 577.700 ;
    END
  END Tile_X5Y6_UI_IN_TT_PROJECT6
  PIN Tile_X5Y6_UI_IN_TT_PROJECT7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 579.820 1076.160 580.220 ;
    END
  END Tile_X5Y6_UI_IN_TT_PROJECT7
  PIN Tile_X5Y6_UO_OUT_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 501.700 1076.160 502.100 ;
    END
  END Tile_X5Y6_UO_OUT_TT_PROJECT0
  PIN Tile_X5Y6_UO_OUT_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 504.220 1076.160 504.620 ;
    END
  END Tile_X5Y6_UO_OUT_TT_PROJECT1
  PIN Tile_X5Y6_UO_OUT_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 506.740 1076.160 507.140 ;
    END
  END Tile_X5Y6_UO_OUT_TT_PROJECT2
  PIN Tile_X5Y6_UO_OUT_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 509.260 1076.160 509.660 ;
    END
  END Tile_X5Y6_UO_OUT_TT_PROJECT3
  PIN Tile_X5Y6_UO_OUT_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.300 511.780 1076.160 512.180 ;
    END
  END Tile_X5Y6_UO_OUT_TT_PROJECT4
  PIN Tile_X5Y6_UO_OUT_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 514.300 1076.160 514.700 ;
    END
  END Tile_X5Y6_UO_OUT_TT_PROJECT5
  PIN Tile_X5Y6_UO_OUT_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 516.820 1076.160 517.220 ;
    END
  END Tile_X5Y6_UO_OUT_TT_PROJECT6
  PIN Tile_X5Y6_UO_OUT_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 519.340 1076.160 519.740 ;
    END
  END Tile_X5Y6_UO_OUT_TT_PROJECT7
  PIN Tile_X5Y7_CLK_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 389.980 1076.160 390.380 ;
    END
  END Tile_X5Y7_CLK_TT_PROJECT
  PIN Tile_X5Y7_ENA_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 387.460 1076.160 387.860 ;
    END
  END Tile_X5Y7_ENA_TT_PROJECT
  PIN Tile_X5Y7_RST_N_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.615900 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.300 392.500 1076.160 392.900 ;
    END
  END Tile_X5Y7_RST_N_TT_PROJECT
  PIN Tile_X5Y7_UIO_IN_TT_PROJECT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 367.300 1076.160 367.700 ;
    END
  END Tile_X5Y7_UIO_IN_TT_PROJECT0
  PIN Tile_X5Y7_UIO_IN_TT_PROJECT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 369.820 1076.160 370.220 ;
    END
  END Tile_X5Y7_UIO_IN_TT_PROJECT1
  PIN Tile_X5Y7_UIO_IN_TT_PROJECT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 372.340 1076.160 372.740 ;
    END
  END Tile_X5Y7_UIO_IN_TT_PROJECT2
  PIN Tile_X5Y7_UIO_IN_TT_PROJECT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 374.860 1076.160 375.260 ;
    END
  END Tile_X5Y7_UIO_IN_TT_PROJECT3
  PIN Tile_X5Y7_UIO_IN_TT_PROJECT4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 377.380 1076.160 377.780 ;
    END
  END Tile_X5Y7_UIO_IN_TT_PROJECT4
  PIN Tile_X5Y7_UIO_IN_TT_PROJECT5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 379.900 1076.160 380.300 ;
    END
  END Tile_X5Y7_UIO_IN_TT_PROJECT5
  PIN Tile_X5Y7_UIO_IN_TT_PROJECT6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 382.420 1076.160 382.820 ;
    END
  END Tile_X5Y7_UIO_IN_TT_PROJECT6
  PIN Tile_X5Y7_UIO_IN_TT_PROJECT7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 384.940 1076.160 385.340 ;
    END
  END Tile_X5Y7_UIO_IN_TT_PROJECT7
  PIN Tile_X5Y7_UIO_OE_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 326.980 1076.160 327.380 ;
    END
  END Tile_X5Y7_UIO_OE_TT_PROJECT0
  PIN Tile_X5Y7_UIO_OE_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 329.500 1076.160 329.900 ;
    END
  END Tile_X5Y7_UIO_OE_TT_PROJECT1
  PIN Tile_X5Y7_UIO_OE_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 332.020 1076.160 332.420 ;
    END
  END Tile_X5Y7_UIO_OE_TT_PROJECT2
  PIN Tile_X5Y7_UIO_OE_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 334.540 1076.160 334.940 ;
    END
  END Tile_X5Y7_UIO_OE_TT_PROJECT3
  PIN Tile_X5Y7_UIO_OE_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 337.060 1076.160 337.460 ;
    END
  END Tile_X5Y7_UIO_OE_TT_PROJECT4
  PIN Tile_X5Y7_UIO_OE_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 339.580 1076.160 339.980 ;
    END
  END Tile_X5Y7_UIO_OE_TT_PROJECT5
  PIN Tile_X5Y7_UIO_OE_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 342.100 1076.160 342.500 ;
    END
  END Tile_X5Y7_UIO_OE_TT_PROJECT6
  PIN Tile_X5Y7_UIO_OE_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 344.620 1076.160 345.020 ;
    END
  END Tile_X5Y7_UIO_OE_TT_PROJECT7
  PIN Tile_X5Y7_UIO_OUT_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 306.820 1076.160 307.220 ;
    END
  END Tile_X5Y7_UIO_OUT_TT_PROJECT0
  PIN Tile_X5Y7_UIO_OUT_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 309.340 1076.160 309.740 ;
    END
  END Tile_X5Y7_UIO_OUT_TT_PROJECT1
  PIN Tile_X5Y7_UIO_OUT_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 311.860 1076.160 312.260 ;
    END
  END Tile_X5Y7_UIO_OUT_TT_PROJECT2
  PIN Tile_X5Y7_UIO_OUT_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 314.380 1076.160 314.780 ;
    END
  END Tile_X5Y7_UIO_OUT_TT_PROJECT3
  PIN Tile_X5Y7_UIO_OUT_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 316.900 1076.160 317.300 ;
    END
  END Tile_X5Y7_UIO_OUT_TT_PROJECT4
  PIN Tile_X5Y7_UIO_OUT_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 319.420 1076.160 319.820 ;
    END
  END Tile_X5Y7_UIO_OUT_TT_PROJECT5
  PIN Tile_X5Y7_UIO_OUT_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 321.940 1076.160 322.340 ;
    END
  END Tile_X5Y7_UIO_OUT_TT_PROJECT6
  PIN Tile_X5Y7_UIO_OUT_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 324.460 1076.160 324.860 ;
    END
  END Tile_X5Y7_UIO_OUT_TT_PROJECT7
  PIN Tile_X5Y7_UI_IN_TT_PROJECT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 347.140 1076.160 347.540 ;
    END
  END Tile_X5Y7_UI_IN_TT_PROJECT0
  PIN Tile_X5Y7_UI_IN_TT_PROJECT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 349.660 1076.160 350.060 ;
    END
  END Tile_X5Y7_UI_IN_TT_PROJECT1
  PIN Tile_X5Y7_UI_IN_TT_PROJECT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 352.180 1076.160 352.580 ;
    END
  END Tile_X5Y7_UI_IN_TT_PROJECT2
  PIN Tile_X5Y7_UI_IN_TT_PROJECT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 354.700 1076.160 355.100 ;
    END
  END Tile_X5Y7_UI_IN_TT_PROJECT3
  PIN Tile_X5Y7_UI_IN_TT_PROJECT4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 357.220 1076.160 357.620 ;
    END
  END Tile_X5Y7_UI_IN_TT_PROJECT4
  PIN Tile_X5Y7_UI_IN_TT_PROJECT5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 359.740 1076.160 360.140 ;
    END
  END Tile_X5Y7_UI_IN_TT_PROJECT5
  PIN Tile_X5Y7_UI_IN_TT_PROJECT6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 362.260 1076.160 362.660 ;
    END
  END Tile_X5Y7_UI_IN_TT_PROJECT6
  PIN Tile_X5Y7_UI_IN_TT_PROJECT7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 364.780 1076.160 365.180 ;
    END
  END Tile_X5Y7_UI_IN_TT_PROJECT7
  PIN Tile_X5Y7_UO_OUT_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 286.660 1076.160 287.060 ;
    END
  END Tile_X5Y7_UO_OUT_TT_PROJECT0
  PIN Tile_X5Y7_UO_OUT_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 289.180 1076.160 289.580 ;
    END
  END Tile_X5Y7_UO_OUT_TT_PROJECT1
  PIN Tile_X5Y7_UO_OUT_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 291.700 1076.160 292.100 ;
    END
  END Tile_X5Y7_UO_OUT_TT_PROJECT2
  PIN Tile_X5Y7_UO_OUT_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 294.220 1076.160 294.620 ;
    END
  END Tile_X5Y7_UO_OUT_TT_PROJECT3
  PIN Tile_X5Y7_UO_OUT_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.300 296.740 1076.160 297.140 ;
    END
  END Tile_X5Y7_UO_OUT_TT_PROJECT4
  PIN Tile_X5Y7_UO_OUT_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 299.260 1076.160 299.660 ;
    END
  END Tile_X5Y7_UO_OUT_TT_PROJECT5
  PIN Tile_X5Y7_UO_OUT_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 301.780 1076.160 302.180 ;
    END
  END Tile_X5Y7_UO_OUT_TT_PROJECT6
  PIN Tile_X5Y7_UO_OUT_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 304.300 1076.160 304.700 ;
    END
  END Tile_X5Y7_UO_OUT_TT_PROJECT7
  PIN Tile_X5Y8_CLK_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 174.940 1076.160 175.340 ;
    END
  END Tile_X5Y8_CLK_TT_PROJECT
  PIN Tile_X5Y8_ENA_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 172.420 1076.160 172.820 ;
    END
  END Tile_X5Y8_ENA_TT_PROJECT
  PIN Tile_X5Y8_RST_N_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.615900 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.300 177.460 1076.160 177.860 ;
    END
  END Tile_X5Y8_RST_N_TT_PROJECT
  PIN Tile_X5Y8_UIO_IN_TT_PROJECT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 152.260 1076.160 152.660 ;
    END
  END Tile_X5Y8_UIO_IN_TT_PROJECT0
  PIN Tile_X5Y8_UIO_IN_TT_PROJECT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 154.780 1076.160 155.180 ;
    END
  END Tile_X5Y8_UIO_IN_TT_PROJECT1
  PIN Tile_X5Y8_UIO_IN_TT_PROJECT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 157.300 1076.160 157.700 ;
    END
  END Tile_X5Y8_UIO_IN_TT_PROJECT2
  PIN Tile_X5Y8_UIO_IN_TT_PROJECT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 159.820 1076.160 160.220 ;
    END
  END Tile_X5Y8_UIO_IN_TT_PROJECT3
  PIN Tile_X5Y8_UIO_IN_TT_PROJECT4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 162.340 1076.160 162.740 ;
    END
  END Tile_X5Y8_UIO_IN_TT_PROJECT4
  PIN Tile_X5Y8_UIO_IN_TT_PROJECT5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 164.860 1076.160 165.260 ;
    END
  END Tile_X5Y8_UIO_IN_TT_PROJECT5
  PIN Tile_X5Y8_UIO_IN_TT_PROJECT6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 167.380 1076.160 167.780 ;
    END
  END Tile_X5Y8_UIO_IN_TT_PROJECT6
  PIN Tile_X5Y8_UIO_IN_TT_PROJECT7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 169.900 1076.160 170.300 ;
    END
  END Tile_X5Y8_UIO_IN_TT_PROJECT7
  PIN Tile_X5Y8_UIO_OE_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 111.940 1076.160 112.340 ;
    END
  END Tile_X5Y8_UIO_OE_TT_PROJECT0
  PIN Tile_X5Y8_UIO_OE_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 114.460 1076.160 114.860 ;
    END
  END Tile_X5Y8_UIO_OE_TT_PROJECT1
  PIN Tile_X5Y8_UIO_OE_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 116.980 1076.160 117.380 ;
    END
  END Tile_X5Y8_UIO_OE_TT_PROJECT2
  PIN Tile_X5Y8_UIO_OE_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 119.500 1076.160 119.900 ;
    END
  END Tile_X5Y8_UIO_OE_TT_PROJECT3
  PIN Tile_X5Y8_UIO_OE_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 122.020 1076.160 122.420 ;
    END
  END Tile_X5Y8_UIO_OE_TT_PROJECT4
  PIN Tile_X5Y8_UIO_OE_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 124.540 1076.160 124.940 ;
    END
  END Tile_X5Y8_UIO_OE_TT_PROJECT5
  PIN Tile_X5Y8_UIO_OE_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 127.060 1076.160 127.460 ;
    END
  END Tile_X5Y8_UIO_OE_TT_PROJECT6
  PIN Tile_X5Y8_UIO_OE_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 129.580 1076.160 129.980 ;
    END
  END Tile_X5Y8_UIO_OE_TT_PROJECT7
  PIN Tile_X5Y8_UIO_OUT_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 91.780 1076.160 92.180 ;
    END
  END Tile_X5Y8_UIO_OUT_TT_PROJECT0
  PIN Tile_X5Y8_UIO_OUT_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 94.300 1076.160 94.700 ;
    END
  END Tile_X5Y8_UIO_OUT_TT_PROJECT1
  PIN Tile_X5Y8_UIO_OUT_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 96.820 1076.160 97.220 ;
    END
  END Tile_X5Y8_UIO_OUT_TT_PROJECT2
  PIN Tile_X5Y8_UIO_OUT_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 99.340 1076.160 99.740 ;
    END
  END Tile_X5Y8_UIO_OUT_TT_PROJECT3
  PIN Tile_X5Y8_UIO_OUT_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 101.860 1076.160 102.260 ;
    END
  END Tile_X5Y8_UIO_OUT_TT_PROJECT4
  PIN Tile_X5Y8_UIO_OUT_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 104.380 1076.160 104.780 ;
    END
  END Tile_X5Y8_UIO_OUT_TT_PROJECT5
  PIN Tile_X5Y8_UIO_OUT_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 106.900 1076.160 107.300 ;
    END
  END Tile_X5Y8_UIO_OUT_TT_PROJECT6
  PIN Tile_X5Y8_UIO_OUT_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 109.420 1076.160 109.820 ;
    END
  END Tile_X5Y8_UIO_OUT_TT_PROJECT7
  PIN Tile_X5Y8_UI_IN_TT_PROJECT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 132.100 1076.160 132.500 ;
    END
  END Tile_X5Y8_UI_IN_TT_PROJECT0
  PIN Tile_X5Y8_UI_IN_TT_PROJECT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 134.620 1076.160 135.020 ;
    END
  END Tile_X5Y8_UI_IN_TT_PROJECT1
  PIN Tile_X5Y8_UI_IN_TT_PROJECT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 137.140 1076.160 137.540 ;
    END
  END Tile_X5Y8_UI_IN_TT_PROJECT2
  PIN Tile_X5Y8_UI_IN_TT_PROJECT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 139.660 1076.160 140.060 ;
    END
  END Tile_X5Y8_UI_IN_TT_PROJECT3
  PIN Tile_X5Y8_UI_IN_TT_PROJECT4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 142.180 1076.160 142.580 ;
    END
  END Tile_X5Y8_UI_IN_TT_PROJECT4
  PIN Tile_X5Y8_UI_IN_TT_PROJECT5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 144.700 1076.160 145.100 ;
    END
  END Tile_X5Y8_UI_IN_TT_PROJECT5
  PIN Tile_X5Y8_UI_IN_TT_PROJECT6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 147.220 1076.160 147.620 ;
    END
  END Tile_X5Y8_UI_IN_TT_PROJECT6
  PIN Tile_X5Y8_UI_IN_TT_PROJECT7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 149.740 1076.160 150.140 ;
    END
  END Tile_X5Y8_UI_IN_TT_PROJECT7
  PIN Tile_X5Y8_UO_OUT_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 71.620 1076.160 72.020 ;
    END
  END Tile_X5Y8_UO_OUT_TT_PROJECT0
  PIN Tile_X5Y8_UO_OUT_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 74.140 1076.160 74.540 ;
    END
  END Tile_X5Y8_UO_OUT_TT_PROJECT1
  PIN Tile_X5Y8_UO_OUT_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 76.660 1076.160 77.060 ;
    END
  END Tile_X5Y8_UO_OUT_TT_PROJECT2
  PIN Tile_X5Y8_UO_OUT_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 79.180 1076.160 79.580 ;
    END
  END Tile_X5Y8_UO_OUT_TT_PROJECT3
  PIN Tile_X5Y8_UO_OUT_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.300 81.700 1076.160 82.100 ;
    END
  END Tile_X5Y8_UO_OUT_TT_PROJECT4
  PIN Tile_X5Y8_UO_OUT_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 84.220 1076.160 84.620 ;
    END
  END Tile_X5Y8_UO_OUT_TT_PROJECT5
  PIN Tile_X5Y8_UO_OUT_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 86.740 1076.160 87.140 ;
    END
  END Tile_X5Y8_UO_OUT_TT_PROJECT6
  PIN Tile_X5Y8_UO_OUT_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 1075.280 89.260 1076.160 89.660 ;
    END
  END Tile_X5Y8_UO_OUT_TT_PROJECT7
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.164600 ;
    PORT
      LAYER Metal2 ;
        RECT 5.560 0.000 5.960 0.480 ;
    END
  END UserCLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER TopMetal1 ;
        RECT 24.940 4.200 27.140 1832.040 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 132.460 4.200 134.660 1832.040 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 208.060 4.200 210.260 1832.040 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 283.660 4.200 285.860 1832.040 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 347.500 4.200 349.700 1832.040 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 423.100 4.200 425.300 1832.040 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 498.700 4.200 500.900 1832.040 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 562.540 4.200 564.740 1832.040 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 638.140 4.200 640.340 1832.040 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 713.740 4.200 715.940 1832.040 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 777.580 4.200 779.780 1832.040 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 853.180 4.200 855.380 1832.040 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 928.780 4.200 930.980 1832.040 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 992.620 4.200 994.820 1832.040 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER TopMetal1 ;
        RECT 18.740 4.200 20.940 1832.040 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 94.340 4.200 96.540 1832.040 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 126.260 4.200 128.460 1832.040 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 201.860 4.200 204.060 1832.040 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 277.460 4.200 279.660 1832.040 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 341.300 4.200 343.500 1832.040 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 416.900 4.200 419.100 1832.040 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 492.500 4.200 494.700 1832.040 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 556.340 4.200 558.540 1832.040 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 631.940 4.200 634.140 1832.040 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 707.540 4.200 709.740 1832.040 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 771.380 4.200 773.580 1832.040 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 846.980 4.200 849.180 1832.040 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 922.580 4.200 924.780 1832.040 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 986.420 4.200 988.620 1832.040 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1062.020 4.200 1064.220 1832.040 ;
    END
  END VPWR
  OBS
      LAYER GatPoly ;
        RECT 6.240 7.830 1069.920 1827.570 ;
      LAYER Metal1 ;
        RECT 6.240 7.760 1070.420 1827.640 ;
      LAYER Metal2 ;
        RECT 0.855 1831.430 122.470 1832.040 ;
        RECT 123.290 1831.430 128.230 1832.040 ;
        RECT 129.050 1831.430 133.990 1832.040 ;
        RECT 134.810 1831.430 139.750 1832.040 ;
        RECT 140.570 1831.430 145.510 1832.040 ;
        RECT 146.330 1831.430 151.270 1832.040 ;
        RECT 152.090 1831.430 157.030 1832.040 ;
        RECT 157.850 1831.430 162.790 1832.040 ;
        RECT 163.610 1831.430 168.550 1832.040 ;
        RECT 169.370 1831.430 174.310 1832.040 ;
        RECT 175.130 1831.430 180.070 1832.040 ;
        RECT 180.890 1831.430 185.830 1832.040 ;
        RECT 186.650 1831.430 337.510 1832.040 ;
        RECT 338.330 1831.430 343.270 1832.040 ;
        RECT 344.090 1831.430 349.030 1832.040 ;
        RECT 349.850 1831.430 354.790 1832.040 ;
        RECT 355.610 1831.430 360.550 1832.040 ;
        RECT 361.370 1831.430 366.310 1832.040 ;
        RECT 367.130 1831.430 372.070 1832.040 ;
        RECT 372.890 1831.430 377.830 1832.040 ;
        RECT 378.650 1831.430 383.590 1832.040 ;
        RECT 384.410 1831.430 389.350 1832.040 ;
        RECT 390.170 1831.430 395.110 1832.040 ;
        RECT 395.930 1831.430 400.870 1832.040 ;
        RECT 401.690 1831.430 552.550 1832.040 ;
        RECT 553.370 1831.430 558.310 1832.040 ;
        RECT 559.130 1831.430 564.070 1832.040 ;
        RECT 564.890 1831.430 569.830 1832.040 ;
        RECT 570.650 1831.430 575.590 1832.040 ;
        RECT 576.410 1831.430 581.350 1832.040 ;
        RECT 582.170 1831.430 587.110 1832.040 ;
        RECT 587.930 1831.430 592.870 1832.040 ;
        RECT 593.690 1831.430 598.630 1832.040 ;
        RECT 599.450 1831.430 604.390 1832.040 ;
        RECT 605.210 1831.430 610.150 1832.040 ;
        RECT 610.970 1831.430 615.910 1832.040 ;
        RECT 616.730 1831.430 767.590 1832.040 ;
        RECT 768.410 1831.430 773.350 1832.040 ;
        RECT 774.170 1831.430 779.110 1832.040 ;
        RECT 779.930 1831.430 784.870 1832.040 ;
        RECT 785.690 1831.430 790.630 1832.040 ;
        RECT 791.450 1831.430 796.390 1832.040 ;
        RECT 797.210 1831.430 802.150 1832.040 ;
        RECT 802.970 1831.430 807.910 1832.040 ;
        RECT 808.730 1831.430 813.670 1832.040 ;
        RECT 814.490 1831.430 819.430 1832.040 ;
        RECT 820.250 1831.430 825.190 1832.040 ;
        RECT 826.010 1831.430 830.950 1832.040 ;
        RECT 831.770 1831.430 1075.305 1832.040 ;
        RECT 0.855 0.690 1075.305 1831.430 ;
        RECT 0.855 0.275 5.350 0.690 ;
        RECT 6.170 0.275 10.150 0.690 ;
        RECT 10.970 0.275 14.950 0.690 ;
        RECT 15.770 0.275 19.750 0.690 ;
        RECT 20.570 0.275 24.550 0.690 ;
        RECT 25.370 0.275 29.350 0.690 ;
        RECT 30.170 0.275 34.150 0.690 ;
        RECT 34.970 0.275 38.950 0.690 ;
        RECT 39.770 0.275 43.750 0.690 ;
        RECT 44.570 0.275 48.550 0.690 ;
        RECT 49.370 0.275 53.350 0.690 ;
        RECT 54.170 0.275 58.150 0.690 ;
        RECT 58.970 0.275 62.950 0.690 ;
        RECT 63.770 0.275 67.750 0.690 ;
        RECT 68.570 0.275 72.550 0.690 ;
        RECT 73.370 0.275 77.350 0.690 ;
        RECT 78.170 0.275 82.150 0.690 ;
        RECT 82.970 0.275 86.950 0.690 ;
        RECT 87.770 0.275 91.750 0.690 ;
        RECT 92.570 0.275 96.550 0.690 ;
        RECT 97.370 0.275 101.350 0.690 ;
        RECT 102.170 0.275 122.470 0.690 ;
        RECT 123.290 0.275 128.230 0.690 ;
        RECT 129.050 0.275 133.990 0.690 ;
        RECT 134.810 0.275 139.750 0.690 ;
        RECT 140.570 0.275 145.510 0.690 ;
        RECT 146.330 0.275 151.270 0.690 ;
        RECT 152.090 0.275 157.030 0.690 ;
        RECT 157.850 0.275 162.790 0.690 ;
        RECT 163.610 0.275 168.550 0.690 ;
        RECT 169.370 0.275 174.310 0.690 ;
        RECT 175.130 0.275 180.070 0.690 ;
        RECT 180.890 0.275 185.830 0.690 ;
        RECT 186.650 0.275 197.350 0.690 ;
        RECT 198.170 0.275 203.110 0.690 ;
        RECT 203.930 0.275 208.870 0.690 ;
        RECT 209.690 0.275 214.630 0.690 ;
        RECT 215.450 0.275 220.390 0.690 ;
        RECT 221.210 0.275 226.150 0.690 ;
        RECT 226.970 0.275 231.910 0.690 ;
        RECT 232.730 0.275 237.670 0.690 ;
        RECT 238.490 0.275 243.430 0.690 ;
        RECT 244.250 0.275 249.190 0.690 ;
        RECT 250.010 0.275 254.950 0.690 ;
        RECT 255.770 0.275 260.710 0.690 ;
        RECT 261.530 0.275 266.470 0.690 ;
        RECT 267.290 0.275 272.230 0.690 ;
        RECT 273.050 0.275 277.990 0.690 ;
        RECT 278.810 0.275 283.750 0.690 ;
        RECT 284.570 0.275 289.510 0.690 ;
        RECT 290.330 0.275 295.270 0.690 ;
        RECT 296.090 0.275 301.030 0.690 ;
        RECT 301.850 0.275 306.790 0.690 ;
        RECT 307.610 0.275 337.510 0.690 ;
        RECT 338.330 0.275 343.270 0.690 ;
        RECT 344.090 0.275 349.030 0.690 ;
        RECT 349.850 0.275 354.790 0.690 ;
        RECT 355.610 0.275 360.550 0.690 ;
        RECT 361.370 0.275 366.310 0.690 ;
        RECT 367.130 0.275 372.070 0.690 ;
        RECT 372.890 0.275 377.830 0.690 ;
        RECT 378.650 0.275 383.590 0.690 ;
        RECT 384.410 0.275 389.350 0.690 ;
        RECT 390.170 0.275 395.110 0.690 ;
        RECT 395.930 0.275 400.870 0.690 ;
        RECT 401.690 0.275 412.390 0.690 ;
        RECT 413.210 0.275 418.150 0.690 ;
        RECT 418.970 0.275 423.910 0.690 ;
        RECT 424.730 0.275 429.670 0.690 ;
        RECT 430.490 0.275 435.430 0.690 ;
        RECT 436.250 0.275 441.190 0.690 ;
        RECT 442.010 0.275 446.950 0.690 ;
        RECT 447.770 0.275 452.710 0.690 ;
        RECT 453.530 0.275 458.470 0.690 ;
        RECT 459.290 0.275 464.230 0.690 ;
        RECT 465.050 0.275 469.990 0.690 ;
        RECT 470.810 0.275 475.750 0.690 ;
        RECT 476.570 0.275 481.510 0.690 ;
        RECT 482.330 0.275 487.270 0.690 ;
        RECT 488.090 0.275 493.030 0.690 ;
        RECT 493.850 0.275 498.790 0.690 ;
        RECT 499.610 0.275 504.550 0.690 ;
        RECT 505.370 0.275 510.310 0.690 ;
        RECT 511.130 0.275 516.070 0.690 ;
        RECT 516.890 0.275 521.830 0.690 ;
        RECT 522.650 0.275 552.550 0.690 ;
        RECT 553.370 0.275 558.310 0.690 ;
        RECT 559.130 0.275 564.070 0.690 ;
        RECT 564.890 0.275 569.830 0.690 ;
        RECT 570.650 0.275 575.590 0.690 ;
        RECT 576.410 0.275 581.350 0.690 ;
        RECT 582.170 0.275 587.110 0.690 ;
        RECT 587.930 0.275 592.870 0.690 ;
        RECT 593.690 0.275 598.630 0.690 ;
        RECT 599.450 0.275 604.390 0.690 ;
        RECT 605.210 0.275 610.150 0.690 ;
        RECT 610.970 0.275 615.910 0.690 ;
        RECT 616.730 0.275 627.430 0.690 ;
        RECT 628.250 0.275 633.190 0.690 ;
        RECT 634.010 0.275 638.950 0.690 ;
        RECT 639.770 0.275 644.710 0.690 ;
        RECT 645.530 0.275 650.470 0.690 ;
        RECT 651.290 0.275 656.230 0.690 ;
        RECT 657.050 0.275 661.990 0.690 ;
        RECT 662.810 0.275 667.750 0.690 ;
        RECT 668.570 0.275 673.510 0.690 ;
        RECT 674.330 0.275 679.270 0.690 ;
        RECT 680.090 0.275 685.030 0.690 ;
        RECT 685.850 0.275 690.790 0.690 ;
        RECT 691.610 0.275 696.550 0.690 ;
        RECT 697.370 0.275 702.310 0.690 ;
        RECT 703.130 0.275 708.070 0.690 ;
        RECT 708.890 0.275 713.830 0.690 ;
        RECT 714.650 0.275 719.590 0.690 ;
        RECT 720.410 0.275 725.350 0.690 ;
        RECT 726.170 0.275 731.110 0.690 ;
        RECT 731.930 0.275 736.870 0.690 ;
        RECT 737.690 0.275 767.590 0.690 ;
        RECT 768.410 0.275 773.350 0.690 ;
        RECT 774.170 0.275 779.110 0.690 ;
        RECT 779.930 0.275 784.870 0.690 ;
        RECT 785.690 0.275 790.630 0.690 ;
        RECT 791.450 0.275 796.390 0.690 ;
        RECT 797.210 0.275 802.150 0.690 ;
        RECT 802.970 0.275 807.910 0.690 ;
        RECT 808.730 0.275 813.670 0.690 ;
        RECT 814.490 0.275 819.430 0.690 ;
        RECT 820.250 0.275 825.190 0.690 ;
        RECT 826.010 0.275 830.950 0.690 ;
        RECT 831.770 0.275 842.470 0.690 ;
        RECT 843.290 0.275 848.230 0.690 ;
        RECT 849.050 0.275 853.990 0.690 ;
        RECT 854.810 0.275 859.750 0.690 ;
        RECT 860.570 0.275 865.510 0.690 ;
        RECT 866.330 0.275 871.270 0.690 ;
        RECT 872.090 0.275 877.030 0.690 ;
        RECT 877.850 0.275 882.790 0.690 ;
        RECT 883.610 0.275 888.550 0.690 ;
        RECT 889.370 0.275 894.310 0.690 ;
        RECT 895.130 0.275 900.070 0.690 ;
        RECT 900.890 0.275 905.830 0.690 ;
        RECT 906.650 0.275 911.590 0.690 ;
        RECT 912.410 0.275 917.350 0.690 ;
        RECT 918.170 0.275 923.110 0.690 ;
        RECT 923.930 0.275 928.870 0.690 ;
        RECT 929.690 0.275 934.630 0.690 ;
        RECT 935.450 0.275 940.390 0.690 ;
        RECT 941.210 0.275 946.150 0.690 ;
        RECT 946.970 0.275 951.910 0.690 ;
        RECT 952.730 0.275 977.830 0.690 ;
        RECT 978.650 0.275 982.630 0.690 ;
        RECT 983.450 0.275 987.430 0.690 ;
        RECT 988.250 0.275 992.230 0.690 ;
        RECT 993.050 0.275 997.030 0.690 ;
        RECT 997.850 0.275 1001.830 0.690 ;
        RECT 1002.650 0.275 1006.630 0.690 ;
        RECT 1007.450 0.275 1011.430 0.690 ;
        RECT 1012.250 0.275 1016.230 0.690 ;
        RECT 1017.050 0.275 1021.030 0.690 ;
        RECT 1021.850 0.275 1025.830 0.690 ;
        RECT 1026.650 0.275 1030.630 0.690 ;
        RECT 1031.450 0.275 1035.430 0.690 ;
        RECT 1036.250 0.275 1040.230 0.690 ;
        RECT 1041.050 0.275 1045.030 0.690 ;
        RECT 1045.850 0.275 1049.830 0.690 ;
        RECT 1050.650 0.275 1054.630 0.690 ;
        RECT 1055.450 0.275 1059.430 0.690 ;
        RECT 1060.250 0.275 1064.230 0.690 ;
        RECT 1065.050 0.275 1069.030 0.690 ;
        RECT 1069.850 0.275 1075.305 0.690 ;
      LAYER Metal3 ;
        RECT 0.580 1831.190 1075.680 1831.720 ;
        RECT 1.090 1830.370 1075.680 1831.190 ;
        RECT 0.580 1829.510 1075.680 1830.370 ;
        RECT 1.090 1828.690 1075.680 1829.510 ;
        RECT 0.580 1827.830 1075.680 1828.690 ;
        RECT 1.090 1827.010 1075.680 1827.830 ;
        RECT 0.580 1826.150 1075.680 1827.010 ;
        RECT 1.090 1825.330 1075.680 1826.150 ;
        RECT 0.580 1824.470 1075.680 1825.330 ;
        RECT 1.090 1823.650 1075.680 1824.470 ;
        RECT 0.580 1822.790 1075.680 1823.650 ;
        RECT 1.090 1821.970 1075.680 1822.790 ;
        RECT 0.580 1821.110 1075.680 1821.970 ;
        RECT 1.090 1820.290 1075.680 1821.110 ;
        RECT 0.580 1819.430 1075.680 1820.290 ;
        RECT 1.090 1818.610 1075.680 1819.430 ;
        RECT 0.580 1817.750 1075.680 1818.610 ;
        RECT 1.090 1816.930 1075.680 1817.750 ;
        RECT 0.580 1816.070 1075.680 1816.930 ;
        RECT 1.090 1815.250 1075.680 1816.070 ;
        RECT 0.580 1814.390 1075.680 1815.250 ;
        RECT 1.090 1813.570 1075.680 1814.390 ;
        RECT 0.580 1812.710 1075.680 1813.570 ;
        RECT 1.090 1811.890 1075.680 1812.710 ;
        RECT 0.580 1811.030 1075.680 1811.890 ;
        RECT 1.090 1810.210 1075.680 1811.030 ;
        RECT 0.580 1809.350 1075.680 1810.210 ;
        RECT 1.090 1808.530 1075.680 1809.350 ;
        RECT 0.580 1807.670 1075.680 1808.530 ;
        RECT 1.090 1806.850 1075.680 1807.670 ;
        RECT 0.580 1805.990 1075.680 1806.850 ;
        RECT 1.090 1805.170 1075.680 1805.990 ;
        RECT 0.580 1804.310 1075.680 1805.170 ;
        RECT 1.090 1803.490 1075.680 1804.310 ;
        RECT 0.580 1802.630 1075.680 1803.490 ;
        RECT 1.090 1801.810 1075.680 1802.630 ;
        RECT 0.580 1800.950 1075.680 1801.810 ;
        RECT 1.090 1800.130 1075.680 1800.950 ;
        RECT 0.580 1799.270 1075.680 1800.130 ;
        RECT 1.090 1798.450 1075.680 1799.270 ;
        RECT 0.580 1797.590 1075.680 1798.450 ;
        RECT 1.090 1796.770 1075.680 1797.590 ;
        RECT 0.580 1795.910 1075.680 1796.770 ;
        RECT 1.090 1795.090 1075.680 1795.910 ;
        RECT 0.580 1794.230 1075.680 1795.090 ;
        RECT 1.090 1793.410 1075.680 1794.230 ;
        RECT 0.580 1792.550 1075.680 1793.410 ;
        RECT 1.090 1791.730 1075.680 1792.550 ;
        RECT 0.580 1790.870 1075.680 1791.730 ;
        RECT 1.090 1790.050 1075.680 1790.870 ;
        RECT 0.580 1789.190 1075.680 1790.050 ;
        RECT 1.090 1788.370 1075.680 1789.190 ;
        RECT 0.580 1787.510 1075.680 1788.370 ;
        RECT 1.090 1786.690 1075.680 1787.510 ;
        RECT 0.580 1785.830 1075.680 1786.690 ;
        RECT 1.090 1785.010 1075.680 1785.830 ;
        RECT 0.580 1784.150 1075.680 1785.010 ;
        RECT 1.090 1783.330 1075.680 1784.150 ;
        RECT 0.580 1782.470 1075.680 1783.330 ;
        RECT 1.090 1781.650 1075.680 1782.470 ;
        RECT 0.580 1780.790 1075.680 1781.650 ;
        RECT 1.090 1779.970 1075.680 1780.790 ;
        RECT 0.580 1779.110 1075.680 1779.970 ;
        RECT 1.090 1778.290 1075.680 1779.110 ;
        RECT 0.580 1763.990 1075.680 1778.290 ;
        RECT 1.090 1763.170 1075.680 1763.990 ;
        RECT 0.580 1761.470 1075.680 1763.170 ;
        RECT 1.090 1760.650 1075.680 1761.470 ;
        RECT 0.580 1758.950 1075.680 1760.650 ;
        RECT 1.090 1758.130 1075.680 1758.950 ;
        RECT 0.580 1756.430 1075.680 1758.130 ;
        RECT 1.090 1755.610 1075.680 1756.430 ;
        RECT 0.580 1753.910 1075.680 1755.610 ;
        RECT 1.090 1753.090 1075.680 1753.910 ;
        RECT 0.580 1751.390 1075.680 1753.090 ;
        RECT 1.090 1750.570 1075.680 1751.390 ;
        RECT 0.580 1748.870 1075.680 1750.570 ;
        RECT 1.090 1748.050 1075.680 1748.870 ;
        RECT 0.580 1746.350 1075.680 1748.050 ;
        RECT 1.090 1745.530 1075.680 1746.350 ;
        RECT 0.580 1743.830 1075.680 1745.530 ;
        RECT 1.090 1743.010 1075.680 1743.830 ;
        RECT 0.580 1741.310 1075.680 1743.010 ;
        RECT 1.090 1740.490 1075.680 1741.310 ;
        RECT 0.580 1738.790 1075.680 1740.490 ;
        RECT 1.090 1737.970 1075.680 1738.790 ;
        RECT 0.580 1736.270 1075.680 1737.970 ;
        RECT 1.090 1735.450 1075.680 1736.270 ;
        RECT 0.580 1733.750 1075.680 1735.450 ;
        RECT 1.090 1732.930 1075.680 1733.750 ;
        RECT 0.580 1731.230 1075.680 1732.930 ;
        RECT 1.090 1730.410 1075.680 1731.230 ;
        RECT 0.580 1728.710 1075.680 1730.410 ;
        RECT 1.090 1727.890 1075.680 1728.710 ;
        RECT 0.580 1726.190 1075.680 1727.890 ;
        RECT 1.090 1725.370 1075.680 1726.190 ;
        RECT 0.580 1723.670 1075.680 1725.370 ;
        RECT 1.090 1722.850 1075.680 1723.670 ;
        RECT 0.580 1721.150 1075.680 1722.850 ;
        RECT 1.090 1720.330 1075.680 1721.150 ;
        RECT 0.580 1718.630 1075.680 1720.330 ;
        RECT 1.090 1717.810 1075.680 1718.630 ;
        RECT 0.580 1716.110 1075.680 1717.810 ;
        RECT 1.090 1715.290 1075.680 1716.110 ;
        RECT 0.580 1713.590 1075.680 1715.290 ;
        RECT 1.090 1712.770 1075.680 1713.590 ;
        RECT 0.580 1711.070 1075.680 1712.770 ;
        RECT 1.090 1710.250 1075.680 1711.070 ;
        RECT 0.580 1708.550 1075.680 1710.250 ;
        RECT 1.090 1707.730 1075.680 1708.550 ;
        RECT 0.580 1706.030 1075.680 1707.730 ;
        RECT 1.090 1705.210 1075.680 1706.030 ;
        RECT 0.580 1703.510 1075.680 1705.210 ;
        RECT 1.090 1702.690 1075.680 1703.510 ;
        RECT 0.580 1700.990 1075.680 1702.690 ;
        RECT 1.090 1700.170 1075.680 1700.990 ;
        RECT 0.580 1698.470 1075.680 1700.170 ;
        RECT 1.090 1697.650 1075.680 1698.470 ;
        RECT 0.580 1695.950 1075.680 1697.650 ;
        RECT 1.070 1695.130 1075.680 1695.950 ;
        RECT 0.580 1693.430 1075.680 1695.130 ;
        RECT 1.090 1692.610 1075.680 1693.430 ;
        RECT 0.580 1690.910 1075.680 1692.610 ;
        RECT 1.090 1690.090 1075.680 1690.910 ;
        RECT 0.580 1688.390 1075.680 1690.090 ;
        RECT 1.090 1687.570 1075.680 1688.390 ;
        RECT 0.580 1685.870 1075.680 1687.570 ;
        RECT 1.090 1685.050 1075.680 1685.870 ;
        RECT 0.580 1683.350 1075.680 1685.050 ;
        RECT 1.070 1682.530 1075.680 1683.350 ;
        RECT 0.580 1680.830 1075.680 1682.530 ;
        RECT 1.090 1680.010 1075.680 1680.830 ;
        RECT 0.580 1678.310 1075.680 1680.010 ;
        RECT 1.090 1677.490 1075.680 1678.310 ;
        RECT 0.580 1675.790 1075.680 1677.490 ;
        RECT 1.090 1674.970 1075.680 1675.790 ;
        RECT 0.580 1673.270 1075.680 1674.970 ;
        RECT 1.090 1672.450 1075.680 1673.270 ;
        RECT 0.580 1670.750 1075.680 1672.450 ;
        RECT 1.090 1669.930 1075.680 1670.750 ;
        RECT 0.580 1668.230 1075.680 1669.930 ;
        RECT 1.090 1667.410 1075.680 1668.230 ;
        RECT 0.580 1665.710 1075.680 1667.410 ;
        RECT 1.090 1664.890 1075.680 1665.710 ;
        RECT 0.580 1663.190 1075.680 1664.890 ;
        RECT 1.090 1662.370 1075.680 1663.190 ;
        RECT 0.580 1660.670 1075.680 1662.370 ;
        RECT 1.090 1659.850 1075.680 1660.670 ;
        RECT 0.580 1658.150 1075.680 1659.850 ;
        RECT 1.090 1657.330 1075.680 1658.150 ;
        RECT 0.580 1655.630 1075.680 1657.330 ;
        RECT 1.090 1654.810 1075.680 1655.630 ;
        RECT 0.580 1653.110 1075.680 1654.810 ;
        RECT 1.070 1652.290 1075.680 1653.110 ;
        RECT 0.580 1650.590 1075.680 1652.290 ;
        RECT 1.090 1649.770 1075.680 1650.590 ;
        RECT 0.580 1648.070 1075.680 1649.770 ;
        RECT 1.090 1647.250 1075.680 1648.070 ;
        RECT 0.580 1645.550 1075.680 1647.250 ;
        RECT 1.090 1644.730 1075.680 1645.550 ;
        RECT 0.580 1643.030 1075.680 1644.730 ;
        RECT 1.090 1642.210 1075.680 1643.030 ;
        RECT 0.580 1640.510 1075.680 1642.210 ;
        RECT 1.090 1639.690 1075.680 1640.510 ;
        RECT 0.580 1637.990 1075.680 1639.690 ;
        RECT 1.090 1637.170 1075.680 1637.990 ;
        RECT 0.580 1635.470 1075.680 1637.170 ;
        RECT 1.090 1634.650 1075.680 1635.470 ;
        RECT 0.580 1632.950 1075.680 1634.650 ;
        RECT 1.090 1632.130 1075.680 1632.950 ;
        RECT 0.580 1630.430 1075.680 1632.130 ;
        RECT 1.090 1629.610 1075.680 1630.430 ;
        RECT 0.580 1627.910 1075.680 1629.610 ;
        RECT 1.090 1627.090 1075.680 1627.910 ;
        RECT 0.580 1625.390 1075.680 1627.090 ;
        RECT 1.090 1624.570 1075.680 1625.390 ;
        RECT 0.580 1622.870 1075.680 1624.570 ;
        RECT 1.090 1622.050 1075.680 1622.870 ;
        RECT 0.580 1620.350 1075.680 1622.050 ;
        RECT 1.090 1619.530 1075.680 1620.350 ;
        RECT 0.580 1617.830 1075.680 1619.530 ;
        RECT 1.090 1617.010 1075.680 1617.830 ;
        RECT 0.580 1615.310 1075.680 1617.010 ;
        RECT 1.090 1614.490 1075.680 1615.310 ;
        RECT 0.580 1612.790 1075.680 1614.490 ;
        RECT 1.090 1611.970 1075.680 1612.790 ;
        RECT 0.580 1610.270 1075.680 1611.970 ;
        RECT 1.090 1609.450 1075.680 1610.270 ;
        RECT 0.580 1607.750 1075.680 1609.450 ;
        RECT 1.090 1606.930 1075.680 1607.750 ;
        RECT 0.580 1605.230 1075.680 1606.930 ;
        RECT 1.090 1604.410 1075.680 1605.230 ;
        RECT 0.580 1603.550 1075.680 1604.410 ;
        RECT 0.580 1602.730 1075.070 1603.550 ;
        RECT 0.580 1602.710 1075.680 1602.730 ;
        RECT 1.090 1601.890 1075.680 1602.710 ;
        RECT 0.580 1601.870 1075.680 1601.890 ;
        RECT 0.580 1601.050 1075.070 1601.870 ;
        RECT 0.580 1600.190 1075.680 1601.050 ;
        RECT 1.090 1599.370 1075.070 1600.190 ;
        RECT 0.580 1598.510 1075.680 1599.370 ;
        RECT 0.580 1597.690 1075.070 1598.510 ;
        RECT 0.580 1597.670 1075.680 1597.690 ;
        RECT 1.090 1596.850 1075.680 1597.670 ;
        RECT 0.580 1596.830 1075.680 1596.850 ;
        RECT 0.580 1596.010 1075.070 1596.830 ;
        RECT 0.580 1595.150 1075.680 1596.010 ;
        RECT 1.090 1594.330 1075.090 1595.150 ;
        RECT 0.580 1593.470 1075.680 1594.330 ;
        RECT 0.580 1592.650 1075.070 1593.470 ;
        RECT 0.580 1592.630 1075.680 1592.650 ;
        RECT 1.090 1591.810 1075.680 1592.630 ;
        RECT 0.580 1591.790 1075.680 1591.810 ;
        RECT 0.580 1590.970 1075.070 1591.790 ;
        RECT 0.580 1590.110 1075.680 1590.970 ;
        RECT 1.090 1589.290 1075.070 1590.110 ;
        RECT 0.580 1588.430 1075.680 1589.290 ;
        RECT 0.580 1587.610 1075.070 1588.430 ;
        RECT 0.580 1587.590 1075.680 1587.610 ;
        RECT 1.090 1586.770 1075.680 1587.590 ;
        RECT 0.580 1586.750 1075.680 1586.770 ;
        RECT 0.580 1585.930 1075.070 1586.750 ;
        RECT 0.580 1585.070 1075.680 1585.930 ;
        RECT 1.090 1584.250 1075.070 1585.070 ;
        RECT 0.580 1583.390 1075.680 1584.250 ;
        RECT 0.580 1582.570 1075.070 1583.390 ;
        RECT 0.580 1582.550 1075.680 1582.570 ;
        RECT 1.090 1581.730 1075.680 1582.550 ;
        RECT 0.580 1581.710 1075.680 1581.730 ;
        RECT 0.580 1580.890 1075.070 1581.710 ;
        RECT 0.580 1580.030 1075.680 1580.890 ;
        RECT 1.090 1579.210 1075.070 1580.030 ;
        RECT 0.580 1578.350 1075.680 1579.210 ;
        RECT 0.580 1577.530 1075.070 1578.350 ;
        RECT 0.580 1577.510 1075.680 1577.530 ;
        RECT 1.090 1576.690 1075.680 1577.510 ;
        RECT 0.580 1576.670 1075.680 1576.690 ;
        RECT 0.580 1575.850 1075.070 1576.670 ;
        RECT 0.580 1574.990 1075.680 1575.850 ;
        RECT 0.580 1574.170 1075.070 1574.990 ;
        RECT 0.580 1573.310 1075.680 1574.170 ;
        RECT 0.580 1572.490 1075.070 1573.310 ;
        RECT 0.580 1571.630 1075.680 1572.490 ;
        RECT 0.580 1570.810 1075.070 1571.630 ;
        RECT 0.580 1569.950 1075.680 1570.810 ;
        RECT 0.580 1569.130 1075.070 1569.950 ;
        RECT 0.580 1568.270 1075.680 1569.130 ;
        RECT 0.580 1567.450 1075.070 1568.270 ;
        RECT 0.580 1566.590 1075.680 1567.450 ;
        RECT 0.580 1565.770 1075.070 1566.590 ;
        RECT 0.580 1564.910 1075.680 1565.770 ;
        RECT 0.580 1564.090 1075.070 1564.910 ;
        RECT 0.580 1563.230 1075.680 1564.090 ;
        RECT 0.580 1562.410 1075.070 1563.230 ;
        RECT 0.580 1561.550 1075.680 1562.410 ;
        RECT 0.580 1560.730 1075.070 1561.550 ;
        RECT 0.580 1559.870 1075.680 1560.730 ;
        RECT 0.580 1559.050 1075.070 1559.870 ;
        RECT 0.580 1558.190 1075.680 1559.050 ;
        RECT 0.580 1557.370 1075.070 1558.190 ;
        RECT 0.580 1556.510 1075.680 1557.370 ;
        RECT 0.580 1555.690 1075.070 1556.510 ;
        RECT 0.580 1554.830 1075.680 1555.690 ;
        RECT 0.580 1554.010 1075.070 1554.830 ;
        RECT 0.580 1553.150 1075.680 1554.010 ;
        RECT 0.580 1552.330 1075.070 1553.150 ;
        RECT 0.580 1551.470 1075.680 1552.330 ;
        RECT 0.580 1550.650 1075.070 1551.470 ;
        RECT 0.580 1549.790 1075.680 1550.650 ;
        RECT 0.580 1548.970 1075.070 1549.790 ;
        RECT 0.580 1548.950 1075.680 1548.970 ;
        RECT 1.090 1548.130 1075.680 1548.950 ;
        RECT 0.580 1548.110 1075.680 1548.130 ;
        RECT 0.580 1547.290 1075.070 1548.110 ;
        RECT 0.580 1546.430 1075.680 1547.290 ;
        RECT 1.090 1545.610 1075.070 1546.430 ;
        RECT 0.580 1544.750 1075.680 1545.610 ;
        RECT 0.580 1543.930 1075.070 1544.750 ;
        RECT 0.580 1543.910 1075.680 1543.930 ;
        RECT 1.090 1543.090 1075.680 1543.910 ;
        RECT 0.580 1543.070 1075.680 1543.090 ;
        RECT 0.580 1542.250 1075.070 1543.070 ;
        RECT 0.580 1541.390 1075.680 1542.250 ;
        RECT 1.090 1540.570 1075.070 1541.390 ;
        RECT 0.580 1539.710 1075.680 1540.570 ;
        RECT 0.580 1538.890 1075.070 1539.710 ;
        RECT 0.580 1538.870 1075.680 1538.890 ;
        RECT 1.090 1538.050 1075.680 1538.870 ;
        RECT 0.580 1538.030 1075.680 1538.050 ;
        RECT 0.580 1537.210 1075.070 1538.030 ;
        RECT 0.580 1536.350 1075.680 1537.210 ;
        RECT 1.090 1535.530 1075.070 1536.350 ;
        RECT 0.580 1534.670 1075.680 1535.530 ;
        RECT 0.580 1533.850 1075.070 1534.670 ;
        RECT 0.580 1533.830 1075.680 1533.850 ;
        RECT 1.090 1533.010 1075.680 1533.830 ;
        RECT 0.580 1532.990 1075.680 1533.010 ;
        RECT 0.580 1532.170 1075.070 1532.990 ;
        RECT 0.580 1531.310 1075.680 1532.170 ;
        RECT 1.090 1530.490 1075.070 1531.310 ;
        RECT 0.580 1529.630 1075.680 1530.490 ;
        RECT 0.580 1528.810 1075.070 1529.630 ;
        RECT 0.580 1528.790 1075.680 1528.810 ;
        RECT 1.090 1527.970 1075.680 1528.790 ;
        RECT 0.580 1527.950 1075.680 1527.970 ;
        RECT 0.580 1527.130 1075.070 1527.950 ;
        RECT 0.580 1526.270 1075.680 1527.130 ;
        RECT 1.090 1525.450 1075.070 1526.270 ;
        RECT 0.580 1524.590 1075.680 1525.450 ;
        RECT 0.580 1523.770 1075.070 1524.590 ;
        RECT 0.580 1523.750 1075.680 1523.770 ;
        RECT 1.090 1522.930 1075.680 1523.750 ;
        RECT 0.580 1522.910 1075.680 1522.930 ;
        RECT 0.580 1522.090 1075.070 1522.910 ;
        RECT 0.580 1521.230 1075.680 1522.090 ;
        RECT 1.090 1520.410 1075.070 1521.230 ;
        RECT 0.580 1519.550 1075.680 1520.410 ;
        RECT 0.580 1518.730 1075.070 1519.550 ;
        RECT 0.580 1518.710 1075.680 1518.730 ;
        RECT 1.090 1517.890 1075.680 1518.710 ;
        RECT 0.580 1517.870 1075.680 1517.890 ;
        RECT 0.580 1517.050 1075.070 1517.870 ;
        RECT 0.580 1516.190 1075.680 1517.050 ;
        RECT 1.090 1515.370 1075.070 1516.190 ;
        RECT 0.580 1514.510 1075.680 1515.370 ;
        RECT 0.580 1513.690 1075.070 1514.510 ;
        RECT 0.580 1513.670 1075.680 1513.690 ;
        RECT 1.090 1512.850 1075.680 1513.670 ;
        RECT 0.580 1512.830 1075.680 1512.850 ;
        RECT 0.580 1512.010 1075.070 1512.830 ;
        RECT 0.580 1511.150 1075.680 1512.010 ;
        RECT 1.090 1510.330 1075.070 1511.150 ;
        RECT 0.580 1509.470 1075.680 1510.330 ;
        RECT 0.580 1508.650 1075.070 1509.470 ;
        RECT 0.580 1508.630 1075.680 1508.650 ;
        RECT 1.090 1507.810 1075.680 1508.630 ;
        RECT 0.580 1507.790 1075.680 1507.810 ;
        RECT 0.580 1506.970 1075.070 1507.790 ;
        RECT 0.580 1506.110 1075.680 1506.970 ;
        RECT 1.090 1505.290 1075.070 1506.110 ;
        RECT 0.580 1504.430 1075.680 1505.290 ;
        RECT 0.580 1503.610 1075.070 1504.430 ;
        RECT 0.580 1503.590 1075.680 1503.610 ;
        RECT 1.090 1502.770 1075.680 1503.590 ;
        RECT 0.580 1502.750 1075.680 1502.770 ;
        RECT 0.580 1501.930 1075.070 1502.750 ;
        RECT 0.580 1501.070 1075.680 1501.930 ;
        RECT 1.090 1500.250 1075.070 1501.070 ;
        RECT 0.580 1499.390 1075.680 1500.250 ;
        RECT 0.580 1498.570 1075.070 1499.390 ;
        RECT 0.580 1498.550 1075.680 1498.570 ;
        RECT 1.090 1497.730 1075.680 1498.550 ;
        RECT 0.580 1497.710 1075.680 1497.730 ;
        RECT 0.580 1496.890 1075.070 1497.710 ;
        RECT 0.580 1496.030 1075.680 1496.890 ;
        RECT 1.090 1495.210 1075.070 1496.030 ;
        RECT 0.580 1494.350 1075.680 1495.210 ;
        RECT 0.580 1493.530 1075.070 1494.350 ;
        RECT 0.580 1493.510 1075.680 1493.530 ;
        RECT 1.090 1492.690 1075.680 1493.510 ;
        RECT 0.580 1492.670 1075.680 1492.690 ;
        RECT 0.580 1491.850 1075.070 1492.670 ;
        RECT 0.580 1490.990 1075.680 1491.850 ;
        RECT 1.090 1490.170 1075.070 1490.990 ;
        RECT 0.580 1489.310 1075.680 1490.170 ;
        RECT 0.580 1488.490 1075.070 1489.310 ;
        RECT 0.580 1488.470 1075.680 1488.490 ;
        RECT 1.090 1487.650 1075.680 1488.470 ;
        RECT 0.580 1487.630 1075.680 1487.650 ;
        RECT 0.580 1486.810 1075.070 1487.630 ;
        RECT 0.580 1485.950 1075.680 1486.810 ;
        RECT 1.090 1485.130 1075.070 1485.950 ;
        RECT 0.580 1484.270 1075.680 1485.130 ;
        RECT 0.580 1483.450 1075.070 1484.270 ;
        RECT 0.580 1483.430 1075.680 1483.450 ;
        RECT 1.090 1482.610 1075.680 1483.430 ;
        RECT 0.580 1482.590 1075.680 1482.610 ;
        RECT 0.580 1481.770 1075.070 1482.590 ;
        RECT 0.580 1480.910 1075.680 1481.770 ;
        RECT 1.070 1480.090 1075.070 1480.910 ;
        RECT 0.580 1479.230 1075.680 1480.090 ;
        RECT 0.580 1478.410 1075.070 1479.230 ;
        RECT 0.580 1478.390 1075.680 1478.410 ;
        RECT 1.090 1477.570 1075.680 1478.390 ;
        RECT 0.580 1477.550 1075.680 1477.570 ;
        RECT 0.580 1476.730 1075.070 1477.550 ;
        RECT 0.580 1475.870 1075.680 1476.730 ;
        RECT 1.090 1475.050 1075.070 1475.870 ;
        RECT 0.580 1474.190 1075.680 1475.050 ;
        RECT 0.580 1473.370 1075.070 1474.190 ;
        RECT 0.580 1473.350 1075.680 1473.370 ;
        RECT 1.090 1472.530 1075.680 1473.350 ;
        RECT 0.580 1472.510 1075.680 1472.530 ;
        RECT 0.580 1471.690 1075.070 1472.510 ;
        RECT 0.580 1470.830 1075.680 1471.690 ;
        RECT 1.090 1470.010 1075.070 1470.830 ;
        RECT 0.580 1469.150 1075.680 1470.010 ;
        RECT 0.580 1468.330 1075.090 1469.150 ;
        RECT 0.580 1468.310 1075.680 1468.330 ;
        RECT 1.070 1467.490 1075.680 1468.310 ;
        RECT 0.580 1467.470 1075.680 1467.490 ;
        RECT 0.580 1466.650 1075.070 1467.470 ;
        RECT 0.580 1465.790 1075.680 1466.650 ;
        RECT 1.090 1464.970 1075.070 1465.790 ;
        RECT 0.580 1464.110 1075.680 1464.970 ;
        RECT 0.580 1463.290 1075.070 1464.110 ;
        RECT 0.580 1463.270 1075.680 1463.290 ;
        RECT 1.090 1462.450 1075.680 1463.270 ;
        RECT 0.580 1462.430 1075.680 1462.450 ;
        RECT 0.580 1461.610 1075.070 1462.430 ;
        RECT 0.580 1460.750 1075.680 1461.610 ;
        RECT 1.090 1459.930 1075.070 1460.750 ;
        RECT 0.580 1459.070 1075.680 1459.930 ;
        RECT 0.580 1458.250 1075.070 1459.070 ;
        RECT 0.580 1458.230 1075.680 1458.250 ;
        RECT 1.090 1457.410 1075.680 1458.230 ;
        RECT 0.580 1457.390 1075.680 1457.410 ;
        RECT 0.580 1456.570 1075.070 1457.390 ;
        RECT 0.580 1455.710 1075.680 1456.570 ;
        RECT 1.090 1454.890 1075.070 1455.710 ;
        RECT 0.580 1454.030 1075.680 1454.890 ;
        RECT 0.580 1453.210 1075.070 1454.030 ;
        RECT 0.580 1453.190 1075.680 1453.210 ;
        RECT 1.090 1452.370 1075.680 1453.190 ;
        RECT 0.580 1452.350 1075.680 1452.370 ;
        RECT 0.580 1451.530 1075.070 1452.350 ;
        RECT 0.580 1450.670 1075.680 1451.530 ;
        RECT 1.090 1449.850 1075.070 1450.670 ;
        RECT 0.580 1448.990 1075.680 1449.850 ;
        RECT 0.580 1448.170 1075.070 1448.990 ;
        RECT 0.580 1448.150 1075.680 1448.170 ;
        RECT 1.090 1447.330 1075.680 1448.150 ;
        RECT 0.580 1447.310 1075.680 1447.330 ;
        RECT 0.580 1446.490 1075.070 1447.310 ;
        RECT 0.580 1445.630 1075.680 1446.490 ;
        RECT 1.090 1444.810 1075.070 1445.630 ;
        RECT 0.580 1443.950 1075.680 1444.810 ;
        RECT 0.580 1443.130 1075.070 1443.950 ;
        RECT 0.580 1443.110 1075.680 1443.130 ;
        RECT 1.090 1442.290 1075.680 1443.110 ;
        RECT 0.580 1442.270 1075.680 1442.290 ;
        RECT 0.580 1441.450 1075.070 1442.270 ;
        RECT 0.580 1440.590 1075.680 1441.450 ;
        RECT 1.090 1439.770 1075.070 1440.590 ;
        RECT 0.580 1438.910 1075.680 1439.770 ;
        RECT 0.580 1438.090 1075.070 1438.910 ;
        RECT 0.580 1438.070 1075.680 1438.090 ;
        RECT 1.070 1437.250 1075.680 1438.070 ;
        RECT 0.580 1437.230 1075.680 1437.250 ;
        RECT 0.580 1436.410 1075.070 1437.230 ;
        RECT 0.580 1435.550 1075.680 1436.410 ;
        RECT 1.090 1434.730 1075.070 1435.550 ;
        RECT 0.580 1433.870 1075.680 1434.730 ;
        RECT 0.580 1433.050 1075.090 1433.870 ;
        RECT 0.580 1433.030 1075.680 1433.050 ;
        RECT 1.090 1432.210 1075.680 1433.030 ;
        RECT 0.580 1432.190 1075.680 1432.210 ;
        RECT 0.580 1431.370 1075.070 1432.190 ;
        RECT 0.580 1430.510 1075.680 1431.370 ;
        RECT 1.090 1429.690 1075.070 1430.510 ;
        RECT 0.580 1428.830 1075.680 1429.690 ;
        RECT 0.580 1428.010 1075.070 1428.830 ;
        RECT 0.580 1427.990 1075.680 1428.010 ;
        RECT 1.090 1427.170 1075.680 1427.990 ;
        RECT 0.580 1427.150 1075.680 1427.170 ;
        RECT 0.580 1426.330 1075.070 1427.150 ;
        RECT 0.580 1425.470 1075.680 1426.330 ;
        RECT 1.090 1424.650 1075.070 1425.470 ;
        RECT 0.580 1423.790 1075.680 1424.650 ;
        RECT 0.580 1422.970 1075.070 1423.790 ;
        RECT 0.580 1422.950 1075.680 1422.970 ;
        RECT 1.090 1422.130 1075.680 1422.950 ;
        RECT 0.580 1422.110 1075.680 1422.130 ;
        RECT 0.580 1421.290 1075.070 1422.110 ;
        RECT 0.580 1420.430 1075.680 1421.290 ;
        RECT 1.090 1419.610 1075.070 1420.430 ;
        RECT 0.580 1418.750 1075.680 1419.610 ;
        RECT 0.580 1417.930 1075.070 1418.750 ;
        RECT 0.580 1417.910 1075.680 1417.930 ;
        RECT 1.090 1417.090 1075.680 1417.910 ;
        RECT 0.580 1417.070 1075.680 1417.090 ;
        RECT 0.580 1416.250 1075.070 1417.070 ;
        RECT 0.580 1415.390 1075.680 1416.250 ;
        RECT 1.090 1414.570 1075.070 1415.390 ;
        RECT 0.580 1412.870 1075.680 1414.570 ;
        RECT 1.090 1412.050 1075.680 1412.870 ;
        RECT 0.580 1410.350 1075.680 1412.050 ;
        RECT 1.090 1409.530 1075.680 1410.350 ;
        RECT 0.580 1407.830 1075.680 1409.530 ;
        RECT 1.090 1407.010 1075.680 1407.830 ;
        RECT 0.580 1405.310 1075.680 1407.010 ;
        RECT 1.090 1404.490 1075.680 1405.310 ;
        RECT 0.580 1402.790 1075.680 1404.490 ;
        RECT 1.090 1401.970 1075.680 1402.790 ;
        RECT 0.580 1400.270 1075.680 1401.970 ;
        RECT 1.090 1399.450 1075.680 1400.270 ;
        RECT 0.580 1397.750 1075.680 1399.450 ;
        RECT 1.090 1396.930 1075.680 1397.750 ;
        RECT 0.580 1395.230 1075.680 1396.930 ;
        RECT 1.090 1394.410 1075.680 1395.230 ;
        RECT 0.580 1392.710 1075.680 1394.410 ;
        RECT 1.090 1391.890 1075.680 1392.710 ;
        RECT 0.580 1390.190 1075.680 1391.890 ;
        RECT 1.090 1389.370 1075.680 1390.190 ;
        RECT 0.580 1387.670 1075.680 1389.370 ;
        RECT 1.090 1386.850 1075.680 1387.670 ;
        RECT 0.580 1385.150 1075.680 1386.850 ;
        RECT 1.090 1384.330 1075.680 1385.150 ;
        RECT 0.580 1382.630 1075.680 1384.330 ;
        RECT 1.090 1381.810 1075.680 1382.630 ;
        RECT 0.580 1380.110 1075.680 1381.810 ;
        RECT 1.090 1379.290 1075.680 1380.110 ;
        RECT 0.580 1377.590 1075.680 1379.290 ;
        RECT 1.090 1376.770 1075.680 1377.590 ;
        RECT 0.580 1375.070 1075.680 1376.770 ;
        RECT 1.090 1374.250 1075.680 1375.070 ;
        RECT 0.580 1372.550 1075.680 1374.250 ;
        RECT 1.090 1371.730 1075.680 1372.550 ;
        RECT 0.580 1370.030 1075.680 1371.730 ;
        RECT 1.090 1369.210 1075.680 1370.030 ;
        RECT 0.580 1367.510 1075.680 1369.210 ;
        RECT 1.090 1366.690 1075.680 1367.510 ;
        RECT 0.580 1364.990 1075.680 1366.690 ;
        RECT 1.090 1364.170 1075.680 1364.990 ;
        RECT 0.580 1362.470 1075.680 1364.170 ;
        RECT 1.090 1361.650 1075.680 1362.470 ;
        RECT 0.580 1333.910 1075.680 1361.650 ;
        RECT 1.090 1333.090 1075.680 1333.910 ;
        RECT 0.580 1331.390 1075.680 1333.090 ;
        RECT 1.090 1330.570 1075.680 1331.390 ;
        RECT 0.580 1328.870 1075.680 1330.570 ;
        RECT 1.090 1328.050 1075.680 1328.870 ;
        RECT 0.580 1326.350 1075.680 1328.050 ;
        RECT 1.090 1325.530 1075.680 1326.350 ;
        RECT 0.580 1323.830 1075.680 1325.530 ;
        RECT 1.090 1323.010 1075.680 1323.830 ;
        RECT 0.580 1321.310 1075.680 1323.010 ;
        RECT 1.090 1320.490 1075.680 1321.310 ;
        RECT 0.580 1318.790 1075.680 1320.490 ;
        RECT 1.090 1317.970 1075.680 1318.790 ;
        RECT 0.580 1316.270 1075.680 1317.970 ;
        RECT 1.090 1315.450 1075.680 1316.270 ;
        RECT 0.580 1313.750 1075.680 1315.450 ;
        RECT 1.090 1312.930 1075.680 1313.750 ;
        RECT 0.580 1311.230 1075.680 1312.930 ;
        RECT 1.090 1310.410 1075.680 1311.230 ;
        RECT 0.580 1308.710 1075.680 1310.410 ;
        RECT 1.090 1307.890 1075.680 1308.710 ;
        RECT 0.580 1306.190 1075.680 1307.890 ;
        RECT 1.090 1305.370 1075.680 1306.190 ;
        RECT 0.580 1303.670 1075.680 1305.370 ;
        RECT 1.090 1302.850 1075.680 1303.670 ;
        RECT 0.580 1301.150 1075.680 1302.850 ;
        RECT 1.090 1300.330 1075.680 1301.150 ;
        RECT 0.580 1298.630 1075.680 1300.330 ;
        RECT 1.090 1297.810 1075.680 1298.630 ;
        RECT 0.580 1296.110 1075.680 1297.810 ;
        RECT 1.090 1295.290 1075.680 1296.110 ;
        RECT 0.580 1293.590 1075.680 1295.290 ;
        RECT 1.090 1292.770 1075.680 1293.590 ;
        RECT 0.580 1291.070 1075.680 1292.770 ;
        RECT 1.090 1290.250 1075.680 1291.070 ;
        RECT 0.580 1288.550 1075.680 1290.250 ;
        RECT 1.090 1287.730 1075.680 1288.550 ;
        RECT 0.580 1286.030 1075.680 1287.730 ;
        RECT 1.090 1285.210 1075.680 1286.030 ;
        RECT 0.580 1283.510 1075.680 1285.210 ;
        RECT 1.090 1282.690 1075.680 1283.510 ;
        RECT 0.580 1280.990 1075.680 1282.690 ;
        RECT 1.090 1280.170 1075.680 1280.990 ;
        RECT 0.580 1278.470 1075.680 1280.170 ;
        RECT 1.090 1277.650 1075.680 1278.470 ;
        RECT 0.580 1275.950 1075.680 1277.650 ;
        RECT 1.090 1275.130 1075.680 1275.950 ;
        RECT 0.580 1273.430 1075.680 1275.130 ;
        RECT 1.090 1272.610 1075.680 1273.430 ;
        RECT 0.580 1270.910 1075.680 1272.610 ;
        RECT 1.090 1270.090 1075.680 1270.910 ;
        RECT 0.580 1268.390 1075.680 1270.090 ;
        RECT 1.090 1267.570 1075.680 1268.390 ;
        RECT 0.580 1265.870 1075.680 1267.570 ;
        RECT 1.070 1265.050 1075.680 1265.870 ;
        RECT 0.580 1263.350 1075.680 1265.050 ;
        RECT 1.090 1262.530 1075.680 1263.350 ;
        RECT 0.580 1260.830 1075.680 1262.530 ;
        RECT 1.090 1260.010 1075.680 1260.830 ;
        RECT 0.580 1258.310 1075.680 1260.010 ;
        RECT 1.090 1257.490 1075.680 1258.310 ;
        RECT 0.580 1255.790 1075.680 1257.490 ;
        RECT 1.090 1254.970 1075.680 1255.790 ;
        RECT 0.580 1253.270 1075.680 1254.970 ;
        RECT 1.070 1252.450 1075.090 1253.270 ;
        RECT 0.580 1250.750 1075.680 1252.450 ;
        RECT 1.090 1249.930 1075.070 1250.750 ;
        RECT 0.580 1248.230 1075.680 1249.930 ;
        RECT 1.090 1247.410 1075.070 1248.230 ;
        RECT 0.580 1245.710 1075.680 1247.410 ;
        RECT 1.090 1244.890 1075.070 1245.710 ;
        RECT 0.580 1243.190 1075.680 1244.890 ;
        RECT 1.090 1242.370 1075.070 1243.190 ;
        RECT 0.580 1240.670 1075.680 1242.370 ;
        RECT 1.090 1239.850 1075.070 1240.670 ;
        RECT 0.580 1238.150 1075.680 1239.850 ;
        RECT 1.090 1237.330 1075.070 1238.150 ;
        RECT 0.580 1235.630 1075.680 1237.330 ;
        RECT 1.090 1234.810 1075.070 1235.630 ;
        RECT 0.580 1233.110 1075.680 1234.810 ;
        RECT 1.090 1232.290 1075.070 1233.110 ;
        RECT 0.580 1230.590 1075.680 1232.290 ;
        RECT 1.090 1229.770 1075.070 1230.590 ;
        RECT 0.580 1228.070 1075.680 1229.770 ;
        RECT 1.090 1227.250 1075.070 1228.070 ;
        RECT 0.580 1225.550 1075.680 1227.250 ;
        RECT 1.090 1224.730 1075.070 1225.550 ;
        RECT 0.580 1223.030 1075.680 1224.730 ;
        RECT 1.070 1222.210 1075.070 1223.030 ;
        RECT 0.580 1220.510 1075.680 1222.210 ;
        RECT 1.090 1219.690 1075.070 1220.510 ;
        RECT 0.580 1217.990 1075.680 1219.690 ;
        RECT 1.090 1217.170 1075.070 1217.990 ;
        RECT 0.580 1215.470 1075.680 1217.170 ;
        RECT 1.090 1214.650 1075.070 1215.470 ;
        RECT 0.580 1212.950 1075.680 1214.650 ;
        RECT 1.090 1212.130 1075.070 1212.950 ;
        RECT 0.580 1210.430 1075.680 1212.130 ;
        RECT 1.090 1209.610 1075.070 1210.430 ;
        RECT 0.580 1207.910 1075.680 1209.610 ;
        RECT 1.090 1207.090 1075.070 1207.910 ;
        RECT 0.580 1205.390 1075.680 1207.090 ;
        RECT 1.090 1204.570 1075.070 1205.390 ;
        RECT 0.580 1202.870 1075.680 1204.570 ;
        RECT 1.090 1202.050 1075.070 1202.870 ;
        RECT 0.580 1200.350 1075.680 1202.050 ;
        RECT 1.090 1199.530 1075.070 1200.350 ;
        RECT 0.580 1197.830 1075.680 1199.530 ;
        RECT 1.090 1197.010 1075.070 1197.830 ;
        RECT 0.580 1195.310 1075.680 1197.010 ;
        RECT 1.090 1194.490 1075.070 1195.310 ;
        RECT 0.580 1192.790 1075.680 1194.490 ;
        RECT 1.090 1191.970 1075.070 1192.790 ;
        RECT 0.580 1190.270 1075.680 1191.970 ;
        RECT 1.090 1189.450 1075.070 1190.270 ;
        RECT 0.580 1187.750 1075.680 1189.450 ;
        RECT 1.090 1186.930 1075.070 1187.750 ;
        RECT 0.580 1185.230 1075.680 1186.930 ;
        RECT 1.090 1184.410 1075.070 1185.230 ;
        RECT 0.580 1182.710 1075.680 1184.410 ;
        RECT 1.090 1181.890 1075.070 1182.710 ;
        RECT 0.580 1180.190 1075.680 1181.890 ;
        RECT 1.090 1179.370 1075.070 1180.190 ;
        RECT 0.580 1177.670 1075.680 1179.370 ;
        RECT 1.090 1176.850 1075.070 1177.670 ;
        RECT 0.580 1175.150 1075.680 1176.850 ;
        RECT 1.090 1174.330 1075.070 1175.150 ;
        RECT 0.580 1172.630 1075.680 1174.330 ;
        RECT 1.090 1171.810 1075.070 1172.630 ;
        RECT 0.580 1170.110 1075.680 1171.810 ;
        RECT 1.090 1169.290 1075.070 1170.110 ;
        RECT 0.580 1167.590 1075.680 1169.290 ;
        RECT 1.090 1166.770 1075.070 1167.590 ;
        RECT 0.580 1165.070 1075.680 1166.770 ;
        RECT 1.090 1164.250 1075.070 1165.070 ;
        RECT 0.580 1162.550 1075.680 1164.250 ;
        RECT 1.090 1161.730 1075.070 1162.550 ;
        RECT 0.580 1160.030 1075.680 1161.730 ;
        RECT 1.090 1159.210 1075.070 1160.030 ;
        RECT 0.580 1157.510 1075.680 1159.210 ;
        RECT 1.090 1156.690 1075.090 1157.510 ;
        RECT 0.580 1154.990 1075.680 1156.690 ;
        RECT 1.090 1154.170 1075.070 1154.990 ;
        RECT 0.580 1152.470 1075.680 1154.170 ;
        RECT 1.090 1151.650 1075.070 1152.470 ;
        RECT 0.580 1149.950 1075.680 1151.650 ;
        RECT 1.090 1149.130 1075.070 1149.950 ;
        RECT 0.580 1147.430 1075.680 1149.130 ;
        RECT 1.090 1146.610 1075.070 1147.430 ;
        RECT 0.580 1118.870 1075.680 1146.610 ;
        RECT 1.090 1118.050 1075.680 1118.870 ;
        RECT 0.580 1116.350 1075.680 1118.050 ;
        RECT 1.090 1115.530 1075.680 1116.350 ;
        RECT 0.580 1113.830 1075.680 1115.530 ;
        RECT 1.090 1113.010 1075.680 1113.830 ;
        RECT 0.580 1111.310 1075.680 1113.010 ;
        RECT 1.090 1110.490 1075.680 1111.310 ;
        RECT 0.580 1108.790 1075.680 1110.490 ;
        RECT 1.090 1107.970 1075.680 1108.790 ;
        RECT 0.580 1106.270 1075.680 1107.970 ;
        RECT 1.090 1105.450 1075.680 1106.270 ;
        RECT 0.580 1103.750 1075.680 1105.450 ;
        RECT 1.090 1102.930 1075.680 1103.750 ;
        RECT 0.580 1101.230 1075.680 1102.930 ;
        RECT 1.090 1100.410 1075.680 1101.230 ;
        RECT 0.580 1098.710 1075.680 1100.410 ;
        RECT 1.090 1097.890 1075.680 1098.710 ;
        RECT 0.580 1096.190 1075.680 1097.890 ;
        RECT 1.090 1095.370 1075.680 1096.190 ;
        RECT 0.580 1093.670 1075.680 1095.370 ;
        RECT 1.090 1092.850 1075.680 1093.670 ;
        RECT 0.580 1091.150 1075.680 1092.850 ;
        RECT 1.090 1090.330 1075.680 1091.150 ;
        RECT 0.580 1088.630 1075.680 1090.330 ;
        RECT 1.090 1087.810 1075.680 1088.630 ;
        RECT 0.580 1086.110 1075.680 1087.810 ;
        RECT 1.090 1085.290 1075.680 1086.110 ;
        RECT 0.580 1083.590 1075.680 1085.290 ;
        RECT 1.090 1082.770 1075.680 1083.590 ;
        RECT 0.580 1081.070 1075.680 1082.770 ;
        RECT 1.090 1080.250 1075.680 1081.070 ;
        RECT 0.580 1078.550 1075.680 1080.250 ;
        RECT 1.090 1077.730 1075.680 1078.550 ;
        RECT 0.580 1076.030 1075.680 1077.730 ;
        RECT 1.090 1075.210 1075.680 1076.030 ;
        RECT 0.580 1073.510 1075.680 1075.210 ;
        RECT 1.090 1072.690 1075.680 1073.510 ;
        RECT 0.580 1070.990 1075.680 1072.690 ;
        RECT 1.090 1070.170 1075.680 1070.990 ;
        RECT 0.580 1068.470 1075.680 1070.170 ;
        RECT 1.090 1067.650 1075.680 1068.470 ;
        RECT 0.580 1065.950 1075.680 1067.650 ;
        RECT 1.090 1065.130 1075.680 1065.950 ;
        RECT 0.580 1063.430 1075.680 1065.130 ;
        RECT 1.090 1062.610 1075.680 1063.430 ;
        RECT 0.580 1060.910 1075.680 1062.610 ;
        RECT 1.090 1060.090 1075.680 1060.910 ;
        RECT 0.580 1058.390 1075.680 1060.090 ;
        RECT 1.090 1057.570 1075.680 1058.390 ;
        RECT 0.580 1055.870 1075.680 1057.570 ;
        RECT 1.090 1055.050 1075.680 1055.870 ;
        RECT 0.580 1053.350 1075.680 1055.050 ;
        RECT 1.090 1052.530 1075.680 1053.350 ;
        RECT 0.580 1050.830 1075.680 1052.530 ;
        RECT 1.070 1050.010 1075.680 1050.830 ;
        RECT 0.580 1048.310 1075.680 1050.010 ;
        RECT 1.090 1047.490 1075.680 1048.310 ;
        RECT 0.580 1045.790 1075.680 1047.490 ;
        RECT 1.090 1044.970 1075.680 1045.790 ;
        RECT 0.580 1043.270 1075.680 1044.970 ;
        RECT 1.090 1042.450 1075.680 1043.270 ;
        RECT 0.580 1040.750 1075.680 1042.450 ;
        RECT 1.090 1039.930 1075.680 1040.750 ;
        RECT 0.580 1038.230 1075.680 1039.930 ;
        RECT 1.070 1037.410 1075.090 1038.230 ;
        RECT 0.580 1035.710 1075.680 1037.410 ;
        RECT 1.090 1034.890 1075.070 1035.710 ;
        RECT 0.580 1033.190 1075.680 1034.890 ;
        RECT 1.090 1032.370 1075.070 1033.190 ;
        RECT 0.580 1030.670 1075.680 1032.370 ;
        RECT 1.090 1029.850 1075.070 1030.670 ;
        RECT 0.580 1028.150 1075.680 1029.850 ;
        RECT 1.090 1027.330 1075.070 1028.150 ;
        RECT 0.580 1025.630 1075.680 1027.330 ;
        RECT 1.090 1024.810 1075.070 1025.630 ;
        RECT 0.580 1023.110 1075.680 1024.810 ;
        RECT 1.090 1022.290 1075.070 1023.110 ;
        RECT 0.580 1020.590 1075.680 1022.290 ;
        RECT 1.090 1019.770 1075.070 1020.590 ;
        RECT 0.580 1018.070 1075.680 1019.770 ;
        RECT 1.090 1017.250 1075.070 1018.070 ;
        RECT 0.580 1015.550 1075.680 1017.250 ;
        RECT 1.090 1014.730 1075.070 1015.550 ;
        RECT 0.580 1013.030 1075.680 1014.730 ;
        RECT 1.090 1012.210 1075.070 1013.030 ;
        RECT 0.580 1010.510 1075.680 1012.210 ;
        RECT 1.090 1009.690 1075.070 1010.510 ;
        RECT 0.580 1007.990 1075.680 1009.690 ;
        RECT 1.070 1007.170 1075.070 1007.990 ;
        RECT 0.580 1005.470 1075.680 1007.170 ;
        RECT 1.090 1004.650 1075.070 1005.470 ;
        RECT 0.580 1002.950 1075.680 1004.650 ;
        RECT 1.090 1002.130 1075.070 1002.950 ;
        RECT 0.580 1000.430 1075.680 1002.130 ;
        RECT 1.090 999.610 1075.070 1000.430 ;
        RECT 0.580 997.910 1075.680 999.610 ;
        RECT 1.090 997.090 1075.070 997.910 ;
        RECT 0.580 995.390 1075.680 997.090 ;
        RECT 1.090 994.570 1075.070 995.390 ;
        RECT 0.580 992.870 1075.680 994.570 ;
        RECT 1.090 992.050 1075.070 992.870 ;
        RECT 0.580 990.350 1075.680 992.050 ;
        RECT 1.090 989.530 1075.070 990.350 ;
        RECT 0.580 987.830 1075.680 989.530 ;
        RECT 1.090 987.010 1075.070 987.830 ;
        RECT 0.580 985.310 1075.680 987.010 ;
        RECT 1.090 984.490 1075.070 985.310 ;
        RECT 0.580 982.790 1075.680 984.490 ;
        RECT 1.090 981.970 1075.070 982.790 ;
        RECT 0.580 980.270 1075.680 981.970 ;
        RECT 1.090 979.450 1075.070 980.270 ;
        RECT 0.580 977.750 1075.680 979.450 ;
        RECT 1.090 976.930 1075.070 977.750 ;
        RECT 0.580 975.230 1075.680 976.930 ;
        RECT 1.090 974.410 1075.070 975.230 ;
        RECT 0.580 972.710 1075.680 974.410 ;
        RECT 1.090 971.890 1075.070 972.710 ;
        RECT 0.580 970.190 1075.680 971.890 ;
        RECT 1.090 969.370 1075.070 970.190 ;
        RECT 0.580 967.670 1075.680 969.370 ;
        RECT 1.090 966.850 1075.070 967.670 ;
        RECT 0.580 965.150 1075.680 966.850 ;
        RECT 1.090 964.330 1075.070 965.150 ;
        RECT 0.580 962.630 1075.680 964.330 ;
        RECT 1.090 961.810 1075.070 962.630 ;
        RECT 0.580 960.110 1075.680 961.810 ;
        RECT 1.090 959.290 1075.070 960.110 ;
        RECT 0.580 957.590 1075.680 959.290 ;
        RECT 1.090 956.770 1075.070 957.590 ;
        RECT 0.580 955.070 1075.680 956.770 ;
        RECT 1.090 954.250 1075.070 955.070 ;
        RECT 0.580 952.550 1075.680 954.250 ;
        RECT 1.090 951.730 1075.070 952.550 ;
        RECT 0.580 950.030 1075.680 951.730 ;
        RECT 1.090 949.210 1075.070 950.030 ;
        RECT 0.580 947.510 1075.680 949.210 ;
        RECT 1.090 946.690 1075.070 947.510 ;
        RECT 0.580 944.990 1075.680 946.690 ;
        RECT 1.090 944.170 1075.070 944.990 ;
        RECT 0.580 942.470 1075.680 944.170 ;
        RECT 1.090 941.650 1075.090 942.470 ;
        RECT 0.580 939.950 1075.680 941.650 ;
        RECT 1.090 939.130 1075.070 939.950 ;
        RECT 0.580 937.430 1075.680 939.130 ;
        RECT 1.090 936.610 1075.070 937.430 ;
        RECT 0.580 934.910 1075.680 936.610 ;
        RECT 1.090 934.090 1075.070 934.910 ;
        RECT 0.580 932.390 1075.680 934.090 ;
        RECT 1.090 931.570 1075.070 932.390 ;
        RECT 0.580 903.830 1075.680 931.570 ;
        RECT 1.090 903.010 1075.680 903.830 ;
        RECT 0.580 901.310 1075.680 903.010 ;
        RECT 1.090 900.490 1075.680 901.310 ;
        RECT 0.580 898.790 1075.680 900.490 ;
        RECT 1.090 897.970 1075.680 898.790 ;
        RECT 0.580 896.270 1075.680 897.970 ;
        RECT 1.090 895.450 1075.680 896.270 ;
        RECT 0.580 893.750 1075.680 895.450 ;
        RECT 1.090 892.930 1075.680 893.750 ;
        RECT 0.580 891.230 1075.680 892.930 ;
        RECT 1.090 890.410 1075.680 891.230 ;
        RECT 0.580 888.710 1075.680 890.410 ;
        RECT 1.090 887.890 1075.680 888.710 ;
        RECT 0.580 886.190 1075.680 887.890 ;
        RECT 1.090 885.370 1075.680 886.190 ;
        RECT 0.580 883.670 1075.680 885.370 ;
        RECT 1.090 882.850 1075.680 883.670 ;
        RECT 0.580 881.150 1075.680 882.850 ;
        RECT 1.090 880.330 1075.680 881.150 ;
        RECT 0.580 878.630 1075.680 880.330 ;
        RECT 1.090 877.810 1075.680 878.630 ;
        RECT 0.580 876.110 1075.680 877.810 ;
        RECT 1.090 875.290 1075.680 876.110 ;
        RECT 0.580 873.590 1075.680 875.290 ;
        RECT 1.090 872.770 1075.680 873.590 ;
        RECT 0.580 871.070 1075.680 872.770 ;
        RECT 1.090 870.250 1075.680 871.070 ;
        RECT 0.580 868.550 1075.680 870.250 ;
        RECT 1.090 867.730 1075.680 868.550 ;
        RECT 0.580 866.030 1075.680 867.730 ;
        RECT 1.090 865.210 1075.680 866.030 ;
        RECT 0.580 863.510 1075.680 865.210 ;
        RECT 1.090 862.690 1075.680 863.510 ;
        RECT 0.580 860.990 1075.680 862.690 ;
        RECT 1.090 860.170 1075.680 860.990 ;
        RECT 0.580 858.470 1075.680 860.170 ;
        RECT 1.090 857.650 1075.680 858.470 ;
        RECT 0.580 855.950 1075.680 857.650 ;
        RECT 1.090 855.130 1075.680 855.950 ;
        RECT 0.580 853.430 1075.680 855.130 ;
        RECT 1.090 852.610 1075.680 853.430 ;
        RECT 0.580 850.910 1075.680 852.610 ;
        RECT 1.090 850.090 1075.680 850.910 ;
        RECT 0.580 848.390 1075.680 850.090 ;
        RECT 1.090 847.570 1075.680 848.390 ;
        RECT 0.580 845.870 1075.680 847.570 ;
        RECT 1.090 845.050 1075.680 845.870 ;
        RECT 0.580 843.350 1075.680 845.050 ;
        RECT 1.090 842.530 1075.680 843.350 ;
        RECT 0.580 840.830 1075.680 842.530 ;
        RECT 1.090 840.010 1075.680 840.830 ;
        RECT 0.580 838.310 1075.680 840.010 ;
        RECT 1.090 837.490 1075.680 838.310 ;
        RECT 0.580 835.790 1075.680 837.490 ;
        RECT 1.070 834.970 1075.680 835.790 ;
        RECT 0.580 833.270 1075.680 834.970 ;
        RECT 1.090 832.450 1075.680 833.270 ;
        RECT 0.580 830.750 1075.680 832.450 ;
        RECT 1.090 829.930 1075.680 830.750 ;
        RECT 0.580 828.230 1075.680 829.930 ;
        RECT 1.090 827.410 1075.680 828.230 ;
        RECT 0.580 825.710 1075.680 827.410 ;
        RECT 1.090 824.890 1075.680 825.710 ;
        RECT 0.580 823.190 1075.680 824.890 ;
        RECT 1.070 822.370 1075.090 823.190 ;
        RECT 0.580 820.670 1075.680 822.370 ;
        RECT 1.090 819.850 1075.070 820.670 ;
        RECT 0.580 818.150 1075.680 819.850 ;
        RECT 1.090 817.330 1075.070 818.150 ;
        RECT 0.580 815.630 1075.680 817.330 ;
        RECT 1.090 814.810 1075.070 815.630 ;
        RECT 0.580 813.110 1075.680 814.810 ;
        RECT 1.090 812.290 1075.070 813.110 ;
        RECT 0.580 810.590 1075.680 812.290 ;
        RECT 1.090 809.770 1075.070 810.590 ;
        RECT 0.580 808.070 1075.680 809.770 ;
        RECT 1.090 807.250 1075.070 808.070 ;
        RECT 0.580 805.550 1075.680 807.250 ;
        RECT 1.090 804.730 1075.070 805.550 ;
        RECT 0.580 803.030 1075.680 804.730 ;
        RECT 1.090 802.210 1075.070 803.030 ;
        RECT 0.580 800.510 1075.680 802.210 ;
        RECT 1.090 799.690 1075.070 800.510 ;
        RECT 0.580 797.990 1075.680 799.690 ;
        RECT 1.090 797.170 1075.070 797.990 ;
        RECT 0.580 795.470 1075.680 797.170 ;
        RECT 1.090 794.650 1075.070 795.470 ;
        RECT 0.580 792.950 1075.680 794.650 ;
        RECT 1.070 792.130 1075.070 792.950 ;
        RECT 0.580 790.430 1075.680 792.130 ;
        RECT 1.090 789.610 1075.070 790.430 ;
        RECT 0.580 787.910 1075.680 789.610 ;
        RECT 1.090 787.090 1075.070 787.910 ;
        RECT 0.580 785.390 1075.680 787.090 ;
        RECT 1.090 784.570 1075.070 785.390 ;
        RECT 0.580 782.870 1075.680 784.570 ;
        RECT 1.090 782.050 1075.070 782.870 ;
        RECT 0.580 780.350 1075.680 782.050 ;
        RECT 1.090 779.530 1075.070 780.350 ;
        RECT 0.580 777.830 1075.680 779.530 ;
        RECT 1.090 777.010 1075.070 777.830 ;
        RECT 0.580 775.310 1075.680 777.010 ;
        RECT 1.090 774.490 1075.070 775.310 ;
        RECT 0.580 772.790 1075.680 774.490 ;
        RECT 1.090 771.970 1075.070 772.790 ;
        RECT 0.580 770.270 1075.680 771.970 ;
        RECT 1.090 769.450 1075.070 770.270 ;
        RECT 0.580 767.750 1075.680 769.450 ;
        RECT 1.090 766.930 1075.070 767.750 ;
        RECT 0.580 765.230 1075.680 766.930 ;
        RECT 1.090 764.410 1075.070 765.230 ;
        RECT 0.580 762.710 1075.680 764.410 ;
        RECT 1.090 761.890 1075.070 762.710 ;
        RECT 0.580 760.190 1075.680 761.890 ;
        RECT 1.090 759.370 1075.070 760.190 ;
        RECT 0.580 757.670 1075.680 759.370 ;
        RECT 1.090 756.850 1075.070 757.670 ;
        RECT 0.580 755.150 1075.680 756.850 ;
        RECT 1.090 754.330 1075.070 755.150 ;
        RECT 0.580 752.630 1075.680 754.330 ;
        RECT 1.090 751.810 1075.070 752.630 ;
        RECT 0.580 750.110 1075.680 751.810 ;
        RECT 1.090 749.290 1075.070 750.110 ;
        RECT 0.580 747.590 1075.680 749.290 ;
        RECT 1.090 746.770 1075.070 747.590 ;
        RECT 0.580 745.070 1075.680 746.770 ;
        RECT 1.090 744.250 1075.070 745.070 ;
        RECT 0.580 742.550 1075.680 744.250 ;
        RECT 1.090 741.730 1075.070 742.550 ;
        RECT 0.580 740.030 1075.680 741.730 ;
        RECT 1.090 739.210 1075.070 740.030 ;
        RECT 0.580 737.510 1075.680 739.210 ;
        RECT 1.090 736.690 1075.070 737.510 ;
        RECT 0.580 734.990 1075.680 736.690 ;
        RECT 1.090 734.170 1075.070 734.990 ;
        RECT 0.580 732.470 1075.680 734.170 ;
        RECT 1.090 731.650 1075.070 732.470 ;
        RECT 0.580 729.950 1075.680 731.650 ;
        RECT 1.090 729.130 1075.070 729.950 ;
        RECT 0.580 727.430 1075.680 729.130 ;
        RECT 1.090 726.610 1075.090 727.430 ;
        RECT 0.580 724.910 1075.680 726.610 ;
        RECT 1.090 724.090 1075.070 724.910 ;
        RECT 0.580 722.390 1075.680 724.090 ;
        RECT 1.090 721.570 1075.070 722.390 ;
        RECT 0.580 719.870 1075.680 721.570 ;
        RECT 1.090 719.050 1075.070 719.870 ;
        RECT 0.580 717.350 1075.680 719.050 ;
        RECT 1.090 716.530 1075.070 717.350 ;
        RECT 0.580 688.790 1075.680 716.530 ;
        RECT 1.090 687.970 1075.680 688.790 ;
        RECT 0.580 686.270 1075.680 687.970 ;
        RECT 1.090 685.450 1075.680 686.270 ;
        RECT 0.580 683.750 1075.680 685.450 ;
        RECT 1.090 682.930 1075.680 683.750 ;
        RECT 0.580 681.230 1075.680 682.930 ;
        RECT 1.090 680.410 1075.680 681.230 ;
        RECT 0.580 678.710 1075.680 680.410 ;
        RECT 1.090 677.890 1075.680 678.710 ;
        RECT 0.580 676.190 1075.680 677.890 ;
        RECT 1.090 675.370 1075.680 676.190 ;
        RECT 0.580 673.670 1075.680 675.370 ;
        RECT 1.090 672.850 1075.680 673.670 ;
        RECT 0.580 671.150 1075.680 672.850 ;
        RECT 1.090 670.330 1075.680 671.150 ;
        RECT 0.580 668.630 1075.680 670.330 ;
        RECT 1.090 667.810 1075.680 668.630 ;
        RECT 0.580 666.110 1075.680 667.810 ;
        RECT 1.090 665.290 1075.680 666.110 ;
        RECT 0.580 663.590 1075.680 665.290 ;
        RECT 1.090 662.770 1075.680 663.590 ;
        RECT 0.580 661.070 1075.680 662.770 ;
        RECT 1.090 660.250 1075.680 661.070 ;
        RECT 0.580 658.550 1075.680 660.250 ;
        RECT 1.090 657.730 1075.680 658.550 ;
        RECT 0.580 656.030 1075.680 657.730 ;
        RECT 1.090 655.210 1075.680 656.030 ;
        RECT 0.580 653.510 1075.680 655.210 ;
        RECT 1.090 652.690 1075.680 653.510 ;
        RECT 0.580 650.990 1075.680 652.690 ;
        RECT 1.090 650.170 1075.680 650.990 ;
        RECT 0.580 648.470 1075.680 650.170 ;
        RECT 1.090 647.650 1075.680 648.470 ;
        RECT 0.580 645.950 1075.680 647.650 ;
        RECT 1.090 645.130 1075.680 645.950 ;
        RECT 0.580 643.430 1075.680 645.130 ;
        RECT 1.090 642.610 1075.680 643.430 ;
        RECT 0.580 640.910 1075.680 642.610 ;
        RECT 1.090 640.090 1075.680 640.910 ;
        RECT 0.580 638.390 1075.680 640.090 ;
        RECT 1.090 637.570 1075.680 638.390 ;
        RECT 0.580 635.870 1075.680 637.570 ;
        RECT 1.090 635.050 1075.680 635.870 ;
        RECT 0.580 633.350 1075.680 635.050 ;
        RECT 1.090 632.530 1075.680 633.350 ;
        RECT 0.580 630.830 1075.680 632.530 ;
        RECT 1.090 630.010 1075.680 630.830 ;
        RECT 0.580 628.310 1075.680 630.010 ;
        RECT 1.090 627.490 1075.680 628.310 ;
        RECT 0.580 625.790 1075.680 627.490 ;
        RECT 1.090 624.970 1075.680 625.790 ;
        RECT 0.580 623.270 1075.680 624.970 ;
        RECT 1.090 622.450 1075.680 623.270 ;
        RECT 0.580 620.750 1075.680 622.450 ;
        RECT 1.070 619.930 1075.680 620.750 ;
        RECT 0.580 618.230 1075.680 619.930 ;
        RECT 1.090 617.410 1075.680 618.230 ;
        RECT 0.580 615.710 1075.680 617.410 ;
        RECT 1.090 614.890 1075.680 615.710 ;
        RECT 0.580 613.190 1075.680 614.890 ;
        RECT 1.090 612.370 1075.680 613.190 ;
        RECT 0.580 610.670 1075.680 612.370 ;
        RECT 1.090 609.850 1075.680 610.670 ;
        RECT 0.580 608.150 1075.680 609.850 ;
        RECT 1.070 607.330 1075.090 608.150 ;
        RECT 0.580 605.630 1075.680 607.330 ;
        RECT 1.090 604.810 1075.070 605.630 ;
        RECT 0.580 603.110 1075.680 604.810 ;
        RECT 1.090 602.290 1075.070 603.110 ;
        RECT 0.580 600.590 1075.680 602.290 ;
        RECT 1.090 599.770 1075.070 600.590 ;
        RECT 0.580 598.070 1075.680 599.770 ;
        RECT 1.090 597.250 1075.070 598.070 ;
        RECT 0.580 595.550 1075.680 597.250 ;
        RECT 1.090 594.730 1075.070 595.550 ;
        RECT 0.580 593.030 1075.680 594.730 ;
        RECT 1.090 592.210 1075.070 593.030 ;
        RECT 0.580 590.510 1075.680 592.210 ;
        RECT 1.090 589.690 1075.070 590.510 ;
        RECT 0.580 587.990 1075.680 589.690 ;
        RECT 1.090 587.170 1075.070 587.990 ;
        RECT 0.580 585.470 1075.680 587.170 ;
        RECT 1.090 584.650 1075.070 585.470 ;
        RECT 0.580 582.950 1075.680 584.650 ;
        RECT 1.090 582.130 1075.070 582.950 ;
        RECT 0.580 580.430 1075.680 582.130 ;
        RECT 1.090 579.610 1075.070 580.430 ;
        RECT 0.580 577.910 1075.680 579.610 ;
        RECT 1.070 577.090 1075.070 577.910 ;
        RECT 0.580 575.390 1075.680 577.090 ;
        RECT 1.090 574.570 1075.070 575.390 ;
        RECT 0.580 572.870 1075.680 574.570 ;
        RECT 1.090 572.050 1075.070 572.870 ;
        RECT 0.580 570.350 1075.680 572.050 ;
        RECT 1.090 569.530 1075.070 570.350 ;
        RECT 0.580 567.830 1075.680 569.530 ;
        RECT 1.090 567.010 1075.070 567.830 ;
        RECT 0.580 565.310 1075.680 567.010 ;
        RECT 1.090 564.490 1075.070 565.310 ;
        RECT 0.580 562.790 1075.680 564.490 ;
        RECT 1.090 561.970 1075.070 562.790 ;
        RECT 0.580 560.270 1075.680 561.970 ;
        RECT 1.090 559.450 1075.070 560.270 ;
        RECT 0.580 557.750 1075.680 559.450 ;
        RECT 1.090 556.930 1075.070 557.750 ;
        RECT 0.580 555.230 1075.680 556.930 ;
        RECT 1.090 554.410 1075.070 555.230 ;
        RECT 0.580 552.710 1075.680 554.410 ;
        RECT 1.090 551.890 1075.070 552.710 ;
        RECT 0.580 550.190 1075.680 551.890 ;
        RECT 1.090 549.370 1075.070 550.190 ;
        RECT 0.580 547.670 1075.680 549.370 ;
        RECT 1.090 546.850 1075.070 547.670 ;
        RECT 0.580 545.150 1075.680 546.850 ;
        RECT 1.090 544.330 1075.070 545.150 ;
        RECT 0.580 542.630 1075.680 544.330 ;
        RECT 1.090 541.810 1075.070 542.630 ;
        RECT 0.580 540.110 1075.680 541.810 ;
        RECT 1.090 539.290 1075.070 540.110 ;
        RECT 0.580 537.590 1075.680 539.290 ;
        RECT 1.090 536.770 1075.070 537.590 ;
        RECT 0.580 535.070 1075.680 536.770 ;
        RECT 1.090 534.250 1075.070 535.070 ;
        RECT 0.580 532.550 1075.680 534.250 ;
        RECT 1.090 531.730 1075.070 532.550 ;
        RECT 0.580 530.030 1075.680 531.730 ;
        RECT 1.090 529.210 1075.070 530.030 ;
        RECT 0.580 527.510 1075.680 529.210 ;
        RECT 1.090 526.690 1075.070 527.510 ;
        RECT 0.580 524.990 1075.680 526.690 ;
        RECT 1.090 524.170 1075.070 524.990 ;
        RECT 0.580 522.470 1075.680 524.170 ;
        RECT 1.090 521.650 1075.070 522.470 ;
        RECT 0.580 519.950 1075.680 521.650 ;
        RECT 1.090 519.130 1075.070 519.950 ;
        RECT 0.580 517.430 1075.680 519.130 ;
        RECT 1.090 516.610 1075.070 517.430 ;
        RECT 0.580 514.910 1075.680 516.610 ;
        RECT 1.090 514.090 1075.070 514.910 ;
        RECT 0.580 512.390 1075.680 514.090 ;
        RECT 1.090 511.570 1075.090 512.390 ;
        RECT 0.580 509.870 1075.680 511.570 ;
        RECT 1.090 509.050 1075.070 509.870 ;
        RECT 0.580 507.350 1075.680 509.050 ;
        RECT 1.090 506.530 1075.070 507.350 ;
        RECT 0.580 504.830 1075.680 506.530 ;
        RECT 1.090 504.010 1075.070 504.830 ;
        RECT 0.580 502.310 1075.680 504.010 ;
        RECT 1.090 501.490 1075.070 502.310 ;
        RECT 0.580 473.750 1075.680 501.490 ;
        RECT 1.090 472.930 1075.680 473.750 ;
        RECT 0.580 471.230 1075.680 472.930 ;
        RECT 1.090 470.410 1075.680 471.230 ;
        RECT 0.580 468.710 1075.680 470.410 ;
        RECT 1.090 467.890 1075.680 468.710 ;
        RECT 0.580 466.190 1075.680 467.890 ;
        RECT 1.090 465.370 1075.680 466.190 ;
        RECT 0.580 463.670 1075.680 465.370 ;
        RECT 1.090 462.850 1075.680 463.670 ;
        RECT 0.580 461.150 1075.680 462.850 ;
        RECT 1.090 460.330 1075.680 461.150 ;
        RECT 0.580 458.630 1075.680 460.330 ;
        RECT 1.090 457.810 1075.680 458.630 ;
        RECT 0.580 456.110 1075.680 457.810 ;
        RECT 1.090 455.290 1075.680 456.110 ;
        RECT 0.580 453.590 1075.680 455.290 ;
        RECT 1.090 452.770 1075.680 453.590 ;
        RECT 0.580 451.070 1075.680 452.770 ;
        RECT 1.090 450.250 1075.680 451.070 ;
        RECT 0.580 448.550 1075.680 450.250 ;
        RECT 1.090 447.730 1075.680 448.550 ;
        RECT 0.580 446.030 1075.680 447.730 ;
        RECT 1.090 445.210 1075.680 446.030 ;
        RECT 0.580 443.510 1075.680 445.210 ;
        RECT 1.090 442.690 1075.680 443.510 ;
        RECT 0.580 440.990 1075.680 442.690 ;
        RECT 1.090 440.170 1075.680 440.990 ;
        RECT 0.580 438.470 1075.680 440.170 ;
        RECT 1.090 437.650 1075.680 438.470 ;
        RECT 0.580 435.950 1075.680 437.650 ;
        RECT 1.090 435.130 1075.680 435.950 ;
        RECT 0.580 433.430 1075.680 435.130 ;
        RECT 1.090 432.610 1075.680 433.430 ;
        RECT 0.580 430.910 1075.680 432.610 ;
        RECT 1.090 430.090 1075.680 430.910 ;
        RECT 0.580 428.390 1075.680 430.090 ;
        RECT 1.090 427.570 1075.680 428.390 ;
        RECT 0.580 425.870 1075.680 427.570 ;
        RECT 1.090 425.050 1075.680 425.870 ;
        RECT 0.580 423.350 1075.680 425.050 ;
        RECT 1.090 422.530 1075.680 423.350 ;
        RECT 0.580 420.830 1075.680 422.530 ;
        RECT 1.090 420.010 1075.680 420.830 ;
        RECT 0.580 418.310 1075.680 420.010 ;
        RECT 1.090 417.490 1075.680 418.310 ;
        RECT 0.580 415.790 1075.680 417.490 ;
        RECT 1.090 414.970 1075.680 415.790 ;
        RECT 0.580 413.270 1075.680 414.970 ;
        RECT 1.090 412.450 1075.680 413.270 ;
        RECT 0.580 410.750 1075.680 412.450 ;
        RECT 1.090 409.930 1075.680 410.750 ;
        RECT 0.580 408.230 1075.680 409.930 ;
        RECT 1.090 407.410 1075.680 408.230 ;
        RECT 0.580 405.710 1075.680 407.410 ;
        RECT 1.070 404.890 1075.680 405.710 ;
        RECT 0.580 403.190 1075.680 404.890 ;
        RECT 1.090 402.370 1075.680 403.190 ;
        RECT 0.580 400.670 1075.680 402.370 ;
        RECT 1.090 399.850 1075.680 400.670 ;
        RECT 0.580 398.150 1075.680 399.850 ;
        RECT 1.090 397.330 1075.680 398.150 ;
        RECT 0.580 395.630 1075.680 397.330 ;
        RECT 1.090 394.810 1075.680 395.630 ;
        RECT 0.580 393.110 1075.680 394.810 ;
        RECT 1.070 392.290 1075.090 393.110 ;
        RECT 0.580 390.590 1075.680 392.290 ;
        RECT 1.090 389.770 1075.070 390.590 ;
        RECT 0.580 388.070 1075.680 389.770 ;
        RECT 1.090 387.250 1075.070 388.070 ;
        RECT 0.580 385.550 1075.680 387.250 ;
        RECT 1.090 384.730 1075.070 385.550 ;
        RECT 0.580 383.030 1075.680 384.730 ;
        RECT 1.090 382.210 1075.070 383.030 ;
        RECT 0.580 380.510 1075.680 382.210 ;
        RECT 1.090 379.690 1075.070 380.510 ;
        RECT 0.580 377.990 1075.680 379.690 ;
        RECT 1.090 377.170 1075.070 377.990 ;
        RECT 0.580 375.470 1075.680 377.170 ;
        RECT 1.090 374.650 1075.070 375.470 ;
        RECT 0.580 372.950 1075.680 374.650 ;
        RECT 1.090 372.130 1075.070 372.950 ;
        RECT 0.580 370.430 1075.680 372.130 ;
        RECT 1.090 369.610 1075.070 370.430 ;
        RECT 0.580 367.910 1075.680 369.610 ;
        RECT 1.090 367.090 1075.070 367.910 ;
        RECT 0.580 365.390 1075.680 367.090 ;
        RECT 1.090 364.570 1075.070 365.390 ;
        RECT 0.580 362.870 1075.680 364.570 ;
        RECT 1.070 362.050 1075.070 362.870 ;
        RECT 0.580 360.350 1075.680 362.050 ;
        RECT 1.090 359.530 1075.070 360.350 ;
        RECT 0.580 357.830 1075.680 359.530 ;
        RECT 1.090 357.010 1075.070 357.830 ;
        RECT 0.580 355.310 1075.680 357.010 ;
        RECT 1.090 354.490 1075.070 355.310 ;
        RECT 0.580 352.790 1075.680 354.490 ;
        RECT 1.090 351.970 1075.070 352.790 ;
        RECT 0.580 350.270 1075.680 351.970 ;
        RECT 1.090 349.450 1075.070 350.270 ;
        RECT 0.580 347.750 1075.680 349.450 ;
        RECT 1.090 346.930 1075.070 347.750 ;
        RECT 0.580 345.230 1075.680 346.930 ;
        RECT 1.090 344.410 1075.070 345.230 ;
        RECT 0.580 342.710 1075.680 344.410 ;
        RECT 1.090 341.890 1075.070 342.710 ;
        RECT 0.580 340.190 1075.680 341.890 ;
        RECT 1.090 339.370 1075.070 340.190 ;
        RECT 0.580 337.670 1075.680 339.370 ;
        RECT 1.090 336.850 1075.070 337.670 ;
        RECT 0.580 335.150 1075.680 336.850 ;
        RECT 1.090 334.330 1075.070 335.150 ;
        RECT 0.580 332.630 1075.680 334.330 ;
        RECT 1.090 331.810 1075.070 332.630 ;
        RECT 0.580 330.110 1075.680 331.810 ;
        RECT 1.090 329.290 1075.070 330.110 ;
        RECT 0.580 327.590 1075.680 329.290 ;
        RECT 1.090 326.770 1075.070 327.590 ;
        RECT 0.580 325.070 1075.680 326.770 ;
        RECT 1.090 324.250 1075.070 325.070 ;
        RECT 0.580 322.550 1075.680 324.250 ;
        RECT 1.090 321.730 1075.070 322.550 ;
        RECT 0.580 320.030 1075.680 321.730 ;
        RECT 1.090 319.210 1075.070 320.030 ;
        RECT 0.580 317.510 1075.680 319.210 ;
        RECT 1.090 316.690 1075.070 317.510 ;
        RECT 0.580 314.990 1075.680 316.690 ;
        RECT 1.090 314.170 1075.070 314.990 ;
        RECT 0.580 312.470 1075.680 314.170 ;
        RECT 1.090 311.650 1075.070 312.470 ;
        RECT 0.580 309.950 1075.680 311.650 ;
        RECT 1.090 309.130 1075.070 309.950 ;
        RECT 0.580 307.430 1075.680 309.130 ;
        RECT 1.090 306.610 1075.070 307.430 ;
        RECT 0.580 304.910 1075.680 306.610 ;
        RECT 1.090 304.090 1075.070 304.910 ;
        RECT 0.580 302.390 1075.680 304.090 ;
        RECT 1.090 301.570 1075.070 302.390 ;
        RECT 0.580 299.870 1075.680 301.570 ;
        RECT 1.090 299.050 1075.070 299.870 ;
        RECT 0.580 297.350 1075.680 299.050 ;
        RECT 1.090 296.530 1075.090 297.350 ;
        RECT 0.580 294.830 1075.680 296.530 ;
        RECT 1.090 294.010 1075.070 294.830 ;
        RECT 0.580 292.310 1075.680 294.010 ;
        RECT 1.090 291.490 1075.070 292.310 ;
        RECT 0.580 289.790 1075.680 291.490 ;
        RECT 1.090 288.970 1075.070 289.790 ;
        RECT 0.580 287.270 1075.680 288.970 ;
        RECT 1.090 286.450 1075.070 287.270 ;
        RECT 0.580 258.710 1075.680 286.450 ;
        RECT 1.090 257.890 1075.680 258.710 ;
        RECT 0.580 256.190 1075.680 257.890 ;
        RECT 1.090 255.370 1075.680 256.190 ;
        RECT 0.580 253.670 1075.680 255.370 ;
        RECT 1.090 252.850 1075.680 253.670 ;
        RECT 0.580 251.150 1075.680 252.850 ;
        RECT 1.090 250.330 1075.680 251.150 ;
        RECT 0.580 248.630 1075.680 250.330 ;
        RECT 1.090 247.810 1075.680 248.630 ;
        RECT 0.580 246.110 1075.680 247.810 ;
        RECT 1.090 245.290 1075.680 246.110 ;
        RECT 0.580 243.590 1075.680 245.290 ;
        RECT 1.090 242.770 1075.680 243.590 ;
        RECT 0.580 241.070 1075.680 242.770 ;
        RECT 1.090 240.250 1075.680 241.070 ;
        RECT 0.580 238.550 1075.680 240.250 ;
        RECT 1.090 237.730 1075.680 238.550 ;
        RECT 0.580 236.030 1075.680 237.730 ;
        RECT 1.090 235.210 1075.680 236.030 ;
        RECT 0.580 233.510 1075.680 235.210 ;
        RECT 1.090 232.690 1075.680 233.510 ;
        RECT 0.580 230.990 1075.680 232.690 ;
        RECT 1.090 230.170 1075.680 230.990 ;
        RECT 0.580 228.470 1075.680 230.170 ;
        RECT 1.090 227.650 1075.680 228.470 ;
        RECT 0.580 225.950 1075.680 227.650 ;
        RECT 1.090 225.130 1075.680 225.950 ;
        RECT 0.580 223.430 1075.680 225.130 ;
        RECT 1.090 222.610 1075.680 223.430 ;
        RECT 0.580 220.910 1075.680 222.610 ;
        RECT 1.090 220.090 1075.680 220.910 ;
        RECT 0.580 218.390 1075.680 220.090 ;
        RECT 1.090 217.570 1075.680 218.390 ;
        RECT 0.580 215.870 1075.680 217.570 ;
        RECT 1.090 215.050 1075.680 215.870 ;
        RECT 0.580 213.350 1075.680 215.050 ;
        RECT 1.090 212.530 1075.680 213.350 ;
        RECT 0.580 210.830 1075.680 212.530 ;
        RECT 1.090 210.010 1075.680 210.830 ;
        RECT 0.580 208.310 1075.680 210.010 ;
        RECT 1.090 207.490 1075.680 208.310 ;
        RECT 0.580 205.790 1075.680 207.490 ;
        RECT 1.090 204.970 1075.680 205.790 ;
        RECT 0.580 203.270 1075.680 204.970 ;
        RECT 1.090 202.450 1075.680 203.270 ;
        RECT 0.580 200.750 1075.680 202.450 ;
        RECT 1.090 199.930 1075.680 200.750 ;
        RECT 0.580 198.230 1075.680 199.930 ;
        RECT 1.090 197.410 1075.680 198.230 ;
        RECT 0.580 195.710 1075.680 197.410 ;
        RECT 1.090 194.890 1075.680 195.710 ;
        RECT 0.580 193.190 1075.680 194.890 ;
        RECT 1.090 192.370 1075.680 193.190 ;
        RECT 0.580 190.670 1075.680 192.370 ;
        RECT 1.070 189.850 1075.680 190.670 ;
        RECT 0.580 188.150 1075.680 189.850 ;
        RECT 1.090 187.330 1075.680 188.150 ;
        RECT 0.580 185.630 1075.680 187.330 ;
        RECT 1.090 184.810 1075.680 185.630 ;
        RECT 0.580 183.110 1075.680 184.810 ;
        RECT 1.090 182.290 1075.680 183.110 ;
        RECT 0.580 180.590 1075.680 182.290 ;
        RECT 1.090 179.770 1075.680 180.590 ;
        RECT 0.580 178.070 1075.680 179.770 ;
        RECT 1.070 177.250 1075.090 178.070 ;
        RECT 0.580 175.550 1075.680 177.250 ;
        RECT 1.090 174.730 1075.070 175.550 ;
        RECT 0.580 173.030 1075.680 174.730 ;
        RECT 1.090 172.210 1075.070 173.030 ;
        RECT 0.580 170.510 1075.680 172.210 ;
        RECT 1.090 169.690 1075.070 170.510 ;
        RECT 0.580 167.990 1075.680 169.690 ;
        RECT 1.090 167.170 1075.070 167.990 ;
        RECT 0.580 165.470 1075.680 167.170 ;
        RECT 1.090 164.650 1075.070 165.470 ;
        RECT 0.580 162.950 1075.680 164.650 ;
        RECT 1.090 162.130 1075.070 162.950 ;
        RECT 0.580 160.430 1075.680 162.130 ;
        RECT 1.090 159.610 1075.070 160.430 ;
        RECT 0.580 157.910 1075.680 159.610 ;
        RECT 1.090 157.090 1075.070 157.910 ;
        RECT 0.580 155.390 1075.680 157.090 ;
        RECT 1.090 154.570 1075.070 155.390 ;
        RECT 0.580 152.870 1075.680 154.570 ;
        RECT 1.090 152.050 1075.070 152.870 ;
        RECT 0.580 150.350 1075.680 152.050 ;
        RECT 1.090 149.530 1075.070 150.350 ;
        RECT 0.580 147.830 1075.680 149.530 ;
        RECT 1.070 147.010 1075.070 147.830 ;
        RECT 0.580 145.310 1075.680 147.010 ;
        RECT 1.090 144.490 1075.070 145.310 ;
        RECT 0.580 142.790 1075.680 144.490 ;
        RECT 1.090 141.970 1075.070 142.790 ;
        RECT 0.580 140.270 1075.680 141.970 ;
        RECT 1.090 139.450 1075.070 140.270 ;
        RECT 0.580 137.750 1075.680 139.450 ;
        RECT 1.090 136.930 1075.070 137.750 ;
        RECT 0.580 135.230 1075.680 136.930 ;
        RECT 1.090 134.410 1075.070 135.230 ;
        RECT 0.580 132.710 1075.680 134.410 ;
        RECT 1.090 131.890 1075.070 132.710 ;
        RECT 0.580 130.190 1075.680 131.890 ;
        RECT 1.090 129.370 1075.070 130.190 ;
        RECT 0.580 127.670 1075.680 129.370 ;
        RECT 1.090 126.850 1075.070 127.670 ;
        RECT 0.580 125.150 1075.680 126.850 ;
        RECT 1.090 124.330 1075.070 125.150 ;
        RECT 0.580 122.630 1075.680 124.330 ;
        RECT 1.090 121.810 1075.070 122.630 ;
        RECT 0.580 120.110 1075.680 121.810 ;
        RECT 1.090 119.290 1075.070 120.110 ;
        RECT 0.580 117.590 1075.680 119.290 ;
        RECT 1.090 116.770 1075.070 117.590 ;
        RECT 0.580 115.070 1075.680 116.770 ;
        RECT 1.090 114.250 1075.070 115.070 ;
        RECT 0.580 112.550 1075.680 114.250 ;
        RECT 1.090 111.730 1075.070 112.550 ;
        RECT 0.580 110.030 1075.680 111.730 ;
        RECT 1.090 109.210 1075.070 110.030 ;
        RECT 0.580 107.510 1075.680 109.210 ;
        RECT 1.090 106.690 1075.070 107.510 ;
        RECT 0.580 104.990 1075.680 106.690 ;
        RECT 1.090 104.170 1075.070 104.990 ;
        RECT 0.580 102.470 1075.680 104.170 ;
        RECT 1.090 101.650 1075.070 102.470 ;
        RECT 0.580 99.950 1075.680 101.650 ;
        RECT 1.090 99.130 1075.070 99.950 ;
        RECT 0.580 97.430 1075.680 99.130 ;
        RECT 1.090 96.610 1075.070 97.430 ;
        RECT 0.580 94.910 1075.680 96.610 ;
        RECT 1.090 94.090 1075.070 94.910 ;
        RECT 0.580 92.390 1075.680 94.090 ;
        RECT 1.090 91.570 1075.070 92.390 ;
        RECT 0.580 89.870 1075.680 91.570 ;
        RECT 1.090 89.050 1075.070 89.870 ;
        RECT 0.580 87.350 1075.680 89.050 ;
        RECT 1.090 86.530 1075.070 87.350 ;
        RECT 0.580 84.830 1075.680 86.530 ;
        RECT 1.090 84.010 1075.070 84.830 ;
        RECT 0.580 82.310 1075.680 84.010 ;
        RECT 1.090 81.490 1075.090 82.310 ;
        RECT 0.580 79.790 1075.680 81.490 ;
        RECT 1.090 78.970 1075.070 79.790 ;
        RECT 0.580 77.270 1075.680 78.970 ;
        RECT 1.090 76.450 1075.070 77.270 ;
        RECT 0.580 74.750 1075.680 76.450 ;
        RECT 1.090 73.930 1075.070 74.750 ;
        RECT 0.580 72.230 1075.680 73.930 ;
        RECT 1.090 71.410 1075.070 72.230 ;
        RECT 0.580 57.110 1075.680 71.410 ;
        RECT 1.090 56.290 1075.680 57.110 ;
        RECT 0.580 55.430 1075.680 56.290 ;
        RECT 1.090 54.610 1075.680 55.430 ;
        RECT 0.580 53.750 1075.680 54.610 ;
        RECT 1.090 52.930 1075.680 53.750 ;
        RECT 0.580 52.070 1075.680 52.930 ;
        RECT 1.090 51.250 1075.680 52.070 ;
        RECT 0.580 50.390 1075.680 51.250 ;
        RECT 1.090 49.570 1075.680 50.390 ;
        RECT 0.580 48.710 1075.680 49.570 ;
        RECT 1.090 47.890 1075.680 48.710 ;
        RECT 0.580 47.030 1075.680 47.890 ;
        RECT 1.090 46.210 1075.680 47.030 ;
        RECT 0.580 45.350 1075.680 46.210 ;
        RECT 1.090 44.530 1075.680 45.350 ;
        RECT 0.580 43.670 1075.680 44.530 ;
        RECT 1.090 42.850 1075.680 43.670 ;
        RECT 0.580 41.990 1075.680 42.850 ;
        RECT 1.090 41.170 1075.680 41.990 ;
        RECT 0.580 40.310 1075.680 41.170 ;
        RECT 1.090 39.490 1075.680 40.310 ;
        RECT 0.580 38.630 1075.680 39.490 ;
        RECT 1.090 37.810 1075.680 38.630 ;
        RECT 0.580 36.950 1075.680 37.810 ;
        RECT 1.090 36.130 1075.680 36.950 ;
        RECT 0.580 35.270 1075.680 36.130 ;
        RECT 1.090 34.450 1075.680 35.270 ;
        RECT 0.580 33.590 1075.680 34.450 ;
        RECT 1.090 32.770 1075.680 33.590 ;
        RECT 0.580 31.910 1075.680 32.770 ;
        RECT 1.090 31.090 1075.680 31.910 ;
        RECT 0.580 30.230 1075.680 31.090 ;
        RECT 1.090 29.410 1075.680 30.230 ;
        RECT 0.580 28.550 1075.680 29.410 ;
        RECT 1.090 27.730 1075.680 28.550 ;
        RECT 0.580 26.870 1075.680 27.730 ;
        RECT 1.090 26.050 1075.680 26.870 ;
        RECT 0.580 25.190 1075.680 26.050 ;
        RECT 1.090 24.370 1075.680 25.190 ;
        RECT 0.580 23.510 1075.680 24.370 ;
        RECT 1.090 22.690 1075.680 23.510 ;
        RECT 0.580 21.830 1075.680 22.690 ;
        RECT 1.090 21.010 1075.680 21.830 ;
        RECT 0.580 20.150 1075.680 21.010 ;
        RECT 1.090 19.330 1075.680 20.150 ;
        RECT 0.580 18.470 1075.680 19.330 ;
        RECT 1.090 17.650 1075.680 18.470 ;
        RECT 0.580 16.790 1075.680 17.650 ;
        RECT 1.090 15.970 1075.680 16.790 ;
        RECT 0.580 15.110 1075.680 15.970 ;
        RECT 1.090 14.290 1075.680 15.110 ;
        RECT 0.580 13.430 1075.680 14.290 ;
        RECT 1.090 12.610 1075.680 13.430 ;
        RECT 0.580 11.750 1075.680 12.610 ;
        RECT 1.090 10.930 1075.680 11.750 ;
        RECT 0.580 10.070 1075.680 10.930 ;
        RECT 1.090 9.250 1075.680 10.070 ;
        RECT 0.580 8.390 1075.680 9.250 ;
        RECT 1.090 7.570 1075.680 8.390 ;
        RECT 0.580 6.710 1075.680 7.570 ;
        RECT 1.090 5.890 1075.680 6.710 ;
        RECT 0.580 5.030 1075.680 5.890 ;
        RECT 1.090 4.210 1075.680 5.030 ;
        RECT 0.580 0.320 1075.680 4.210 ;
      LAYER Metal4 ;
        RECT 0.860 4.895 1075.300 1829.245 ;
      LAYER Metal5 ;
        RECT 1.295 6.620 1074.865 1827.730 ;
      LAYER TopMetal1 ;
        RECT 60.580 4.200 92.700 1832.040 ;
        RECT 98.180 4.200 124.620 1832.040 ;
        RECT 130.100 4.200 130.820 1832.040 ;
        RECT 136.300 4.200 200.220 1832.040 ;
        RECT 205.700 4.200 206.420 1832.040 ;
        RECT 211.900 4.200 275.820 1832.040 ;
        RECT 281.300 4.200 282.020 1832.040 ;
        RECT 287.500 4.200 339.660 1832.040 ;
        RECT 345.140 4.200 345.860 1832.040 ;
        RECT 351.340 4.200 415.260 1832.040 ;
        RECT 420.740 4.200 421.460 1832.040 ;
        RECT 426.940 4.200 490.860 1832.040 ;
        RECT 496.340 4.200 497.060 1832.040 ;
        RECT 502.540 4.200 554.700 1832.040 ;
        RECT 560.180 4.200 560.900 1832.040 ;
        RECT 566.380 4.200 630.300 1832.040 ;
        RECT 635.780 4.200 636.500 1832.040 ;
        RECT 641.980 4.200 705.900 1832.040 ;
        RECT 711.380 4.200 712.100 1832.040 ;
        RECT 717.580 4.200 769.740 1832.040 ;
        RECT 775.220 4.200 775.940 1832.040 ;
        RECT 781.420 4.200 845.340 1832.040 ;
        RECT 850.820 4.200 851.540 1832.040 ;
        RECT 857.020 4.200 920.940 1832.040 ;
        RECT 926.420 4.200 927.140 1832.040 ;
        RECT 932.620 4.200 984.780 1832.040 ;
        RECT 990.260 4.200 990.980 1832.040 ;
        RECT 996.460 4.200 1060.380 1832.040 ;
        RECT 1065.860 4.200 1070.420 1832.040 ;
  END
END eFPGA
END LIBRARY

