module heichips25_example_large (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net25;

 sg13g2_and2_1 _29_ (.A(net1),
    .B(net9),
    .X(_00_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _30_ (.A(net2),
    .B(net10),
    .X(_01_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _31_ (.B(net10),
    .A(net2),
    .X(_02_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _32_ (.B(_02_),
    .A(_00_),
    .X(net18),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _33_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_01_),
    .Y(_03_),
    .A2(_02_),
    .A1(_00_));
 sg13g2_and2_1 _34_ (.A(net3),
    .B(net11),
    .X(_04_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _35_ (.Y(_05_),
    .A(net3),
    .B(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _36_ (.A(_03_),
    .B(_05_),
    .Y(_06_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _37_ (.B(_05_),
    .A(_03_),
    .X(net19),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _38_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_07_),
    .B(net12),
    .A(net4));
 sg13g2_and2_1 _39_ (.A(net4),
    .B(net12),
    .X(_08_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _40_ (.B(net12),
    .A(net4),
    .X(_09_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _41_ (.A(_04_),
    .B(_06_),
    .Y(_10_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _42_ (.Y(net20),
    .A(_09_),
    .B(_10_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _43_ (.Y(_11_),
    .B(_09_),
    .A_N(_05_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _44_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04_),
    .A2(_07_),
    .Y(_12_),
    .B1(_08_));
 sg13g2_o21ai_1 _45_ (.B1(_12_),
    .VDD(VPWR),
    .Y(_13_),
    .VSS(VGND),
    .A1(_03_),
    .A2(_11_));
 sg13g2_nand2_1 _46_ (.Y(_14_),
    .A(net5),
    .B(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _47_ (.B(net13),
    .A(net5),
    .X(_15_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _48_ (.VDD(VPWR),
    .Y(_16_),
    .A(_15_),
    .VSS(VGND));
 sg13g2_nand2_1 _49_ (.Y(_17_),
    .A(_13_),
    .B(_15_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _50_ (.Y(net21),
    .A(_13_),
    .B(_16_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _51_ (.A(net6),
    .B(net14),
    .Y(_18_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _52_ (.Y(_19_),
    .A(net6),
    .B(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _53_ (.Y(_20_),
    .A(_14_),
    .B(_17_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _54_ (.Y(net22),
    .A(_19_),
    .B(_20_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _55_ (.A(_16_),
    .B(_19_),
    .Y(_21_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _56_ (.A(_14_),
    .B(_18_),
    .Y(_22_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _57_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_21_),
    .C1(_22_),
    .B1(_13_),
    .A1(net6),
    .Y(_23_),
    .A2(net14));
 sg13g2_nand2_1 _58_ (.Y(_24_),
    .A(net7),
    .B(net15),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _59_ (.A(net7),
    .B(net15),
    .Y(_25_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _60_ (.B(net15),
    .A(net7),
    .X(_26_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _61_ (.Y(net23),
    .A(_23_),
    .B(_26_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _62_ (.B1(_24_),
    .VDD(VPWR),
    .Y(_27_),
    .VSS(VGND),
    .A1(_23_),
    .A2(_25_));
 sg13g2_xnor2_1 _63_ (.Y(_28_),
    .A(net8),
    .B(net16),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _64_ (.Y(net24),
    .A(_27_),
    .B(_28_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _65_ (.B(net9),
    .A(net1),
    .X(net17),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo heichips25_example_large_26 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net26));
 sg13g2_tielo heichips25_example_large_27 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net27));
 sg13g2_tielo heichips25_example_large_28 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net28));
 sg13g2_tielo heichips25_example_large_29 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net29));
 sg13g2_tielo heichips25_example_large_30 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net30));
 sg13g2_tielo heichips25_example_large_31 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net31));
 sg13g2_tielo heichips25_example_large_32 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net32));
 sg13g2_tielo heichips25_example_large_33 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net33));
 sg13g2_tielo heichips25_example_large_34 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net34));
 sg13g2_tielo heichips25_example_large_35 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net35));
 sg13g2_tielo heichips25_example_large_36 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net36));
 sg13g2_tielo heichips25_example_large_37 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net37));
 sg13g2_tielo heichips25_example_large_38 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net38));
 sg13g2_tielo heichips25_example_large_39 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net39));
 sg13g2_tielo heichips25_example_large_40 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net40));
 sg13g2_decap_8 FILLER_0_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input9 (.A(uio_in[0]),
    .X(net9),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input10 (.A(uio_in[1]),
    .X(net10),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input11 (.A(uio_in[2]),
    .X(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input12 (.A(uio_in[3]),
    .X(net12),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input13 (.A(uio_in[4]),
    .X(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input14 (.A(uio_in[5]),
    .X(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input15 (.A(uio_in[6]),
    .X(net15),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input16 (.A(uio_in[7]),
    .X(net16),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo heichips25_example_large_25 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net25));
 sg13g2_decap_8 FILLER_0_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_58_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_59_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_59_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_60_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_60_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_60_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_60_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_60_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_13 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_61_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_68_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_68_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_68_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_69_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_69_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_69_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_71_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_71_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_73_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_73_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_73_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_74_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_74_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_74_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_75_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_76_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_79_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_79_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_81_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_81_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_83_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_86_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_86_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_88_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_90_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_5 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_95_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_98_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_98_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_1022 (.VDD(VPWR),
    .VSS(VGND));
 assign uio_oe[0] = net25;
 assign uio_oe[1] = net26;
 assign uio_oe[2] = net27;
 assign uio_oe[3] = net28;
 assign uio_oe[4] = net29;
 assign uio_oe[5] = net30;
 assign uio_oe[6] = net31;
 assign uio_oe[7] = net32;
 assign uio_out[0] = net33;
 assign uio_out[1] = net34;
 assign uio_out[2] = net35;
 assign uio_out[3] = net36;
 assign uio_out[4] = net37;
 assign uio_out[5] = net38;
 assign uio_out[6] = net39;
 assign uio_out[7] = net40;
endmodule
