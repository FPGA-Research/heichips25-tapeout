magic
tech ihp-sg13g2
magscale 1 2
timestamp 1752760856
<< metal1 >>
rect 1152 9848 20452 9872
rect 1152 9808 4928 9848
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 5296 9808 20048 9848
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20416 9808 20452 9848
rect 1152 9784 20452 9808
rect 19371 9680 19413 9689
rect 19371 9640 19372 9680
rect 19412 9640 19413 9680
rect 19371 9631 19413 9640
rect 19171 9428 19229 9429
rect 19171 9388 19180 9428
rect 19220 9388 19229 9428
rect 19171 9387 19229 9388
rect 1152 9092 20352 9116
rect 1152 9052 3688 9092
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 4056 9052 18808 9092
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 19176 9052 20352 9092
rect 1152 9028 20352 9052
rect 11403 8924 11445 8933
rect 11403 8884 11404 8924
rect 11444 8884 11445 8924
rect 11403 8875 11445 8884
rect 2187 8840 2229 8849
rect 2187 8800 2188 8840
rect 2228 8800 2229 8840
rect 2187 8791 2229 8800
rect 4395 8840 4437 8849
rect 4395 8800 4396 8840
rect 4436 8800 4437 8840
rect 4395 8791 4437 8800
rect 5163 8840 5205 8849
rect 5163 8800 5164 8840
rect 5204 8800 5205 8840
rect 5163 8791 5205 8800
rect 5643 8840 5685 8849
rect 5643 8800 5644 8840
rect 5684 8800 5685 8840
rect 5643 8791 5685 8800
rect 7083 8840 7125 8849
rect 7083 8800 7084 8840
rect 7124 8800 7125 8840
rect 7083 8791 7125 8800
rect 7467 8840 7509 8849
rect 7467 8800 7468 8840
rect 7508 8800 7509 8840
rect 7467 8791 7509 8800
rect 8043 8840 8085 8849
rect 8043 8800 8044 8840
rect 8084 8800 8085 8840
rect 8043 8791 8085 8800
rect 10059 8840 10101 8849
rect 10059 8800 10060 8840
rect 10100 8800 10101 8840
rect 10059 8791 10101 8800
rect 10635 8840 10677 8849
rect 10635 8800 10636 8840
rect 10676 8800 10677 8840
rect 10635 8791 10677 8800
rect 11019 8840 11061 8849
rect 11019 8800 11020 8840
rect 11060 8800 11061 8840
rect 11019 8791 11061 8800
rect 16299 8840 16341 8849
rect 16299 8800 16300 8840
rect 16340 8800 16341 8840
rect 16299 8791 16341 8800
rect 16491 8840 16533 8849
rect 16491 8800 16492 8840
rect 16532 8800 16533 8840
rect 16491 8791 16533 8800
rect 17067 8840 17109 8849
rect 17067 8800 17068 8840
rect 17108 8800 17109 8840
rect 17067 8791 17109 8800
rect 18987 8840 19029 8849
rect 18987 8800 18988 8840
rect 19028 8800 19029 8840
rect 18987 8791 19029 8800
rect 19371 8840 19413 8849
rect 19371 8800 19372 8840
rect 19412 8800 19413 8840
rect 19371 8791 19413 8800
rect 19755 8840 19797 8849
rect 19755 8800 19756 8840
rect 19796 8800 19797 8840
rect 19755 8791 19797 8800
rect 1795 8756 1853 8757
rect 1795 8716 1804 8756
rect 1844 8716 1853 8756
rect 1795 8715 1853 8716
rect 2371 8756 2429 8757
rect 2371 8716 2380 8756
rect 2420 8716 2429 8756
rect 2371 8715 2429 8716
rect 2755 8756 2813 8757
rect 2755 8716 2764 8756
rect 2804 8716 2813 8756
rect 2755 8715 2813 8716
rect 4579 8756 4637 8757
rect 4579 8716 4588 8756
rect 4628 8716 4637 8756
rect 4579 8715 4637 8716
rect 4963 8756 5021 8757
rect 4963 8716 4972 8756
rect 5012 8716 5021 8756
rect 4963 8715 5021 8716
rect 5347 8756 5405 8757
rect 5347 8716 5356 8756
rect 5396 8716 5405 8756
rect 5347 8715 5405 8716
rect 5827 8756 5885 8757
rect 5827 8716 5836 8756
rect 5876 8716 5885 8756
rect 5827 8715 5885 8716
rect 6307 8756 6365 8757
rect 6307 8716 6316 8756
rect 6356 8716 6365 8756
rect 6307 8715 6365 8716
rect 7267 8756 7325 8757
rect 7267 8716 7276 8756
rect 7316 8716 7325 8756
rect 7267 8715 7325 8716
rect 7651 8756 7709 8757
rect 7651 8716 7660 8756
rect 7700 8716 7709 8756
rect 7651 8715 7709 8716
rect 8227 8756 8285 8757
rect 8227 8716 8236 8756
rect 8276 8716 8285 8756
rect 8227 8715 8285 8716
rect 10243 8756 10301 8757
rect 10243 8716 10252 8756
rect 10292 8716 10301 8756
rect 10243 8715 10301 8716
rect 10819 8756 10877 8757
rect 10819 8716 10828 8756
rect 10868 8716 10877 8756
rect 10819 8715 10877 8716
rect 11203 8756 11261 8757
rect 11203 8716 11212 8756
rect 11252 8716 11261 8756
rect 11203 8715 11261 8716
rect 11587 8756 11645 8757
rect 11587 8716 11596 8756
rect 11636 8716 11645 8756
rect 11587 8715 11645 8716
rect 11971 8756 12029 8757
rect 11971 8716 11980 8756
rect 12020 8716 12029 8756
rect 11971 8715 12029 8716
rect 14467 8756 14525 8757
rect 14467 8716 14476 8756
rect 14516 8716 14525 8756
rect 14467 8715 14525 8716
rect 14851 8756 14909 8757
rect 14851 8716 14860 8756
rect 14900 8716 14909 8756
rect 14851 8715 14909 8716
rect 15427 8756 15485 8757
rect 15427 8716 15436 8756
rect 15476 8716 15485 8756
rect 15427 8715 15485 8716
rect 16099 8756 16157 8757
rect 16099 8716 16108 8756
rect 16148 8716 16157 8756
rect 16099 8715 16157 8716
rect 16675 8756 16733 8757
rect 16675 8716 16684 8756
rect 16724 8716 16733 8756
rect 16675 8715 16733 8716
rect 17251 8756 17309 8757
rect 17251 8716 17260 8756
rect 17300 8716 17309 8756
rect 17251 8715 17309 8716
rect 17731 8756 17789 8757
rect 17731 8716 17740 8756
rect 17780 8716 17789 8756
rect 17731 8715 17789 8716
rect 18787 8756 18845 8757
rect 18787 8716 18796 8756
rect 18836 8716 18845 8756
rect 18787 8715 18845 8716
rect 19171 8756 19229 8757
rect 19171 8716 19180 8756
rect 19220 8716 19229 8756
rect 19171 8715 19229 8716
rect 19555 8756 19613 8757
rect 19555 8716 19564 8756
rect 19604 8716 19613 8756
rect 19555 8715 19613 8716
rect 1995 8504 2037 8513
rect 1995 8464 1996 8504
rect 2036 8464 2037 8504
rect 1995 8455 2037 8464
rect 2571 8504 2613 8513
rect 2571 8464 2572 8504
rect 2612 8464 2613 8504
rect 2571 8455 2613 8464
rect 4779 8504 4821 8513
rect 4779 8464 4780 8504
rect 4820 8464 4821 8504
rect 4779 8455 4821 8464
rect 6123 8504 6165 8513
rect 6123 8464 6124 8504
rect 6164 8464 6165 8504
rect 6123 8455 6165 8464
rect 11787 8504 11829 8513
rect 11787 8464 11788 8504
rect 11828 8464 11829 8504
rect 11787 8455 11829 8464
rect 14283 8504 14325 8513
rect 14283 8464 14284 8504
rect 14324 8464 14325 8504
rect 14283 8455 14325 8464
rect 14667 8504 14709 8513
rect 14667 8464 14668 8504
rect 14708 8464 14709 8504
rect 14667 8455 14709 8464
rect 15243 8504 15285 8513
rect 15243 8464 15244 8504
rect 15284 8464 15285 8504
rect 15243 8455 15285 8464
rect 17931 8504 17973 8513
rect 17931 8464 17932 8504
rect 17972 8464 17973 8504
rect 17931 8455 17973 8464
rect 1152 8336 20452 8360
rect 1152 8296 4928 8336
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 5296 8296 20048 8336
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20416 8296 20452 8336
rect 1152 8272 20452 8296
rect 2091 8168 2133 8177
rect 2091 8128 2092 8168
rect 2132 8128 2133 8168
rect 2091 8119 2133 8128
rect 2763 8168 2805 8177
rect 2763 8128 2764 8168
rect 2804 8128 2805 8168
rect 2763 8119 2805 8128
rect 3339 8168 3381 8177
rect 3339 8128 3340 8168
rect 3380 8128 3381 8168
rect 3339 8119 3381 8128
rect 4107 8168 4149 8177
rect 4107 8128 4108 8168
rect 4148 8128 4149 8168
rect 4107 8119 4149 8128
rect 7083 8168 7125 8177
rect 7083 8128 7084 8168
rect 7124 8128 7125 8168
rect 7083 8119 7125 8128
rect 7659 8168 7701 8177
rect 7659 8128 7660 8168
rect 7700 8128 7701 8168
rect 7659 8119 7701 8128
rect 8043 8168 8085 8177
rect 8043 8128 8044 8168
rect 8084 8128 8085 8168
rect 8043 8119 8085 8128
rect 8427 8168 8469 8177
rect 8427 8128 8428 8168
rect 8468 8128 8469 8168
rect 8427 8119 8469 8128
rect 9579 8168 9621 8177
rect 9579 8128 9580 8168
rect 9620 8128 9621 8168
rect 9579 8119 9621 8128
rect 9963 8168 10005 8177
rect 9963 8128 9964 8168
rect 10004 8128 10005 8168
rect 9963 8119 10005 8128
rect 11403 8168 11445 8177
rect 11403 8128 11404 8168
rect 11444 8128 11445 8168
rect 11403 8119 11445 8128
rect 13227 8168 13269 8177
rect 13227 8128 13228 8168
rect 13268 8128 13269 8168
rect 13227 8119 13269 8128
rect 13707 8168 13749 8177
rect 13707 8128 13708 8168
rect 13748 8128 13749 8168
rect 13707 8119 13749 8128
rect 17163 8168 17205 8177
rect 17163 8128 17164 8168
rect 17204 8128 17205 8168
rect 17163 8119 17205 8128
rect 19371 8168 19413 8177
rect 19371 8128 19372 8168
rect 19412 8128 19413 8168
rect 19371 8119 19413 8128
rect 1891 7916 1949 7917
rect 1891 7876 1900 7916
rect 1940 7876 1949 7916
rect 1891 7875 1949 7876
rect 2563 7916 2621 7917
rect 2563 7876 2572 7916
rect 2612 7876 2621 7916
rect 2563 7875 2621 7876
rect 3523 7916 3581 7917
rect 3523 7876 3532 7916
rect 3572 7876 3581 7916
rect 3523 7875 3581 7876
rect 4291 7916 4349 7917
rect 4291 7876 4300 7916
rect 4340 7876 4349 7916
rect 4291 7875 4349 7876
rect 7267 7916 7325 7917
rect 7267 7876 7276 7916
rect 7316 7876 7325 7916
rect 7267 7875 7325 7876
rect 7843 7916 7901 7917
rect 7843 7876 7852 7916
rect 7892 7876 7901 7916
rect 7843 7875 7901 7876
rect 8227 7916 8285 7917
rect 8227 7876 8236 7916
rect 8276 7876 8285 7916
rect 8227 7875 8285 7876
rect 8611 7916 8669 7917
rect 8611 7876 8620 7916
rect 8660 7876 8669 7916
rect 8611 7875 8669 7876
rect 9763 7916 9821 7917
rect 9763 7876 9772 7916
rect 9812 7876 9821 7916
rect 9763 7875 9821 7876
rect 10147 7916 10205 7917
rect 10147 7876 10156 7916
rect 10196 7876 10205 7916
rect 10147 7875 10205 7876
rect 11587 7916 11645 7917
rect 11587 7876 11596 7916
rect 11636 7876 11645 7916
rect 11587 7875 11645 7876
rect 12931 7916 12989 7917
rect 12931 7876 12940 7916
rect 12980 7876 12989 7916
rect 12931 7875 12989 7876
rect 13411 7916 13469 7917
rect 13411 7876 13420 7916
rect 13460 7876 13469 7916
rect 13411 7875 13469 7876
rect 13891 7916 13949 7917
rect 13891 7876 13900 7916
rect 13940 7876 13949 7916
rect 13891 7875 13949 7876
rect 16195 7916 16253 7917
rect 16195 7876 16204 7916
rect 16244 7876 16253 7916
rect 16195 7875 16253 7876
rect 16963 7916 17021 7917
rect 16963 7876 16972 7916
rect 17012 7876 17021 7916
rect 16963 7875 17021 7876
rect 19171 7916 19229 7917
rect 19171 7876 19180 7916
rect 19220 7876 19229 7916
rect 19171 7875 19229 7876
rect 16395 7832 16437 7841
rect 16395 7792 16396 7832
rect 16436 7792 16437 7832
rect 16395 7783 16437 7792
rect 12747 7748 12789 7757
rect 12747 7708 12748 7748
rect 12788 7708 12789 7748
rect 12747 7699 12789 7708
rect 1152 7580 20352 7604
rect 1152 7540 3688 7580
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 4056 7540 18808 7580
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 19176 7540 20352 7580
rect 1152 7516 20352 7540
rect 2091 7412 2133 7421
rect 2091 7372 2092 7412
rect 2132 7372 2133 7412
rect 2091 7363 2133 7372
rect 1891 7244 1949 7245
rect 1891 7204 1900 7244
rect 1940 7204 1949 7244
rect 1891 7203 1949 7204
rect 1152 6824 20452 6848
rect 1152 6784 4928 6824
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 5296 6784 20048 6824
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20416 6784 20452 6824
rect 1152 6760 20452 6784
rect 16491 6656 16533 6665
rect 16491 6616 16492 6656
rect 16532 6616 16533 6656
rect 16491 6607 16533 6616
rect 17931 6656 17973 6665
rect 17931 6616 17932 6656
rect 17972 6616 17973 6656
rect 17931 6607 17973 6616
rect 19179 6656 19221 6665
rect 19179 6616 19180 6656
rect 19220 6616 19221 6656
rect 19179 6607 19221 6616
rect 19563 6656 19605 6665
rect 19563 6616 19564 6656
rect 19604 6616 19605 6656
rect 19563 6607 19605 6616
rect 1987 6404 2045 6405
rect 1987 6364 1996 6404
rect 2036 6364 2045 6404
rect 1987 6363 2045 6364
rect 16291 6404 16349 6405
rect 16291 6364 16300 6404
rect 16340 6364 16349 6404
rect 16291 6363 16349 6364
rect 17731 6404 17789 6405
rect 17731 6364 17740 6404
rect 17780 6364 17789 6404
rect 17731 6363 17789 6364
rect 18979 6404 19037 6405
rect 18979 6364 18988 6404
rect 19028 6364 19037 6404
rect 18979 6363 19037 6364
rect 19363 6404 19421 6405
rect 19363 6364 19372 6404
rect 19412 6364 19421 6404
rect 19363 6363 19421 6364
rect 2187 6236 2229 6245
rect 2187 6196 2188 6236
rect 2228 6196 2229 6236
rect 2187 6187 2229 6196
rect 1152 6068 20352 6092
rect 1152 6028 3688 6068
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 4056 6028 18808 6068
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 19176 6028 20352 6068
rect 1152 6004 20352 6028
rect 16971 5900 17013 5909
rect 16971 5860 16972 5900
rect 17012 5860 17013 5900
rect 16971 5851 17013 5860
rect 18699 5900 18741 5909
rect 18699 5860 18700 5900
rect 18740 5860 18741 5900
rect 18699 5851 18741 5860
rect 19563 5900 19605 5909
rect 19563 5860 19564 5900
rect 19604 5860 19605 5900
rect 19563 5851 19605 5860
rect 12163 5732 12221 5733
rect 12163 5692 12172 5732
rect 12212 5692 12221 5732
rect 12163 5691 12221 5692
rect 16771 5732 16829 5733
rect 16771 5692 16780 5732
rect 16820 5692 16829 5732
rect 16771 5691 16829 5692
rect 18499 5732 18557 5733
rect 18499 5692 18508 5732
rect 18548 5692 18557 5732
rect 18499 5691 18557 5692
rect 19363 5732 19421 5733
rect 19363 5692 19372 5732
rect 19412 5692 19421 5732
rect 19363 5691 19421 5692
rect 12363 5480 12405 5489
rect 12363 5440 12364 5480
rect 12404 5440 12405 5480
rect 12363 5431 12405 5440
rect 1152 5312 20452 5336
rect 1152 5272 4928 5312
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 5296 5272 20048 5312
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20416 5272 20452 5312
rect 1152 5248 20452 5272
rect 2275 4892 2333 4893
rect 2275 4852 2284 4892
rect 2324 4852 2333 4892
rect 2275 4851 2333 4852
rect 9475 4892 9533 4893
rect 9475 4852 9484 4892
rect 9524 4852 9533 4892
rect 9475 4851 9533 4852
rect 2475 4808 2517 4817
rect 2475 4768 2476 4808
rect 2516 4768 2517 4808
rect 2475 4759 2517 4768
rect 9675 4808 9717 4817
rect 9675 4768 9676 4808
rect 9716 4768 9717 4808
rect 9675 4759 9717 4768
rect 1152 4556 20352 4580
rect 1152 4516 3688 4556
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 4056 4516 18808 4556
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 19176 4516 20352 4556
rect 1152 4492 20352 4516
rect 19275 4388 19317 4397
rect 19275 4348 19276 4388
rect 19316 4348 19317 4388
rect 19275 4339 19317 4348
rect 1891 4220 1949 4221
rect 1891 4180 1900 4220
rect 1940 4180 1949 4220
rect 1891 4179 1949 4180
rect 2275 4220 2333 4221
rect 2275 4180 2284 4220
rect 2324 4180 2333 4220
rect 2275 4179 2333 4180
rect 2659 4220 2717 4221
rect 2659 4180 2668 4220
rect 2708 4180 2717 4220
rect 2659 4179 2717 4180
rect 9763 4220 9821 4221
rect 9763 4180 9772 4220
rect 9812 4180 9821 4220
rect 9763 4179 9821 4180
rect 12931 4220 12989 4221
rect 12931 4180 12940 4220
rect 12980 4180 12989 4220
rect 12931 4179 12989 4180
rect 19075 4220 19133 4221
rect 19075 4180 19084 4220
rect 19124 4180 19133 4220
rect 19075 4179 19133 4180
rect 19459 4220 19517 4221
rect 19459 4180 19468 4220
rect 19508 4180 19517 4220
rect 19459 4179 19517 4180
rect 2091 3968 2133 3977
rect 2091 3928 2092 3968
rect 2132 3928 2133 3968
rect 2091 3919 2133 3928
rect 2475 3968 2517 3977
rect 2475 3928 2476 3968
rect 2516 3928 2517 3968
rect 2475 3919 2517 3928
rect 2859 3968 2901 3977
rect 2859 3928 2860 3968
rect 2900 3928 2901 3968
rect 2859 3919 2901 3928
rect 9963 3968 10005 3977
rect 9963 3928 9964 3968
rect 10004 3928 10005 3968
rect 9963 3919 10005 3928
rect 13131 3968 13173 3977
rect 13131 3928 13132 3968
rect 13172 3928 13173 3968
rect 13131 3919 13173 3928
rect 19659 3968 19701 3977
rect 19659 3928 19660 3968
rect 19700 3928 19701 3968
rect 19659 3919 19701 3928
rect 1152 3800 20452 3824
rect 1152 3760 4928 3800
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 5296 3760 20048 3800
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20416 3760 20452 3800
rect 1152 3736 20452 3760
rect 2179 3380 2237 3381
rect 2179 3340 2188 3380
rect 2228 3340 2237 3380
rect 2179 3339 2237 3340
rect 2379 3212 2421 3221
rect 2379 3172 2380 3212
rect 2420 3172 2421 3212
rect 2379 3163 2421 3172
rect 1152 3044 20352 3068
rect 1152 3004 3688 3044
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 4056 3004 18808 3044
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 19176 3004 20352 3044
rect 1152 2980 20352 3004
rect 14667 2792 14709 2801
rect 14667 2752 14668 2792
rect 14708 2752 14709 2792
rect 14667 2743 14709 2752
rect 14467 2708 14525 2709
rect 14467 2668 14476 2708
rect 14516 2668 14525 2708
rect 14467 2667 14525 2668
rect 1152 2288 20452 2312
rect 1152 2248 4928 2288
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 5296 2248 20048 2288
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20416 2248 20452 2288
rect 1152 2224 20452 2248
rect 3435 2120 3477 2129
rect 3435 2080 3436 2120
rect 3476 2080 3477 2120
rect 3435 2071 3477 2080
rect 4107 2120 4149 2129
rect 4107 2080 4108 2120
rect 4148 2080 4149 2120
rect 4107 2071 4149 2080
rect 5835 2120 5877 2129
rect 5835 2080 5836 2120
rect 5876 2080 5877 2120
rect 5835 2071 5877 2080
rect 6603 2120 6645 2129
rect 6603 2080 6604 2120
rect 6644 2080 6645 2120
rect 6603 2071 6645 2080
rect 9963 2120 10005 2129
rect 9963 2080 9964 2120
rect 10004 2080 10005 2120
rect 9963 2071 10005 2080
rect 10731 2120 10773 2129
rect 10731 2080 10732 2120
rect 10772 2080 10773 2120
rect 10731 2071 10773 2080
rect 12075 2120 12117 2129
rect 12075 2080 12076 2120
rect 12116 2080 12117 2120
rect 12075 2071 12117 2080
rect 13227 2120 13269 2129
rect 13227 2080 13228 2120
rect 13268 2080 13269 2120
rect 13227 2071 13269 2080
rect 14571 2120 14613 2129
rect 14571 2080 14572 2120
rect 14612 2080 14613 2120
rect 14571 2071 14613 2080
rect 15339 2120 15381 2129
rect 15339 2080 15340 2120
rect 15380 2080 15381 2120
rect 15339 2071 15381 2080
rect 15915 2120 15957 2129
rect 15915 2080 15916 2120
rect 15956 2080 15957 2120
rect 15915 2071 15957 2080
rect 16395 2120 16437 2129
rect 16395 2080 16396 2120
rect 16436 2080 16437 2120
rect 16395 2071 16437 2080
rect 17643 2120 17685 2129
rect 17643 2080 17644 2120
rect 17684 2080 17685 2120
rect 17643 2071 17685 2080
rect 18027 2120 18069 2129
rect 18027 2080 18028 2120
rect 18068 2080 18069 2120
rect 18027 2071 18069 2080
rect 19275 2120 19317 2129
rect 19275 2080 19276 2120
rect 19316 2080 19317 2120
rect 19275 2071 19317 2080
rect 19851 2120 19893 2129
rect 19851 2080 19852 2120
rect 19892 2080 19893 2120
rect 19851 2071 19893 2080
rect 1507 1868 1565 1869
rect 1507 1828 1516 1868
rect 1556 1828 1565 1868
rect 1507 1827 1565 1828
rect 1891 1868 1949 1869
rect 1891 1828 1900 1868
rect 1940 1828 1949 1868
rect 1891 1827 1949 1828
rect 2275 1868 2333 1869
rect 2275 1828 2284 1868
rect 2324 1828 2333 1868
rect 2275 1827 2333 1828
rect 3235 1868 3293 1869
rect 3235 1828 3244 1868
rect 3284 1828 3293 1868
rect 3235 1827 3293 1828
rect 3907 1868 3965 1869
rect 3907 1828 3916 1868
rect 3956 1828 3965 1868
rect 3907 1827 3965 1828
rect 4291 1868 4349 1869
rect 4291 1828 4300 1868
rect 4340 1828 4349 1868
rect 4291 1827 4349 1828
rect 4675 1868 4733 1869
rect 4675 1828 4684 1868
rect 4724 1828 4733 1868
rect 4675 1827 4733 1828
rect 5635 1868 5693 1869
rect 5635 1828 5644 1868
rect 5684 1828 5693 1868
rect 5635 1827 5693 1828
rect 6019 1868 6077 1869
rect 6019 1828 6028 1868
rect 6068 1828 6077 1868
rect 6019 1827 6077 1828
rect 6403 1868 6461 1869
rect 6403 1828 6412 1868
rect 6452 1828 6461 1868
rect 6403 1827 6461 1828
rect 8323 1868 8381 1869
rect 8323 1828 8332 1868
rect 8372 1828 8381 1868
rect 8323 1827 8381 1828
rect 9763 1868 9821 1869
rect 9763 1828 9772 1868
rect 9812 1828 9821 1868
rect 9763 1827 9821 1828
rect 10531 1868 10589 1869
rect 10531 1828 10540 1868
rect 10580 1828 10589 1868
rect 10531 1827 10589 1828
rect 11875 1868 11933 1869
rect 11875 1828 11884 1868
rect 11924 1828 11933 1868
rect 11875 1827 11933 1828
rect 13027 1868 13085 1869
rect 13027 1828 13036 1868
rect 13076 1828 13085 1868
rect 13027 1827 13085 1828
rect 14371 1868 14429 1869
rect 14371 1828 14380 1868
rect 14420 1828 14429 1868
rect 14371 1827 14429 1828
rect 15139 1868 15197 1869
rect 15139 1828 15148 1868
rect 15188 1828 15197 1868
rect 15139 1827 15197 1828
rect 15715 1868 15773 1869
rect 15715 1828 15724 1868
rect 15764 1828 15773 1868
rect 15715 1827 15773 1828
rect 16195 1868 16253 1869
rect 16195 1828 16204 1868
rect 16244 1828 16253 1868
rect 16195 1827 16253 1828
rect 17443 1868 17501 1869
rect 17443 1828 17452 1868
rect 17492 1828 17501 1868
rect 17443 1827 17501 1828
rect 17827 1868 17885 1869
rect 17827 1828 17836 1868
rect 17876 1828 17885 1868
rect 17827 1827 17885 1828
rect 19075 1868 19133 1869
rect 19075 1828 19084 1868
rect 19124 1828 19133 1868
rect 19075 1827 19133 1828
rect 19459 1868 19517 1869
rect 19459 1828 19468 1868
rect 19508 1828 19517 1868
rect 19459 1827 19517 1828
rect 20035 1868 20093 1869
rect 20035 1828 20044 1868
rect 20084 1828 20093 1868
rect 20035 1827 20093 1828
rect 19659 1784 19701 1793
rect 19659 1744 19660 1784
rect 19700 1744 19701 1784
rect 19659 1735 19701 1744
rect 1707 1700 1749 1709
rect 1707 1660 1708 1700
rect 1748 1660 1749 1700
rect 1707 1651 1749 1660
rect 2091 1700 2133 1709
rect 2091 1660 2092 1700
rect 2132 1660 2133 1700
rect 2091 1651 2133 1660
rect 2475 1700 2517 1709
rect 2475 1660 2476 1700
rect 2516 1660 2517 1700
rect 2475 1651 2517 1660
rect 4491 1700 4533 1709
rect 4491 1660 4492 1700
rect 4532 1660 4533 1700
rect 4491 1651 4533 1660
rect 4875 1700 4917 1709
rect 4875 1660 4876 1700
rect 4916 1660 4917 1700
rect 4875 1651 4917 1660
rect 6219 1700 6261 1709
rect 6219 1660 6220 1700
rect 6260 1660 6261 1700
rect 6219 1651 6261 1660
rect 8523 1700 8565 1709
rect 8523 1660 8524 1700
rect 8564 1660 8565 1700
rect 8523 1651 8565 1660
rect 1152 1532 20352 1556
rect 1152 1492 3688 1532
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 4056 1492 18808 1532
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 19176 1492 20352 1532
rect 1152 1468 20352 1492
rect 1152 776 20452 800
rect 1152 736 4928 776
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 5296 736 20048 776
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20416 736 20452 776
rect 1152 712 20452 736
<< via1 >>
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 19372 9640 19412 9680
rect 19180 9388 19220 9428
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 11404 8884 11444 8924
rect 2188 8800 2228 8840
rect 4396 8800 4436 8840
rect 5164 8800 5204 8840
rect 5644 8800 5684 8840
rect 7084 8800 7124 8840
rect 7468 8800 7508 8840
rect 8044 8800 8084 8840
rect 10060 8800 10100 8840
rect 10636 8800 10676 8840
rect 11020 8800 11060 8840
rect 16300 8800 16340 8840
rect 16492 8800 16532 8840
rect 17068 8800 17108 8840
rect 18988 8800 19028 8840
rect 19372 8800 19412 8840
rect 19756 8800 19796 8840
rect 1804 8716 1844 8756
rect 2380 8716 2420 8756
rect 2764 8716 2804 8756
rect 4588 8716 4628 8756
rect 4972 8716 5012 8756
rect 5356 8716 5396 8756
rect 5836 8716 5876 8756
rect 6316 8716 6356 8756
rect 7276 8716 7316 8756
rect 7660 8716 7700 8756
rect 8236 8716 8276 8756
rect 10252 8716 10292 8756
rect 10828 8716 10868 8756
rect 11212 8716 11252 8756
rect 11596 8716 11636 8756
rect 11980 8716 12020 8756
rect 14476 8716 14516 8756
rect 14860 8716 14900 8756
rect 15436 8716 15476 8756
rect 16108 8716 16148 8756
rect 16684 8716 16724 8756
rect 17260 8716 17300 8756
rect 17740 8716 17780 8756
rect 18796 8716 18836 8756
rect 19180 8716 19220 8756
rect 19564 8716 19604 8756
rect 1996 8464 2036 8504
rect 2572 8464 2612 8504
rect 4780 8464 4820 8504
rect 6124 8464 6164 8504
rect 11788 8464 11828 8504
rect 14284 8464 14324 8504
rect 14668 8464 14708 8504
rect 15244 8464 15284 8504
rect 17932 8464 17972 8504
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 2092 8128 2132 8168
rect 2764 8128 2804 8168
rect 3340 8128 3380 8168
rect 4108 8128 4148 8168
rect 7084 8128 7124 8168
rect 7660 8128 7700 8168
rect 8044 8128 8084 8168
rect 8428 8128 8468 8168
rect 9580 8128 9620 8168
rect 9964 8128 10004 8168
rect 11404 8128 11444 8168
rect 13228 8128 13268 8168
rect 13708 8128 13748 8168
rect 17164 8128 17204 8168
rect 19372 8128 19412 8168
rect 1900 7876 1940 7916
rect 2572 7876 2612 7916
rect 3532 7876 3572 7916
rect 4300 7876 4340 7916
rect 7276 7876 7316 7916
rect 7852 7876 7892 7916
rect 8236 7876 8276 7916
rect 8620 7876 8660 7916
rect 9772 7876 9812 7916
rect 10156 7876 10196 7916
rect 11596 7876 11636 7916
rect 12940 7876 12980 7916
rect 13420 7876 13460 7916
rect 13900 7876 13940 7916
rect 16204 7876 16244 7916
rect 16972 7876 17012 7916
rect 19180 7876 19220 7916
rect 16396 7792 16436 7832
rect 12748 7708 12788 7748
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 2092 7372 2132 7412
rect 1900 7204 1940 7244
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 16492 6616 16532 6656
rect 17932 6616 17972 6656
rect 19180 6616 19220 6656
rect 19564 6616 19604 6656
rect 1996 6364 2036 6404
rect 16300 6364 16340 6404
rect 17740 6364 17780 6404
rect 18988 6364 19028 6404
rect 19372 6364 19412 6404
rect 2188 6196 2228 6236
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 16972 5860 17012 5900
rect 18700 5860 18740 5900
rect 19564 5860 19604 5900
rect 12172 5692 12212 5732
rect 16780 5692 16820 5732
rect 18508 5692 18548 5732
rect 19372 5692 19412 5732
rect 12364 5440 12404 5480
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 2284 4852 2324 4892
rect 9484 4852 9524 4892
rect 2476 4768 2516 4808
rect 9676 4768 9716 4808
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 19276 4348 19316 4388
rect 1900 4180 1940 4220
rect 2284 4180 2324 4220
rect 2668 4180 2708 4220
rect 9772 4180 9812 4220
rect 12940 4180 12980 4220
rect 19084 4180 19124 4220
rect 19468 4180 19508 4220
rect 2092 3928 2132 3968
rect 2476 3928 2516 3968
rect 2860 3928 2900 3968
rect 9964 3928 10004 3968
rect 13132 3928 13172 3968
rect 19660 3928 19700 3968
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 2188 3340 2228 3380
rect 2380 3172 2420 3212
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 14668 2752 14708 2792
rect 14476 2668 14516 2708
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 3436 2080 3476 2120
rect 4108 2080 4148 2120
rect 5836 2080 5876 2120
rect 6604 2080 6644 2120
rect 9964 2080 10004 2120
rect 10732 2080 10772 2120
rect 12076 2080 12116 2120
rect 13228 2080 13268 2120
rect 14572 2080 14612 2120
rect 15340 2080 15380 2120
rect 15916 2080 15956 2120
rect 16396 2080 16436 2120
rect 17644 2080 17684 2120
rect 18028 2080 18068 2120
rect 19276 2080 19316 2120
rect 19852 2080 19892 2120
rect 1516 1828 1556 1868
rect 1900 1828 1940 1868
rect 2284 1828 2324 1868
rect 3244 1828 3284 1868
rect 3916 1828 3956 1868
rect 4300 1828 4340 1868
rect 4684 1828 4724 1868
rect 5644 1828 5684 1868
rect 6028 1828 6068 1868
rect 6412 1828 6452 1868
rect 8332 1828 8372 1868
rect 9772 1828 9812 1868
rect 10540 1828 10580 1868
rect 11884 1828 11924 1868
rect 13036 1828 13076 1868
rect 14380 1828 14420 1868
rect 15148 1828 15188 1868
rect 15724 1828 15764 1868
rect 16204 1828 16244 1868
rect 17452 1828 17492 1868
rect 17836 1828 17876 1868
rect 19084 1828 19124 1868
rect 19468 1828 19508 1868
rect 20044 1828 20084 1868
rect 19660 1744 19700 1784
rect 1708 1660 1748 1700
rect 2092 1660 2132 1700
rect 2476 1660 2516 1700
rect 4492 1660 4532 1700
rect 4876 1660 4916 1700
rect 6220 1660 6260 1700
rect 8524 1660 8564 1700
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
<< metal2 >>
rect 1784 10672 1864 10752
rect 1976 10672 2056 10752
rect 2168 10672 2248 10752
rect 2360 10672 2440 10752
rect 2552 10672 2632 10752
rect 2744 10672 2824 10752
rect 2936 10672 3016 10752
rect 3128 10672 3208 10752
rect 3320 10672 3400 10752
rect 3512 10672 3592 10752
rect 3704 10672 3784 10752
rect 3896 10672 3976 10752
rect 4088 10672 4168 10752
rect 4280 10672 4360 10752
rect 4472 10672 4552 10752
rect 4664 10672 4744 10752
rect 4856 10672 4936 10752
rect 5048 10672 5128 10752
rect 5240 10672 5320 10752
rect 5432 10672 5512 10752
rect 5624 10672 5704 10752
rect 5816 10688 5896 10752
rect 5816 10672 5836 10688
rect 1611 9176 1653 9185
rect 1611 9136 1612 9176
rect 1652 9136 1653 9176
rect 1611 9127 1653 9136
rect 1612 7925 1652 9127
rect 1804 9008 1844 10672
rect 1708 8968 1844 9008
rect 1708 8513 1748 8968
rect 1996 8840 2036 10672
rect 2188 9008 2228 10672
rect 2188 8968 2324 9008
rect 2188 8840 2228 8849
rect 1996 8800 2188 8840
rect 2188 8791 2228 8800
rect 1804 8756 1844 8765
rect 1707 8504 1749 8513
rect 1707 8464 1708 8504
rect 1748 8464 1749 8504
rect 1707 8455 1749 8464
rect 1611 7916 1653 7925
rect 1611 7876 1612 7916
rect 1652 7876 1653 7916
rect 1611 7867 1653 7876
rect 1804 7085 1844 8716
rect 1899 8672 1941 8681
rect 1899 8632 1900 8672
rect 1940 8632 1941 8672
rect 1899 8623 1941 8632
rect 1900 8084 1940 8623
rect 1996 8504 2036 8513
rect 2284 8504 2324 8968
rect 2380 8924 2420 10672
rect 2380 8884 2516 8924
rect 2036 8464 2324 8504
rect 2380 8756 2420 8765
rect 1996 8455 2036 8464
rect 2091 8168 2133 8177
rect 2091 8128 2092 8168
rect 2132 8128 2133 8168
rect 2091 8119 2133 8128
rect 1900 8044 2036 8084
rect 1899 7916 1941 7925
rect 1899 7876 1900 7916
rect 1940 7876 1941 7916
rect 1899 7867 1941 7876
rect 1900 7782 1940 7867
rect 1996 7412 2036 8044
rect 2092 8034 2132 8119
rect 2092 7412 2132 7421
rect 1996 7372 2092 7412
rect 2092 7363 2132 7372
rect 1899 7244 1941 7253
rect 1899 7204 1900 7244
rect 1940 7204 1941 7244
rect 1899 7195 1941 7204
rect 1900 7110 1940 7195
rect 1803 7076 1845 7085
rect 1803 7036 1804 7076
rect 1844 7036 1845 7076
rect 1803 7027 1845 7036
rect 2380 6917 2420 8716
rect 2476 8177 2516 8884
rect 2572 8681 2612 10672
rect 2764 8924 2804 10672
rect 2859 10268 2901 10277
rect 2859 10228 2860 10268
rect 2900 10228 2901 10268
rect 2859 10219 2901 10228
rect 2668 8884 2804 8924
rect 2571 8672 2613 8681
rect 2571 8632 2572 8672
rect 2612 8632 2613 8672
rect 2571 8623 2613 8632
rect 2571 8504 2613 8513
rect 2571 8464 2572 8504
rect 2612 8464 2613 8504
rect 2571 8455 2613 8464
rect 2572 8370 2612 8455
rect 2475 8168 2517 8177
rect 2475 8128 2476 8168
rect 2516 8128 2517 8168
rect 2668 8168 2708 8884
rect 2764 8756 2804 8765
rect 2860 8756 2900 10219
rect 2804 8716 2900 8756
rect 2764 8707 2804 8716
rect 2764 8168 2804 8177
rect 2668 8128 2764 8168
rect 2475 8119 2517 8128
rect 2764 8119 2804 8128
rect 2956 8000 2996 10672
rect 3148 8177 3188 10672
rect 3340 9680 3380 10672
rect 3435 10352 3477 10361
rect 3435 10312 3436 10352
rect 3476 10312 3477 10352
rect 3435 10303 3477 10312
rect 3244 9640 3380 9680
rect 3244 8513 3284 9640
rect 3243 8504 3285 8513
rect 3243 8464 3244 8504
rect 3284 8464 3285 8504
rect 3243 8455 3285 8464
rect 3147 8168 3189 8177
rect 3147 8128 3148 8168
rect 3188 8128 3189 8168
rect 3147 8119 3189 8128
rect 3340 8168 3380 8177
rect 3340 8000 3380 8128
rect 2956 7960 3380 8000
rect 2572 7916 2612 7925
rect 3436 7916 3476 10303
rect 3532 8849 3572 10672
rect 3724 10613 3764 10672
rect 3723 10604 3765 10613
rect 3723 10564 3724 10604
rect 3764 10564 3765 10604
rect 3723 10555 3765 10564
rect 3916 9269 3956 10672
rect 3915 9260 3957 9269
rect 3915 9220 3916 9260
rect 3956 9220 3957 9260
rect 3915 9211 3957 9220
rect 3688 9092 4056 9101
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 3688 9043 4056 9052
rect 3531 8840 3573 8849
rect 3531 8800 3532 8840
rect 3572 8800 3573 8840
rect 3531 8791 3573 8800
rect 4108 8765 4148 10672
rect 4203 9596 4245 9605
rect 4203 9556 4204 9596
rect 4244 9556 4245 9596
rect 4203 9547 4245 9556
rect 4107 8756 4149 8765
rect 4107 8716 4108 8756
rect 4148 8716 4149 8756
rect 4107 8707 4149 8716
rect 4107 8168 4149 8177
rect 4107 8128 4108 8168
rect 4148 8128 4149 8168
rect 4107 8119 4149 8128
rect 4108 8034 4148 8119
rect 3532 7916 3572 7925
rect 3436 7876 3532 7916
rect 4204 7916 4244 9547
rect 4300 8681 4340 10672
rect 4395 8840 4437 8849
rect 4395 8800 4396 8840
rect 4436 8800 4437 8840
rect 4395 8791 4437 8800
rect 4396 8706 4436 8791
rect 4299 8672 4341 8681
rect 4299 8632 4300 8672
rect 4340 8632 4341 8672
rect 4299 8623 4341 8632
rect 4492 8597 4532 10672
rect 4588 8756 4628 8765
rect 4491 8588 4533 8597
rect 4491 8548 4492 8588
rect 4532 8548 4533 8588
rect 4491 8539 4533 8548
rect 4588 8177 4628 8716
rect 4684 8261 4724 10672
rect 4876 10025 4916 10672
rect 5068 10193 5108 10672
rect 5067 10184 5109 10193
rect 5067 10144 5068 10184
rect 5108 10144 5109 10184
rect 5067 10135 5109 10144
rect 5260 10109 5300 10672
rect 5355 10436 5397 10445
rect 5355 10396 5356 10436
rect 5396 10396 5397 10436
rect 5355 10387 5397 10396
rect 5259 10100 5301 10109
rect 5259 10060 5260 10100
rect 5300 10060 5301 10100
rect 5259 10051 5301 10060
rect 4875 10016 4917 10025
rect 4875 9976 4876 10016
rect 4916 9976 4917 10016
rect 4875 9967 4917 9976
rect 4928 9848 5296 9857
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 4928 9799 5296 9808
rect 4971 9680 5013 9689
rect 4971 9640 4972 9680
rect 5012 9640 5013 9680
rect 4971 9631 5013 9640
rect 4972 8756 5012 9631
rect 5164 8840 5204 8851
rect 5164 8765 5204 8800
rect 4972 8707 5012 8716
rect 5163 8756 5205 8765
rect 5163 8716 5164 8756
rect 5204 8716 5205 8756
rect 5163 8707 5205 8716
rect 5356 8756 5396 10387
rect 5452 9185 5492 10672
rect 5547 10184 5589 10193
rect 5547 10144 5548 10184
rect 5588 10144 5589 10184
rect 5547 10135 5589 10144
rect 5451 9176 5493 9185
rect 5451 9136 5452 9176
rect 5492 9136 5493 9176
rect 5451 9127 5493 9136
rect 5548 8765 5588 10135
rect 5644 9848 5684 10672
rect 5835 10648 5836 10672
rect 5876 10672 5896 10688
rect 6008 10672 6088 10752
rect 6200 10672 6280 10752
rect 6392 10672 6472 10752
rect 6584 10672 6664 10752
rect 6776 10672 6856 10752
rect 6968 10672 7048 10752
rect 7160 10672 7240 10752
rect 7352 10672 7432 10752
rect 7544 10672 7624 10752
rect 7736 10672 7816 10752
rect 7928 10672 8008 10752
rect 8120 10672 8200 10752
rect 8312 10672 8392 10752
rect 8504 10672 8584 10752
rect 8696 10672 8776 10752
rect 8888 10672 8968 10752
rect 9080 10672 9160 10752
rect 9272 10672 9352 10752
rect 9464 10672 9544 10752
rect 9656 10672 9736 10752
rect 9848 10672 9928 10752
rect 10040 10672 10120 10752
rect 10232 10688 10312 10752
rect 10166 10672 10312 10688
rect 10424 10672 10504 10752
rect 10616 10672 10696 10752
rect 10808 10672 10888 10752
rect 11000 10672 11080 10752
rect 11192 10672 11272 10752
rect 11384 10672 11464 10752
rect 11576 10672 11656 10752
rect 11768 10672 11848 10752
rect 11960 10672 12040 10752
rect 12152 10672 12232 10752
rect 12344 10672 12424 10752
rect 12536 10672 12616 10752
rect 12728 10672 12808 10752
rect 12920 10672 13000 10752
rect 13112 10672 13192 10752
rect 13304 10672 13384 10752
rect 13496 10672 13576 10752
rect 13688 10672 13768 10752
rect 13880 10672 13960 10752
rect 14072 10672 14152 10752
rect 14264 10672 14344 10752
rect 14456 10672 14536 10752
rect 14648 10672 14728 10752
rect 14840 10672 14920 10752
rect 15032 10672 15112 10752
rect 15224 10672 15304 10752
rect 15416 10672 15496 10752
rect 15608 10672 15688 10752
rect 15800 10672 15880 10752
rect 15992 10672 16072 10752
rect 16184 10672 16264 10752
rect 16376 10672 16456 10752
rect 16568 10672 16648 10752
rect 16760 10672 16840 10752
rect 16952 10672 17032 10752
rect 17144 10672 17224 10752
rect 17336 10672 17416 10752
rect 17528 10672 17608 10752
rect 17720 10672 17800 10752
rect 17912 10672 17992 10752
rect 18104 10672 18184 10752
rect 18296 10672 18376 10752
rect 18488 10672 18568 10752
rect 18680 10672 18760 10752
rect 18872 10672 18952 10752
rect 19064 10672 19144 10752
rect 19256 10672 19336 10752
rect 19448 10688 19528 10752
rect 19660 10697 19892 10732
rect 19448 10672 19468 10688
rect 5876 10648 5877 10672
rect 5835 10639 5877 10648
rect 5835 9932 5877 9941
rect 5835 9892 5836 9932
rect 5876 9892 5877 9932
rect 5835 9883 5877 9892
rect 5644 9808 5780 9848
rect 5740 8933 5780 9808
rect 5739 8924 5781 8933
rect 5739 8884 5740 8924
rect 5780 8884 5781 8924
rect 5739 8875 5781 8884
rect 5644 8840 5684 8849
rect 5356 8707 5396 8716
rect 5547 8756 5589 8765
rect 5547 8716 5548 8756
rect 5588 8716 5589 8756
rect 5547 8707 5589 8716
rect 5644 8681 5684 8800
rect 5836 8756 5876 9883
rect 5836 8707 5876 8716
rect 5643 8672 5685 8681
rect 5643 8632 5644 8672
rect 5684 8632 5685 8672
rect 5643 8623 5685 8632
rect 4779 8504 4821 8513
rect 4779 8464 4780 8504
rect 4820 8464 4821 8504
rect 4779 8455 4821 8464
rect 4780 8370 4820 8455
rect 4928 8336 5296 8345
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 4928 8287 5296 8296
rect 4683 8252 4725 8261
rect 4683 8212 4684 8252
rect 4724 8212 4725 8252
rect 4683 8203 4725 8212
rect 4587 8168 4629 8177
rect 4587 8128 4588 8168
rect 4628 8128 4629 8168
rect 4587 8119 4629 8128
rect 4300 7916 4340 7925
rect 4204 7876 4300 7916
rect 2572 7001 2612 7876
rect 3532 7867 3572 7876
rect 4300 7867 4340 7876
rect 3688 7580 4056 7589
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 3688 7531 4056 7540
rect 6028 7505 6068 10672
rect 6123 8588 6165 8597
rect 6123 8548 6124 8588
rect 6164 8548 6165 8588
rect 6123 8539 6165 8548
rect 6124 8504 6164 8539
rect 6124 8453 6164 8464
rect 6027 7496 6069 7505
rect 6027 7456 6028 7496
rect 6068 7456 6069 7496
rect 6027 7447 6069 7456
rect 2571 6992 2613 7001
rect 2571 6952 2572 6992
rect 2612 6952 2613 6992
rect 2571 6943 2613 6952
rect 2379 6908 2421 6917
rect 2379 6868 2380 6908
rect 2420 6868 2421 6908
rect 2379 6859 2421 6868
rect 4928 6824 5296 6833
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 4928 6775 5296 6784
rect 1227 6488 1269 6497
rect 1227 6448 1228 6488
rect 1268 6448 1269 6488
rect 1227 6439 1269 6448
rect 1228 5993 1268 6439
rect 1996 6404 2036 6413
rect 1996 6161 2036 6364
rect 6220 6245 6260 10672
rect 6316 8756 6356 8765
rect 6316 8345 6356 8716
rect 6315 8336 6357 8345
rect 6315 8296 6316 8336
rect 6356 8296 6357 8336
rect 6315 8287 6357 8296
rect 6412 7421 6452 10672
rect 6604 10529 6644 10672
rect 6603 10520 6645 10529
rect 6603 10480 6604 10520
rect 6644 10480 6645 10520
rect 6603 10471 6645 10480
rect 6796 10193 6836 10672
rect 6795 10184 6837 10193
rect 6795 10144 6796 10184
rect 6836 10144 6837 10184
rect 6795 10135 6837 10144
rect 6411 7412 6453 7421
rect 6411 7372 6412 7412
rect 6452 7372 6453 7412
rect 6411 7363 6453 7372
rect 6988 7337 7028 10672
rect 7083 10016 7125 10025
rect 7083 9976 7084 10016
rect 7124 9976 7125 10016
rect 7083 9967 7125 9976
rect 7084 8840 7124 9967
rect 7084 8791 7124 8800
rect 7180 8513 7220 10672
rect 7275 8756 7317 8765
rect 7275 8716 7276 8756
rect 7316 8716 7317 8756
rect 7275 8707 7317 8716
rect 7276 8622 7316 8707
rect 7372 8597 7412 10672
rect 7564 9521 7604 10672
rect 7659 9764 7701 9773
rect 7659 9724 7660 9764
rect 7700 9724 7701 9764
rect 7659 9715 7701 9724
rect 7563 9512 7605 9521
rect 7563 9472 7564 9512
rect 7604 9472 7605 9512
rect 7563 9463 7605 9472
rect 7467 8840 7509 8849
rect 7467 8800 7468 8840
rect 7508 8800 7509 8840
rect 7467 8791 7509 8800
rect 7468 8706 7508 8791
rect 7660 8756 7700 9715
rect 7660 8707 7700 8716
rect 7371 8588 7413 8597
rect 7371 8548 7372 8588
rect 7412 8548 7413 8588
rect 7371 8539 7413 8548
rect 7179 8504 7221 8513
rect 7179 8464 7180 8504
rect 7220 8464 7221 8504
rect 7179 8455 7221 8464
rect 7083 8252 7125 8261
rect 7083 8212 7084 8252
rect 7124 8212 7125 8252
rect 7083 8203 7125 8212
rect 7084 8168 7124 8203
rect 7084 8117 7124 8128
rect 7660 8168 7700 8177
rect 7756 8168 7796 10672
rect 7851 9428 7893 9437
rect 7851 9388 7852 9428
rect 7892 9388 7893 9428
rect 7851 9379 7893 9388
rect 7700 8128 7796 8168
rect 7660 8119 7700 8128
rect 7275 7916 7317 7925
rect 7275 7876 7276 7916
rect 7316 7876 7317 7916
rect 7275 7867 7317 7876
rect 7852 7916 7892 9379
rect 7948 8168 7988 10672
rect 8043 9260 8085 9269
rect 8043 9220 8044 9260
rect 8084 9220 8085 9260
rect 8043 9211 8085 9220
rect 8044 8840 8084 9211
rect 8044 8791 8084 8800
rect 8140 8177 8180 10672
rect 8235 8756 8277 8765
rect 8235 8716 8236 8756
rect 8276 8716 8277 8756
rect 8235 8707 8277 8716
rect 8236 8622 8276 8707
rect 8332 8261 8372 10672
rect 8427 10604 8469 10613
rect 8427 10564 8428 10604
rect 8468 10564 8469 10604
rect 8427 10555 8469 10564
rect 8331 8252 8373 8261
rect 8331 8212 8332 8252
rect 8372 8212 8373 8252
rect 8331 8203 8373 8212
rect 8044 8168 8084 8177
rect 7948 8128 8044 8168
rect 8044 8119 8084 8128
rect 8139 8168 8181 8177
rect 8139 8128 8140 8168
rect 8180 8128 8181 8168
rect 8139 8119 8181 8128
rect 8428 8168 8468 10555
rect 8524 8849 8564 10672
rect 8619 9344 8661 9353
rect 8619 9304 8620 9344
rect 8660 9304 8661 9344
rect 8619 9295 8661 9304
rect 8523 8840 8565 8849
rect 8523 8800 8524 8840
rect 8564 8800 8565 8840
rect 8523 8791 8565 8800
rect 8620 8672 8660 9295
rect 8716 9101 8756 10672
rect 8715 9092 8757 9101
rect 8715 9052 8716 9092
rect 8756 9052 8757 9092
rect 8715 9043 8757 9052
rect 8428 8119 8468 8128
rect 8524 8632 8660 8672
rect 7852 7867 7892 7876
rect 8236 7916 8276 7925
rect 8524 7916 8564 8632
rect 8276 7876 8564 7916
rect 8619 7916 8661 7925
rect 8619 7876 8620 7916
rect 8660 7876 8661 7916
rect 8236 7867 8276 7876
rect 8619 7867 8661 7876
rect 7276 7782 7316 7867
rect 8620 7782 8660 7867
rect 6987 7328 7029 7337
rect 6987 7288 6988 7328
rect 7028 7288 7029 7328
rect 6987 7279 7029 7288
rect 8908 7085 8948 10672
rect 8907 7076 8949 7085
rect 8907 7036 8908 7076
rect 8948 7036 8949 7076
rect 8907 7027 8949 7036
rect 9100 6917 9140 10672
rect 9292 10277 9332 10672
rect 9291 10268 9333 10277
rect 9291 10228 9292 10268
rect 9332 10228 9333 10268
rect 9291 10219 9333 10228
rect 9484 8765 9524 10672
rect 9483 8756 9525 8765
rect 9483 8716 9484 8756
rect 9524 8716 9525 8756
rect 9483 8707 9525 8716
rect 9483 8420 9525 8429
rect 9483 8380 9484 8420
rect 9524 8380 9525 8420
rect 9483 8371 9525 8380
rect 9099 6908 9141 6917
rect 9099 6868 9100 6908
rect 9140 6868 9141 6908
rect 9099 6859 9141 6868
rect 9484 6320 9524 8371
rect 9579 8168 9621 8177
rect 9579 8128 9580 8168
rect 9620 8128 9621 8168
rect 9579 8119 9621 8128
rect 9580 8034 9620 8119
rect 9676 7925 9716 10672
rect 9771 9848 9813 9857
rect 9771 9808 9772 9848
rect 9812 9808 9813 9848
rect 9771 9799 9813 9808
rect 9675 7916 9717 7925
rect 9675 7876 9676 7916
rect 9716 7876 9717 7916
rect 9675 7867 9717 7876
rect 9772 7916 9812 9799
rect 9868 8093 9908 10672
rect 10060 9689 10100 10672
rect 10166 10648 10292 10672
rect 10166 10604 10206 10648
rect 10156 10564 10206 10604
rect 10059 9680 10101 9689
rect 10059 9640 10060 9680
rect 10100 9640 10101 9680
rect 10059 9631 10101 9640
rect 10156 9605 10196 10564
rect 10444 10361 10484 10672
rect 10443 10352 10485 10361
rect 10443 10312 10444 10352
rect 10484 10312 10485 10352
rect 10443 10303 10485 10312
rect 10251 9680 10293 9689
rect 10251 9640 10252 9680
rect 10292 9640 10293 9680
rect 10251 9631 10293 9640
rect 10155 9596 10197 9605
rect 10155 9556 10156 9596
rect 10196 9556 10197 9596
rect 10155 9547 10197 9556
rect 10155 9260 10197 9269
rect 10155 9220 10156 9260
rect 10196 9220 10197 9260
rect 10155 9211 10197 9220
rect 10059 9176 10101 9185
rect 10059 9136 10060 9176
rect 10100 9136 10101 9176
rect 10059 9127 10101 9136
rect 9963 9092 10005 9101
rect 9963 9052 9964 9092
rect 10004 9052 10005 9092
rect 9963 9043 10005 9052
rect 9964 8420 10004 9043
rect 10060 8840 10100 9127
rect 10060 8791 10100 8800
rect 9964 8380 10100 8420
rect 9963 8252 10005 8261
rect 9963 8212 9964 8252
rect 10004 8212 10005 8252
rect 9963 8203 10005 8212
rect 9964 8168 10004 8203
rect 9964 8117 10004 8128
rect 9867 8084 9909 8093
rect 9867 8044 9868 8084
rect 9908 8044 9909 8084
rect 9867 8035 9909 8044
rect 9772 7867 9812 7876
rect 10060 6320 10100 8380
rect 10156 7916 10196 9211
rect 10252 8756 10292 9631
rect 10636 9008 10676 10672
rect 10828 10520 10868 10672
rect 10252 8707 10292 8716
rect 10540 8968 10676 9008
rect 10732 10480 10868 10520
rect 10156 7867 10196 7876
rect 10540 7001 10580 8968
rect 10635 8840 10677 8849
rect 10635 8800 10636 8840
rect 10676 8800 10677 8840
rect 10635 8791 10677 8800
rect 10636 8706 10676 8791
rect 10732 7253 10772 10480
rect 11020 9689 11060 10672
rect 11212 9764 11252 10672
rect 11404 9773 11444 10672
rect 11499 10100 11541 10109
rect 11499 10060 11500 10100
rect 11540 10060 11541 10100
rect 11499 10051 11541 10060
rect 11403 9764 11445 9773
rect 11212 9724 11348 9764
rect 11019 9680 11061 9689
rect 11019 9640 11020 9680
rect 11060 9640 11061 9680
rect 11019 9631 11061 9640
rect 11211 9596 11253 9605
rect 11211 9556 11212 9596
rect 11252 9556 11253 9596
rect 11211 9547 11253 9556
rect 11019 9512 11061 9521
rect 11019 9472 11020 9512
rect 11060 9472 11061 9512
rect 11019 9463 11061 9472
rect 11020 8840 11060 9463
rect 11020 8791 11060 8800
rect 10827 8756 10869 8765
rect 10827 8716 10828 8756
rect 10868 8716 10869 8756
rect 10827 8707 10869 8716
rect 11212 8756 11252 9547
rect 11308 8756 11348 9724
rect 11403 9724 11404 9764
rect 11444 9724 11445 9764
rect 11403 9715 11445 9724
rect 11404 8924 11444 8933
rect 11500 8924 11540 10051
rect 11596 9764 11636 10672
rect 11596 9724 11732 9764
rect 11444 8884 11540 8924
rect 11404 8875 11444 8884
rect 11596 8756 11636 8765
rect 11308 8716 11596 8756
rect 11212 8707 11252 8716
rect 11596 8707 11636 8716
rect 10828 8622 10868 8707
rect 11692 8681 11732 9724
rect 11788 8849 11828 10672
rect 11980 10648 12030 10672
rect 11990 10520 12030 10648
rect 11884 10480 12030 10520
rect 11787 8840 11829 8849
rect 11787 8800 11788 8840
rect 11828 8800 11829 8840
rect 11787 8791 11829 8800
rect 11691 8672 11733 8681
rect 11691 8632 11692 8672
rect 11732 8632 11733 8672
rect 11691 8623 11733 8632
rect 11403 8588 11445 8597
rect 11403 8548 11404 8588
rect 11444 8548 11445 8588
rect 11403 8539 11445 8548
rect 11595 8588 11637 8597
rect 11595 8548 11596 8588
rect 11636 8548 11637 8588
rect 11595 8539 11637 8548
rect 11404 8168 11444 8539
rect 11404 8119 11444 8128
rect 11596 7916 11636 8539
rect 11787 8504 11829 8513
rect 11787 8464 11788 8504
rect 11828 8464 11829 8504
rect 11787 8455 11829 8464
rect 11788 8370 11828 8455
rect 11884 8345 11924 10480
rect 12172 9941 12212 10672
rect 12364 10445 12404 10672
rect 12363 10436 12405 10445
rect 12363 10396 12364 10436
rect 12404 10396 12405 10436
rect 12363 10387 12405 10396
rect 12171 9932 12213 9941
rect 12171 9892 12172 9932
rect 12212 9892 12213 9932
rect 12171 9883 12213 9892
rect 11979 9764 12021 9773
rect 11979 9724 11980 9764
rect 12020 9724 12021 9764
rect 11979 9715 12021 9724
rect 11980 8756 12020 9715
rect 12075 8840 12117 8849
rect 12075 8800 12076 8840
rect 12116 8800 12117 8840
rect 12075 8791 12117 8800
rect 11980 8707 12020 8716
rect 11883 8336 11925 8345
rect 11883 8296 11884 8336
rect 11924 8296 11925 8336
rect 11883 8287 11925 8296
rect 12076 8009 12116 8791
rect 12556 8765 12596 10672
rect 12748 9269 12788 10672
rect 12940 9857 12980 10672
rect 12939 9848 12981 9857
rect 12939 9808 12940 9848
rect 12980 9808 12981 9848
rect 12939 9799 12981 9808
rect 13132 9353 13172 10672
rect 13227 10184 13269 10193
rect 13227 10144 13228 10184
rect 13268 10144 13269 10184
rect 13227 10135 13269 10144
rect 13131 9344 13173 9353
rect 13131 9304 13132 9344
rect 13172 9304 13173 9344
rect 13131 9295 13173 9304
rect 12747 9260 12789 9269
rect 12747 9220 12748 9260
rect 12788 9220 12789 9260
rect 12747 9211 12789 9220
rect 12555 8756 12597 8765
rect 12555 8716 12556 8756
rect 12596 8716 12597 8756
rect 12555 8707 12597 8716
rect 13228 8168 13268 10135
rect 13324 9437 13364 10672
rect 13516 9605 13556 10672
rect 13611 10520 13653 10529
rect 13611 10480 13612 10520
rect 13652 10480 13653 10520
rect 13611 10471 13653 10480
rect 13515 9596 13557 9605
rect 13515 9556 13516 9596
rect 13556 9556 13557 9596
rect 13515 9547 13557 9556
rect 13323 9428 13365 9437
rect 13323 9388 13324 9428
rect 13364 9388 13365 9428
rect 13323 9379 13365 9388
rect 13419 8840 13461 8849
rect 13419 8800 13420 8840
rect 13460 8800 13461 8840
rect 13419 8791 13461 8800
rect 13228 8119 13268 8128
rect 13323 8168 13365 8177
rect 13323 8128 13324 8168
rect 13364 8128 13365 8168
rect 13323 8119 13365 8128
rect 12075 8000 12117 8009
rect 12075 7960 12076 8000
rect 12116 7960 12117 8000
rect 12075 7951 12117 7960
rect 11596 7867 11636 7876
rect 12939 7916 12981 7925
rect 12939 7876 12940 7916
rect 12980 7876 12981 7916
rect 12939 7867 12981 7876
rect 12940 7782 12980 7867
rect 12748 7748 12788 7757
rect 10827 7580 10869 7589
rect 10827 7540 10828 7580
rect 10868 7540 10869 7580
rect 10827 7531 10869 7540
rect 10731 7244 10773 7253
rect 10731 7204 10732 7244
rect 10772 7204 10773 7244
rect 10731 7195 10773 7204
rect 10539 6992 10581 7001
rect 10539 6952 10540 6992
rect 10580 6952 10581 6992
rect 10539 6943 10581 6952
rect 9484 6280 9620 6320
rect 2187 6236 2229 6245
rect 2187 6196 2188 6236
rect 2228 6196 2229 6236
rect 2187 6187 2229 6196
rect 6219 6236 6261 6245
rect 6219 6196 6220 6236
rect 6260 6196 6261 6236
rect 6219 6187 6261 6196
rect 1995 6152 2037 6161
rect 1995 6112 1996 6152
rect 2036 6112 2037 6152
rect 1995 6103 2037 6112
rect 2188 6102 2228 6187
rect 3688 6068 4056 6077
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 3688 6019 4056 6028
rect 1227 5984 1269 5993
rect 1227 5944 1228 5984
rect 1268 5944 1269 5984
rect 1227 5935 1269 5944
rect 459 5816 501 5825
rect 459 5776 460 5816
rect 500 5776 501 5816
rect 459 5767 501 5776
rect 460 4229 500 5767
rect 6603 5648 6645 5657
rect 6603 5608 6604 5648
rect 6644 5608 6645 5648
rect 6603 5599 6645 5608
rect 4928 5312 5296 5321
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 4928 5263 5296 5272
rect 2283 5144 2325 5153
rect 2283 5104 2284 5144
rect 2324 5104 2325 5144
rect 2283 5095 2325 5104
rect 2475 5144 2517 5153
rect 2475 5104 2476 5144
rect 2516 5104 2517 5144
rect 2475 5095 2517 5104
rect 2284 4892 2324 5095
rect 2284 4843 2324 4852
rect 2476 4808 2516 5095
rect 2476 4759 2516 4768
rect 2283 4724 2325 4733
rect 2283 4684 2284 4724
rect 2324 4684 2325 4724
rect 2283 4675 2325 4684
rect 459 4220 501 4229
rect 459 4180 460 4220
rect 500 4180 501 4220
rect 459 4171 501 4180
rect 1900 4220 1940 4229
rect 1900 3137 1940 4180
rect 2284 4220 2324 4675
rect 3688 4556 4056 4565
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 3688 4507 4056 4516
rect 2667 4472 2709 4481
rect 2667 4432 2668 4472
rect 2708 4432 2709 4472
rect 2667 4423 2709 4432
rect 2284 4171 2324 4180
rect 2668 4220 2708 4423
rect 5835 4388 5877 4397
rect 5835 4348 5836 4388
rect 5876 4348 5877 4388
rect 5835 4339 5877 4348
rect 2668 4171 2708 4180
rect 2092 3968 2132 3977
rect 2092 3305 2132 3928
rect 2475 3968 2517 3977
rect 2475 3928 2476 3968
rect 2516 3928 2517 3968
rect 2475 3919 2517 3928
rect 2860 3968 2900 3977
rect 2900 3928 3188 3968
rect 2860 3919 2900 3928
rect 2476 3834 2516 3919
rect 3148 3884 3188 3928
rect 3243 3884 3285 3893
rect 3148 3844 3244 3884
rect 3284 3844 3285 3884
rect 3243 3835 3285 3844
rect 4928 3800 5296 3809
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 4928 3751 5296 3760
rect 2188 3380 2228 3389
rect 2091 3296 2133 3305
rect 2091 3256 2092 3296
rect 2132 3256 2133 3296
rect 2091 3247 2133 3256
rect 1899 3128 1941 3137
rect 1899 3088 1900 3128
rect 1940 3088 1941 3128
rect 1899 3079 1941 3088
rect 2188 2465 2228 3340
rect 2380 3212 2420 3221
rect 2380 2969 2420 3172
rect 3435 3128 3477 3137
rect 3435 3088 3436 3128
rect 3476 3088 3477 3128
rect 3435 3079 3477 3088
rect 2379 2960 2421 2969
rect 2379 2920 2380 2960
rect 2420 2920 2421 2960
rect 2379 2911 2421 2920
rect 2187 2456 2229 2465
rect 2187 2416 2188 2456
rect 2228 2416 2229 2456
rect 2187 2407 2229 2416
rect 3436 2120 3476 3079
rect 3688 3044 4056 3053
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 3688 2995 4056 3004
rect 4928 2288 5296 2297
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 4928 2239 5296 2248
rect 4107 2204 4149 2213
rect 4107 2164 4108 2204
rect 4148 2164 4149 2204
rect 4107 2155 4149 2164
rect 3436 2071 3476 2080
rect 4108 2120 4148 2155
rect 4108 2069 4148 2080
rect 5836 2120 5876 4339
rect 5836 2071 5876 2080
rect 6027 2120 6069 2129
rect 6027 2080 6028 2120
rect 6068 2080 6069 2120
rect 6027 2071 6069 2080
rect 6604 2120 6644 5599
rect 9483 4892 9525 4901
rect 9483 4852 9484 4892
rect 9524 4852 9525 4892
rect 9483 4843 9525 4852
rect 9484 4758 9524 4843
rect 9580 4808 9620 6280
rect 9868 6280 10100 6320
rect 9676 4808 9716 4817
rect 9580 4768 9676 4808
rect 9676 4759 9716 4768
rect 9772 4220 9812 4229
rect 9772 3473 9812 4180
rect 9771 3464 9813 3473
rect 9771 3424 9772 3464
rect 9812 3424 9813 3464
rect 9771 3415 9813 3424
rect 6987 3380 7029 3389
rect 6987 3340 6988 3380
rect 7028 3340 7029 3380
rect 6987 3331 7029 3340
rect 6988 2213 7028 3331
rect 6987 2204 7029 2213
rect 6987 2164 6988 2204
rect 7028 2164 7029 2204
rect 6987 2155 7029 2164
rect 9868 2120 9908 6280
rect 9964 3968 10004 3977
rect 9964 3473 10004 3928
rect 9963 3464 10005 3473
rect 9963 3424 9964 3464
rect 10004 3424 10005 3464
rect 9963 3415 10005 3424
rect 10059 2624 10101 2633
rect 10059 2584 10060 2624
rect 10100 2584 10101 2624
rect 10059 2575 10101 2584
rect 9964 2120 10004 2129
rect 9868 2080 9964 2120
rect 6604 2071 6644 2080
rect 9964 2071 10004 2080
rect 1035 1868 1077 1877
rect 1035 1828 1036 1868
rect 1076 1828 1077 1868
rect 1035 1819 1077 1828
rect 1516 1868 1556 1877
rect 1036 80 1076 1819
rect 1516 449 1556 1828
rect 1900 1868 1940 1877
rect 1708 1700 1748 1709
rect 1708 449 1748 1660
rect 1515 440 1557 449
rect 1515 400 1516 440
rect 1556 400 1557 440
rect 1515 391 1557 400
rect 1707 440 1749 449
rect 1707 400 1708 440
rect 1748 400 1749 440
rect 1707 391 1749 400
rect 1900 197 1940 1828
rect 2284 1868 2324 1877
rect 2091 1700 2133 1709
rect 2091 1660 2092 1700
rect 2132 1660 2133 1700
rect 2091 1651 2133 1660
rect 2092 1566 2132 1651
rect 2284 1457 2324 1828
rect 3243 1868 3285 1877
rect 3243 1828 3244 1868
rect 3284 1828 3285 1868
rect 3243 1819 3285 1828
rect 3916 1868 3956 1877
rect 4300 1868 4340 1877
rect 3956 1828 4244 1868
rect 3916 1819 3956 1828
rect 3244 1734 3284 1819
rect 2476 1700 2516 1709
rect 2476 1457 2516 1660
rect 3531 1700 3573 1709
rect 3531 1660 3532 1700
rect 3572 1660 3573 1700
rect 3531 1651 3573 1660
rect 2283 1448 2325 1457
rect 2283 1408 2284 1448
rect 2324 1408 2325 1448
rect 2283 1399 2325 1408
rect 2475 1448 2517 1457
rect 2475 1408 2476 1448
rect 2516 1408 2517 1448
rect 2475 1399 2517 1408
rect 2955 1280 2997 1289
rect 2955 1240 2956 1280
rect 2996 1240 2997 1280
rect 2955 1231 2997 1240
rect 1995 944 2037 953
rect 1995 904 1996 944
rect 2036 904 2037 944
rect 1995 895 2037 904
rect 1899 188 1941 197
rect 1899 148 1900 188
rect 1940 148 1941 188
rect 1899 139 1941 148
rect 1996 80 2036 895
rect 2956 80 2996 1231
rect 3532 113 3572 1651
rect 3688 1532 4056 1541
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 3688 1483 4056 1492
rect 3915 1364 3957 1373
rect 3915 1324 3916 1364
rect 3956 1324 3957 1364
rect 3915 1315 3957 1324
rect 3531 104 3573 113
rect 1016 0 1096 80
rect 1976 0 2056 80
rect 2936 0 3016 80
rect 3531 64 3532 104
rect 3572 64 3573 104
rect 3916 80 3956 1315
rect 4204 953 4244 1828
rect 4300 1289 4340 1828
rect 4684 1868 4724 1877
rect 4491 1700 4533 1709
rect 4491 1660 4492 1700
rect 4532 1660 4533 1700
rect 4491 1651 4533 1660
rect 4492 1566 4532 1651
rect 4299 1280 4341 1289
rect 4299 1240 4300 1280
rect 4340 1240 4341 1280
rect 4299 1231 4341 1240
rect 4203 944 4245 953
rect 4203 904 4204 944
rect 4244 904 4245 944
rect 4203 895 4245 904
rect 4684 785 4724 1828
rect 5644 1868 5684 1877
rect 4876 1700 4916 1709
rect 4876 953 4916 1660
rect 5644 1373 5684 1828
rect 6028 1868 6068 2071
rect 6028 1819 6068 1828
rect 6412 1868 6452 1877
rect 6220 1700 6260 1709
rect 6220 1541 6260 1660
rect 6219 1532 6261 1541
rect 6219 1492 6220 1532
rect 6260 1492 6261 1532
rect 6219 1483 6261 1492
rect 5643 1364 5685 1373
rect 5643 1324 5644 1364
rect 5684 1324 5685 1364
rect 5643 1315 5685 1324
rect 4875 944 4917 953
rect 4875 904 4876 944
rect 4916 904 4917 944
rect 4875 895 4917 904
rect 4683 776 4725 785
rect 4683 736 4684 776
rect 4724 736 4725 776
rect 4683 727 4725 736
rect 4928 776 5296 785
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 4928 727 5296 736
rect 6412 365 6452 1828
rect 8332 1868 8372 1877
rect 8332 1121 8372 1828
rect 8715 1868 8757 1877
rect 8715 1828 8716 1868
rect 8756 1828 8757 1868
rect 8715 1819 8757 1828
rect 9771 1868 9813 1877
rect 9771 1828 9772 1868
rect 9812 1828 9813 1868
rect 9771 1819 9813 1828
rect 8524 1700 8564 1709
rect 8524 1121 8564 1660
rect 8331 1112 8373 1121
rect 8331 1072 8332 1112
rect 8372 1072 8373 1112
rect 8331 1063 8373 1072
rect 8523 1112 8565 1121
rect 8523 1072 8524 1112
rect 8564 1072 8565 1112
rect 8523 1063 8565 1072
rect 4875 356 4917 365
rect 4875 316 4876 356
rect 4916 316 4917 356
rect 4875 307 4917 316
rect 6411 356 6453 365
rect 6411 316 6412 356
rect 6452 316 6453 356
rect 6411 307 6453 316
rect 7755 356 7797 365
rect 7755 316 7756 356
rect 7796 316 7797 356
rect 7755 307 7797 316
rect 4876 80 4916 307
rect 6795 272 6837 281
rect 6795 232 6796 272
rect 6836 232 6837 272
rect 6795 223 6837 232
rect 5835 188 5877 197
rect 5835 148 5836 188
rect 5876 148 5877 188
rect 5835 139 5877 148
rect 5836 80 5876 139
rect 6796 80 6836 223
rect 7756 80 7796 307
rect 8716 80 8756 1819
rect 9772 1734 9812 1819
rect 10060 1709 10100 2575
rect 10732 2120 10772 2129
rect 10828 2120 10868 7531
rect 12748 7337 12788 7708
rect 12747 7328 12789 7337
rect 12747 7288 12748 7328
rect 12788 7288 12789 7328
rect 12747 7279 12789 7288
rect 12172 5732 12212 5741
rect 12172 5489 12212 5692
rect 12171 5480 12213 5489
rect 12171 5440 12172 5480
rect 12212 5440 12213 5480
rect 12171 5431 12213 5440
rect 12363 5480 12405 5489
rect 12363 5440 12364 5480
rect 12404 5440 12405 5480
rect 12363 5431 12405 5440
rect 12364 5346 12404 5431
rect 12940 4220 12980 4229
rect 12843 4136 12885 4145
rect 12940 4136 12980 4180
rect 12843 4096 12844 4136
rect 12884 4096 12980 4136
rect 13131 4136 13173 4145
rect 13131 4096 13132 4136
rect 13172 4096 13173 4136
rect 12843 4087 12885 4096
rect 13131 4087 13173 4096
rect 13132 3968 13172 4087
rect 13132 3919 13172 3928
rect 12075 3800 12117 3809
rect 12075 3760 12076 3800
rect 12116 3760 12117 3800
rect 12075 3751 12117 3760
rect 10772 2080 10868 2120
rect 12076 2120 12116 3751
rect 10732 2071 10772 2080
rect 12076 2071 12116 2080
rect 13228 2120 13268 2129
rect 13324 2120 13364 8119
rect 13420 7916 13460 8791
rect 13612 8168 13652 10471
rect 13708 8597 13748 10672
rect 13900 9773 13940 10672
rect 13899 9764 13941 9773
rect 13899 9724 13900 9764
rect 13940 9724 13941 9764
rect 13899 9715 13941 9724
rect 13707 8588 13749 8597
rect 13707 8548 13708 8588
rect 13748 8548 13749 8588
rect 13707 8539 13749 8548
rect 13708 8168 13748 8177
rect 13612 8128 13708 8168
rect 13708 8119 13748 8128
rect 14092 7925 14132 10672
rect 14284 8849 14324 10672
rect 14476 9344 14516 10672
rect 14380 9304 14516 9344
rect 14283 8840 14325 8849
rect 14283 8800 14284 8840
rect 14324 8800 14325 8840
rect 14283 8791 14325 8800
rect 14380 8672 14420 9304
rect 14476 8756 14516 8765
rect 14668 8756 14708 10672
rect 14516 8716 14708 8756
rect 14860 8756 14900 10672
rect 15052 8765 15092 10672
rect 15244 8849 15284 10672
rect 15436 9764 15476 10672
rect 15340 9724 15476 9764
rect 15243 8840 15285 8849
rect 15243 8800 15244 8840
rect 15284 8800 15285 8840
rect 15243 8791 15285 8800
rect 14476 8707 14516 8716
rect 14860 8707 14900 8716
rect 15051 8756 15093 8765
rect 15051 8716 15052 8756
rect 15092 8716 15093 8756
rect 15051 8707 15093 8716
rect 15340 8681 15380 9724
rect 15531 8924 15573 8933
rect 15531 8884 15532 8924
rect 15572 8884 15573 8924
rect 15531 8875 15573 8884
rect 15435 8756 15477 8765
rect 15435 8716 15436 8756
rect 15476 8716 15477 8756
rect 15435 8707 15477 8716
rect 14188 8632 14420 8672
rect 15339 8672 15381 8681
rect 15339 8632 15340 8672
rect 15380 8632 15381 8672
rect 13420 7867 13460 7876
rect 13900 7916 13940 7925
rect 14091 7916 14133 7925
rect 13940 7876 14036 7916
rect 13900 7867 13940 7876
rect 13996 7748 14036 7876
rect 14091 7876 14092 7916
rect 14132 7876 14133 7916
rect 14091 7867 14133 7876
rect 14188 7748 14228 8632
rect 15339 8623 15381 8632
rect 15436 8622 15476 8707
rect 13996 7708 14228 7748
rect 14284 8504 14324 8513
rect 14284 7421 14324 8464
rect 14668 8504 14708 8513
rect 14283 7412 14325 7421
rect 14283 7372 14284 7412
rect 14324 7372 14325 7412
rect 14283 7363 14325 7372
rect 14571 6572 14613 6581
rect 14571 6532 14572 6572
rect 14612 6532 14613 6572
rect 14571 6523 14613 6532
rect 14475 2708 14517 2717
rect 14475 2668 14476 2708
rect 14516 2668 14517 2708
rect 14475 2659 14517 2668
rect 14476 2574 14516 2659
rect 14572 2456 14612 6523
rect 14668 6245 14708 8464
rect 15244 8504 15284 8513
rect 14763 8336 14805 8345
rect 14763 8296 14764 8336
rect 14804 8296 14805 8336
rect 14763 8287 14805 8296
rect 14667 6236 14709 6245
rect 14667 6196 14668 6236
rect 14708 6196 14709 6236
rect 14667 6187 14709 6196
rect 14668 2792 14708 2801
rect 14668 2633 14708 2752
rect 14667 2624 14709 2633
rect 14667 2584 14668 2624
rect 14708 2584 14709 2624
rect 14667 2575 14709 2584
rect 13268 2080 13364 2120
rect 14476 2416 14612 2456
rect 13228 2071 13268 2080
rect 10540 1868 10580 1877
rect 10059 1700 10101 1709
rect 10059 1660 10060 1700
rect 10100 1660 10101 1700
rect 10059 1651 10101 1660
rect 10540 1289 10580 1828
rect 10635 1868 10677 1877
rect 10635 1828 10636 1868
rect 10676 1828 10677 1868
rect 10635 1819 10677 1828
rect 11883 1868 11925 1877
rect 11883 1828 11884 1868
rect 11924 1828 11925 1868
rect 11883 1819 11925 1828
rect 13036 1868 13076 1877
rect 9675 1280 9717 1289
rect 9675 1240 9676 1280
rect 9716 1240 9717 1280
rect 9675 1231 9717 1240
rect 10539 1280 10581 1289
rect 10539 1240 10540 1280
rect 10580 1240 10581 1280
rect 10539 1231 10581 1240
rect 9676 80 9716 1231
rect 10636 80 10676 1819
rect 11884 1734 11924 1819
rect 13036 1289 13076 1828
rect 13515 1868 13557 1877
rect 13515 1828 13516 1868
rect 13556 1828 13557 1868
rect 13515 1819 13557 1828
rect 14379 1868 14421 1877
rect 14379 1828 14380 1868
rect 14420 1828 14421 1868
rect 14379 1819 14421 1828
rect 11595 1280 11637 1289
rect 11595 1240 11596 1280
rect 11636 1240 11637 1280
rect 11595 1231 11637 1240
rect 13035 1280 13077 1289
rect 13035 1240 13036 1280
rect 13076 1240 13077 1280
rect 13035 1231 13077 1240
rect 11596 80 11636 1231
rect 12555 776 12597 785
rect 12555 736 12556 776
rect 12596 736 12597 776
rect 12555 727 12597 736
rect 12556 80 12596 727
rect 13516 80 13556 1819
rect 14380 1734 14420 1819
rect 14476 80 14516 2416
rect 14572 2120 14612 2129
rect 14764 2120 14804 8287
rect 15244 7505 15284 8464
rect 15243 7496 15285 7505
rect 15243 7456 15244 7496
rect 15284 7456 15285 7496
rect 15243 7447 15285 7456
rect 15339 7412 15381 7421
rect 15339 7372 15340 7412
rect 15380 7372 15381 7412
rect 15339 7363 15381 7372
rect 14612 2080 14804 2120
rect 15340 2120 15380 7363
rect 15532 2717 15572 8875
rect 15628 3137 15668 10672
rect 15723 8504 15765 8513
rect 15723 8464 15724 8504
rect 15764 8464 15765 8504
rect 15723 8455 15765 8464
rect 15724 4397 15764 8455
rect 15723 4388 15765 4397
rect 15723 4348 15724 4388
rect 15764 4348 15765 4388
rect 15723 4339 15765 4348
rect 15820 3389 15860 10672
rect 16012 8933 16052 10672
rect 16011 8924 16053 8933
rect 16011 8884 16012 8924
rect 16052 8884 16053 8924
rect 16011 8875 16053 8884
rect 16108 8756 16148 8765
rect 16012 8716 16108 8756
rect 15915 6236 15957 6245
rect 15915 6196 15916 6236
rect 15956 6196 15957 6236
rect 15915 6187 15957 6196
rect 15819 3380 15861 3389
rect 15819 3340 15820 3380
rect 15860 3340 15861 3380
rect 15819 3331 15861 3340
rect 15627 3128 15669 3137
rect 15627 3088 15628 3128
rect 15668 3088 15669 3128
rect 15627 3079 15669 3088
rect 15531 2708 15573 2717
rect 15531 2668 15532 2708
rect 15572 2668 15573 2708
rect 15531 2659 15573 2668
rect 14572 2071 14612 2080
rect 15340 2071 15380 2080
rect 15916 2120 15956 6187
rect 16012 2549 16052 8716
rect 16108 8707 16148 8716
rect 16204 8513 16244 10672
rect 16299 9344 16341 9353
rect 16299 9304 16300 9344
rect 16340 9304 16341 9344
rect 16299 9295 16341 9304
rect 16300 8840 16340 9295
rect 16300 8791 16340 8800
rect 16396 8513 16436 10672
rect 16491 10604 16533 10613
rect 16491 10564 16492 10604
rect 16532 10564 16533 10604
rect 16491 10555 16533 10564
rect 16492 8840 16532 10555
rect 16492 8791 16532 8800
rect 16203 8504 16245 8513
rect 16203 8464 16204 8504
rect 16244 8464 16245 8504
rect 16203 8455 16245 8464
rect 16395 8504 16437 8513
rect 16395 8464 16396 8504
rect 16436 8464 16437 8504
rect 16395 8455 16437 8464
rect 16204 7916 16244 7925
rect 16204 6581 16244 7876
rect 16396 7841 16436 7926
rect 16395 7832 16437 7841
rect 16395 7792 16396 7832
rect 16436 7792 16437 7832
rect 16395 7783 16437 7792
rect 16491 7664 16533 7673
rect 16491 7624 16492 7664
rect 16532 7624 16533 7664
rect 16491 7615 16533 7624
rect 16395 7580 16437 7589
rect 16395 7540 16396 7580
rect 16436 7540 16437 7580
rect 16395 7531 16437 7540
rect 16203 6572 16245 6581
rect 16203 6532 16204 6572
rect 16244 6532 16245 6572
rect 16203 6523 16245 6532
rect 16300 6404 16340 6413
rect 16300 6320 16340 6364
rect 16108 6280 16340 6320
rect 16011 2540 16053 2549
rect 16011 2500 16012 2540
rect 16052 2500 16053 2540
rect 16011 2491 16053 2500
rect 15916 2071 15956 2080
rect 15148 1868 15188 1877
rect 15148 197 15188 1828
rect 15724 1868 15764 1877
rect 15724 281 15764 1828
rect 15723 272 15765 281
rect 15723 232 15724 272
rect 15764 232 15765 272
rect 15723 223 15765 232
rect 15147 188 15189 197
rect 15147 148 15148 188
rect 15188 148 15189 188
rect 15147 139 15189 148
rect 15436 148 15668 188
rect 15436 80 15476 148
rect 15628 104 15668 148
rect 3531 55 3573 64
rect 3896 0 3976 80
rect 4856 0 4936 80
rect 5816 0 5896 80
rect 6776 0 6856 80
rect 7736 0 7816 80
rect 8696 0 8776 80
rect 9656 0 9736 80
rect 10616 0 10696 80
rect 11576 0 11656 80
rect 12536 0 12616 80
rect 13496 0 13576 80
rect 14456 0 14536 80
rect 15416 0 15496 80
rect 15628 64 15764 104
rect 15724 60 15764 64
rect 16108 60 16148 6280
rect 16396 2120 16436 7531
rect 16492 6656 16532 7615
rect 16588 7421 16628 10672
rect 16683 8756 16725 8765
rect 16683 8716 16684 8756
rect 16724 8716 16725 8756
rect 16683 8707 16725 8716
rect 16684 8622 16724 8707
rect 16587 7412 16629 7421
rect 16587 7372 16588 7412
rect 16628 7372 16629 7412
rect 16587 7363 16629 7372
rect 16492 6607 16532 6616
rect 16780 6329 16820 10672
rect 16972 8504 17012 10672
rect 17164 9269 17204 10672
rect 17163 9260 17205 9269
rect 17163 9220 17164 9260
rect 17204 9220 17205 9260
rect 17163 9211 17205 9220
rect 17163 8924 17205 8933
rect 17163 8884 17164 8924
rect 17204 8884 17205 8924
rect 17163 8875 17205 8884
rect 17067 8840 17109 8849
rect 17067 8800 17068 8840
rect 17108 8800 17109 8840
rect 17067 8791 17109 8800
rect 17068 8706 17108 8791
rect 16876 8464 17012 8504
rect 17067 8504 17109 8513
rect 17067 8464 17068 8504
rect 17108 8464 17109 8504
rect 16876 7589 16916 8464
rect 17067 8455 17109 8464
rect 17068 8000 17108 8455
rect 17164 8168 17204 8875
rect 17259 8756 17301 8765
rect 17259 8716 17260 8756
rect 17300 8716 17301 8756
rect 17259 8707 17301 8716
rect 17260 8622 17300 8707
rect 17164 8119 17204 8128
rect 17068 7960 17204 8000
rect 16972 7916 17012 7925
rect 16875 7580 16917 7589
rect 16875 7540 16876 7580
rect 16916 7540 16917 7580
rect 16875 7531 16917 7540
rect 16779 6320 16821 6329
rect 16972 6320 17012 7876
rect 17067 7664 17109 7673
rect 17067 7624 17068 7664
rect 17108 7624 17109 7664
rect 17067 7615 17109 7624
rect 16779 6280 16780 6320
rect 16820 6280 16821 6320
rect 16779 6271 16821 6280
rect 16876 6280 17012 6320
rect 16779 5900 16821 5909
rect 16779 5860 16780 5900
rect 16820 5860 16821 5900
rect 16779 5851 16821 5860
rect 16780 5732 16820 5851
rect 16780 5683 16820 5692
rect 16396 2071 16436 2080
rect 16204 1868 16244 1877
rect 16204 365 16244 1828
rect 16203 356 16245 365
rect 16203 316 16204 356
rect 16244 316 16245 356
rect 16203 307 16245 316
rect 16396 148 16724 188
rect 16396 80 16436 148
rect 15724 20 16148 60
rect 16376 0 16456 80
rect 16684 60 16724 148
rect 16876 60 16916 6280
rect 16972 5900 17012 5909
rect 17068 5900 17108 7615
rect 17012 5860 17108 5900
rect 16972 5851 17012 5860
rect 17164 5657 17204 7960
rect 17356 7925 17396 10672
rect 17355 7916 17397 7925
rect 17355 7876 17356 7916
rect 17396 7876 17397 7916
rect 17355 7867 17397 7876
rect 17163 5648 17205 5657
rect 17163 5608 17164 5648
rect 17204 5608 17205 5648
rect 17163 5599 17205 5608
rect 17548 3809 17588 10672
rect 17740 9269 17780 10672
rect 17739 9260 17781 9269
rect 17739 9220 17740 9260
rect 17780 9220 17781 9260
rect 17739 9211 17781 9220
rect 17932 9101 17972 10672
rect 18124 9512 18164 10672
rect 18124 9472 18260 9512
rect 18123 9260 18165 9269
rect 18123 9220 18124 9260
rect 18164 9220 18165 9260
rect 18123 9211 18165 9220
rect 17643 9092 17685 9101
rect 17643 9052 17644 9092
rect 17684 9052 17685 9092
rect 17643 9043 17685 9052
rect 17931 9092 17973 9101
rect 17931 9052 17932 9092
rect 17972 9052 17973 9092
rect 17931 9043 17973 9052
rect 17547 3800 17589 3809
rect 17547 3760 17548 3800
rect 17588 3760 17589 3800
rect 17547 3751 17589 3760
rect 17355 2540 17397 2549
rect 17355 2500 17356 2540
rect 17396 2500 17397 2540
rect 17355 2491 17397 2500
rect 17356 80 17396 2491
rect 17644 2120 17684 9043
rect 18027 8840 18069 8849
rect 17932 8800 18028 8840
rect 18068 8800 18069 8840
rect 17739 8756 17781 8765
rect 17739 8716 17740 8756
rect 17780 8716 17781 8756
rect 17739 8707 17781 8716
rect 17740 8622 17780 8707
rect 17932 8504 17972 8800
rect 18027 8791 18069 8800
rect 17932 8455 17972 8464
rect 17931 8168 17973 8177
rect 17931 8128 17932 8168
rect 17972 8128 17973 8168
rect 17931 8119 17973 8128
rect 17932 6656 17972 8119
rect 17932 6607 17972 6616
rect 17740 6413 17780 6498
rect 17739 6404 17781 6413
rect 17739 6364 17740 6404
rect 17780 6364 17781 6404
rect 17739 6355 17781 6364
rect 18124 6320 18164 9211
rect 18220 8345 18260 9472
rect 18219 8336 18261 8345
rect 18219 8296 18220 8336
rect 18260 8296 18261 8336
rect 18219 8287 18261 8296
rect 18316 7841 18356 10672
rect 18315 7832 18357 7841
rect 18315 7792 18316 7832
rect 18356 7792 18357 7832
rect 18315 7783 18357 7792
rect 18508 7589 18548 10672
rect 18700 8933 18740 10672
rect 18892 9353 18932 10672
rect 18891 9344 18933 9353
rect 18891 9304 18892 9344
rect 18932 9304 18933 9344
rect 18891 9295 18933 9304
rect 19084 9269 19124 10672
rect 19276 9689 19316 10672
rect 19467 10648 19468 10672
rect 19508 10672 19528 10688
rect 19659 10692 19892 10697
rect 19659 10688 19701 10692
rect 19508 10648 19509 10672
rect 19467 10639 19509 10648
rect 19659 10648 19660 10688
rect 19700 10648 19701 10688
rect 19659 10639 19701 10648
rect 19371 10520 19413 10529
rect 19371 10480 19372 10520
rect 19412 10480 19413 10520
rect 19371 10471 19413 10480
rect 19275 9680 19317 9689
rect 19275 9640 19276 9680
rect 19316 9640 19317 9680
rect 19275 9631 19317 9640
rect 19372 9680 19412 10471
rect 19467 10184 19509 10193
rect 19467 10144 19468 10184
rect 19508 10144 19509 10184
rect 19467 10135 19509 10144
rect 19372 9631 19412 9640
rect 19275 9512 19317 9521
rect 19275 9472 19276 9512
rect 19316 9472 19317 9512
rect 19275 9463 19317 9472
rect 19179 9428 19221 9437
rect 19179 9388 19180 9428
rect 19220 9388 19221 9428
rect 19179 9379 19221 9388
rect 19180 9294 19220 9379
rect 19083 9260 19125 9269
rect 19083 9220 19084 9260
rect 19124 9220 19125 9260
rect 19083 9211 19125 9220
rect 18808 9092 19176 9101
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 18808 9043 19176 9052
rect 18699 8924 18741 8933
rect 19276 8924 19316 9463
rect 19371 9176 19413 9185
rect 19371 9136 19372 9176
rect 19412 9136 19413 9176
rect 19371 9127 19413 9136
rect 18699 8884 18700 8924
rect 18740 8884 18741 8924
rect 18699 8875 18741 8884
rect 18988 8884 19316 8924
rect 18988 8840 19028 8884
rect 18988 8791 19028 8800
rect 19372 8840 19412 9127
rect 19372 8791 19412 8800
rect 18795 8756 18837 8765
rect 18795 8716 18796 8756
rect 18836 8716 18837 8756
rect 18795 8707 18837 8716
rect 19180 8756 19220 8765
rect 18796 8622 18836 8707
rect 19180 8093 19220 8716
rect 19372 8168 19412 8177
rect 19468 8168 19508 10135
rect 19755 9764 19797 9773
rect 19755 9724 19756 9764
rect 19796 9724 19797 9764
rect 19755 9715 19797 9724
rect 19756 8840 19796 9715
rect 19756 8791 19796 8800
rect 19564 8756 19604 8765
rect 19564 8261 19604 8716
rect 19563 8252 19605 8261
rect 19563 8212 19564 8252
rect 19604 8212 19605 8252
rect 19563 8203 19605 8212
rect 19412 8128 19508 8168
rect 19372 8119 19412 8128
rect 19179 8084 19221 8093
rect 19179 8044 19180 8084
rect 19220 8044 19221 8084
rect 19179 8035 19221 8044
rect 19179 7916 19221 7925
rect 19179 7876 19180 7916
rect 19220 7876 19221 7916
rect 19179 7867 19221 7876
rect 19180 7782 19220 7867
rect 18507 7580 18549 7589
rect 18507 7540 18508 7580
rect 18548 7540 18549 7580
rect 18507 7531 18549 7540
rect 18808 7580 19176 7589
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 18808 7531 19176 7540
rect 18699 7496 18741 7505
rect 18699 7456 18700 7496
rect 18740 7456 18741 7496
rect 18699 7447 18741 7456
rect 17644 2071 17684 2080
rect 18028 6280 18164 6320
rect 18028 2120 18068 6280
rect 18700 5900 18740 7447
rect 19371 7160 19413 7169
rect 19371 7120 19372 7160
rect 19412 7120 19413 7160
rect 19371 7111 19413 7120
rect 19563 7160 19605 7169
rect 19563 7120 19564 7160
rect 19604 7120 19605 7160
rect 19563 7111 19605 7120
rect 18987 6740 19029 6749
rect 18987 6700 18988 6740
rect 19028 6700 19029 6740
rect 18987 6691 19029 6700
rect 19179 6740 19221 6749
rect 19179 6700 19180 6740
rect 19220 6700 19221 6740
rect 19179 6691 19221 6700
rect 18988 6404 19028 6691
rect 19180 6656 19220 6691
rect 19180 6605 19220 6616
rect 18988 6355 19028 6364
rect 19372 6404 19412 7111
rect 19564 6656 19604 7111
rect 19564 6607 19604 6616
rect 19659 6488 19701 6497
rect 19659 6448 19660 6488
rect 19700 6448 19701 6488
rect 19659 6439 19701 6448
rect 19372 6355 19412 6364
rect 19660 6320 19700 6439
rect 19564 6280 19700 6320
rect 18808 6068 19176 6077
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 18808 6019 19176 6028
rect 19371 5984 19413 5993
rect 19371 5944 19372 5984
rect 19412 5944 19413 5984
rect 19371 5935 19413 5944
rect 18700 5851 18740 5860
rect 19275 5816 19317 5825
rect 19275 5776 19276 5816
rect 19316 5776 19317 5816
rect 19275 5767 19317 5776
rect 18507 5732 18549 5741
rect 18507 5692 18508 5732
rect 18548 5692 18549 5732
rect 18507 5683 18549 5692
rect 18508 5598 18548 5683
rect 18315 4808 18357 4817
rect 18315 4768 18316 4808
rect 18356 4768 18357 4808
rect 18315 4759 18357 4768
rect 18219 4472 18261 4481
rect 18219 4432 18220 4472
rect 18260 4432 18261 4472
rect 18219 4423 18261 4432
rect 18220 3893 18260 4423
rect 18316 4061 18356 4759
rect 18808 4556 19176 4565
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 18808 4507 19176 4516
rect 19276 4388 19316 5767
rect 19372 5732 19412 5935
rect 19564 5900 19604 6280
rect 19564 5851 19604 5860
rect 19372 5683 19412 5692
rect 19276 4339 19316 4348
rect 19083 4220 19125 4229
rect 19083 4180 19084 4220
rect 19124 4180 19125 4220
rect 19083 4171 19125 4180
rect 19468 4220 19508 4229
rect 19084 4086 19124 4171
rect 18315 4052 18357 4061
rect 18315 4012 18316 4052
rect 18356 4012 18357 4052
rect 18315 4003 18357 4012
rect 19468 3977 19508 4180
rect 19467 3968 19509 3977
rect 19467 3928 19468 3968
rect 19508 3928 19509 3968
rect 19467 3919 19509 3928
rect 19659 3968 19701 3977
rect 19659 3928 19660 3968
rect 19700 3928 19701 3968
rect 19659 3919 19701 3928
rect 18219 3884 18261 3893
rect 18219 3844 18220 3884
rect 18260 3844 18261 3884
rect 18219 3835 18261 3844
rect 19660 3834 19700 3919
rect 18808 3044 19176 3053
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 18808 2995 19176 3004
rect 18028 2071 18068 2080
rect 19275 2120 19317 2129
rect 19275 2080 19276 2120
rect 19316 2080 19317 2120
rect 19275 2071 19317 2080
rect 19852 2120 19892 10692
rect 20048 9848 20416 9857
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20048 9799 20416 9808
rect 19947 9680 19989 9689
rect 19947 9640 19948 9680
rect 19988 9640 19989 9680
rect 19947 9631 19989 9640
rect 19948 2129 19988 9631
rect 20048 8336 20416 8345
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20048 8287 20416 8296
rect 20048 6824 20416 6833
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20048 6775 20416 6784
rect 20048 5312 20416 5321
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20048 5263 20416 5272
rect 20048 3800 20416 3809
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20048 3751 20416 3760
rect 20139 2960 20181 2969
rect 20139 2920 20140 2960
rect 20180 2920 20181 2960
rect 20139 2911 20181 2920
rect 20140 2465 20180 2911
rect 20139 2456 20181 2465
rect 20139 2416 20140 2456
rect 20180 2416 20181 2456
rect 20139 2407 20181 2416
rect 20048 2288 20416 2297
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20048 2239 20416 2248
rect 19852 2071 19892 2080
rect 19947 2120 19989 2129
rect 19947 2080 19948 2120
rect 19988 2080 19989 2120
rect 19947 2071 19989 2080
rect 21387 2120 21429 2129
rect 21387 2080 21388 2120
rect 21428 2080 21429 2120
rect 21387 2071 21429 2080
rect 19276 1986 19316 2071
rect 17452 1868 17492 1877
rect 17452 785 17492 1828
rect 17836 1868 17876 1877
rect 17451 776 17493 785
rect 17451 736 17452 776
rect 17492 736 17493 776
rect 17451 727 17493 736
rect 16684 20 16916 60
rect 17336 0 17416 80
rect 17836 60 17876 1828
rect 19084 1868 19124 1877
rect 19467 1868 19509 1877
rect 20044 1868 20084 1877
rect 19124 1828 19412 1868
rect 19084 1819 19124 1828
rect 18808 1532 19176 1541
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 18808 1483 19176 1492
rect 19372 944 19412 1828
rect 19467 1828 19468 1868
rect 19508 1828 19509 1868
rect 19467 1819 19509 1828
rect 19948 1828 20044 1868
rect 19468 1734 19508 1819
rect 19659 1784 19701 1793
rect 19659 1744 19660 1784
rect 19700 1744 19701 1784
rect 19659 1735 19701 1744
rect 19660 1650 19700 1735
rect 19276 904 19412 944
rect 18124 148 18356 188
rect 18124 60 18164 148
rect 18316 80 18356 148
rect 19276 80 19316 904
rect 17836 20 18164 60
rect 18296 0 18376 80
rect 19256 0 19336 80
rect 19948 60 19988 1828
rect 20044 1819 20084 1828
rect 21388 1625 21428 2071
rect 21387 1616 21429 1625
rect 21387 1576 21388 1616
rect 21428 1576 21429 1616
rect 21387 1567 21429 1576
rect 20048 776 20416 785
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20048 727 20416 736
rect 20044 80 20276 104
rect 20044 64 20296 80
rect 20044 60 20084 64
rect 19948 20 20084 60
rect 20216 0 20296 64
<< via2 >>
rect 1612 9136 1652 9176
rect 1708 8464 1748 8504
rect 1612 7876 1652 7916
rect 1900 8632 1940 8672
rect 2092 8128 2132 8168
rect 1900 7876 1940 7916
rect 1900 7204 1940 7244
rect 1804 7036 1844 7076
rect 2860 10228 2900 10268
rect 2572 8632 2612 8672
rect 2572 8464 2612 8504
rect 2476 8128 2516 8168
rect 3436 10312 3476 10352
rect 3244 8464 3284 8504
rect 3148 8128 3188 8168
rect 3724 10564 3764 10604
rect 3916 9220 3956 9260
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 3532 8800 3572 8840
rect 4204 9556 4244 9596
rect 4108 8716 4148 8756
rect 4108 8128 4148 8168
rect 4396 8800 4436 8840
rect 4300 8632 4340 8672
rect 4492 8548 4532 8588
rect 5068 10144 5108 10184
rect 5356 10396 5396 10436
rect 5260 10060 5300 10100
rect 4876 9976 4916 10016
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 4972 9640 5012 9680
rect 5164 8716 5204 8756
rect 5548 10144 5588 10184
rect 5452 9136 5492 9176
rect 5836 10648 5876 10688
rect 5836 9892 5876 9932
rect 5740 8884 5780 8924
rect 5548 8716 5588 8756
rect 5644 8632 5684 8672
rect 4780 8464 4820 8504
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 4684 8212 4724 8252
rect 4588 8128 4628 8168
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 6124 8548 6164 8588
rect 6028 7456 6068 7496
rect 2572 6952 2612 6992
rect 2380 6868 2420 6908
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 1228 6448 1268 6488
rect 6316 8296 6356 8336
rect 6604 10480 6644 10520
rect 6796 10144 6836 10184
rect 6412 7372 6452 7412
rect 7084 9976 7124 10016
rect 7276 8716 7316 8756
rect 7660 9724 7700 9764
rect 7564 9472 7604 9512
rect 7468 8800 7508 8840
rect 7372 8548 7412 8588
rect 7180 8464 7220 8504
rect 7084 8212 7124 8252
rect 7852 9388 7892 9428
rect 7276 7876 7316 7916
rect 8044 9220 8084 9260
rect 8236 8716 8276 8756
rect 8428 10564 8468 10604
rect 8332 8212 8372 8252
rect 8140 8128 8180 8168
rect 8620 9304 8660 9344
rect 8524 8800 8564 8840
rect 8716 9052 8756 9092
rect 8620 7876 8660 7916
rect 6988 7288 7028 7328
rect 8908 7036 8948 7076
rect 9292 10228 9332 10268
rect 9484 8716 9524 8756
rect 9484 8380 9524 8420
rect 9100 6868 9140 6908
rect 9580 8128 9620 8168
rect 9772 9808 9812 9848
rect 9676 7876 9716 7916
rect 10060 9640 10100 9680
rect 10444 10312 10484 10352
rect 10252 9640 10292 9680
rect 10156 9556 10196 9596
rect 10156 9220 10196 9260
rect 10060 9136 10100 9176
rect 9964 9052 10004 9092
rect 9964 8212 10004 8252
rect 9868 8044 9908 8084
rect 10636 8800 10676 8840
rect 11500 10060 11540 10100
rect 11020 9640 11060 9680
rect 11212 9556 11252 9596
rect 11020 9472 11060 9512
rect 10828 8716 10868 8756
rect 11404 9724 11444 9764
rect 11788 8800 11828 8840
rect 11692 8632 11732 8672
rect 11404 8548 11444 8588
rect 11596 8548 11636 8588
rect 11788 8464 11828 8504
rect 12364 10396 12404 10436
rect 12172 9892 12212 9932
rect 11980 9724 12020 9764
rect 12076 8800 12116 8840
rect 11884 8296 11924 8336
rect 12940 9808 12980 9848
rect 13228 10144 13268 10184
rect 13132 9304 13172 9344
rect 12748 9220 12788 9260
rect 12556 8716 12596 8756
rect 13612 10480 13652 10520
rect 13516 9556 13556 9596
rect 13324 9388 13364 9428
rect 13420 8800 13460 8840
rect 13324 8128 13364 8168
rect 12076 7960 12116 8000
rect 12940 7876 12980 7916
rect 10828 7540 10868 7580
rect 10732 7204 10772 7244
rect 10540 6952 10580 6992
rect 2188 6196 2228 6236
rect 6220 6196 6260 6236
rect 1996 6112 2036 6152
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 1228 5944 1268 5984
rect 460 5776 500 5816
rect 6604 5608 6644 5648
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 2284 5104 2324 5144
rect 2476 5104 2516 5144
rect 2284 4684 2324 4724
rect 460 4180 500 4220
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 2668 4432 2708 4472
rect 5836 4348 5876 4388
rect 2476 3928 2516 3968
rect 3244 3844 3284 3884
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 2092 3256 2132 3296
rect 1900 3088 1940 3128
rect 3436 3088 3476 3128
rect 2380 2920 2420 2960
rect 2188 2416 2228 2456
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 4108 2164 4148 2204
rect 6028 2080 6068 2120
rect 9484 4852 9524 4892
rect 9772 3424 9812 3464
rect 6988 3340 7028 3380
rect 6988 2164 7028 2204
rect 9964 3424 10004 3464
rect 10060 2584 10100 2624
rect 1036 1828 1076 1868
rect 1516 400 1556 440
rect 1708 400 1748 440
rect 2092 1660 2132 1700
rect 3244 1828 3284 1868
rect 3532 1660 3572 1700
rect 2284 1408 2324 1448
rect 2476 1408 2516 1448
rect 2956 1240 2996 1280
rect 1996 904 2036 944
rect 1900 148 1940 188
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 3916 1324 3956 1364
rect 3532 64 3572 104
rect 4492 1660 4532 1700
rect 4300 1240 4340 1280
rect 4204 904 4244 944
rect 6220 1492 6260 1532
rect 5644 1324 5684 1364
rect 4876 904 4916 944
rect 4684 736 4724 776
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 8716 1828 8756 1868
rect 9772 1828 9812 1868
rect 8332 1072 8372 1112
rect 8524 1072 8564 1112
rect 4876 316 4916 356
rect 6412 316 6452 356
rect 7756 316 7796 356
rect 6796 232 6836 272
rect 5836 148 5876 188
rect 12748 7288 12788 7328
rect 12172 5440 12212 5480
rect 12364 5440 12404 5480
rect 12844 4096 12884 4136
rect 13132 4096 13172 4136
rect 12076 3760 12116 3800
rect 13900 9724 13940 9764
rect 13708 8548 13748 8588
rect 14284 8800 14324 8840
rect 15244 8800 15284 8840
rect 15052 8716 15092 8756
rect 15532 8884 15572 8924
rect 15436 8716 15476 8756
rect 15340 8632 15380 8672
rect 14092 7876 14132 7916
rect 14284 7372 14324 7412
rect 14572 6532 14612 6572
rect 14476 2668 14516 2708
rect 14764 8296 14804 8336
rect 14668 6196 14708 6236
rect 14668 2584 14708 2624
rect 10060 1660 10100 1700
rect 10636 1828 10676 1868
rect 11884 1828 11924 1868
rect 9676 1240 9716 1280
rect 10540 1240 10580 1280
rect 13516 1828 13556 1868
rect 14380 1828 14420 1868
rect 11596 1240 11636 1280
rect 13036 1240 13076 1280
rect 12556 736 12596 776
rect 15244 7456 15284 7496
rect 15340 7372 15380 7412
rect 15724 8464 15764 8504
rect 15724 4348 15764 4388
rect 16012 8884 16052 8924
rect 15916 6196 15956 6236
rect 15820 3340 15860 3380
rect 15628 3088 15668 3128
rect 15532 2668 15572 2708
rect 16300 9304 16340 9344
rect 16492 10564 16532 10604
rect 16204 8464 16244 8504
rect 16396 8464 16436 8504
rect 16396 7792 16436 7832
rect 16492 7624 16532 7664
rect 16396 7540 16436 7580
rect 16204 6532 16244 6572
rect 16012 2500 16052 2540
rect 15724 232 15764 272
rect 15148 148 15188 188
rect 16684 8716 16724 8756
rect 16588 7372 16628 7412
rect 17164 9220 17204 9260
rect 17164 8884 17204 8924
rect 17068 8800 17108 8840
rect 17068 8464 17108 8504
rect 17260 8716 17300 8756
rect 16876 7540 16916 7580
rect 17068 7624 17108 7664
rect 16780 6280 16820 6320
rect 16780 5860 16820 5900
rect 16204 316 16244 356
rect 17356 7876 17396 7916
rect 17164 5608 17204 5648
rect 17740 9220 17780 9260
rect 18124 9220 18164 9260
rect 17644 9052 17684 9092
rect 17932 9052 17972 9092
rect 17548 3760 17588 3800
rect 17356 2500 17396 2540
rect 18028 8800 18068 8840
rect 17740 8716 17780 8756
rect 17932 8128 17972 8168
rect 17740 6364 17780 6404
rect 18220 8296 18260 8336
rect 18316 7792 18356 7832
rect 18892 9304 18932 9344
rect 19468 10648 19508 10688
rect 19660 10648 19700 10688
rect 19372 10480 19412 10520
rect 19276 9640 19316 9680
rect 19468 10144 19508 10184
rect 19276 9472 19316 9512
rect 19180 9388 19220 9428
rect 19084 9220 19124 9260
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 19372 9136 19412 9176
rect 18700 8884 18740 8924
rect 18796 8716 18836 8756
rect 19756 9724 19796 9764
rect 19564 8212 19604 8252
rect 19180 8044 19220 8084
rect 19180 7876 19220 7916
rect 18508 7540 18548 7580
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 18700 7456 18740 7496
rect 19372 7120 19412 7160
rect 19564 7120 19604 7160
rect 18988 6700 19028 6740
rect 19180 6700 19220 6740
rect 19660 6448 19700 6488
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 19372 5944 19412 5984
rect 19276 5776 19316 5816
rect 18508 5692 18548 5732
rect 18316 4768 18356 4808
rect 18220 4432 18260 4472
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 19084 4180 19124 4220
rect 18316 4012 18356 4052
rect 19468 3928 19508 3968
rect 19660 3928 19700 3968
rect 18220 3844 18260 3884
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 19276 2080 19316 2120
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 19948 9640 19988 9680
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 20140 2920 20180 2960
rect 20140 2416 20180 2456
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 19948 2080 19988 2120
rect 21388 2080 21428 2120
rect 17452 736 17492 776
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 19468 1828 19508 1868
rect 19660 1744 19700 1784
rect 21388 1576 21428 1616
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
<< metal3 >>
rect 5827 10648 5836 10688
rect 5876 10648 15140 10688
rect 19459 10648 19468 10688
rect 19508 10648 19660 10688
rect 19700 10648 19709 10688
rect 15100 10604 15140 10648
rect 3715 10564 3724 10604
rect 3764 10564 8428 10604
rect 8468 10564 8477 10604
rect 15100 10564 16492 10604
rect 16532 10564 16541 10604
rect 0 10520 80 10540
rect 547 10520 605 10521
rect 21424 10520 21504 10540
rect 0 10480 556 10520
rect 596 10480 605 10520
rect 6595 10480 6604 10520
rect 6644 10480 13612 10520
rect 13652 10480 13661 10520
rect 19363 10480 19372 10520
rect 19412 10480 21504 10520
rect 0 10460 80 10480
rect 547 10479 605 10480
rect 21424 10460 21504 10480
rect 5347 10396 5356 10436
rect 5396 10396 12364 10436
rect 12404 10396 12413 10436
rect 3427 10312 3436 10352
rect 3476 10312 10444 10352
rect 10484 10312 10493 10352
rect 2851 10228 2860 10268
rect 2900 10228 9292 10268
rect 9332 10228 9341 10268
rect 0 10184 80 10204
rect 1123 10184 1181 10185
rect 21424 10184 21504 10204
rect 0 10144 1132 10184
rect 1172 10144 1181 10184
rect 5059 10144 5068 10184
rect 5108 10144 5548 10184
rect 5588 10144 5597 10184
rect 6787 10144 6796 10184
rect 6836 10144 13228 10184
rect 13268 10144 13277 10184
rect 19459 10144 19468 10184
rect 19508 10144 21504 10184
rect 0 10124 80 10144
rect 1123 10143 1181 10144
rect 21424 10124 21504 10144
rect 5251 10060 5260 10100
rect 5300 10060 11500 10100
rect 11540 10060 11549 10100
rect 4867 9976 4876 10016
rect 4916 9976 7084 10016
rect 7124 9976 7133 10016
rect 5827 9892 5836 9932
rect 5876 9892 12172 9932
rect 12212 9892 12221 9932
rect 0 9848 80 9868
rect 643 9848 701 9849
rect 21424 9848 21504 9868
rect 0 9808 652 9848
rect 692 9808 701 9848
rect 4919 9808 4928 9848
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 5296 9808 5305 9848
rect 9763 9808 9772 9848
rect 9812 9808 12940 9848
rect 12980 9808 12989 9848
rect 20039 9808 20048 9848
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20416 9808 20425 9848
rect 20524 9808 21504 9848
rect 0 9788 80 9808
rect 643 9807 701 9808
rect 20524 9764 20564 9808
rect 21424 9788 21504 9808
rect 7651 9724 7660 9764
rect 7700 9724 11404 9764
rect 11444 9724 11453 9764
rect 11971 9724 11980 9764
rect 12020 9724 13900 9764
rect 13940 9724 13949 9764
rect 19747 9724 19756 9764
rect 19796 9724 20564 9764
rect 4963 9640 4972 9680
rect 5012 9640 10060 9680
rect 10100 9640 10109 9680
rect 10243 9640 10252 9680
rect 10292 9640 11020 9680
rect 11060 9640 11069 9680
rect 19267 9640 19276 9680
rect 19316 9640 19948 9680
rect 19988 9640 19997 9680
rect 4195 9556 4204 9596
rect 4244 9556 10156 9596
rect 10196 9556 10205 9596
rect 11203 9556 11212 9596
rect 11252 9556 13516 9596
rect 13556 9556 13565 9596
rect 0 9512 80 9532
rect 5059 9512 5117 9513
rect 21424 9512 21504 9532
rect 0 9472 5068 9512
rect 5108 9472 5117 9512
rect 7555 9472 7564 9512
rect 7604 9472 11020 9512
rect 11060 9472 11069 9512
rect 19267 9472 19276 9512
rect 19316 9472 21504 9512
rect 0 9452 80 9472
rect 5059 9471 5117 9472
rect 21424 9452 21504 9472
rect 16867 9428 16925 9429
rect 7843 9388 7852 9428
rect 7892 9388 13324 9428
rect 13364 9388 13373 9428
rect 16867 9388 16876 9428
rect 16916 9388 19180 9428
rect 19220 9388 19229 9428
rect 16867 9387 16925 9388
rect 8611 9304 8620 9344
rect 8660 9304 13132 9344
rect 13172 9304 13181 9344
rect 16291 9304 16300 9344
rect 16340 9304 18892 9344
rect 18932 9304 18941 9344
rect 17635 9260 17693 9261
rect 3907 9220 3916 9260
rect 3956 9220 8044 9260
rect 8084 9220 8093 9260
rect 10147 9220 10156 9260
rect 10196 9220 12748 9260
rect 12788 9220 12797 9260
rect 15100 9220 17164 9260
rect 17204 9220 17213 9260
rect 17635 9220 17644 9260
rect 17684 9220 17740 9260
rect 17780 9220 17789 9260
rect 18115 9220 18124 9260
rect 18164 9220 19084 9260
rect 19124 9220 19133 9260
rect 0 9176 80 9196
rect 355 9176 413 9177
rect 0 9136 364 9176
rect 404 9136 413 9176
rect 1603 9136 1612 9176
rect 1652 9136 4148 9176
rect 5443 9136 5452 9176
rect 5492 9136 10060 9176
rect 10100 9136 10109 9176
rect 0 9116 80 9136
rect 355 9135 413 9136
rect 4108 9092 4148 9136
rect 15100 9092 15140 9220
rect 17635 9219 17693 9220
rect 21424 9176 21504 9196
rect 19363 9136 19372 9176
rect 19412 9136 21504 9176
rect 21424 9116 21504 9136
rect 3679 9052 3688 9092
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 4056 9052 4065 9092
rect 4108 9052 8716 9092
rect 8756 9052 8765 9092
rect 9955 9052 9964 9092
rect 10004 9052 15140 9092
rect 17635 9052 17644 9092
rect 17684 9052 17932 9092
rect 17972 9052 17981 9092
rect 18799 9052 18808 9092
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 19176 9052 19185 9092
rect 7075 9008 7133 9009
rect 172 8968 7084 9008
rect 7124 8968 7133 9008
rect 0 8840 80 8860
rect 172 8840 212 8968
rect 7075 8967 7133 8968
rect 8707 8924 8765 8925
rect 5731 8884 5740 8924
rect 5780 8884 8716 8924
rect 8756 8884 8765 8924
rect 15523 8884 15532 8924
rect 15572 8884 16012 8924
rect 16052 8884 16061 8924
rect 17155 8884 17164 8924
rect 17204 8884 18700 8924
rect 18740 8884 18749 8924
rect 8707 8883 8765 8884
rect 16291 8840 16349 8841
rect 17731 8840 17789 8841
rect 21424 8840 21504 8860
rect 0 8800 212 8840
rect 3523 8800 3532 8840
rect 3572 8800 4396 8840
rect 4436 8800 4445 8840
rect 6280 8800 7468 8840
rect 7508 8800 7517 8840
rect 8515 8800 8524 8840
rect 8564 8800 10636 8840
rect 10676 8800 10685 8840
rect 11779 8800 11788 8840
rect 11828 8800 12076 8840
rect 12116 8800 12125 8840
rect 13411 8800 13420 8840
rect 13460 8800 14284 8840
rect 14324 8800 14333 8840
rect 15235 8800 15244 8840
rect 15284 8800 15572 8840
rect 0 8780 80 8800
rect 6280 8756 6320 8800
rect 15532 8756 15572 8800
rect 16291 8800 16300 8840
rect 16340 8800 17068 8840
rect 17108 8800 17117 8840
rect 17731 8800 17740 8840
rect 17780 8800 17791 8840
rect 18019 8800 18028 8840
rect 18068 8800 21504 8840
rect 16291 8799 16349 8800
rect 17731 8799 17789 8800
rect 17740 8756 17780 8799
rect 21424 8780 21504 8800
rect 18787 8756 18845 8757
rect 4099 8716 4108 8756
rect 4148 8716 5164 8756
rect 5204 8716 5213 8756
rect 5539 8716 5548 8756
rect 5588 8716 6320 8756
rect 7267 8716 7276 8756
rect 7316 8716 7325 8756
rect 8227 8716 8236 8756
rect 8276 8716 9484 8756
rect 9524 8716 9533 8756
rect 10819 8716 10828 8756
rect 10868 8716 12556 8756
rect 12596 8716 12605 8756
rect 15043 8716 15052 8756
rect 15092 8716 15436 8756
rect 15476 8716 15485 8756
rect 15532 8716 16684 8756
rect 16724 8716 16733 8756
rect 17251 8716 17260 8756
rect 17300 8716 17309 8756
rect 17731 8716 17740 8756
rect 17780 8716 17789 8756
rect 18702 8716 18796 8756
rect 18836 8716 18845 8756
rect 7276 8672 7316 8716
rect 17260 8672 17300 8716
rect 18787 8715 18845 8716
rect 1891 8632 1900 8672
rect 1940 8632 2572 8672
rect 2612 8632 2621 8672
rect 4291 8632 4300 8672
rect 4340 8632 5644 8672
rect 5684 8632 5693 8672
rect 7276 8632 11692 8672
rect 11732 8632 11741 8672
rect 15331 8632 15340 8672
rect 15380 8632 17300 8672
rect 4483 8548 4492 8588
rect 4532 8548 6124 8588
rect 6164 8548 6173 8588
rect 7363 8548 7372 8588
rect 7412 8548 11404 8588
rect 11444 8548 11453 8588
rect 11587 8548 11596 8588
rect 11636 8548 13708 8588
rect 13748 8548 13757 8588
rect 0 8504 80 8524
rect 21424 8504 21504 8524
rect 0 8464 1652 8504
rect 1699 8464 1708 8504
rect 1748 8464 2572 8504
rect 2612 8464 2621 8504
rect 3235 8464 3244 8504
rect 3284 8464 4780 8504
rect 4820 8464 4829 8504
rect 7171 8464 7180 8504
rect 7220 8464 11788 8504
rect 11828 8464 11837 8504
rect 15715 8464 15724 8504
rect 15764 8464 16204 8504
rect 16244 8464 16253 8504
rect 16387 8464 16396 8504
rect 16436 8464 17068 8504
rect 17108 8464 17117 8504
rect 18604 8464 21504 8504
rect 0 8444 80 8464
rect 0 8168 80 8188
rect 1507 8168 1565 8169
rect 0 8128 1516 8168
rect 1556 8128 1565 8168
rect 0 8108 80 8128
rect 1507 8127 1565 8128
rect 1612 8084 1652 8464
rect 18604 8420 18644 8464
rect 21424 8444 21504 8464
rect 9475 8380 9484 8420
rect 9524 8380 18644 8420
rect 4919 8296 4928 8336
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 5296 8296 5305 8336
rect 6307 8296 6316 8336
rect 6356 8296 11884 8336
rect 11924 8296 11933 8336
rect 14755 8296 14764 8336
rect 14804 8296 18220 8336
rect 18260 8296 18269 8336
rect 20039 8296 20048 8336
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20416 8296 20425 8336
rect 12739 8252 12797 8253
rect 4675 8212 4684 8252
rect 4724 8212 7084 8252
rect 7124 8212 7133 8252
rect 8323 8212 8332 8252
rect 8372 8212 9964 8252
rect 10004 8212 10013 8252
rect 12739 8212 12748 8252
rect 12788 8212 19564 8252
rect 19604 8212 19613 8252
rect 12739 8211 12797 8212
rect 17635 8168 17693 8169
rect 21424 8168 21504 8188
rect 2083 8128 2092 8168
rect 2132 8128 2476 8168
rect 2516 8128 2525 8168
rect 3139 8128 3148 8168
rect 3188 8128 4108 8168
rect 4148 8128 4157 8168
rect 4579 8128 4588 8168
rect 4628 8128 8084 8168
rect 8131 8128 8140 8168
rect 8180 8128 9580 8168
rect 9620 8128 9629 8168
rect 13315 8128 13324 8168
rect 13364 8128 17644 8168
rect 17684 8128 17693 8168
rect 17923 8128 17932 8168
rect 17972 8128 21504 8168
rect 7651 8084 7709 8085
rect 1612 8044 7660 8084
rect 7700 8044 7709 8084
rect 8044 8084 8084 8128
rect 17635 8127 17693 8128
rect 21424 8108 21504 8128
rect 17155 8084 17213 8085
rect 8044 8044 9868 8084
rect 9908 8044 9917 8084
rect 17155 8044 17164 8084
rect 17204 8044 19180 8084
rect 19220 8044 19229 8084
rect 7651 8043 7709 8044
rect 17155 8043 17213 8044
rect 12643 8000 12701 8001
rect 7276 7960 12076 8000
rect 12116 7960 12125 8000
rect 12643 7960 12652 8000
rect 12692 7960 19220 8000
rect 7276 7916 7316 7960
rect 12643 7959 12701 7960
rect 19180 7916 19220 7960
rect 1603 7876 1612 7916
rect 1652 7876 1900 7916
rect 1940 7876 1949 7916
rect 7267 7876 7276 7916
rect 7316 7876 7325 7916
rect 8611 7876 8620 7916
rect 8660 7876 9676 7916
rect 9716 7876 9725 7916
rect 12931 7876 12940 7916
rect 12980 7876 14092 7916
rect 14132 7876 14141 7916
rect 16204 7876 17356 7916
rect 17396 7876 17405 7916
rect 19171 7876 19180 7916
rect 19220 7876 19229 7916
rect 0 7832 80 7852
rect 7555 7832 7613 7833
rect 0 7792 7564 7832
rect 7604 7792 7613 7832
rect 0 7772 80 7792
rect 7555 7791 7613 7792
rect 16204 7580 16244 7876
rect 21424 7832 21504 7852
rect 16387 7792 16396 7832
rect 16436 7792 18316 7832
rect 18356 7792 18365 7832
rect 21292 7792 21504 7832
rect 21292 7664 21332 7792
rect 21424 7772 21504 7792
rect 16483 7624 16492 7664
rect 16532 7624 17012 7664
rect 17059 7624 17068 7664
rect 17108 7624 21332 7664
rect 16972 7580 17012 7624
rect 3679 7540 3688 7580
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 4056 7540 4065 7580
rect 10819 7540 10828 7580
rect 10868 7540 16244 7580
rect 16387 7540 16396 7580
rect 16436 7540 16876 7580
rect 16916 7540 16925 7580
rect 16972 7540 18508 7580
rect 18548 7540 18557 7580
rect 18799 7540 18808 7580
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 19176 7540 19185 7580
rect 0 7496 80 7516
rect 4387 7496 4445 7497
rect 21424 7496 21504 7516
rect 0 7456 4396 7496
rect 4436 7456 4445 7496
rect 6019 7456 6028 7496
rect 6068 7456 15244 7496
rect 15284 7456 15293 7496
rect 18691 7456 18700 7496
rect 18740 7456 21504 7496
rect 0 7436 80 7456
rect 4387 7455 4445 7456
rect 21424 7436 21504 7456
rect 6403 7372 6412 7412
rect 6452 7372 14284 7412
rect 14324 7372 14333 7412
rect 15331 7372 15340 7412
rect 15380 7372 16588 7412
rect 16628 7372 16637 7412
rect 6979 7288 6988 7328
rect 7028 7288 12748 7328
rect 12788 7288 12797 7328
rect 1891 7204 1900 7244
rect 1940 7204 10732 7244
rect 10772 7204 10781 7244
rect 0 7160 80 7180
rect 21424 7160 21504 7180
rect 0 7120 19372 7160
rect 19412 7120 19421 7160
rect 19555 7120 19564 7160
rect 19604 7120 21504 7160
rect 0 7100 80 7120
rect 21424 7100 21504 7120
rect 1795 7036 1804 7076
rect 1844 7036 8908 7076
rect 8948 7036 8957 7076
rect 2563 6952 2572 6992
rect 2612 6952 10540 6992
rect 10580 6952 10589 6992
rect 2371 6868 2380 6908
rect 2420 6868 9100 6908
rect 9140 6868 9149 6908
rect 0 6824 80 6844
rect 21424 6824 21504 6844
rect 0 6784 3188 6824
rect 4919 6784 4928 6824
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 5296 6784 5305 6824
rect 20039 6784 20048 6824
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20416 6784 20425 6824
rect 20524 6784 21504 6824
rect 0 6764 80 6784
rect 3148 6740 3188 6784
rect 20524 6740 20564 6784
rect 21424 6764 21504 6784
rect 3148 6700 18988 6740
rect 19028 6700 19037 6740
rect 19171 6700 19180 6740
rect 19220 6700 20564 6740
rect 14563 6532 14572 6572
rect 14612 6532 16204 6572
rect 16244 6532 16253 6572
rect 0 6488 80 6508
rect 21424 6488 21504 6508
rect 0 6448 1228 6488
rect 1268 6448 1277 6488
rect 19651 6448 19660 6488
rect 19700 6448 21504 6488
rect 0 6428 80 6448
rect 21424 6428 21504 6448
rect 1507 6404 1565 6405
rect 1507 6364 1516 6404
rect 1556 6364 17740 6404
rect 17780 6364 17789 6404
rect 1507 6363 1565 6364
rect 16740 6280 16780 6320
rect 16820 6280 16829 6320
rect 16780 6236 16820 6280
rect 2179 6196 2188 6236
rect 2228 6196 2237 6236
rect 6211 6196 6220 6236
rect 6260 6196 14668 6236
rect 14708 6196 14717 6236
rect 15907 6196 15916 6236
rect 15956 6196 16820 6236
rect 0 6152 80 6172
rect 2188 6152 2228 6196
rect 21424 6152 21504 6172
rect 0 6112 1996 6152
rect 2036 6112 2045 6152
rect 2188 6112 21504 6152
rect 0 6092 80 6112
rect 21424 6092 21504 6112
rect 3679 6028 3688 6068
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 4056 6028 4065 6068
rect 18799 6028 18808 6068
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 19176 6028 19185 6068
rect 1219 5944 1228 5984
rect 1268 5944 19372 5984
rect 19412 5944 19421 5984
rect 7555 5900 7613 5901
rect 7555 5860 7564 5900
rect 7604 5860 16780 5900
rect 16820 5860 16829 5900
rect 7555 5859 7613 5860
rect 0 5816 80 5836
rect 4387 5816 4445 5817
rect 21424 5816 21504 5836
rect 0 5776 460 5816
rect 500 5776 509 5816
rect 4387 5776 4396 5816
rect 4436 5776 6320 5816
rect 19267 5776 19276 5816
rect 19316 5776 21504 5816
rect 0 5756 80 5776
rect 4387 5775 4445 5776
rect 6280 5732 6320 5776
rect 21424 5756 21504 5776
rect 6280 5692 18508 5732
rect 18548 5692 18557 5732
rect 6595 5608 6604 5648
rect 6644 5608 17164 5648
rect 17204 5608 17213 5648
rect 0 5480 80 5500
rect 21424 5480 21504 5500
rect 0 5440 12172 5480
rect 12212 5440 12221 5480
rect 12355 5440 12364 5480
rect 12404 5440 21504 5480
rect 0 5420 80 5440
rect 21424 5420 21504 5440
rect 4919 5272 4928 5312
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 5296 5272 5305 5312
rect 20039 5272 20048 5312
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20416 5272 20425 5312
rect 0 5144 80 5164
rect 21424 5144 21504 5164
rect 0 5104 2284 5144
rect 2324 5104 2333 5144
rect 2467 5104 2476 5144
rect 2516 5104 21504 5144
rect 0 5084 80 5104
rect 21424 5084 21504 5104
rect 7651 4892 7709 4893
rect 7651 4852 7660 4892
rect 7700 4852 9484 4892
rect 9524 4852 9533 4892
rect 7651 4851 7709 4852
rect 0 4808 80 4828
rect 21424 4808 21504 4828
rect 0 4768 2324 4808
rect 18307 4768 18316 4808
rect 18356 4768 21504 4808
rect 0 4748 80 4768
rect 2284 4724 2324 4768
rect 21424 4748 21504 4768
rect 2275 4684 2284 4724
rect 2324 4684 2333 4724
rect 3679 4516 3688 4556
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 4056 4516 4065 4556
rect 18799 4516 18808 4556
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 19176 4516 19185 4556
rect 0 4472 80 4492
rect 21424 4472 21504 4492
rect 0 4432 2668 4472
rect 2708 4432 2717 4472
rect 18211 4432 18220 4472
rect 18260 4432 21504 4472
rect 0 4412 80 4432
rect 21424 4412 21504 4432
rect 5827 4348 5836 4388
rect 5876 4348 15724 4388
rect 15764 4348 15773 4388
rect 451 4180 460 4220
rect 500 4180 19084 4220
rect 19124 4180 19133 4220
rect 0 4136 80 4156
rect 21424 4136 21504 4156
rect 0 4096 12844 4136
rect 12884 4096 12893 4136
rect 13123 4096 13132 4136
rect 13172 4096 21504 4136
rect 0 4076 80 4096
rect 21424 4076 21504 4096
rect 2476 4012 18316 4052
rect 18356 4012 18365 4052
rect 2476 3968 2516 4012
rect 2467 3928 2476 3968
rect 2516 3928 2525 3968
rect 3148 3928 19468 3968
rect 19508 3928 19517 3968
rect 19651 3928 19660 3968
rect 19700 3928 21428 3968
rect 0 3800 80 3820
rect 3148 3800 3188 3928
rect 3235 3844 3244 3884
rect 3284 3844 18220 3884
rect 18260 3844 18269 3884
rect 21388 3820 21428 3928
rect 0 3760 3188 3800
rect 4919 3760 4928 3800
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 5296 3760 5305 3800
rect 12067 3760 12076 3800
rect 12116 3760 17548 3800
rect 17588 3760 17597 3800
rect 20039 3760 20048 3800
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20416 3760 20425 3800
rect 21388 3760 21504 3820
rect 0 3740 80 3760
rect 21424 3740 21504 3760
rect 0 3464 80 3484
rect 21424 3464 21504 3484
rect 0 3424 9772 3464
rect 9812 3424 9821 3464
rect 9955 3424 9964 3464
rect 10004 3424 21504 3464
rect 0 3404 80 3424
rect 21424 3404 21504 3424
rect 6979 3340 6988 3380
rect 7028 3340 15820 3380
rect 15860 3340 15869 3380
rect 2083 3256 2092 3296
rect 2132 3256 21332 3296
rect 0 3128 80 3148
rect 21292 3128 21332 3256
rect 21424 3128 21504 3148
rect 0 3088 1900 3128
rect 1940 3088 1949 3128
rect 3427 3088 3436 3128
rect 3476 3088 15628 3128
rect 15668 3088 15677 3128
rect 21292 3088 21504 3128
rect 0 3068 80 3088
rect 21424 3068 21504 3088
rect 3679 3004 3688 3044
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 4056 3004 4065 3044
rect 18799 3004 18808 3044
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 19176 3004 19185 3044
rect 2371 2920 2380 2960
rect 2420 2920 20140 2960
rect 20180 2920 20189 2960
rect 0 2792 80 2812
rect 21424 2792 21504 2812
rect 0 2752 6320 2792
rect 0 2732 80 2752
rect 6280 2708 6320 2752
rect 19852 2752 21504 2792
rect 6280 2668 14476 2708
rect 14516 2668 14525 2708
rect 14572 2668 15532 2708
rect 15572 2668 15581 2708
rect 14572 2624 14612 2668
rect 19852 2624 19892 2752
rect 21424 2732 21504 2752
rect 10051 2584 10060 2624
rect 10100 2584 14612 2624
rect 14659 2584 14668 2624
rect 14708 2584 19892 2624
rect 16003 2500 16012 2540
rect 16052 2500 17356 2540
rect 17396 2500 17405 2540
rect 0 2456 80 2476
rect 21424 2456 21504 2476
rect 0 2416 2188 2456
rect 2228 2416 2237 2456
rect 20131 2416 20140 2456
rect 20180 2416 21504 2456
rect 0 2396 80 2416
rect 21424 2396 21504 2416
rect 4919 2248 4928 2288
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 5296 2248 5305 2288
rect 20039 2248 20048 2288
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20416 2248 20425 2288
rect 4099 2164 4108 2204
rect 4148 2164 6988 2204
rect 7028 2164 7037 2204
rect 0 2120 80 2140
rect 21424 2120 21504 2140
rect 0 2080 6028 2120
rect 6068 2080 6077 2120
rect 19267 2080 19276 2120
rect 19316 2080 19948 2120
rect 19988 2080 19997 2120
rect 21379 2080 21388 2120
rect 21428 2080 21504 2120
rect 0 2060 80 2080
rect 21424 2060 21504 2080
rect 1027 1828 1036 1868
rect 1076 1828 3244 1868
rect 3284 1828 3293 1868
rect 8707 1828 8716 1868
rect 8756 1828 9772 1868
rect 9812 1828 9821 1868
rect 10627 1828 10636 1868
rect 10676 1828 11884 1868
rect 11924 1828 11933 1868
rect 13507 1828 13516 1868
rect 13556 1828 14380 1868
rect 14420 1828 14429 1868
rect 15100 1828 19468 1868
rect 19508 1828 19517 1868
rect 0 1784 80 1804
rect 15100 1784 15140 1828
rect 21424 1784 21504 1804
rect 0 1744 15140 1784
rect 19651 1744 19660 1784
rect 19700 1744 21504 1784
rect 0 1724 80 1744
rect 21424 1724 21504 1744
rect 2083 1660 2092 1700
rect 2132 1660 3532 1700
rect 3572 1660 3581 1700
rect 4483 1660 4492 1700
rect 4532 1660 10060 1700
rect 10100 1660 10109 1700
rect 6280 1576 21388 1616
rect 21428 1576 21437 1616
rect 6280 1532 6320 1576
rect 3679 1492 3688 1532
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 4056 1492 4065 1532
rect 6211 1492 6220 1532
rect 6260 1492 6320 1532
rect 18799 1492 18808 1532
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 19176 1492 19185 1532
rect 0 1448 80 1468
rect 21424 1448 21504 1468
rect 0 1408 2284 1448
rect 2324 1408 2333 1448
rect 2467 1408 2476 1448
rect 2516 1408 21504 1448
rect 0 1388 80 1408
rect 21424 1388 21504 1408
rect 3907 1324 3916 1364
rect 3956 1324 5644 1364
rect 5684 1324 5693 1364
rect 2947 1240 2956 1280
rect 2996 1240 4300 1280
rect 4340 1240 4349 1280
rect 9667 1240 9676 1280
rect 9716 1240 10540 1280
rect 10580 1240 10589 1280
rect 11587 1240 11596 1280
rect 11636 1240 13036 1280
rect 13076 1240 13085 1280
rect 0 1112 80 1132
rect 21424 1112 21504 1132
rect 0 1072 8332 1112
rect 8372 1072 8381 1112
rect 8515 1072 8524 1112
rect 8564 1072 21504 1112
rect 0 1052 80 1072
rect 21424 1052 21504 1072
rect 1987 904 1996 944
rect 2036 904 4204 944
rect 4244 904 4253 944
rect 4867 904 4876 944
rect 4916 904 6320 944
rect 6280 860 6320 904
rect 6280 820 20564 860
rect 0 776 80 796
rect 20524 776 20564 820
rect 21424 776 21504 796
rect 0 736 4684 776
rect 4724 736 4733 776
rect 4919 736 4928 776
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 5296 736 5305 776
rect 12547 736 12556 776
rect 12596 736 17452 776
rect 17492 736 17501 776
rect 20039 736 20048 776
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20416 736 20425 776
rect 20524 736 21504 776
rect 0 716 80 736
rect 21424 716 21504 736
rect 0 440 80 460
rect 21424 440 21504 460
rect 0 400 1516 440
rect 1556 400 1565 440
rect 1699 400 1708 440
rect 1748 400 21504 440
rect 0 380 80 400
rect 21424 380 21504 400
rect 4867 316 4876 356
rect 4916 316 6412 356
rect 6452 316 6461 356
rect 7747 316 7756 356
rect 7796 316 16204 356
rect 16244 316 16253 356
rect 6787 232 6796 272
rect 6836 232 15724 272
rect 15764 232 15773 272
rect 1891 148 1900 188
rect 1940 148 1949 188
rect 5827 148 5836 188
rect 5876 148 15148 188
rect 15188 148 15197 188
rect 0 104 80 124
rect 1900 104 1940 148
rect 21424 104 21504 124
rect 0 64 1940 104
rect 3523 64 3532 104
rect 3572 64 21504 104
rect 0 44 80 64
rect 21424 44 21504 64
<< via3 >>
rect 556 10480 596 10520
rect 1132 10144 1172 10184
rect 652 9808 692 9848
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 5068 9472 5108 9512
rect 16876 9388 16916 9428
rect 17644 9220 17684 9260
rect 364 9136 404 9176
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 7084 8968 7124 9008
rect 8716 8884 8756 8924
rect 16300 8800 16340 8840
rect 17740 8800 17780 8840
rect 18796 8716 18836 8756
rect 1516 8128 1556 8168
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 12748 8212 12788 8252
rect 17644 8128 17684 8168
rect 7660 8044 7700 8084
rect 17164 8044 17204 8084
rect 12652 7960 12692 8000
rect 7564 7792 7604 7832
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 4396 7456 4436 7496
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 1516 6364 1556 6404
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 7564 5860 7604 5900
rect 4396 5776 4436 5816
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 7660 4852 7700 4892
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
<< metal4 >>
rect 556 10520 596 10529
rect 364 9176 404 9185
rect 364 7169 404 9136
rect 556 7421 596 10480
rect 1132 10184 1172 10193
rect 652 9848 692 9857
rect 555 7412 597 7421
rect 555 7372 556 7412
rect 596 7372 597 7412
rect 555 7363 597 7372
rect 652 7253 692 9808
rect 1132 7337 1172 10144
rect 4928 9848 5296 9857
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 4928 9799 5296 9808
rect 20048 9848 20416 9857
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20048 9799 20416 9808
rect 7083 9764 7125 9773
rect 7083 9724 7084 9764
rect 7124 9724 7125 9764
rect 7083 9715 7125 9724
rect 17739 9764 17781 9773
rect 17739 9724 17740 9764
rect 17780 9724 17781 9764
rect 17739 9715 17781 9724
rect 5068 9512 5108 9521
rect 3688 9092 4056 9101
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 3688 9043 4056 9052
rect 5068 8765 5108 9472
rect 7084 9008 7124 9715
rect 7084 8959 7124 8968
rect 16876 9428 16916 9437
rect 8715 8924 8757 8933
rect 8715 8884 8716 8924
rect 8756 8884 8757 8924
rect 8715 8875 8757 8884
rect 16299 8924 16341 8933
rect 16299 8884 16300 8924
rect 16340 8884 16341 8924
rect 16299 8875 16341 8884
rect 8716 8790 8756 8875
rect 16300 8840 16340 8875
rect 16300 8789 16340 8800
rect 5067 8756 5109 8765
rect 5067 8716 5068 8756
rect 5108 8716 5109 8756
rect 5067 8707 5109 8716
rect 4928 8336 5296 8345
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 4928 8287 5296 8296
rect 12748 8252 12788 8261
rect 1516 8168 1556 8177
rect 1131 7328 1173 7337
rect 1131 7288 1132 7328
rect 1172 7288 1173 7328
rect 1131 7279 1173 7288
rect 651 7244 693 7253
rect 651 7204 652 7244
rect 692 7204 693 7244
rect 651 7195 693 7204
rect 363 7160 405 7169
rect 363 7120 364 7160
rect 404 7120 405 7160
rect 363 7111 405 7120
rect 1516 6404 1556 8128
rect 7660 8084 7700 8093
rect 7564 7832 7604 7841
rect 3688 7580 4056 7589
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 3688 7531 4056 7540
rect 1516 6355 1556 6364
rect 4396 7496 4436 7505
rect 3688 6068 4056 6077
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 3688 6019 4056 6028
rect 4396 5816 4436 7456
rect 4928 6824 5296 6833
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 4928 6775 5296 6784
rect 7564 5900 7604 7792
rect 7564 5851 7604 5860
rect 4396 5767 4436 5776
rect 4928 5312 5296 5321
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 4928 5263 5296 5272
rect 7660 4892 7700 8044
rect 12652 8000 12692 8009
rect 12652 7337 12692 7960
rect 12651 7328 12693 7337
rect 12651 7288 12652 7328
rect 12692 7288 12693 7328
rect 12651 7279 12693 7288
rect 12748 7253 12788 8212
rect 16876 7421 16916 9388
rect 17644 9260 17684 9269
rect 17644 8168 17684 9220
rect 17740 8840 17780 9715
rect 18808 9092 19176 9101
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 18808 9043 19176 9052
rect 17740 8791 17780 8800
rect 18795 8756 18837 8765
rect 18795 8716 18796 8756
rect 18836 8716 18837 8756
rect 18795 8707 18837 8716
rect 18796 8622 18836 8707
rect 20048 8336 20416 8345
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20048 8287 20416 8296
rect 17644 8119 17684 8128
rect 17164 8084 17204 8093
rect 16875 7412 16917 7421
rect 16875 7372 16876 7412
rect 16916 7372 16917 7412
rect 16875 7363 16917 7372
rect 12747 7244 12789 7253
rect 12747 7204 12748 7244
rect 12788 7204 12789 7244
rect 12747 7195 12789 7204
rect 17164 7169 17204 8044
rect 18808 7580 19176 7589
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 18808 7531 19176 7540
rect 17163 7160 17205 7169
rect 17163 7120 17164 7160
rect 17204 7120 17205 7160
rect 17163 7111 17205 7120
rect 20048 6824 20416 6833
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20048 6775 20416 6784
rect 18808 6068 19176 6077
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 18808 6019 19176 6028
rect 20048 5312 20416 5321
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20048 5263 20416 5272
rect 7660 4843 7700 4852
rect 3688 4556 4056 4565
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 3688 4507 4056 4516
rect 18808 4556 19176 4565
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 18808 4507 19176 4516
rect 4928 3800 5296 3809
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 4928 3751 5296 3760
rect 20048 3800 20416 3809
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20048 3751 20416 3760
rect 3688 3044 4056 3053
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 3688 2995 4056 3004
rect 18808 3044 19176 3053
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 18808 2995 19176 3004
rect 4928 2288 5296 2297
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 4928 2239 5296 2248
rect 20048 2288 20416 2297
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20048 2239 20416 2248
rect 3688 1532 4056 1541
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 3688 1483 4056 1492
rect 18808 1532 19176 1541
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 18808 1483 19176 1492
rect 4928 776 5296 785
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 4928 727 5296 736
rect 20048 776 20416 785
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20048 727 20416 736
<< via4 >>
rect 556 7372 596 7412
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 7084 9724 7124 9764
rect 17740 9724 17780 9764
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 8716 8884 8756 8924
rect 16300 8884 16340 8924
rect 5068 8716 5108 8756
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 1132 7288 1172 7328
rect 652 7204 692 7244
rect 364 7120 404 7160
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 12652 7288 12692 7328
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 18796 8716 18836 8756
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 16876 7372 16916 7412
rect 12748 7204 12788 7244
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 17164 7120 17204 7160
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
<< metal5 >>
rect 4919 9871 5305 9890
rect 4919 9848 4985 9871
rect 5071 9848 5153 9871
rect 5239 9848 5305 9871
rect 4919 9808 4928 9848
rect 4968 9808 4985 9848
rect 5071 9808 5092 9848
rect 5132 9808 5153 9848
rect 5239 9808 5256 9848
rect 5296 9808 5305 9848
rect 4919 9785 4985 9808
rect 5071 9785 5153 9808
rect 5239 9785 5305 9808
rect 4919 9766 5305 9785
rect 20039 9871 20425 9890
rect 20039 9848 20105 9871
rect 20191 9848 20273 9871
rect 20359 9848 20425 9871
rect 20039 9808 20048 9848
rect 20088 9808 20105 9848
rect 20191 9808 20212 9848
rect 20252 9808 20273 9848
rect 20359 9808 20376 9848
rect 20416 9808 20425 9848
rect 20039 9785 20105 9808
rect 20191 9785 20273 9808
rect 20359 9785 20425 9808
rect 20039 9766 20425 9785
rect 7075 9724 7084 9764
rect 7124 9724 17740 9764
rect 17780 9724 17789 9764
rect 3679 9115 4065 9134
rect 3679 9092 3745 9115
rect 3831 9092 3913 9115
rect 3999 9092 4065 9115
rect 3679 9052 3688 9092
rect 3728 9052 3745 9092
rect 3831 9052 3852 9092
rect 3892 9052 3913 9092
rect 3999 9052 4016 9092
rect 4056 9052 4065 9092
rect 3679 9029 3745 9052
rect 3831 9029 3913 9052
rect 3999 9029 4065 9052
rect 3679 9010 4065 9029
rect 18799 9115 19185 9134
rect 18799 9092 18865 9115
rect 18951 9092 19033 9115
rect 19119 9092 19185 9115
rect 18799 9052 18808 9092
rect 18848 9052 18865 9092
rect 18951 9052 18972 9092
rect 19012 9052 19033 9092
rect 19119 9052 19136 9092
rect 19176 9052 19185 9092
rect 18799 9029 18865 9052
rect 18951 9029 19033 9052
rect 19119 9029 19185 9052
rect 18799 9010 19185 9029
rect 8707 8884 8716 8924
rect 8756 8884 16300 8924
rect 16340 8884 16349 8924
rect 5059 8716 5068 8756
rect 5108 8716 18796 8756
rect 18836 8716 18845 8756
rect 4919 8359 5305 8378
rect 4919 8336 4985 8359
rect 5071 8336 5153 8359
rect 5239 8336 5305 8359
rect 4919 8296 4928 8336
rect 4968 8296 4985 8336
rect 5071 8296 5092 8336
rect 5132 8296 5153 8336
rect 5239 8296 5256 8336
rect 5296 8296 5305 8336
rect 4919 8273 4985 8296
rect 5071 8273 5153 8296
rect 5239 8273 5305 8296
rect 4919 8254 5305 8273
rect 20039 8359 20425 8378
rect 20039 8336 20105 8359
rect 20191 8336 20273 8359
rect 20359 8336 20425 8359
rect 20039 8296 20048 8336
rect 20088 8296 20105 8336
rect 20191 8296 20212 8336
rect 20252 8296 20273 8336
rect 20359 8296 20376 8336
rect 20416 8296 20425 8336
rect 20039 8273 20105 8296
rect 20191 8273 20273 8296
rect 20359 8273 20425 8296
rect 20039 8254 20425 8273
rect 3679 7603 4065 7622
rect 3679 7580 3745 7603
rect 3831 7580 3913 7603
rect 3999 7580 4065 7603
rect 3679 7540 3688 7580
rect 3728 7540 3745 7580
rect 3831 7540 3852 7580
rect 3892 7540 3913 7580
rect 3999 7540 4016 7580
rect 4056 7540 4065 7580
rect 3679 7517 3745 7540
rect 3831 7517 3913 7540
rect 3999 7517 4065 7540
rect 3679 7498 4065 7517
rect 18799 7603 19185 7622
rect 18799 7580 18865 7603
rect 18951 7580 19033 7603
rect 19119 7580 19185 7603
rect 18799 7540 18808 7580
rect 18848 7540 18865 7580
rect 18951 7540 18972 7580
rect 19012 7540 19033 7580
rect 19119 7540 19136 7580
rect 19176 7540 19185 7580
rect 18799 7517 18865 7540
rect 18951 7517 19033 7540
rect 19119 7517 19185 7540
rect 18799 7498 19185 7517
rect 547 7372 556 7412
rect 596 7372 16876 7412
rect 16916 7372 16925 7412
rect 1123 7288 1132 7328
rect 1172 7288 12652 7328
rect 12692 7288 12701 7328
rect 643 7204 652 7244
rect 692 7204 12748 7244
rect 12788 7204 12797 7244
rect 355 7120 364 7160
rect 404 7120 17164 7160
rect 17204 7120 17213 7160
rect 4919 6847 5305 6866
rect 4919 6824 4985 6847
rect 5071 6824 5153 6847
rect 5239 6824 5305 6847
rect 4919 6784 4928 6824
rect 4968 6784 4985 6824
rect 5071 6784 5092 6824
rect 5132 6784 5153 6824
rect 5239 6784 5256 6824
rect 5296 6784 5305 6824
rect 4919 6761 4985 6784
rect 5071 6761 5153 6784
rect 5239 6761 5305 6784
rect 4919 6742 5305 6761
rect 20039 6847 20425 6866
rect 20039 6824 20105 6847
rect 20191 6824 20273 6847
rect 20359 6824 20425 6847
rect 20039 6784 20048 6824
rect 20088 6784 20105 6824
rect 20191 6784 20212 6824
rect 20252 6784 20273 6824
rect 20359 6784 20376 6824
rect 20416 6784 20425 6824
rect 20039 6761 20105 6784
rect 20191 6761 20273 6784
rect 20359 6761 20425 6784
rect 20039 6742 20425 6761
rect 3679 6091 4065 6110
rect 3679 6068 3745 6091
rect 3831 6068 3913 6091
rect 3999 6068 4065 6091
rect 3679 6028 3688 6068
rect 3728 6028 3745 6068
rect 3831 6028 3852 6068
rect 3892 6028 3913 6068
rect 3999 6028 4016 6068
rect 4056 6028 4065 6068
rect 3679 6005 3745 6028
rect 3831 6005 3913 6028
rect 3999 6005 4065 6028
rect 3679 5986 4065 6005
rect 18799 6091 19185 6110
rect 18799 6068 18865 6091
rect 18951 6068 19033 6091
rect 19119 6068 19185 6091
rect 18799 6028 18808 6068
rect 18848 6028 18865 6068
rect 18951 6028 18972 6068
rect 19012 6028 19033 6068
rect 19119 6028 19136 6068
rect 19176 6028 19185 6068
rect 18799 6005 18865 6028
rect 18951 6005 19033 6028
rect 19119 6005 19185 6028
rect 18799 5986 19185 6005
rect 4919 5335 5305 5354
rect 4919 5312 4985 5335
rect 5071 5312 5153 5335
rect 5239 5312 5305 5335
rect 4919 5272 4928 5312
rect 4968 5272 4985 5312
rect 5071 5272 5092 5312
rect 5132 5272 5153 5312
rect 5239 5272 5256 5312
rect 5296 5272 5305 5312
rect 4919 5249 4985 5272
rect 5071 5249 5153 5272
rect 5239 5249 5305 5272
rect 4919 5230 5305 5249
rect 20039 5335 20425 5354
rect 20039 5312 20105 5335
rect 20191 5312 20273 5335
rect 20359 5312 20425 5335
rect 20039 5272 20048 5312
rect 20088 5272 20105 5312
rect 20191 5272 20212 5312
rect 20252 5272 20273 5312
rect 20359 5272 20376 5312
rect 20416 5272 20425 5312
rect 20039 5249 20105 5272
rect 20191 5249 20273 5272
rect 20359 5249 20425 5272
rect 20039 5230 20425 5249
rect 3679 4579 4065 4598
rect 3679 4556 3745 4579
rect 3831 4556 3913 4579
rect 3999 4556 4065 4579
rect 3679 4516 3688 4556
rect 3728 4516 3745 4556
rect 3831 4516 3852 4556
rect 3892 4516 3913 4556
rect 3999 4516 4016 4556
rect 4056 4516 4065 4556
rect 3679 4493 3745 4516
rect 3831 4493 3913 4516
rect 3999 4493 4065 4516
rect 3679 4474 4065 4493
rect 18799 4579 19185 4598
rect 18799 4556 18865 4579
rect 18951 4556 19033 4579
rect 19119 4556 19185 4579
rect 18799 4516 18808 4556
rect 18848 4516 18865 4556
rect 18951 4516 18972 4556
rect 19012 4516 19033 4556
rect 19119 4516 19136 4556
rect 19176 4516 19185 4556
rect 18799 4493 18865 4516
rect 18951 4493 19033 4516
rect 19119 4493 19185 4516
rect 18799 4474 19185 4493
rect 4919 3823 5305 3842
rect 4919 3800 4985 3823
rect 5071 3800 5153 3823
rect 5239 3800 5305 3823
rect 4919 3760 4928 3800
rect 4968 3760 4985 3800
rect 5071 3760 5092 3800
rect 5132 3760 5153 3800
rect 5239 3760 5256 3800
rect 5296 3760 5305 3800
rect 4919 3737 4985 3760
rect 5071 3737 5153 3760
rect 5239 3737 5305 3760
rect 4919 3718 5305 3737
rect 20039 3823 20425 3842
rect 20039 3800 20105 3823
rect 20191 3800 20273 3823
rect 20359 3800 20425 3823
rect 20039 3760 20048 3800
rect 20088 3760 20105 3800
rect 20191 3760 20212 3800
rect 20252 3760 20273 3800
rect 20359 3760 20376 3800
rect 20416 3760 20425 3800
rect 20039 3737 20105 3760
rect 20191 3737 20273 3760
rect 20359 3737 20425 3760
rect 20039 3718 20425 3737
rect 3679 3067 4065 3086
rect 3679 3044 3745 3067
rect 3831 3044 3913 3067
rect 3999 3044 4065 3067
rect 3679 3004 3688 3044
rect 3728 3004 3745 3044
rect 3831 3004 3852 3044
rect 3892 3004 3913 3044
rect 3999 3004 4016 3044
rect 4056 3004 4065 3044
rect 3679 2981 3745 3004
rect 3831 2981 3913 3004
rect 3999 2981 4065 3004
rect 3679 2962 4065 2981
rect 18799 3067 19185 3086
rect 18799 3044 18865 3067
rect 18951 3044 19033 3067
rect 19119 3044 19185 3067
rect 18799 3004 18808 3044
rect 18848 3004 18865 3044
rect 18951 3004 18972 3044
rect 19012 3004 19033 3044
rect 19119 3004 19136 3044
rect 19176 3004 19185 3044
rect 18799 2981 18865 3004
rect 18951 2981 19033 3004
rect 19119 2981 19185 3004
rect 18799 2962 19185 2981
rect 4919 2311 5305 2330
rect 4919 2288 4985 2311
rect 5071 2288 5153 2311
rect 5239 2288 5305 2311
rect 4919 2248 4928 2288
rect 4968 2248 4985 2288
rect 5071 2248 5092 2288
rect 5132 2248 5153 2288
rect 5239 2248 5256 2288
rect 5296 2248 5305 2288
rect 4919 2225 4985 2248
rect 5071 2225 5153 2248
rect 5239 2225 5305 2248
rect 4919 2206 5305 2225
rect 20039 2311 20425 2330
rect 20039 2288 20105 2311
rect 20191 2288 20273 2311
rect 20359 2288 20425 2311
rect 20039 2248 20048 2288
rect 20088 2248 20105 2288
rect 20191 2248 20212 2288
rect 20252 2248 20273 2288
rect 20359 2248 20376 2288
rect 20416 2248 20425 2288
rect 20039 2225 20105 2248
rect 20191 2225 20273 2248
rect 20359 2225 20425 2248
rect 20039 2206 20425 2225
rect 3679 1555 4065 1574
rect 3679 1532 3745 1555
rect 3831 1532 3913 1555
rect 3999 1532 4065 1555
rect 3679 1492 3688 1532
rect 3728 1492 3745 1532
rect 3831 1492 3852 1532
rect 3892 1492 3913 1532
rect 3999 1492 4016 1532
rect 4056 1492 4065 1532
rect 3679 1469 3745 1492
rect 3831 1469 3913 1492
rect 3999 1469 4065 1492
rect 3679 1450 4065 1469
rect 18799 1555 19185 1574
rect 18799 1532 18865 1555
rect 18951 1532 19033 1555
rect 19119 1532 19185 1555
rect 18799 1492 18808 1532
rect 18848 1492 18865 1532
rect 18951 1492 18972 1532
rect 19012 1492 19033 1532
rect 19119 1492 19136 1532
rect 19176 1492 19185 1532
rect 18799 1469 18865 1492
rect 18951 1469 19033 1492
rect 19119 1469 19185 1492
rect 18799 1450 19185 1469
rect 4919 799 5305 818
rect 4919 776 4985 799
rect 5071 776 5153 799
rect 5239 776 5305 799
rect 4919 736 4928 776
rect 4968 736 4985 776
rect 5071 736 5092 776
rect 5132 736 5153 776
rect 5239 736 5256 776
rect 5296 736 5305 776
rect 4919 713 4985 736
rect 5071 713 5153 736
rect 5239 713 5305 736
rect 4919 694 5305 713
rect 20039 799 20425 818
rect 20039 776 20105 799
rect 20191 776 20273 799
rect 20359 776 20425 799
rect 20039 736 20048 776
rect 20088 736 20105 776
rect 20191 736 20212 776
rect 20252 736 20273 776
rect 20359 736 20376 776
rect 20416 736 20425 776
rect 20039 713 20105 736
rect 20191 713 20273 736
rect 20359 713 20425 736
rect 20039 694 20425 713
<< via5 >>
rect 4985 9848 5071 9871
rect 5153 9848 5239 9871
rect 4985 9808 5010 9848
rect 5010 9808 5050 9848
rect 5050 9808 5071 9848
rect 5153 9808 5174 9848
rect 5174 9808 5214 9848
rect 5214 9808 5239 9848
rect 4985 9785 5071 9808
rect 5153 9785 5239 9808
rect 20105 9848 20191 9871
rect 20273 9848 20359 9871
rect 20105 9808 20130 9848
rect 20130 9808 20170 9848
rect 20170 9808 20191 9848
rect 20273 9808 20294 9848
rect 20294 9808 20334 9848
rect 20334 9808 20359 9848
rect 20105 9785 20191 9808
rect 20273 9785 20359 9808
rect 3745 9092 3831 9115
rect 3913 9092 3999 9115
rect 3745 9052 3770 9092
rect 3770 9052 3810 9092
rect 3810 9052 3831 9092
rect 3913 9052 3934 9092
rect 3934 9052 3974 9092
rect 3974 9052 3999 9092
rect 3745 9029 3831 9052
rect 3913 9029 3999 9052
rect 18865 9092 18951 9115
rect 19033 9092 19119 9115
rect 18865 9052 18890 9092
rect 18890 9052 18930 9092
rect 18930 9052 18951 9092
rect 19033 9052 19054 9092
rect 19054 9052 19094 9092
rect 19094 9052 19119 9092
rect 18865 9029 18951 9052
rect 19033 9029 19119 9052
rect 4985 8336 5071 8359
rect 5153 8336 5239 8359
rect 4985 8296 5010 8336
rect 5010 8296 5050 8336
rect 5050 8296 5071 8336
rect 5153 8296 5174 8336
rect 5174 8296 5214 8336
rect 5214 8296 5239 8336
rect 4985 8273 5071 8296
rect 5153 8273 5239 8296
rect 20105 8336 20191 8359
rect 20273 8336 20359 8359
rect 20105 8296 20130 8336
rect 20130 8296 20170 8336
rect 20170 8296 20191 8336
rect 20273 8296 20294 8336
rect 20294 8296 20334 8336
rect 20334 8296 20359 8336
rect 20105 8273 20191 8296
rect 20273 8273 20359 8296
rect 3745 7580 3831 7603
rect 3913 7580 3999 7603
rect 3745 7540 3770 7580
rect 3770 7540 3810 7580
rect 3810 7540 3831 7580
rect 3913 7540 3934 7580
rect 3934 7540 3974 7580
rect 3974 7540 3999 7580
rect 3745 7517 3831 7540
rect 3913 7517 3999 7540
rect 18865 7580 18951 7603
rect 19033 7580 19119 7603
rect 18865 7540 18890 7580
rect 18890 7540 18930 7580
rect 18930 7540 18951 7580
rect 19033 7540 19054 7580
rect 19054 7540 19094 7580
rect 19094 7540 19119 7580
rect 18865 7517 18951 7540
rect 19033 7517 19119 7540
rect 4985 6824 5071 6847
rect 5153 6824 5239 6847
rect 4985 6784 5010 6824
rect 5010 6784 5050 6824
rect 5050 6784 5071 6824
rect 5153 6784 5174 6824
rect 5174 6784 5214 6824
rect 5214 6784 5239 6824
rect 4985 6761 5071 6784
rect 5153 6761 5239 6784
rect 20105 6824 20191 6847
rect 20273 6824 20359 6847
rect 20105 6784 20130 6824
rect 20130 6784 20170 6824
rect 20170 6784 20191 6824
rect 20273 6784 20294 6824
rect 20294 6784 20334 6824
rect 20334 6784 20359 6824
rect 20105 6761 20191 6784
rect 20273 6761 20359 6784
rect 3745 6068 3831 6091
rect 3913 6068 3999 6091
rect 3745 6028 3770 6068
rect 3770 6028 3810 6068
rect 3810 6028 3831 6068
rect 3913 6028 3934 6068
rect 3934 6028 3974 6068
rect 3974 6028 3999 6068
rect 3745 6005 3831 6028
rect 3913 6005 3999 6028
rect 18865 6068 18951 6091
rect 19033 6068 19119 6091
rect 18865 6028 18890 6068
rect 18890 6028 18930 6068
rect 18930 6028 18951 6068
rect 19033 6028 19054 6068
rect 19054 6028 19094 6068
rect 19094 6028 19119 6068
rect 18865 6005 18951 6028
rect 19033 6005 19119 6028
rect 4985 5312 5071 5335
rect 5153 5312 5239 5335
rect 4985 5272 5010 5312
rect 5010 5272 5050 5312
rect 5050 5272 5071 5312
rect 5153 5272 5174 5312
rect 5174 5272 5214 5312
rect 5214 5272 5239 5312
rect 4985 5249 5071 5272
rect 5153 5249 5239 5272
rect 20105 5312 20191 5335
rect 20273 5312 20359 5335
rect 20105 5272 20130 5312
rect 20130 5272 20170 5312
rect 20170 5272 20191 5312
rect 20273 5272 20294 5312
rect 20294 5272 20334 5312
rect 20334 5272 20359 5312
rect 20105 5249 20191 5272
rect 20273 5249 20359 5272
rect 3745 4556 3831 4579
rect 3913 4556 3999 4579
rect 3745 4516 3770 4556
rect 3770 4516 3810 4556
rect 3810 4516 3831 4556
rect 3913 4516 3934 4556
rect 3934 4516 3974 4556
rect 3974 4516 3999 4556
rect 3745 4493 3831 4516
rect 3913 4493 3999 4516
rect 18865 4556 18951 4579
rect 19033 4556 19119 4579
rect 18865 4516 18890 4556
rect 18890 4516 18930 4556
rect 18930 4516 18951 4556
rect 19033 4516 19054 4556
rect 19054 4516 19094 4556
rect 19094 4516 19119 4556
rect 18865 4493 18951 4516
rect 19033 4493 19119 4516
rect 4985 3800 5071 3823
rect 5153 3800 5239 3823
rect 4985 3760 5010 3800
rect 5010 3760 5050 3800
rect 5050 3760 5071 3800
rect 5153 3760 5174 3800
rect 5174 3760 5214 3800
rect 5214 3760 5239 3800
rect 4985 3737 5071 3760
rect 5153 3737 5239 3760
rect 20105 3800 20191 3823
rect 20273 3800 20359 3823
rect 20105 3760 20130 3800
rect 20130 3760 20170 3800
rect 20170 3760 20191 3800
rect 20273 3760 20294 3800
rect 20294 3760 20334 3800
rect 20334 3760 20359 3800
rect 20105 3737 20191 3760
rect 20273 3737 20359 3760
rect 3745 3044 3831 3067
rect 3913 3044 3999 3067
rect 3745 3004 3770 3044
rect 3770 3004 3810 3044
rect 3810 3004 3831 3044
rect 3913 3004 3934 3044
rect 3934 3004 3974 3044
rect 3974 3004 3999 3044
rect 3745 2981 3831 3004
rect 3913 2981 3999 3004
rect 18865 3044 18951 3067
rect 19033 3044 19119 3067
rect 18865 3004 18890 3044
rect 18890 3004 18930 3044
rect 18930 3004 18951 3044
rect 19033 3004 19054 3044
rect 19054 3004 19094 3044
rect 19094 3004 19119 3044
rect 18865 2981 18951 3004
rect 19033 2981 19119 3004
rect 4985 2288 5071 2311
rect 5153 2288 5239 2311
rect 4985 2248 5010 2288
rect 5010 2248 5050 2288
rect 5050 2248 5071 2288
rect 5153 2248 5174 2288
rect 5174 2248 5214 2288
rect 5214 2248 5239 2288
rect 4985 2225 5071 2248
rect 5153 2225 5239 2248
rect 20105 2288 20191 2311
rect 20273 2288 20359 2311
rect 20105 2248 20130 2288
rect 20130 2248 20170 2288
rect 20170 2248 20191 2288
rect 20273 2248 20294 2288
rect 20294 2248 20334 2288
rect 20334 2248 20359 2288
rect 20105 2225 20191 2248
rect 20273 2225 20359 2248
rect 3745 1532 3831 1555
rect 3913 1532 3999 1555
rect 3745 1492 3770 1532
rect 3770 1492 3810 1532
rect 3810 1492 3831 1532
rect 3913 1492 3934 1532
rect 3934 1492 3974 1532
rect 3974 1492 3999 1532
rect 3745 1469 3831 1492
rect 3913 1469 3999 1492
rect 18865 1532 18951 1555
rect 19033 1532 19119 1555
rect 18865 1492 18890 1532
rect 18890 1492 18930 1532
rect 18930 1492 18951 1532
rect 19033 1492 19054 1532
rect 19054 1492 19094 1532
rect 19094 1492 19119 1532
rect 18865 1469 18951 1492
rect 19033 1469 19119 1492
rect 4985 776 5071 799
rect 5153 776 5239 799
rect 4985 736 5010 776
rect 5010 736 5050 776
rect 5050 736 5071 776
rect 5153 736 5174 776
rect 5174 736 5214 776
rect 5214 736 5239 776
rect 4985 713 5071 736
rect 5153 713 5239 736
rect 20105 776 20191 799
rect 20273 776 20359 799
rect 20105 736 20130 776
rect 20130 736 20170 776
rect 20170 736 20191 776
rect 20273 736 20294 776
rect 20294 736 20334 776
rect 20334 736 20359 776
rect 20105 713 20191 736
rect 20273 713 20359 736
<< metal6 >>
rect 3652 9115 4092 10752
rect 3652 9029 3745 9115
rect 3831 9029 3913 9115
rect 3999 9029 4092 9115
rect 3652 7603 4092 9029
rect 3652 7517 3745 7603
rect 3831 7517 3913 7603
rect 3999 7517 4092 7603
rect 3652 6091 4092 7517
rect 3652 6005 3745 6091
rect 3831 6005 3913 6091
rect 3999 6005 4092 6091
rect 3652 4579 4092 6005
rect 3652 4493 3745 4579
rect 3831 4493 3913 4579
rect 3999 4493 4092 4579
rect 3652 3067 4092 4493
rect 3652 2981 3745 3067
rect 3831 2981 3913 3067
rect 3999 2981 4092 3067
rect 3652 1555 4092 2981
rect 3652 1469 3745 1555
rect 3831 1469 3913 1555
rect 3999 1469 4092 1555
rect 3652 0 4092 1469
rect 4892 9871 5332 10752
rect 4892 9785 4985 9871
rect 5071 9785 5153 9871
rect 5239 9785 5332 9871
rect 4892 8359 5332 9785
rect 4892 8273 4985 8359
rect 5071 8273 5153 8359
rect 5239 8273 5332 8359
rect 4892 6847 5332 8273
rect 4892 6761 4985 6847
rect 5071 6761 5153 6847
rect 5239 6761 5332 6847
rect 4892 5335 5332 6761
rect 4892 5249 4985 5335
rect 5071 5249 5153 5335
rect 5239 5249 5332 5335
rect 4892 3823 5332 5249
rect 4892 3737 4985 3823
rect 5071 3737 5153 3823
rect 5239 3737 5332 3823
rect 4892 2311 5332 3737
rect 4892 2225 4985 2311
rect 5071 2225 5153 2311
rect 5239 2225 5332 2311
rect 4892 799 5332 2225
rect 4892 713 4985 799
rect 5071 713 5153 799
rect 5239 713 5332 799
rect 4892 0 5332 713
rect 18772 9115 19212 10752
rect 18772 9029 18865 9115
rect 18951 9029 19033 9115
rect 19119 9029 19212 9115
rect 18772 7603 19212 9029
rect 18772 7517 18865 7603
rect 18951 7517 19033 7603
rect 19119 7517 19212 7603
rect 18772 6091 19212 7517
rect 18772 6005 18865 6091
rect 18951 6005 19033 6091
rect 19119 6005 19212 6091
rect 18772 4579 19212 6005
rect 18772 4493 18865 4579
rect 18951 4493 19033 4579
rect 19119 4493 19212 4579
rect 18772 3067 19212 4493
rect 18772 2981 18865 3067
rect 18951 2981 19033 3067
rect 19119 2981 19212 3067
rect 18772 1555 19212 2981
rect 18772 1469 18865 1555
rect 18951 1469 19033 1555
rect 19119 1469 19212 1555
rect 18772 0 19212 1469
rect 20012 9871 20452 10752
rect 20012 9785 20105 9871
rect 20191 9785 20273 9871
rect 20359 9785 20452 9871
rect 20012 8359 20452 9785
rect 20012 8273 20105 8359
rect 20191 8273 20273 8359
rect 20359 8273 20452 8359
rect 20012 6847 20452 8273
rect 20012 6761 20105 6847
rect 20191 6761 20273 6847
rect 20359 6761 20452 6847
rect 20012 5335 20452 6761
rect 20012 5249 20105 5335
rect 20191 5249 20273 5335
rect 20359 5249 20452 5335
rect 20012 3823 20452 5249
rect 20012 3737 20105 3823
rect 20191 3737 20273 3823
rect 20359 3737 20452 3823
rect 20012 2311 20452 3737
rect 20012 2225 20105 2311
rect 20191 2225 20273 2311
rect 20359 2225 20452 2311
rect 20012 799 20452 2225
rect 20012 713 20105 799
rect 20191 713 20273 799
rect 20359 713 20452 799
rect 20012 0 20452 713
use sg13g2_buf_1  _00_
timestamp 1676381911
transform 1 0 1824 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _01_
timestamp 1676381911
transform 1 0 1440 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _02_
timestamp 1676381911
transform 1 0 4608 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _03_
timestamp 1676381911
transform 1 0 8256 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _04_
timestamp 1676381911
transform 1 0 2208 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _05_
timestamp 1676381911
transform 1 0 19392 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _06_
timestamp 1676381911
transform 1 0 5952 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _07_
timestamp 1676381911
transform 1 0 2112 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _08_
timestamp 1676381911
transform 1 0 14400 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _09_
timestamp 1676381911
transform 1 0 1824 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _10_
timestamp 1676381911
transform 1 0 9696 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _11_
timestamp 1676381911
transform 1 0 19392 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _12_
timestamp 1676381911
transform 1 0 12864 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _13_
timestamp 1676381911
transform 1 0 2592 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _14_
timestamp 1676381911
transform 1 0 2208 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _15_
timestamp 1676381911
transform 1 0 2208 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _16_
timestamp 1676381911
transform 1 0 12096 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _17_
timestamp 1676381911
transform 1 0 19008 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _18_
timestamp 1676381911
transform 1 0 1920 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _19_
timestamp 1676381911
transform 1 0 19296 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _20_
timestamp 1676381911
transform 1 0 18912 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _21_
timestamp 1676381911
transform 1 0 19296 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _22_
timestamp 1676381911
transform 1 0 18432 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _23_
timestamp 1676381911
transform 1 0 16704 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _24_
timestamp 1676381911
transform 1 0 17664 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _25_
timestamp 1676381911
transform 1 0 9408 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _26_
timestamp 1676381911
transform 1 0 17664 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _27_
timestamp 1676381911
transform 1 0 19104 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _28_
timestamp 1676381911
transform 1 0 18720 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _29_
timestamp 1676381911
transform 1 0 19488 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _30_
timestamp 1676381911
transform 1 0 19104 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _31_
timestamp 1676381911
transform 1 0 19104 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _32_
timestamp 1676381911
transform 1 0 3840 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _33_
timestamp 1676381911
transform 1 0 4224 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _34_
timestamp 1676381911
transform 1 0 5568 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _35_
timestamp 1676381911
transform 1 0 6336 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _36_
timestamp 1676381911
transform 1 0 15072 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _37_
timestamp 1676381911
transform 1 0 15648 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _38_
timestamp 1676381911
transform 1 0 16128 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _39_
timestamp 1676381911
transform 1 0 9696 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _40_
timestamp 1676381911
transform 1 0 10464 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _41_
timestamp 1676381911
transform 1 0 11808 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _42_
timestamp 1676381911
transform 1 0 12960 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _43_
timestamp 1676381911
transform 1 0 17376 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _44_
timestamp 1676381911
transform 1 0 14304 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _45_
timestamp 1676381911
transform 1 0 16128 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _46_
timestamp 1676381911
transform 1 0 16224 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _47_
timestamp 1676381911
transform 1 0 16896 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _48_
timestamp 1676381911
transform 1 0 16032 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _49_
timestamp 1676381911
transform 1 0 17760 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _50_
timestamp 1676381911
transform 1 0 19008 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _51_
timestamp 1676381911
transform -1 0 20160 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _52_
timestamp 1676381911
transform -1 0 2880 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _53_
timestamp 1676381911
transform -1 0 2496 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _54_
timestamp 1676381911
transform 1 0 1728 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _55_
timestamp 1676381911
transform 1 0 1824 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _56_
timestamp 1676381911
transform 1 0 1824 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _57_
timestamp 1676381911
transform 1 0 2496 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _58_
timestamp 1676381911
transform -1 0 3648 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _59_
timestamp 1676381911
transform -1 0 4416 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _60_
timestamp 1676381911
transform -1 0 5088 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _61_
timestamp 1676381911
transform -1 0 4704 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _62_
timestamp 1676381911
transform -1 0 8736 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _63_
timestamp 1676381911
transform -1 0 8352 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _64_
timestamp 1676381911
transform -1 0 5472 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _65_
timestamp 1676381911
transform -1 0 5952 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _66_
timestamp 1676381911
transform -1 0 6432 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _67_
timestamp 1676381911
transform -1 0 7392 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _68_
timestamp 1676381911
transform -1 0 7392 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _69_
timestamp 1676381911
transform -1 0 7776 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _70_
timestamp 1676381911
transform -1 0 11712 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _71_
timestamp 1676381911
transform -1 0 10368 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _72_
timestamp 1676381911
transform -1 0 17376 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _73_
timestamp 1676381911
transform -1 0 16800 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _74_
timestamp 1676381911
transform -1 0 15552 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _75_
timestamp 1676381911
transform -1 0 14976 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _76_
timestamp 1676381911
transform -1 0 14592 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _77_
timestamp 1676381911
transform -1 0 14016 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _78_
timestamp 1676381911
transform -1 0 13536 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _79_
timestamp 1676381911
transform -1 0 13056 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _80_
timestamp 1676381911
transform -1 0 12096 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _81_
timestamp 1676381911
transform -1 0 11712 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _82_
timestamp 1676381911
transform -1 0 11328 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _83_
timestamp 1676381911
transform -1 0 7968 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _84_
timestamp 1676381911
transform -1 0 8352 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _85_
timestamp 1676381911
transform -1 0 9888 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _86_
timestamp 1676381911
transform -1 0 10272 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _87_
timestamp 1676381911
transform -1 0 10944 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _88_
timestamp 1676381911
transform 1 0 3168 0 -1 2268
box -48 -56 432 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1679581782
transform 1 0 1152 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1679581782
transform 1 0 1824 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1679581782
transform 1 0 2496 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_21
timestamp 1679581782
transform 1 0 3168 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_28
timestamp 1679581782
transform 1 0 3840 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_35
timestamp 1679581782
transform 1 0 4512 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_42
timestamp 1679581782
transform 1 0 5184 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_49
timestamp 1679581782
transform 1 0 5856 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_56
timestamp 1679581782
transform 1 0 6528 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_63
timestamp 1679581782
transform 1 0 7200 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_70
timestamp 1679581782
transform 1 0 7872 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_77
timestamp 1679581782
transform 1 0 8544 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_84
timestamp 1679581782
transform 1 0 9216 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_91
timestamp 1679581782
transform 1 0 9888 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_98
timestamp 1679581782
transform 1 0 10560 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_105
timestamp 1679581782
transform 1 0 11232 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_112
timestamp 1679581782
transform 1 0 11904 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_119
timestamp 1679581782
transform 1 0 12576 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_126
timestamp 1679581782
transform 1 0 13248 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_133
timestamp 1679581782
transform 1 0 13920 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_140
timestamp 1679581782
transform 1 0 14592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_147
timestamp 1679581782
transform 1 0 15264 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_154
timestamp 1679581782
transform 1 0 15936 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_161
timestamp 1679581782
transform 1 0 16608 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_168
timestamp 1679581782
transform 1 0 17280 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_175
timestamp 1679581782
transform 1 0 17952 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_182
timestamp 1679581782
transform 1 0 18624 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_189
timestamp 1679581782
transform 1 0 19296 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_196
timestamp 1679577901
transform 1 0 19968 0 1 756
box -48 -56 432 834
use sg13g2_fill_2  FILLER_1_0
timestamp 1677580104
transform 1 0 1152 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_2
timestamp 1677579658
transform 1 0 1344 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_1_15
timestamp 1679577901
transform 1 0 2592 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_1_19
timestamp 1677580104
transform 1 0 2976 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_1_25
timestamp 1677580104
transform 1 0 3552 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_27
timestamp 1677579658
transform 1 0 3744 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_1_40
timestamp 1679577901
transform 1 0 4992 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_1_44
timestamp 1677580104
transform 1 0 5376 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_58
timestamp 1679581782
transform 1 0 6720 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_65
timestamp 1679581782
transform 1 0 7392 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_72
timestamp 1677580104
transform 1 0 8064 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_78
timestamp 1679581782
transform 1 0 8640 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_85
timestamp 1679577901
transform 1 0 9312 0 -1 2268
box -48 -56 432 834
use sg13g2_decap_4  FILLER_1_93
timestamp 1679577901
transform 1 0 10080 0 -1 2268
box -48 -56 432 834
use sg13g2_decap_8  FILLER_1_101
timestamp 1679581782
transform 1 0 10848 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_108
timestamp 1677580104
transform 1 0 11520 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_110
timestamp 1677579658
transform 1 0 11712 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_115
timestamp 1679581782
transform 1 0 12192 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_1_122
timestamp 1677579658
transform 1 0 12864 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_127
timestamp 1679581782
transform 1 0 13344 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_134
timestamp 1677580104
transform 1 0 14016 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_136
timestamp 1677579658
transform 1 0 14208 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_1_141
timestamp 1679577901
transform 1 0 14688 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_1_149
timestamp 1677580104
transform 1 0 15456 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_155
timestamp 1677579658
transform 1 0 16032 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_160
timestamp 1679581782
transform 1 0 16512 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_167
timestamp 1677580104
transform 1 0 17184 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_177
timestamp 1679581782
transform 1 0 18144 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_184
timestamp 1677580104
transform 1 0 18816 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_1_198
timestamp 1677580104
transform 1 0 20160 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_0
timestamp 1679581782
transform 1 0 1152 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_7
timestamp 1679581782
transform 1 0 1824 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_14
timestamp 1679581782
transform 1 0 2496 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_21
timestamp 1679581782
transform 1 0 3168 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_28
timestamp 1679581782
transform 1 0 3840 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_35
timestamp 1679581782
transform 1 0 4512 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_42
timestamp 1679581782
transform 1 0 5184 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_49
timestamp 1679581782
transform 1 0 5856 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_56
timestamp 1679581782
transform 1 0 6528 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_63
timestamp 1679581782
transform 1 0 7200 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_70
timestamp 1679581782
transform 1 0 7872 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_77
timestamp 1679581782
transform 1 0 8544 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_84
timestamp 1679581782
transform 1 0 9216 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_91
timestamp 1679581782
transform 1 0 9888 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_98
timestamp 1679581782
transform 1 0 10560 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_105
timestamp 1679581782
transform 1 0 11232 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_112
timestamp 1679581782
transform 1 0 11904 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_119
timestamp 1679581782
transform 1 0 12576 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_126
timestamp 1679581782
transform 1 0 13248 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_133
timestamp 1679577901
transform 1 0 13920 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_137
timestamp 1677579658
transform 1 0 14304 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_142
timestamp 1679581782
transform 1 0 14784 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_149
timestamp 1679581782
transform 1 0 15456 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_156
timestamp 1679581782
transform 1 0 16128 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_163
timestamp 1679581782
transform 1 0 16800 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_170
timestamp 1679581782
transform 1 0 17472 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_177
timestamp 1679581782
transform 1 0 18144 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_184
timestamp 1679581782
transform 1 0 18816 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_191
timestamp 1679581782
transform 1 0 19488 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_198
timestamp 1677580104
transform 1 0 20160 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_0
timestamp 1679581782
transform 1 0 1152 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_7
timestamp 1677580104
transform 1 0 1824 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_9
timestamp 1677579658
transform 1 0 2016 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_14
timestamp 1679581782
transform 1 0 2496 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_21
timestamp 1679581782
transform 1 0 3168 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_28
timestamp 1679581782
transform 1 0 3840 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_35
timestamp 1679581782
transform 1 0 4512 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_42
timestamp 1679581782
transform 1 0 5184 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_49
timestamp 1679581782
transform 1 0 5856 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_56
timestamp 1679581782
transform 1 0 6528 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_63
timestamp 1679581782
transform 1 0 7200 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_70
timestamp 1679581782
transform 1 0 7872 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_77
timestamp 1679581782
transform 1 0 8544 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_84
timestamp 1679581782
transform 1 0 9216 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_91
timestamp 1679581782
transform 1 0 9888 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_98
timestamp 1679581782
transform 1 0 10560 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_105
timestamp 1679581782
transform 1 0 11232 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_112
timestamp 1679581782
transform 1 0 11904 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_119
timestamp 1679581782
transform 1 0 12576 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_126
timestamp 1679581782
transform 1 0 13248 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_133
timestamp 1679581782
transform 1 0 13920 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_140
timestamp 1679581782
transform 1 0 14592 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_147
timestamp 1679581782
transform 1 0 15264 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_154
timestamp 1679581782
transform 1 0 15936 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_161
timestamp 1679581782
transform 1 0 16608 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_168
timestamp 1679581782
transform 1 0 17280 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_175
timestamp 1679581782
transform 1 0 17952 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_182
timestamp 1679581782
transform 1 0 18624 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_189
timestamp 1679581782
transform 1 0 19296 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_196
timestamp 1679577901
transform 1 0 19968 0 -1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_4_0
timestamp 1679581782
transform 1 0 1152 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_19
timestamp 1679581782
transform 1 0 2976 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_26
timestamp 1679581782
transform 1 0 3648 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_33
timestamp 1679581782
transform 1 0 4320 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_40
timestamp 1679581782
transform 1 0 4992 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_47
timestamp 1679581782
transform 1 0 5664 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_54
timestamp 1679581782
transform 1 0 6336 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_61
timestamp 1679581782
transform 1 0 7008 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_68
timestamp 1679581782
transform 1 0 7680 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_75
timestamp 1679581782
transform 1 0 8352 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_82
timestamp 1679581782
transform 1 0 9024 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_93
timestamp 1679581782
transform 1 0 10080 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_100
timestamp 1679581782
transform 1 0 10752 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_107
timestamp 1679581782
transform 1 0 11424 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_114
timestamp 1679581782
transform 1 0 12096 0 1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_121
timestamp 1677579658
transform 1 0 12768 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_126
timestamp 1679581782
transform 1 0 13248 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_133
timestamp 1679581782
transform 1 0 13920 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_140
timestamp 1679581782
transform 1 0 14592 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_147
timestamp 1679581782
transform 1 0 15264 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_154
timestamp 1679581782
transform 1 0 15936 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_161
timestamp 1679581782
transform 1 0 16608 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_168
timestamp 1679581782
transform 1 0 17280 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_175
timestamp 1679581782
transform 1 0 17952 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_182
timestamp 1679577901
transform 1 0 18624 0 1 3780
box -48 -56 432 834
use sg13g2_decap_4  FILLER_4_194
timestamp 1679577901
transform 1 0 19776 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_198
timestamp 1677580104
transform 1 0 20160 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_0
timestamp 1679581782
transform 1 0 1152 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_7
timestamp 1679577901
transform 1 0 1824 0 -1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_5_15
timestamp 1679581782
transform 1 0 2592 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_22
timestamp 1679581782
transform 1 0 3264 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_29
timestamp 1679581782
transform 1 0 3936 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_36
timestamp 1679581782
transform 1 0 4608 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_43
timestamp 1679581782
transform 1 0 5280 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_50
timestamp 1679581782
transform 1 0 5952 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_57
timestamp 1679581782
transform 1 0 6624 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_64
timestamp 1679581782
transform 1 0 7296 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_71
timestamp 1679581782
transform 1 0 7968 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_78
timestamp 1679581782
transform 1 0 8640 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_85
timestamp 1677579658
transform 1 0 9312 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_90
timestamp 1679581782
transform 1 0 9792 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_97
timestamp 1679581782
transform 1 0 10464 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_104
timestamp 1679581782
transform 1 0 11136 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_111
timestamp 1679581782
transform 1 0 11808 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_118
timestamp 1679581782
transform 1 0 12480 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_125
timestamp 1679581782
transform 1 0 13152 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_132
timestamp 1679581782
transform 1 0 13824 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_139
timestamp 1679581782
transform 1 0 14496 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_146
timestamp 1679581782
transform 1 0 15168 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_153
timestamp 1679581782
transform 1 0 15840 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_160
timestamp 1679581782
transform 1 0 16512 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_167
timestamp 1679581782
transform 1 0 17184 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_174
timestamp 1679581782
transform 1 0 17856 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_181
timestamp 1679581782
transform 1 0 18528 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_188
timestamp 1679581782
transform 1 0 19200 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_195
timestamp 1679577901
transform 1 0 19872 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_199
timestamp 1677579658
transform 1 0 20256 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_0
timestamp 1679581782
transform 1 0 1152 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_7
timestamp 1679581782
transform 1 0 1824 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_14
timestamp 1679581782
transform 1 0 2496 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_21
timestamp 1679581782
transform 1 0 3168 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_28
timestamp 1679581782
transform 1 0 3840 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_35
timestamp 1679581782
transform 1 0 4512 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_42
timestamp 1679581782
transform 1 0 5184 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_49
timestamp 1679581782
transform 1 0 5856 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_56
timestamp 1679581782
transform 1 0 6528 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_63
timestamp 1679581782
transform 1 0 7200 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_70
timestamp 1679581782
transform 1 0 7872 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_77
timestamp 1679581782
transform 1 0 8544 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_84
timestamp 1679581782
transform 1 0 9216 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_91
timestamp 1679581782
transform 1 0 9888 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_98
timestamp 1679581782
transform 1 0 10560 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_105
timestamp 1679581782
transform 1 0 11232 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_112
timestamp 1677580104
transform 1 0 11904 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_118
timestamp 1679581782
transform 1 0 12480 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_125
timestamp 1679581782
transform 1 0 13152 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_132
timestamp 1679581782
transform 1 0 13824 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_139
timestamp 1679581782
transform 1 0 14496 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_146
timestamp 1679581782
transform 1 0 15168 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_153
timestamp 1679581782
transform 1 0 15840 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_160
timestamp 1677580104
transform 1 0 16512 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_166
timestamp 1679581782
transform 1 0 17088 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_173
timestamp 1679581782
transform 1 0 17760 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_184
timestamp 1679577901
transform 1 0 18816 0 1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_188
timestamp 1677579658
transform 1 0 19200 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_193
timestamp 1679581782
transform 1 0 19680 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_0
timestamp 1679581782
transform 1 0 1152 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_7
timestamp 1677579658
transform 1 0 1824 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_12
timestamp 1679581782
transform 1 0 2304 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_19
timestamp 1679581782
transform 1 0 2976 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_26
timestamp 1679581782
transform 1 0 3648 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_33
timestamp 1679581782
transform 1 0 4320 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_40
timestamp 1679581782
transform 1 0 4992 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_47
timestamp 1679581782
transform 1 0 5664 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_54
timestamp 1679581782
transform 1 0 6336 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_61
timestamp 1679581782
transform 1 0 7008 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_68
timestamp 1679581782
transform 1 0 7680 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_75
timestamp 1679581782
transform 1 0 8352 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_82
timestamp 1679581782
transform 1 0 9024 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_89
timestamp 1679581782
transform 1 0 9696 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_96
timestamp 1679581782
transform 1 0 10368 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_103
timestamp 1679581782
transform 1 0 11040 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_110
timestamp 1679581782
transform 1 0 11712 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_117
timestamp 1679581782
transform 1 0 12384 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_124
timestamp 1679581782
transform 1 0 13056 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_131
timestamp 1679581782
transform 1 0 13728 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_138
timestamp 1679581782
transform 1 0 14400 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_145
timestamp 1679581782
transform 1 0 15072 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_152
timestamp 1679577901
transform 1 0 15744 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_156
timestamp 1677579658
transform 1 0 16128 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_161
timestamp 1679581782
transform 1 0 16608 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_168
timestamp 1679577901
transform 1 0 17280 0 -1 6804
box -48 -56 432 834
use sg13g2_decap_8  FILLER_7_176
timestamp 1679581782
transform 1 0 18048 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_183
timestamp 1677580104
transform 1 0 18720 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_193
timestamp 1679581782
transform 1 0 19680 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_0
timestamp 1679581782
transform 1 0 1152 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_11
timestamp 1679581782
transform 1 0 2208 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_18
timestamp 1679581782
transform 1 0 2880 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_25
timestamp 1679581782
transform 1 0 3552 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_32
timestamp 1679581782
transform 1 0 4224 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_39
timestamp 1679581782
transform 1 0 4896 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_46
timestamp 1679581782
transform 1 0 5568 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_53
timestamp 1679581782
transform 1 0 6240 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_60
timestamp 1679581782
transform 1 0 6912 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_67
timestamp 1679581782
transform 1 0 7584 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_74
timestamp 1679581782
transform 1 0 8256 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_81
timestamp 1679581782
transform 1 0 8928 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_88
timestamp 1679581782
transform 1 0 9600 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_95
timestamp 1679581782
transform 1 0 10272 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_102
timestamp 1679581782
transform 1 0 10944 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_109
timestamp 1679581782
transform 1 0 11616 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_116
timestamp 1679581782
transform 1 0 12288 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_123
timestamp 1679581782
transform 1 0 12960 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_130
timestamp 1679581782
transform 1 0 13632 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_137
timestamp 1679581782
transform 1 0 14304 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_144
timestamp 1679581782
transform 1 0 14976 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_151
timestamp 1679581782
transform 1 0 15648 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_158
timestamp 1679581782
transform 1 0 16320 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_165
timestamp 1679581782
transform 1 0 16992 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_172
timestamp 1679581782
transform 1 0 17664 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_179
timestamp 1679581782
transform 1 0 18336 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_186
timestamp 1679581782
transform 1 0 19008 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_193
timestamp 1679581782
transform 1 0 19680 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_0
timestamp 1679581782
transform 1 0 1152 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_11
timestamp 1677580104
transform 1 0 2208 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_13
timestamp 1677579658
transform 1 0 2400 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_18
timestamp 1679577901
transform 1 0 2880 0 -1 8316
box -48 -56 432 834
use sg13g2_decap_4  FILLER_9_26
timestamp 1679577901
transform 1 0 3648 0 -1 8316
box -48 -56 432 834
use sg13g2_decap_8  FILLER_9_34
timestamp 1679581782
transform 1 0 4416 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_41
timestamp 1679581782
transform 1 0 5088 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_48
timestamp 1679581782
transform 1 0 5760 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_55
timestamp 1679577901
transform 1 0 6432 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_59
timestamp 1677580104
transform 1 0 6816 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_65
timestamp 1677580104
transform 1 0 7392 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_79
timestamp 1679581782
transform 1 0 8736 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_86
timestamp 1677579658
transform 1 0 9408 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_95
timestamp 1679581782
transform 1 0 10272 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_102
timestamp 1679577901
transform 1 0 10944 0 -1 8316
box -48 -56 432 834
use sg13g2_decap_8  FILLER_9_110
timestamp 1679581782
transform 1 0 11712 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_117
timestamp 1677580104
transform 1 0 12384 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_119
timestamp 1677579658
transform 1 0 12576 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_124
timestamp 1677579658
transform 1 0 13056 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_129
timestamp 1677579658
transform 1 0 13536 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_134
timestamp 1679581782
transform 1 0 14016 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_141
timestamp 1679581782
transform 1 0 14688 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_148
timestamp 1679581782
transform 1 0 15360 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_155
timestamp 1677579658
transform 1 0 16032 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_160
timestamp 1679577901
transform 1 0 16512 0 -1 8316
box -48 -56 432 834
use sg13g2_decap_8  FILLER_9_168
timestamp 1679581782
transform 1 0 17280 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_175
timestamp 1679581782
transform 1 0 17952 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_182
timestamp 1679577901
transform 1 0 18624 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_186
timestamp 1677579658
transform 1 0 19008 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_191
timestamp 1679581782
transform 1 0 19488 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_198
timestamp 1677580104
transform 1 0 20160 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_4  FILLER_10_0
timestamp 1679577901
transform 1 0 1152 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_4
timestamp 1677580104
transform 1 0 1536 0 1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_18
timestamp 1679581782
transform 1 0 2880 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_25
timestamp 1679581782
transform 1 0 3552 0 1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_32
timestamp 1677579658
transform 1 0 4224 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_45
timestamp 1677579658
transform 1 0 5472 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_50
timestamp 1677579658
transform 1 0 5952 0 1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_10_55
timestamp 1679577901
transform 1 0 6432 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_59
timestamp 1677580104
transform 1 0 6816 0 1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_69
timestamp 1677580104
transform 1 0 7776 0 1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_75
timestamp 1679581782
transform 1 0 8352 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_82
timestamp 1679581782
transform 1 0 9024 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_89
timestamp 1677580104
transform 1 0 9696 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_91
timestamp 1677579658
transform 1 0 9888 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_96
timestamp 1677580104
transform 1 0 10368 0 1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_114
timestamp 1679581782
transform 1 0 12096 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_121
timestamp 1679581782
transform 1 0 12768 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_128
timestamp 1679581782
transform 1 0 13440 0 1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_135
timestamp 1677579658
transform 1 0 14112 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_144
timestamp 1677580104
transform 1 0 14976 0 1 8316
box -48 -56 240 834
use sg13g2_decap_4  FILLER_10_150
timestamp 1679577901
transform 1 0 15552 0 1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_154
timestamp 1677579658
transform 1 0 15936 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_163
timestamp 1677580104
transform 1 0 16800 0 1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_169
timestamp 1677580104
transform 1 0 17376 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_171
timestamp 1677579658
transform 1 0 17568 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_176
timestamp 1679581782
transform 1 0 18048 0 1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_195
timestamp 1679577901
transform 1 0 19872 0 1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_199
timestamp 1677579658
transform 1 0 20256 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_0
timestamp 1679581782
transform 1 0 1152 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_7
timestamp 1679581782
transform 1 0 1824 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_14
timestamp 1679581782
transform 1 0 2496 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_21
timestamp 1679581782
transform 1 0 3168 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_28
timestamp 1679581782
transform 1 0 3840 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_35
timestamp 1679581782
transform 1 0 4512 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_42
timestamp 1679581782
transform 1 0 5184 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_49
timestamp 1679581782
transform 1 0 5856 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_56
timestamp 1679581782
transform 1 0 6528 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_63
timestamp 1679581782
transform 1 0 7200 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_70
timestamp 1679581782
transform 1 0 7872 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_77
timestamp 1679581782
transform 1 0 8544 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_84
timestamp 1679581782
transform 1 0 9216 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_91
timestamp 1679581782
transform 1 0 9888 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_98
timestamp 1679581782
transform 1 0 10560 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_105
timestamp 1679581782
transform 1 0 11232 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_112
timestamp 1679581782
transform 1 0 11904 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_119
timestamp 1679581782
transform 1 0 12576 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_126
timestamp 1679581782
transform 1 0 13248 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_133
timestamp 1679581782
transform 1 0 13920 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_140
timestamp 1679581782
transform 1 0 14592 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_147
timestamp 1679581782
transform 1 0 15264 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_154
timestamp 1679581782
transform 1 0 15936 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_161
timestamp 1679581782
transform 1 0 16608 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_168
timestamp 1679581782
transform 1 0 17280 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_175
timestamp 1679581782
transform 1 0 17952 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_182
timestamp 1679577901
transform 1 0 18624 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_11_186
timestamp 1677579658
transform 1 0 19008 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_191
timestamp 1679581782
transform 1 0 19488 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_198
timestamp 1677580104
transform 1 0 20160 0 -1 9828
box -48 -56 240 834
<< labels >>
flabel metal3 s 0 44 80 124 0 FreeSans 320 0 0 0 FrameData[0]
port 0 nsew signal input
flabel metal3 s 0 3404 80 3484 0 FreeSans 320 0 0 0 FrameData[10]
port 1 nsew signal input
flabel metal3 s 0 3740 80 3820 0 FreeSans 320 0 0 0 FrameData[11]
port 2 nsew signal input
flabel metal3 s 0 4076 80 4156 0 FreeSans 320 0 0 0 FrameData[12]
port 3 nsew signal input
flabel metal3 s 0 4412 80 4492 0 FreeSans 320 0 0 0 FrameData[13]
port 4 nsew signal input
flabel metal3 s 0 4748 80 4828 0 FreeSans 320 0 0 0 FrameData[14]
port 5 nsew signal input
flabel metal3 s 0 5084 80 5164 0 FreeSans 320 0 0 0 FrameData[15]
port 6 nsew signal input
flabel metal3 s 0 5420 80 5500 0 FreeSans 320 0 0 0 FrameData[16]
port 7 nsew signal input
flabel metal3 s 0 5756 80 5836 0 FreeSans 320 0 0 0 FrameData[17]
port 8 nsew signal input
flabel metal3 s 0 6092 80 6172 0 FreeSans 320 0 0 0 FrameData[18]
port 9 nsew signal input
flabel metal3 s 0 6428 80 6508 0 FreeSans 320 0 0 0 FrameData[19]
port 10 nsew signal input
flabel metal3 s 0 380 80 460 0 FreeSans 320 0 0 0 FrameData[1]
port 11 nsew signal input
flabel metal3 s 0 6764 80 6844 0 FreeSans 320 0 0 0 FrameData[20]
port 12 nsew signal input
flabel metal3 s 0 7100 80 7180 0 FreeSans 320 0 0 0 FrameData[21]
port 13 nsew signal input
flabel metal3 s 0 7436 80 7516 0 FreeSans 320 0 0 0 FrameData[22]
port 14 nsew signal input
flabel metal3 s 0 7772 80 7852 0 FreeSans 320 0 0 0 FrameData[23]
port 15 nsew signal input
flabel metal3 s 0 8108 80 8188 0 FreeSans 320 0 0 0 FrameData[24]
port 16 nsew signal input
flabel metal3 s 0 8444 80 8524 0 FreeSans 320 0 0 0 FrameData[25]
port 17 nsew signal input
flabel metal3 s 0 8780 80 8860 0 FreeSans 320 0 0 0 FrameData[26]
port 18 nsew signal input
flabel metal3 s 0 9116 80 9196 0 FreeSans 320 0 0 0 FrameData[27]
port 19 nsew signal input
flabel metal3 s 0 9452 80 9532 0 FreeSans 320 0 0 0 FrameData[28]
port 20 nsew signal input
flabel metal3 s 0 9788 80 9868 0 FreeSans 320 0 0 0 FrameData[29]
port 21 nsew signal input
flabel metal3 s 0 716 80 796 0 FreeSans 320 0 0 0 FrameData[2]
port 22 nsew signal input
flabel metal3 s 0 10124 80 10204 0 FreeSans 320 0 0 0 FrameData[30]
port 23 nsew signal input
flabel metal3 s 0 10460 80 10540 0 FreeSans 320 0 0 0 FrameData[31]
port 24 nsew signal input
flabel metal3 s 0 1052 80 1132 0 FreeSans 320 0 0 0 FrameData[3]
port 25 nsew signal input
flabel metal3 s 0 1388 80 1468 0 FreeSans 320 0 0 0 FrameData[4]
port 26 nsew signal input
flabel metal3 s 0 1724 80 1804 0 FreeSans 320 0 0 0 FrameData[5]
port 27 nsew signal input
flabel metal3 s 0 2060 80 2140 0 FreeSans 320 0 0 0 FrameData[6]
port 28 nsew signal input
flabel metal3 s 0 2396 80 2476 0 FreeSans 320 0 0 0 FrameData[7]
port 29 nsew signal input
flabel metal3 s 0 2732 80 2812 0 FreeSans 320 0 0 0 FrameData[8]
port 30 nsew signal input
flabel metal3 s 0 3068 80 3148 0 FreeSans 320 0 0 0 FrameData[9]
port 31 nsew signal input
flabel metal3 s 21424 44 21504 124 0 FreeSans 320 0 0 0 FrameData_O[0]
port 32 nsew signal output
flabel metal3 s 21424 3404 21504 3484 0 FreeSans 320 0 0 0 FrameData_O[10]
port 33 nsew signal output
flabel metal3 s 21424 3740 21504 3820 0 FreeSans 320 0 0 0 FrameData_O[11]
port 34 nsew signal output
flabel metal3 s 21424 4076 21504 4156 0 FreeSans 320 0 0 0 FrameData_O[12]
port 35 nsew signal output
flabel metal3 s 21424 4412 21504 4492 0 FreeSans 320 0 0 0 FrameData_O[13]
port 36 nsew signal output
flabel metal3 s 21424 4748 21504 4828 0 FreeSans 320 0 0 0 FrameData_O[14]
port 37 nsew signal output
flabel metal3 s 21424 5084 21504 5164 0 FreeSans 320 0 0 0 FrameData_O[15]
port 38 nsew signal output
flabel metal3 s 21424 5420 21504 5500 0 FreeSans 320 0 0 0 FrameData_O[16]
port 39 nsew signal output
flabel metal3 s 21424 5756 21504 5836 0 FreeSans 320 0 0 0 FrameData_O[17]
port 40 nsew signal output
flabel metal3 s 21424 6092 21504 6172 0 FreeSans 320 0 0 0 FrameData_O[18]
port 41 nsew signal output
flabel metal3 s 21424 6428 21504 6508 0 FreeSans 320 0 0 0 FrameData_O[19]
port 42 nsew signal output
flabel metal3 s 21424 380 21504 460 0 FreeSans 320 0 0 0 FrameData_O[1]
port 43 nsew signal output
flabel metal3 s 21424 6764 21504 6844 0 FreeSans 320 0 0 0 FrameData_O[20]
port 44 nsew signal output
flabel metal3 s 21424 7100 21504 7180 0 FreeSans 320 0 0 0 FrameData_O[21]
port 45 nsew signal output
flabel metal3 s 21424 7436 21504 7516 0 FreeSans 320 0 0 0 FrameData_O[22]
port 46 nsew signal output
flabel metal3 s 21424 7772 21504 7852 0 FreeSans 320 0 0 0 FrameData_O[23]
port 47 nsew signal output
flabel metal3 s 21424 8108 21504 8188 0 FreeSans 320 0 0 0 FrameData_O[24]
port 48 nsew signal output
flabel metal3 s 21424 8444 21504 8524 0 FreeSans 320 0 0 0 FrameData_O[25]
port 49 nsew signal output
flabel metal3 s 21424 8780 21504 8860 0 FreeSans 320 0 0 0 FrameData_O[26]
port 50 nsew signal output
flabel metal3 s 21424 9116 21504 9196 0 FreeSans 320 0 0 0 FrameData_O[27]
port 51 nsew signal output
flabel metal3 s 21424 9452 21504 9532 0 FreeSans 320 0 0 0 FrameData_O[28]
port 52 nsew signal output
flabel metal3 s 21424 9788 21504 9868 0 FreeSans 320 0 0 0 FrameData_O[29]
port 53 nsew signal output
flabel metal3 s 21424 716 21504 796 0 FreeSans 320 0 0 0 FrameData_O[2]
port 54 nsew signal output
flabel metal3 s 21424 10124 21504 10204 0 FreeSans 320 0 0 0 FrameData_O[30]
port 55 nsew signal output
flabel metal3 s 21424 10460 21504 10540 0 FreeSans 320 0 0 0 FrameData_O[31]
port 56 nsew signal output
flabel metal3 s 21424 1052 21504 1132 0 FreeSans 320 0 0 0 FrameData_O[3]
port 57 nsew signal output
flabel metal3 s 21424 1388 21504 1468 0 FreeSans 320 0 0 0 FrameData_O[4]
port 58 nsew signal output
flabel metal3 s 21424 1724 21504 1804 0 FreeSans 320 0 0 0 FrameData_O[5]
port 59 nsew signal output
flabel metal3 s 21424 2060 21504 2140 0 FreeSans 320 0 0 0 FrameData_O[6]
port 60 nsew signal output
flabel metal3 s 21424 2396 21504 2476 0 FreeSans 320 0 0 0 FrameData_O[7]
port 61 nsew signal output
flabel metal3 s 21424 2732 21504 2812 0 FreeSans 320 0 0 0 FrameData_O[8]
port 62 nsew signal output
flabel metal3 s 21424 3068 21504 3148 0 FreeSans 320 0 0 0 FrameData_O[9]
port 63 nsew signal output
flabel metal2 s 1976 0 2056 80 0 FreeSans 320 0 0 0 FrameStrobe[0]
port 64 nsew signal input
flabel metal2 s 11576 0 11656 80 0 FreeSans 320 0 0 0 FrameStrobe[10]
port 65 nsew signal input
flabel metal2 s 12536 0 12616 80 0 FreeSans 320 0 0 0 FrameStrobe[11]
port 66 nsew signal input
flabel metal2 s 13496 0 13576 80 0 FreeSans 320 0 0 0 FrameStrobe[12]
port 67 nsew signal input
flabel metal2 s 14456 0 14536 80 0 FreeSans 320 0 0 0 FrameStrobe[13]
port 68 nsew signal input
flabel metal2 s 15416 0 15496 80 0 FreeSans 320 0 0 0 FrameStrobe[14]
port 69 nsew signal input
flabel metal2 s 16376 0 16456 80 0 FreeSans 320 0 0 0 FrameStrobe[15]
port 70 nsew signal input
flabel metal2 s 17336 0 17416 80 0 FreeSans 320 0 0 0 FrameStrobe[16]
port 71 nsew signal input
flabel metal2 s 18296 0 18376 80 0 FreeSans 320 0 0 0 FrameStrobe[17]
port 72 nsew signal input
flabel metal2 s 19256 0 19336 80 0 FreeSans 320 0 0 0 FrameStrobe[18]
port 73 nsew signal input
flabel metal2 s 20216 0 20296 80 0 FreeSans 320 0 0 0 FrameStrobe[19]
port 74 nsew signal input
flabel metal2 s 2936 0 3016 80 0 FreeSans 320 0 0 0 FrameStrobe[1]
port 75 nsew signal input
flabel metal2 s 3896 0 3976 80 0 FreeSans 320 0 0 0 FrameStrobe[2]
port 76 nsew signal input
flabel metal2 s 4856 0 4936 80 0 FreeSans 320 0 0 0 FrameStrobe[3]
port 77 nsew signal input
flabel metal2 s 5816 0 5896 80 0 FreeSans 320 0 0 0 FrameStrobe[4]
port 78 nsew signal input
flabel metal2 s 6776 0 6856 80 0 FreeSans 320 0 0 0 FrameStrobe[5]
port 79 nsew signal input
flabel metal2 s 7736 0 7816 80 0 FreeSans 320 0 0 0 FrameStrobe[6]
port 80 nsew signal input
flabel metal2 s 8696 0 8776 80 0 FreeSans 320 0 0 0 FrameStrobe[7]
port 81 nsew signal input
flabel metal2 s 9656 0 9736 80 0 FreeSans 320 0 0 0 FrameStrobe[8]
port 82 nsew signal input
flabel metal2 s 10616 0 10696 80 0 FreeSans 320 0 0 0 FrameStrobe[9]
port 83 nsew signal input
flabel metal2 s 15800 10672 15880 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[0]
port 84 nsew signal output
flabel metal2 s 17720 10672 17800 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[10]
port 85 nsew signal output
flabel metal2 s 17912 10672 17992 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[11]
port 86 nsew signal output
flabel metal2 s 18104 10672 18184 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[12]
port 87 nsew signal output
flabel metal2 s 18296 10672 18376 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[13]
port 88 nsew signal output
flabel metal2 s 18488 10672 18568 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[14]
port 89 nsew signal output
flabel metal2 s 18680 10672 18760 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[15]
port 90 nsew signal output
flabel metal2 s 18872 10672 18952 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[16]
port 91 nsew signal output
flabel metal2 s 19064 10672 19144 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[17]
port 92 nsew signal output
flabel metal2 s 19256 10672 19336 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[18]
port 93 nsew signal output
flabel metal2 s 19448 10672 19528 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[19]
port 94 nsew signal output
flabel metal2 s 15992 10672 16072 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[1]
port 95 nsew signal output
flabel metal2 s 16184 10672 16264 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[2]
port 96 nsew signal output
flabel metal2 s 16376 10672 16456 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[3]
port 97 nsew signal output
flabel metal2 s 16568 10672 16648 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[4]
port 98 nsew signal output
flabel metal2 s 16760 10672 16840 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[5]
port 99 nsew signal output
flabel metal2 s 16952 10672 17032 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[6]
port 100 nsew signal output
flabel metal2 s 17144 10672 17224 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[7]
port 101 nsew signal output
flabel metal2 s 17336 10672 17416 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[8]
port 102 nsew signal output
flabel metal2 s 17528 10672 17608 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[9]
port 103 nsew signal output
flabel metal2 s 1784 10672 1864 10752 0 FreeSans 320 0 0 0 N1BEG[0]
port 104 nsew signal output
flabel metal2 s 1976 10672 2056 10752 0 FreeSans 320 0 0 0 N1BEG[1]
port 105 nsew signal output
flabel metal2 s 2168 10672 2248 10752 0 FreeSans 320 0 0 0 N1BEG[2]
port 106 nsew signal output
flabel metal2 s 2360 10672 2440 10752 0 FreeSans 320 0 0 0 N1BEG[3]
port 107 nsew signal output
flabel metal2 s 2552 10672 2632 10752 0 FreeSans 320 0 0 0 N2BEG[0]
port 108 nsew signal output
flabel metal2 s 2744 10672 2824 10752 0 FreeSans 320 0 0 0 N2BEG[1]
port 109 nsew signal output
flabel metal2 s 2936 10672 3016 10752 0 FreeSans 320 0 0 0 N2BEG[2]
port 110 nsew signal output
flabel metal2 s 3128 10672 3208 10752 0 FreeSans 320 0 0 0 N2BEG[3]
port 111 nsew signal output
flabel metal2 s 3320 10672 3400 10752 0 FreeSans 320 0 0 0 N2BEG[4]
port 112 nsew signal output
flabel metal2 s 3512 10672 3592 10752 0 FreeSans 320 0 0 0 N2BEG[5]
port 113 nsew signal output
flabel metal2 s 3704 10672 3784 10752 0 FreeSans 320 0 0 0 N2BEG[6]
port 114 nsew signal output
flabel metal2 s 3896 10672 3976 10752 0 FreeSans 320 0 0 0 N2BEG[7]
port 115 nsew signal output
flabel metal2 s 4088 10672 4168 10752 0 FreeSans 320 0 0 0 N2BEGb[0]
port 116 nsew signal output
flabel metal2 s 4280 10672 4360 10752 0 FreeSans 320 0 0 0 N2BEGb[1]
port 117 nsew signal output
flabel metal2 s 4472 10672 4552 10752 0 FreeSans 320 0 0 0 N2BEGb[2]
port 118 nsew signal output
flabel metal2 s 4664 10672 4744 10752 0 FreeSans 320 0 0 0 N2BEGb[3]
port 119 nsew signal output
flabel metal2 s 4856 10672 4936 10752 0 FreeSans 320 0 0 0 N2BEGb[4]
port 120 nsew signal output
flabel metal2 s 5048 10672 5128 10752 0 FreeSans 320 0 0 0 N2BEGb[5]
port 121 nsew signal output
flabel metal2 s 5240 10672 5320 10752 0 FreeSans 320 0 0 0 N2BEGb[6]
port 122 nsew signal output
flabel metal2 s 5432 10672 5512 10752 0 FreeSans 320 0 0 0 N2BEGb[7]
port 123 nsew signal output
flabel metal2 s 5624 10672 5704 10752 0 FreeSans 320 0 0 0 N4BEG[0]
port 124 nsew signal output
flabel metal2 s 7544 10672 7624 10752 0 FreeSans 320 0 0 0 N4BEG[10]
port 125 nsew signal output
flabel metal2 s 7736 10672 7816 10752 0 FreeSans 320 0 0 0 N4BEG[11]
port 126 nsew signal output
flabel metal2 s 7928 10672 8008 10752 0 FreeSans 320 0 0 0 N4BEG[12]
port 127 nsew signal output
flabel metal2 s 8120 10672 8200 10752 0 FreeSans 320 0 0 0 N4BEG[13]
port 128 nsew signal output
flabel metal2 s 8312 10672 8392 10752 0 FreeSans 320 0 0 0 N4BEG[14]
port 129 nsew signal output
flabel metal2 s 8504 10672 8584 10752 0 FreeSans 320 0 0 0 N4BEG[15]
port 130 nsew signal output
flabel metal2 s 5816 10672 5896 10752 0 FreeSans 320 0 0 0 N4BEG[1]
port 131 nsew signal output
flabel metal2 s 6008 10672 6088 10752 0 FreeSans 320 0 0 0 N4BEG[2]
port 132 nsew signal output
flabel metal2 s 6200 10672 6280 10752 0 FreeSans 320 0 0 0 N4BEG[3]
port 133 nsew signal output
flabel metal2 s 6392 10672 6472 10752 0 FreeSans 320 0 0 0 N4BEG[4]
port 134 nsew signal output
flabel metal2 s 6584 10672 6664 10752 0 FreeSans 320 0 0 0 N4BEG[5]
port 135 nsew signal output
flabel metal2 s 6776 10672 6856 10752 0 FreeSans 320 0 0 0 N4BEG[6]
port 136 nsew signal output
flabel metal2 s 6968 10672 7048 10752 0 FreeSans 320 0 0 0 N4BEG[7]
port 137 nsew signal output
flabel metal2 s 7160 10672 7240 10752 0 FreeSans 320 0 0 0 N4BEG[8]
port 138 nsew signal output
flabel metal2 s 7352 10672 7432 10752 0 FreeSans 320 0 0 0 N4BEG[9]
port 139 nsew signal output
flabel metal2 s 8696 10672 8776 10752 0 FreeSans 320 0 0 0 S1END[0]
port 140 nsew signal input
flabel metal2 s 8888 10672 8968 10752 0 FreeSans 320 0 0 0 S1END[1]
port 141 nsew signal input
flabel metal2 s 9080 10672 9160 10752 0 FreeSans 320 0 0 0 S1END[2]
port 142 nsew signal input
flabel metal2 s 9272 10672 9352 10752 0 FreeSans 320 0 0 0 S1END[3]
port 143 nsew signal input
flabel metal2 s 11000 10672 11080 10752 0 FreeSans 320 0 0 0 S2END[0]
port 144 nsew signal input
flabel metal2 s 11192 10672 11272 10752 0 FreeSans 320 0 0 0 S2END[1]
port 145 nsew signal input
flabel metal2 s 11384 10672 11464 10752 0 FreeSans 320 0 0 0 S2END[2]
port 146 nsew signal input
flabel metal2 s 11576 10672 11656 10752 0 FreeSans 320 0 0 0 S2END[3]
port 147 nsew signal input
flabel metal2 s 11768 10672 11848 10752 0 FreeSans 320 0 0 0 S2END[4]
port 148 nsew signal input
flabel metal2 s 11960 10672 12040 10752 0 FreeSans 320 0 0 0 S2END[5]
port 149 nsew signal input
flabel metal2 s 12152 10672 12232 10752 0 FreeSans 320 0 0 0 S2END[6]
port 150 nsew signal input
flabel metal2 s 12344 10672 12424 10752 0 FreeSans 320 0 0 0 S2END[7]
port 151 nsew signal input
flabel metal2 s 9464 10672 9544 10752 0 FreeSans 320 0 0 0 S2MID[0]
port 152 nsew signal input
flabel metal2 s 9656 10672 9736 10752 0 FreeSans 320 0 0 0 S2MID[1]
port 153 nsew signal input
flabel metal2 s 9848 10672 9928 10752 0 FreeSans 320 0 0 0 S2MID[2]
port 154 nsew signal input
flabel metal2 s 10040 10672 10120 10752 0 FreeSans 320 0 0 0 S2MID[3]
port 155 nsew signal input
flabel metal2 s 10232 10672 10312 10752 0 FreeSans 320 0 0 0 S2MID[4]
port 156 nsew signal input
flabel metal2 s 10424 10672 10504 10752 0 FreeSans 320 0 0 0 S2MID[5]
port 157 nsew signal input
flabel metal2 s 10616 10672 10696 10752 0 FreeSans 320 0 0 0 S2MID[6]
port 158 nsew signal input
flabel metal2 s 10808 10672 10888 10752 0 FreeSans 320 0 0 0 S2MID[7]
port 159 nsew signal input
flabel metal2 s 12536 10672 12616 10752 0 FreeSans 320 0 0 0 S4END[0]
port 160 nsew signal input
flabel metal2 s 14456 10672 14536 10752 0 FreeSans 320 0 0 0 S4END[10]
port 161 nsew signal input
flabel metal2 s 14648 10672 14728 10752 0 FreeSans 320 0 0 0 S4END[11]
port 162 nsew signal input
flabel metal2 s 14840 10672 14920 10752 0 FreeSans 320 0 0 0 S4END[12]
port 163 nsew signal input
flabel metal2 s 15032 10672 15112 10752 0 FreeSans 320 0 0 0 S4END[13]
port 164 nsew signal input
flabel metal2 s 15224 10672 15304 10752 0 FreeSans 320 0 0 0 S4END[14]
port 165 nsew signal input
flabel metal2 s 15416 10672 15496 10752 0 FreeSans 320 0 0 0 S4END[15]
port 166 nsew signal input
flabel metal2 s 12728 10672 12808 10752 0 FreeSans 320 0 0 0 S4END[1]
port 167 nsew signal input
flabel metal2 s 12920 10672 13000 10752 0 FreeSans 320 0 0 0 S4END[2]
port 168 nsew signal input
flabel metal2 s 13112 10672 13192 10752 0 FreeSans 320 0 0 0 S4END[3]
port 169 nsew signal input
flabel metal2 s 13304 10672 13384 10752 0 FreeSans 320 0 0 0 S4END[4]
port 170 nsew signal input
flabel metal2 s 13496 10672 13576 10752 0 FreeSans 320 0 0 0 S4END[5]
port 171 nsew signal input
flabel metal2 s 13688 10672 13768 10752 0 FreeSans 320 0 0 0 S4END[6]
port 172 nsew signal input
flabel metal2 s 13880 10672 13960 10752 0 FreeSans 320 0 0 0 S4END[7]
port 173 nsew signal input
flabel metal2 s 14072 10672 14152 10752 0 FreeSans 320 0 0 0 S4END[8]
port 174 nsew signal input
flabel metal2 s 14264 10672 14344 10752 0 FreeSans 320 0 0 0 S4END[9]
port 175 nsew signal input
flabel metal2 s 1016 0 1096 80 0 FreeSans 320 0 0 0 UserCLK
port 176 nsew signal input
flabel metal2 s 15608 10672 15688 10752 0 FreeSans 320 0 0 0 UserCLKo
port 177 nsew signal output
flabel metal6 s 4892 0 5332 10752 0 FreeSans 2624 90 0 0 VGND
port 178 nsew ground bidirectional
flabel metal6 s 4892 0 5332 328 0 FreeSans 2624 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal6 s 4892 10424 5332 10752 0 FreeSans 2624 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal6 s 20012 0 20452 10752 0 FreeSans 2624 90 0 0 VGND
port 178 nsew ground bidirectional
flabel metal6 s 20012 0 20452 328 0 FreeSans 2624 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal6 s 20012 10424 20452 10752 0 FreeSans 2624 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal6 s 3652 0 4092 10752 0 FreeSans 2624 90 0 0 VPWR
port 179 nsew power bidirectional
flabel metal6 s 3652 0 4092 328 0 FreeSans 2624 0 0 0 VPWR
port 179 nsew power bidirectional
flabel metal6 s 3652 10424 4092 10752 0 FreeSans 2624 0 0 0 VPWR
port 179 nsew power bidirectional
flabel metal6 s 18772 0 19212 10752 0 FreeSans 2624 90 0 0 VPWR
port 179 nsew power bidirectional
flabel metal6 s 18772 0 19212 328 0 FreeSans 2624 0 0 0 VPWR
port 179 nsew power bidirectional
flabel metal6 s 18772 10424 19212 10752 0 FreeSans 2624 0 0 0 VPWR
port 179 nsew power bidirectional
rlabel metal1 10802 9828 10802 9828 0 VGND
rlabel metal1 10752 9072 10752 9072 0 VPWR
rlabel metal3 990 84 990 84 0 FrameData[0]
rlabel metal2 9792 3822 9792 3822 0 FrameData[10]
rlabel metal3 1614 3780 1614 3780 0 FrameData[11]
rlabel metal2 12912 4116 12912 4116 0 FrameData[12]
rlabel metal3 1374 4452 1374 4452 0 FrameData[13]
rlabel metal3 1182 4788 1182 4788 0 FrameData[14]
rlabel metal3 1182 5124 1182 5124 0 FrameData[15]
rlabel metal2 12192 5586 12192 5586 0 FrameData[16]
rlabel metal3 270 5796 270 5796 0 FrameData[17]
rlabel metal3 1038 6132 1038 6132 0 FrameData[18]
rlabel metal2 19392 5838 19392 5838 0 FrameData[19]
rlabel metal3 798 420 798 420 0 FrameData[1]
rlabel metal3 1614 6804 1614 6804 0 FrameData[20]
rlabel metal2 19392 6762 19392 6762 0 FrameData[21]
rlabel metal3 2238 7476 2238 7476 0 FrameData[22]
rlabel metal2 16800 5796 16800 5796 0 FrameData[23]
rlabel metal3 798 8148 798 8148 0 FrameData[24]
rlabel metal3 846 8484 846 8484 0 FrameData[25]
rlabel metal3 126 8820 126 8820 0 FrameData[26]
rlabel metal3 222 9156 222 9156 0 FrameData[27]
rlabel metal3 2574 9492 2574 9492 0 FrameData[28]
rlabel metal3 366 9828 366 9828 0 FrameData[29]
rlabel metal3 2382 756 2382 756 0 FrameData[2]
rlabel metal3 606 10164 606 10164 0 FrameData[30]
rlabel metal3 318 10500 318 10500 0 FrameData[31]
rlabel metal2 8352 1470 8352 1470 0 FrameData[3]
rlabel metal3 1182 1428 1182 1428 0 FrameData[4]
rlabel metal3 17304 1848 17304 1848 0 FrameData[5]
rlabel metal3 3054 2100 3054 2100 0 FrameData[6]
rlabel metal3 1134 2436 1134 2436 0 FrameData[7]
rlabel metal3 3180 2772 3180 2772 0 FrameData[8]
rlabel metal3 990 3108 990 3108 0 FrameData[9]
rlabel metal2 3552 882 3552 882 0 FrameData_O[0]
rlabel metal2 9984 3696 9984 3696 0 FrameData_O[10]
rlabel metal3 21426 3780 21426 3780 0 FrameData_O[11]
rlabel metal2 13152 4032 13152 4032 0 FrameData_O[12]
rlabel metal2 3216 3864 3216 3864 0 FrameData_O[13]
rlabel metal3 2496 3990 2496 3990 0 FrameData_O[14]
rlabel metal2 2496 4956 2496 4956 0 FrameData_O[15]
rlabel metal3 16914 5460 16914 5460 0 FrameData_O[16]
rlabel metal2 19296 5082 19296 5082 0 FrameData_O[17]
rlabel metal3 2208 6174 2208 6174 0 FrameData_O[18]
rlabel metal2 19584 6090 19584 6090 0 FrameData_O[19]
rlabel metal2 1728 1050 1728 1050 0 FrameData_O[1]
rlabel metal2 19200 6678 19200 6678 0 FrameData_O[20]
rlabel metal2 19584 6888 19584 6888 0 FrameData_O[21]
rlabel metal3 20082 7476 20082 7476 0 FrameData_O[22]
rlabel metal2 17040 5880 17040 5880 0 FrameData_O[23]
rlabel metal2 17952 7392 17952 7392 0 FrameData_O[24]
rlabel metal3 20034 8484 20034 8484 0 FrameData_O[25]
rlabel metal3 19746 8820 19746 8820 0 FrameData_O[26]
rlabel metal2 19392 8988 19392 8988 0 FrameData_O[27]
rlabel metal2 19008 8862 19008 8862 0 FrameData_O[28]
rlabel metal2 19776 9282 19776 9282 0 FrameData_O[29]
rlabel metal2 4896 1302 4896 1302 0 FrameData_O[2]
rlabel metal2 19440 8148 19440 8148 0 FrameData_O[30]
rlabel metal2 19392 10080 19392 10080 0 FrameData_O[31]
rlabel metal2 8544 1386 8544 1386 0 FrameData_O[3]
rlabel metal2 2496 1554 2496 1554 0 FrameData_O[4]
rlabel metal3 20562 1764 20562 1764 0 FrameData_O[5]
rlabel metal2 6240 1596 6240 1596 0 FrameData_O[6]
rlabel metal2 2400 3066 2400 3066 0 FrameData_O[7]
rlabel metal3 20658 2772 20658 2772 0 FrameData_O[8]
rlabel metal2 2112 3612 2112 3612 0 FrameData_O[9]
rlabel metal2 2016 492 2016 492 0 FrameStrobe[0]
rlabel metal2 11616 660 11616 660 0 FrameStrobe[10]
rlabel metal2 17472 1302 17472 1302 0 FrameStrobe[11]
rlabel metal2 13536 954 13536 954 0 FrameStrobe[12]
rlabel metal2 16224 7224 16224 7224 0 FrameStrobe[13]
rlabel metal2 15456 114 15456 114 0 FrameStrobe[14]
rlabel metal2 16416 114 16416 114 0 FrameStrobe[15]
rlabel metal2 17376 1290 17376 1290 0 FrameStrobe[16]
rlabel metal2 18336 114 18336 114 0 FrameStrobe[17]
rlabel metal2 19296 492 19296 492 0 FrameStrobe[18]
rlabel metal2 20256 72 20256 72 0 FrameStrobe[19]
rlabel metal2 2976 660 2976 660 0 FrameStrobe[1]
rlabel metal2 3936 702 3936 702 0 FrameStrobe[2]
rlabel metal2 4896 198 4896 198 0 FrameStrobe[3]
rlabel metal2 5856 114 5856 114 0 FrameStrobe[4]
rlabel metal2 15744 1050 15744 1050 0 FrameStrobe[5]
rlabel metal2 16224 1092 16224 1092 0 FrameStrobe[6]
rlabel metal2 8736 954 8736 954 0 FrameStrobe[7]
rlabel metal2 9696 660 9696 660 0 FrameStrobe[8]
rlabel metal2 10656 954 10656 954 0 FrameStrobe[9]
rlabel metal2 4128 2142 4128 2142 0 FrameStrobe_O[0]
rlabel metal2 17760 9966 17760 9966 0 FrameStrobe_O[10]
rlabel metal2 17952 9882 17952 9882 0 FrameStrobe_O[11]
rlabel metal2 18144 10092 18144 10092 0 FrameStrobe_O[12]
rlabel metal3 17376 7812 17376 7812 0 FrameStrobe_O[13]
rlabel metal2 16512 7140 16512 7140 0 FrameStrobe_O[14]
rlabel metal2 17184 8526 17184 8526 0 FrameStrobe_O[15]
rlabel metal2 16320 9072 16320 9072 0 FrameStrobe_O[16]
rlabel metal2 18048 4200 18048 4200 0 FrameStrobe_O[17]
rlabel metal3 19632 2100 19632 2100 0 FrameStrobe_O[18]
rlabel via2 19488 10680 19488 10680 0 FrameStrobe_O[19]
rlabel metal2 16032 9798 16032 9798 0 FrameStrobe_O[1]
rlabel metal2 5856 3234 5856 3234 0 FrameStrobe_O[2]
rlabel metal2 16416 9588 16416 9588 0 FrameStrobe_O[3]
rlabel metal2 16608 9042 16608 9042 0 FrameStrobe_O[4]
rlabel metal2 15936 4158 15936 4158 0 FrameStrobe_O[5]
rlabel metal2 16992 9588 16992 9588 0 FrameStrobe_O[6]
rlabel metal2 17184 9966 17184 9966 0 FrameStrobe_O[7]
rlabel metal2 17376 9294 17376 9294 0 FrameStrobe_O[8]
rlabel metal2 17568 7236 17568 7236 0 FrameStrobe_O[9]
rlabel metal3 2160 8484 2160 8484 0 N1BEG[0]
rlabel metal2 2112 8820 2112 8820 0 N1BEG[1]
rlabel metal2 2160 8484 2160 8484 0 N1BEG[2]
rlabel metal3 2304 8148 2304 8148 0 N1BEG[3]
rlabel metal2 2064 7392 2064 7392 0 N2BEG[0]
rlabel metal2 2736 8148 2736 8148 0 N2BEG[1]
rlabel metal2 3360 8064 3360 8064 0 N2BEG[2]
rlabel metal3 3648 8148 3648 8148 0 N2BEG[3]
rlabel metal3 4032 8484 4032 8484 0 N2BEG[4]
rlabel metal3 3984 8820 3984 8820 0 N2BEG[5]
rlabel metal2 3744 10638 3744 10638 0 N2BEG[6]
rlabel metal2 3936 9966 3936 9966 0 N2BEG[7]
rlabel metal2 5184 8778 5184 8778 0 N2BEGb[0]
rlabel metal2 5664 8736 5664 8736 0 N2BEGb[1]
rlabel metal2 6144 8526 6144 8526 0 N2BEGb[2]
rlabel metal2 4704 9462 4704 9462 0 N2BEGb[3]
rlabel metal2 4896 10344 4896 10344 0 N2BEGb[4]
rlabel metal2 5088 10428 5088 10428 0 N2BEGb[5]
rlabel metal2 5280 10386 5280 10386 0 N2BEGb[6]
rlabel metal2 5472 9924 5472 9924 0 N2BEGb[7]
rlabel metal2 5664 10260 5664 10260 0 N4BEG[0]
rlabel metal2 11040 9156 11040 9156 0 N4BEG[10]
rlabel metal2 7728 8148 7728 8148 0 N4BEG[11]
rlabel metal2 8016 8148 8016 8148 0 N4BEG[12]
rlabel metal3 8880 8148 8880 8148 0 N4BEG[13]
rlabel metal2 9984 8190 9984 8190 0 N4BEG[14]
rlabel metal3 9600 8820 9600 8820 0 N4BEG[15]
rlabel via2 5856 10680 5856 10680 0 N4BEG[1]
rlabel metal2 6048 9084 6048 9084 0 N4BEG[2]
rlabel metal2 6240 8454 6240 8454 0 N4BEG[3]
rlabel metal2 14304 7938 14304 7938 0 N4BEG[4]
rlabel metal2 13680 8148 13680 8148 0 N4BEG[5]
rlabel metal2 13248 9156 13248 9156 0 N4BEG[6]
rlabel metal2 12768 7518 12768 7518 0 N4BEG[7]
rlabel metal3 9504 8484 9504 8484 0 N4BEG[8]
rlabel metal2 11424 8358 11424 8358 0 N4BEG[9]
rlabel metal3 4128 9114 4128 9114 0 S1END[0]
rlabel metal2 1824 7896 1824 7896 0 S1END[1]
rlabel metal2 2400 7812 2400 7812 0 S1END[2]
rlabel metal2 2880 9492 2880 9492 0 S1END[3]
rlabel metal2 11040 10176 11040 10176 0 S2END[0]
rlabel metal2 11232 10218 11232 10218 0 S2END[1]
rlabel metal2 11424 10218 11424 10218 0 S2END[2]
rlabel metal2 11616 10218 11616 10218 0 S2END[3]
rlabel metal2 11808 9756 11808 9756 0 S2END[4]
rlabel metal2 12000 10680 12000 10680 0 S2END[5]
rlabel metal2 5856 9324 5856 9324 0 S2END[6]
rlabel metal2 5376 9576 5376 9576 0 S2END[7]
rlabel metal2 9504 9714 9504 9714 0 S2MID[0]
rlabel metal2 9696 9294 9696 9294 0 S2MID[1]
rlabel metal2 4608 8442 4608 8442 0 S2MID[2]
rlabel metal2 4992 9198 4992 9198 0 S2MID[3]
rlabel metal2 4224 8736 4224 8736 0 S2MID[4]
rlabel metal2 3456 9114 3456 9114 0 S2MID[5]
rlabel metal2 2592 7434 2592 7434 0 S2MID[6]
rlabel metal2 10848 10596 10848 10596 0 S2MID[7]
rlabel metal2 12576 9714 12576 9714 0 S4END[0]
rlabel metal2 14496 10008 14496 10008 0 S4END[10]
rlabel metal2 14688 9714 14688 9714 0 S4END[11]
rlabel metal2 14880 9714 14880 9714 0 S4END[12]
rlabel metal2 15072 9714 15072 9714 0 S4END[13]
rlabel metal2 15264 9756 15264 9756 0 S4END[14]
rlabel metal2 15456 10218 15456 10218 0 S4END[15]
rlabel metal2 12768 9966 12768 9966 0 S4END[1]
rlabel metal2 12960 10260 12960 10260 0 S4END[2]
rlabel metal2 13152 10008 13152 10008 0 S4END[3]
rlabel metal2 13344 10050 13344 10050 0 S4END[4]
rlabel metal2 13536 10134 13536 10134 0 S4END[5]
rlabel metal2 13728 9630 13728 9630 0 S4END[6]
rlabel metal2 13920 10218 13920 10218 0 S4END[7]
rlabel metal2 14112 9294 14112 9294 0 S4END[8]
rlabel metal2 14304 9756 14304 9756 0 S4END[9]
rlabel metal2 1056 954 1056 954 0 UserCLK
rlabel metal2 3456 2604 3456 2604 0 UserCLKo
<< properties >>
string FIXED_BBOX 0 0 21504 10752
<< end >>
