magic
tech ihp-sg13g2
magscale 1 2
timestamp 1755182808
<< metal1 >>
rect 1152 84692 20352 84716
rect 1152 84652 3688 84692
rect 3728 84652 3770 84692
rect 3810 84652 3852 84692
rect 3892 84652 3934 84692
rect 3974 84652 4016 84692
rect 4056 84652 18808 84692
rect 18848 84652 18890 84692
rect 18930 84652 18972 84692
rect 19012 84652 19054 84692
rect 19094 84652 19136 84692
rect 19176 84652 20352 84692
rect 1152 84628 20352 84652
rect 3051 84440 3093 84449
rect 3051 84400 3052 84440
rect 3092 84400 3093 84440
rect 3051 84391 3093 84400
rect 3435 84440 3477 84449
rect 3435 84400 3436 84440
rect 3476 84400 3477 84440
rect 3435 84391 3477 84400
rect 3235 84356 3293 84357
rect 3235 84316 3244 84356
rect 3284 84316 3293 84356
rect 3235 84315 3293 84316
rect 3619 84356 3677 84357
rect 3619 84316 3628 84356
rect 3668 84316 3677 84356
rect 3619 84315 3677 84316
rect 18115 84104 18173 84105
rect 18115 84064 18124 84104
rect 18164 84064 18173 84104
rect 18115 84063 18173 84064
rect 18499 84104 18557 84105
rect 18499 84064 18508 84104
rect 18548 84064 18557 84104
rect 18499 84063 18557 84064
rect 18987 84104 19029 84113
rect 18987 84064 18988 84104
rect 19028 84064 19029 84104
rect 18987 84055 19029 84064
rect 19267 84104 19325 84105
rect 19267 84064 19276 84104
rect 19316 84064 19325 84104
rect 19267 84063 19325 84064
rect 1152 83936 20452 83960
rect 1152 83896 4928 83936
rect 4968 83896 5010 83936
rect 5050 83896 5092 83936
rect 5132 83896 5174 83936
rect 5214 83896 5256 83936
rect 5296 83896 20048 83936
rect 20088 83896 20130 83936
rect 20170 83896 20212 83936
rect 20252 83896 20294 83936
rect 20334 83896 20376 83936
rect 20416 83896 20452 83936
rect 1152 83872 20452 83896
rect 1899 83768 1941 83777
rect 1899 83728 1900 83768
rect 1940 83728 1941 83768
rect 1899 83719 1941 83728
rect 2283 83768 2325 83777
rect 2283 83728 2284 83768
rect 2324 83728 2325 83768
rect 2283 83719 2325 83728
rect 2667 83768 2709 83777
rect 2667 83728 2668 83768
rect 2708 83728 2709 83768
rect 2667 83719 2709 83728
rect 3051 83768 3093 83777
rect 3051 83728 3052 83768
rect 3092 83728 3093 83768
rect 3051 83719 3093 83728
rect 3435 83768 3477 83777
rect 3435 83728 3436 83768
rect 3476 83728 3477 83768
rect 3435 83719 3477 83728
rect 3819 83768 3861 83777
rect 3819 83728 3820 83768
rect 3860 83728 3861 83768
rect 3819 83719 3861 83728
rect 4203 83768 4245 83777
rect 4203 83728 4204 83768
rect 4244 83728 4245 83768
rect 4203 83719 4245 83728
rect 5355 83768 5397 83777
rect 5355 83728 5356 83768
rect 5396 83728 5397 83768
rect 5355 83719 5397 83728
rect 5547 83768 5589 83777
rect 5547 83728 5548 83768
rect 5588 83728 5589 83768
rect 5547 83719 5589 83728
rect 6219 83768 6261 83777
rect 6219 83728 6220 83768
rect 6260 83728 6261 83768
rect 6219 83719 6261 83728
rect 6411 83768 6453 83777
rect 6411 83728 6412 83768
rect 6452 83728 6453 83768
rect 6411 83719 6453 83728
rect 6987 83768 7029 83777
rect 6987 83728 6988 83768
rect 7028 83728 7029 83768
rect 6987 83719 7029 83728
rect 7563 83768 7605 83777
rect 7563 83728 7564 83768
rect 7604 83728 7605 83768
rect 7563 83719 7605 83728
rect 8427 83768 8469 83777
rect 8427 83728 8428 83768
rect 8468 83728 8469 83768
rect 8427 83719 8469 83728
rect 8811 83768 8853 83777
rect 8811 83728 8812 83768
rect 8852 83728 8853 83768
rect 8811 83719 8853 83728
rect 9579 83768 9621 83777
rect 9579 83728 9580 83768
rect 9620 83728 9621 83768
rect 9579 83719 9621 83728
rect 10059 83768 10101 83777
rect 10059 83728 10060 83768
rect 10100 83728 10101 83768
rect 10059 83719 10101 83728
rect 10443 83768 10485 83777
rect 10443 83728 10444 83768
rect 10484 83728 10485 83768
rect 10443 83719 10485 83728
rect 11307 83768 11349 83777
rect 11307 83728 11308 83768
rect 11348 83728 11349 83768
rect 11307 83719 11349 83728
rect 15723 83768 15765 83777
rect 15723 83728 15724 83768
rect 15764 83728 15765 83768
rect 15723 83719 15765 83728
rect 16779 83768 16821 83777
rect 16779 83728 16780 83768
rect 16820 83728 16821 83768
rect 16779 83719 16821 83728
rect 17355 83768 17397 83777
rect 17355 83728 17356 83768
rect 17396 83728 17397 83768
rect 17355 83719 17397 83728
rect 17739 83768 17781 83777
rect 17739 83728 17740 83768
rect 17780 83728 17781 83768
rect 17739 83719 17781 83728
rect 18891 83768 18933 83777
rect 18891 83728 18892 83768
rect 18932 83728 18933 83768
rect 18891 83719 18933 83728
rect 19659 83768 19701 83777
rect 19659 83728 19660 83768
rect 19700 83728 19701 83768
rect 19659 83719 19701 83728
rect 20043 83768 20085 83777
rect 20043 83728 20044 83768
rect 20084 83728 20085 83768
rect 20043 83719 20085 83728
rect 1699 83516 1757 83517
rect 1699 83476 1708 83516
rect 1748 83476 1757 83516
rect 1699 83475 1757 83476
rect 2083 83516 2141 83517
rect 2083 83476 2092 83516
rect 2132 83476 2141 83516
rect 2083 83475 2141 83476
rect 2467 83516 2525 83517
rect 2467 83476 2476 83516
rect 2516 83476 2525 83516
rect 2467 83475 2525 83476
rect 2851 83516 2909 83517
rect 2851 83476 2860 83516
rect 2900 83476 2909 83516
rect 2851 83475 2909 83476
rect 3235 83516 3293 83517
rect 3235 83476 3244 83516
rect 3284 83476 3293 83516
rect 3235 83475 3293 83476
rect 3619 83516 3677 83517
rect 3619 83476 3628 83516
rect 3668 83476 3677 83516
rect 3619 83475 3677 83476
rect 4003 83516 4061 83517
rect 4003 83476 4012 83516
rect 4052 83476 4061 83516
rect 4003 83475 4061 83476
rect 4387 83516 4445 83517
rect 4387 83476 4396 83516
rect 4436 83476 4445 83516
rect 4387 83475 4445 83476
rect 4963 83516 5021 83517
rect 4963 83476 4972 83516
rect 5012 83476 5021 83516
rect 4963 83475 5021 83476
rect 5155 83516 5213 83517
rect 5155 83476 5164 83516
rect 5204 83476 5213 83516
rect 5155 83475 5213 83476
rect 5731 83516 5789 83517
rect 5731 83476 5740 83516
rect 5780 83476 5789 83516
rect 5731 83475 5789 83476
rect 6019 83516 6077 83517
rect 6019 83476 6028 83516
rect 6068 83476 6077 83516
rect 6019 83475 6077 83476
rect 6595 83516 6653 83517
rect 6595 83476 6604 83516
rect 6644 83476 6653 83516
rect 6595 83475 6653 83476
rect 6787 83516 6845 83517
rect 6787 83476 6796 83516
rect 6836 83476 6845 83516
rect 6787 83475 6845 83476
rect 7171 83516 7229 83517
rect 7171 83476 7180 83516
rect 7220 83476 7229 83516
rect 7171 83475 7229 83476
rect 7747 83516 7805 83517
rect 7747 83476 7756 83516
rect 7796 83476 7805 83516
rect 7747 83475 7805 83476
rect 8131 83516 8189 83517
rect 8131 83476 8140 83516
rect 8180 83476 8189 83516
rect 8131 83475 8189 83476
rect 8611 83516 8669 83517
rect 8611 83476 8620 83516
rect 8660 83476 8669 83516
rect 8611 83475 8669 83476
rect 8995 83516 9053 83517
rect 8995 83476 9004 83516
rect 9044 83476 9053 83516
rect 8995 83475 9053 83476
rect 9763 83516 9821 83517
rect 9763 83476 9772 83516
rect 9812 83476 9821 83516
rect 9763 83475 9821 83476
rect 10243 83516 10301 83517
rect 10243 83476 10252 83516
rect 10292 83476 10301 83516
rect 10243 83475 10301 83476
rect 10627 83516 10685 83517
rect 10627 83476 10636 83516
rect 10676 83476 10685 83516
rect 10627 83475 10685 83476
rect 11491 83516 11549 83517
rect 11491 83476 11500 83516
rect 11540 83476 11549 83516
rect 11491 83475 11549 83476
rect 13315 83516 13373 83517
rect 13315 83476 13324 83516
rect 13364 83476 13373 83516
rect 13315 83475 13373 83476
rect 13699 83516 13757 83517
rect 13699 83476 13708 83516
rect 13748 83476 13757 83516
rect 13699 83475 13757 83476
rect 14083 83516 14141 83517
rect 14083 83476 14092 83516
rect 14132 83476 14141 83516
rect 14083 83475 14141 83476
rect 14467 83516 14525 83517
rect 14467 83476 14476 83516
rect 14516 83476 14525 83516
rect 14467 83475 14525 83476
rect 14851 83516 14909 83517
rect 14851 83476 14860 83516
rect 14900 83476 14909 83516
rect 14851 83475 14909 83476
rect 15235 83516 15293 83517
rect 15235 83476 15244 83516
rect 15284 83476 15293 83516
rect 15235 83475 15293 83476
rect 15907 83516 15965 83517
rect 15907 83476 15916 83516
rect 15956 83476 15965 83516
rect 15907 83475 15965 83476
rect 16579 83516 16637 83517
rect 16579 83476 16588 83516
rect 16628 83476 16637 83516
rect 16579 83475 16637 83476
rect 17155 83516 17213 83517
rect 17155 83476 17164 83516
rect 17204 83476 17213 83516
rect 17155 83475 17213 83476
rect 17539 83516 17597 83517
rect 17539 83476 17548 83516
rect 17588 83476 17597 83516
rect 17539 83475 17597 83476
rect 17923 83516 17981 83517
rect 17923 83476 17932 83516
rect 17972 83476 17981 83516
rect 17923 83475 17981 83476
rect 18307 83516 18365 83517
rect 18307 83476 18316 83516
rect 18356 83476 18365 83516
rect 18307 83475 18365 83476
rect 18691 83516 18749 83517
rect 18691 83476 18700 83516
rect 18740 83476 18749 83516
rect 18691 83475 18749 83476
rect 19075 83516 19133 83517
rect 19075 83476 19084 83516
rect 19124 83476 19133 83516
rect 19075 83475 19133 83476
rect 19459 83516 19517 83517
rect 19459 83476 19468 83516
rect 19508 83476 19517 83516
rect 19459 83475 19517 83476
rect 19843 83516 19901 83517
rect 19843 83476 19852 83516
rect 19892 83476 19901 83516
rect 19843 83475 19901 83476
rect 20227 83516 20285 83517
rect 20227 83476 20236 83516
rect 20276 83476 20285 83516
rect 20227 83475 20285 83476
rect 4587 83432 4629 83441
rect 4587 83392 4588 83432
rect 4628 83392 4629 83432
rect 4587 83383 4629 83392
rect 7371 83432 7413 83441
rect 7371 83392 7372 83432
rect 7412 83392 7413 83432
rect 7371 83383 7413 83392
rect 4779 83348 4821 83357
rect 4779 83308 4780 83348
rect 4820 83308 4821 83348
rect 4779 83299 4821 83308
rect 7947 83348 7989 83357
rect 7947 83308 7948 83348
rect 7988 83308 7989 83348
rect 7947 83299 7989 83308
rect 13131 83348 13173 83357
rect 13131 83308 13132 83348
rect 13172 83308 13173 83348
rect 13131 83299 13173 83308
rect 13515 83348 13557 83357
rect 13515 83308 13516 83348
rect 13556 83308 13557 83348
rect 13515 83299 13557 83308
rect 13899 83348 13941 83357
rect 13899 83308 13900 83348
rect 13940 83308 13941 83348
rect 13899 83299 13941 83308
rect 14283 83348 14325 83357
rect 14283 83308 14284 83348
rect 14324 83308 14325 83348
rect 14283 83299 14325 83308
rect 14667 83348 14709 83357
rect 14667 83308 14668 83348
rect 14708 83308 14709 83348
rect 14667 83299 14709 83308
rect 15051 83348 15093 83357
rect 15051 83308 15052 83348
rect 15092 83308 15093 83348
rect 15051 83299 15093 83308
rect 16971 83348 17013 83357
rect 16971 83308 16972 83348
rect 17012 83308 17013 83348
rect 16971 83299 17013 83308
rect 18123 83348 18165 83357
rect 18123 83308 18124 83348
rect 18164 83308 18165 83348
rect 18123 83299 18165 83308
rect 18507 83348 18549 83357
rect 18507 83308 18508 83348
rect 18548 83308 18549 83348
rect 18507 83299 18549 83308
rect 19275 83348 19317 83357
rect 19275 83308 19276 83348
rect 19316 83308 19317 83348
rect 19275 83299 19317 83308
rect 1152 83180 20352 83204
rect 1152 83140 3688 83180
rect 3728 83140 3770 83180
rect 3810 83140 3852 83180
rect 3892 83140 3934 83180
rect 3974 83140 4016 83180
rect 4056 83140 18808 83180
rect 18848 83140 18890 83180
rect 18930 83140 18972 83180
rect 19012 83140 19054 83180
rect 19094 83140 19136 83180
rect 19176 83140 20352 83180
rect 1152 83116 20352 83140
rect 3627 83012 3669 83021
rect 3627 82972 3628 83012
rect 3668 82972 3669 83012
rect 3627 82963 3669 82972
rect 7467 83012 7509 83021
rect 7467 82972 7468 83012
rect 7508 82972 7509 83012
rect 7467 82963 7509 82972
rect 18219 83012 18261 83021
rect 18219 82972 18220 83012
rect 18260 82972 18261 83012
rect 18219 82963 18261 82972
rect 18603 83012 18645 83021
rect 18603 82972 18604 83012
rect 18644 82972 18645 83012
rect 18603 82963 18645 82972
rect 18987 83012 19029 83021
rect 18987 82972 18988 83012
rect 19028 82972 19029 83012
rect 18987 82963 19029 82972
rect 17451 82928 17493 82937
rect 17451 82888 17452 82928
rect 17492 82888 17493 82928
rect 17451 82879 17493 82888
rect 17835 82928 17877 82937
rect 17835 82888 17836 82928
rect 17876 82888 17877 82928
rect 17835 82879 17877 82888
rect 19371 82928 19413 82937
rect 19371 82888 19372 82928
rect 19412 82888 19413 82928
rect 19371 82879 19413 82888
rect 19755 82928 19797 82937
rect 19755 82888 19756 82928
rect 19796 82888 19797 82928
rect 19755 82879 19797 82888
rect 20139 82928 20181 82937
rect 20139 82888 20140 82928
rect 20180 82888 20181 82928
rect 20139 82879 20181 82888
rect 3811 82844 3869 82845
rect 3811 82804 3820 82844
rect 3860 82804 3869 82844
rect 3811 82803 3869 82804
rect 7267 82844 7325 82845
rect 7267 82804 7276 82844
rect 7316 82804 7325 82844
rect 7267 82803 7325 82804
rect 14371 82844 14429 82845
rect 14371 82804 14380 82844
rect 14420 82804 14429 82844
rect 14371 82803 14429 82804
rect 14755 82844 14813 82845
rect 14755 82804 14764 82844
rect 14804 82804 14813 82844
rect 14755 82803 14813 82804
rect 18019 82844 18077 82845
rect 18019 82804 18028 82844
rect 18068 82804 18077 82844
rect 18019 82803 18077 82804
rect 18403 82844 18461 82845
rect 18403 82804 18412 82844
rect 18452 82804 18461 82844
rect 18403 82803 18461 82804
rect 18787 82844 18845 82845
rect 18787 82804 18796 82844
rect 18836 82804 18845 82844
rect 18787 82803 18845 82804
rect 19171 82844 19229 82845
rect 19171 82804 19180 82844
rect 19220 82804 19229 82844
rect 19171 82803 19229 82804
rect 1891 82760 1949 82761
rect 1891 82720 1900 82760
rect 1940 82720 1949 82760
rect 1891 82719 1949 82720
rect 3139 82760 3197 82761
rect 3139 82720 3148 82760
rect 3188 82720 3197 82760
rect 3139 82719 3197 82720
rect 4099 82760 4157 82761
rect 4099 82720 4108 82760
rect 4148 82720 4157 82760
rect 4099 82719 4157 82720
rect 5347 82760 5405 82761
rect 5347 82720 5356 82760
rect 5396 82720 5405 82760
rect 5347 82719 5405 82720
rect 3339 82592 3381 82601
rect 3339 82552 3340 82592
rect 3380 82552 3381 82592
rect 3339 82543 3381 82552
rect 5547 82592 5589 82601
rect 5547 82552 5548 82592
rect 5588 82552 5589 82592
rect 5547 82543 5589 82552
rect 14187 82592 14229 82601
rect 14187 82552 14188 82592
rect 14228 82552 14229 82592
rect 14187 82543 14229 82552
rect 14571 82592 14613 82601
rect 14571 82552 14572 82592
rect 14612 82552 14613 82592
rect 14571 82543 14613 82552
rect 17347 82592 17405 82593
rect 17347 82552 17356 82592
rect 17396 82552 17405 82592
rect 17347 82551 17405 82552
rect 17731 82592 17789 82593
rect 17731 82552 17740 82592
rect 17780 82552 17789 82592
rect 17731 82551 17789 82552
rect 19651 82592 19709 82593
rect 19651 82552 19660 82592
rect 19700 82552 19709 82592
rect 19651 82551 19709 82552
rect 20035 82592 20093 82593
rect 20035 82552 20044 82592
rect 20084 82552 20093 82592
rect 20035 82551 20093 82552
rect 1152 82424 20452 82448
rect 1152 82384 4928 82424
rect 4968 82384 5010 82424
rect 5050 82384 5092 82424
rect 5132 82384 5174 82424
rect 5214 82384 5256 82424
rect 5296 82384 20048 82424
rect 20088 82384 20130 82424
rect 20170 82384 20212 82424
rect 20252 82384 20294 82424
rect 20334 82384 20376 82424
rect 20416 82384 20452 82424
rect 1152 82360 20452 82384
rect 18019 82256 18077 82257
rect 18019 82216 18028 82256
rect 18068 82216 18077 82256
rect 18019 82215 18077 82216
rect 18403 82256 18461 82257
rect 18403 82216 18412 82256
rect 18452 82216 18461 82256
rect 18403 82215 18461 82216
rect 19171 82256 19229 82257
rect 19171 82216 19180 82256
rect 19220 82216 19229 82256
rect 19171 82215 19229 82216
rect 1219 82088 1277 82089
rect 1219 82048 1228 82088
rect 1268 82048 1277 82088
rect 1219 82047 1277 82048
rect 2467 82088 2525 82089
rect 2467 82048 2476 82088
rect 2516 82048 2525 82088
rect 2467 82047 2525 82048
rect 3715 82088 3773 82089
rect 3715 82048 3724 82088
rect 3764 82048 3773 82088
rect 3715 82047 3773 82048
rect 4963 82088 5021 82089
rect 4963 82048 4972 82088
rect 5012 82048 5021 82088
rect 4963 82047 5021 82048
rect 18795 82004 18837 82013
rect 18795 81964 18796 82004
rect 18836 81964 18837 82004
rect 18795 81955 18837 81964
rect 18123 81920 18165 81929
rect 18123 81880 18124 81920
rect 18164 81880 18165 81920
rect 18123 81871 18165 81880
rect 18507 81920 18549 81929
rect 18507 81880 18508 81920
rect 18548 81880 18549 81920
rect 18507 81871 18549 81880
rect 19275 81920 19317 81929
rect 19275 81880 19276 81920
rect 19316 81880 19317 81920
rect 19275 81871 19317 81880
rect 2667 81836 2709 81845
rect 2667 81796 2668 81836
rect 2708 81796 2709 81836
rect 2667 81787 2709 81796
rect 5163 81836 5205 81845
rect 5163 81796 5164 81836
rect 5204 81796 5205 81836
rect 5163 81787 5205 81796
rect 1152 81668 20352 81692
rect 1152 81628 3688 81668
rect 3728 81628 3770 81668
rect 3810 81628 3852 81668
rect 3892 81628 3934 81668
rect 3974 81628 4016 81668
rect 4056 81628 18808 81668
rect 18848 81628 18890 81668
rect 18930 81628 18972 81668
rect 19012 81628 19054 81668
rect 19094 81628 19136 81668
rect 19176 81628 20352 81668
rect 1152 81604 20352 81628
rect 15819 81500 15861 81509
rect 15819 81460 15820 81500
rect 15860 81460 15861 81500
rect 15819 81451 15861 81460
rect 15619 81332 15677 81333
rect 15619 81292 15628 81332
rect 15668 81292 15677 81332
rect 15619 81291 15677 81292
rect 1411 81248 1469 81249
rect 1411 81208 1420 81248
rect 1460 81208 1469 81248
rect 1411 81207 1469 81208
rect 2659 81248 2717 81249
rect 2659 81208 2668 81248
rect 2708 81208 2717 81248
rect 2659 81207 2717 81208
rect 2851 81248 2909 81249
rect 2851 81208 2860 81248
rect 2900 81208 2909 81248
rect 2851 81207 2909 81208
rect 4099 81248 4157 81249
rect 4099 81208 4108 81248
rect 4148 81208 4157 81248
rect 4099 81207 4157 81208
rect 4483 81248 4541 81249
rect 4483 81208 4492 81248
rect 4532 81208 4541 81248
rect 4483 81207 4541 81208
rect 5731 81248 5789 81249
rect 5731 81208 5740 81248
rect 5780 81208 5789 81248
rect 5731 81207 5789 81208
rect 6115 81248 6173 81249
rect 6115 81208 6124 81248
rect 6164 81208 6173 81248
rect 6115 81207 6173 81208
rect 7363 81248 7421 81249
rect 7363 81208 7372 81248
rect 7412 81208 7421 81248
rect 7363 81207 7421 81208
rect 1227 81164 1269 81173
rect 1227 81124 1228 81164
rect 1268 81124 1269 81164
rect 1227 81115 1269 81124
rect 4299 81080 4341 81089
rect 4299 81040 4300 81080
rect 4340 81040 4341 81080
rect 4299 81031 4341 81040
rect 5931 81080 5973 81089
rect 5931 81040 5932 81080
rect 5972 81040 5973 81080
rect 5931 81031 5973 81040
rect 7563 81080 7605 81089
rect 7563 81040 7564 81080
rect 7604 81040 7605 81080
rect 7563 81031 7605 81040
rect 1152 80912 20452 80936
rect 1152 80872 4928 80912
rect 4968 80872 5010 80912
rect 5050 80872 5092 80912
rect 5132 80872 5174 80912
rect 5214 80872 5256 80912
rect 5296 80872 20048 80912
rect 20088 80872 20130 80912
rect 20170 80872 20212 80912
rect 20252 80872 20294 80912
rect 20334 80872 20376 80912
rect 20416 80872 20452 80912
rect 1152 80848 20452 80872
rect 7179 80660 7221 80669
rect 7179 80620 7180 80660
rect 7220 80620 7221 80660
rect 7179 80611 7221 80620
rect 1603 80576 1661 80577
rect 1603 80536 1612 80576
rect 1652 80536 1661 80576
rect 1603 80535 1661 80536
rect 2851 80576 2909 80577
rect 2851 80536 2860 80576
rect 2900 80536 2909 80576
rect 2851 80535 2909 80536
rect 3715 80576 3773 80577
rect 3715 80536 3724 80576
rect 3764 80536 3773 80576
rect 3715 80535 3773 80536
rect 4963 80576 5021 80577
rect 4963 80536 4972 80576
rect 5012 80536 5021 80576
rect 4963 80535 5021 80536
rect 5451 80576 5493 80585
rect 5451 80536 5452 80576
rect 5492 80536 5493 80576
rect 5451 80527 5493 80536
rect 5547 80576 5589 80585
rect 5547 80536 5548 80576
rect 5588 80536 5589 80576
rect 5547 80527 5589 80536
rect 6499 80576 6557 80577
rect 6499 80536 6508 80576
rect 6548 80536 6557 80576
rect 6499 80535 6557 80536
rect 6987 80571 7029 80580
rect 6987 80531 6988 80571
rect 7028 80531 7029 80571
rect 6987 80522 7029 80531
rect 5931 80492 5973 80501
rect 5931 80452 5932 80492
rect 5972 80452 5973 80492
rect 5931 80443 5973 80452
rect 6027 80492 6069 80501
rect 6027 80452 6028 80492
rect 6068 80452 6069 80492
rect 6027 80443 6069 80452
rect 3051 80324 3093 80333
rect 3051 80284 3052 80324
rect 3092 80284 3093 80324
rect 3051 80275 3093 80284
rect 5163 80324 5205 80333
rect 5163 80284 5164 80324
rect 5204 80284 5205 80324
rect 5163 80275 5205 80284
rect 1152 80156 20352 80180
rect 1152 80116 3688 80156
rect 3728 80116 3770 80156
rect 3810 80116 3852 80156
rect 3892 80116 3934 80156
rect 3974 80116 4016 80156
rect 4056 80116 18808 80156
rect 18848 80116 18890 80156
rect 18930 80116 18972 80156
rect 19012 80116 19054 80156
rect 19094 80116 19136 80156
rect 19176 80116 20352 80156
rect 1152 80092 20352 80116
rect 16011 79988 16053 79997
rect 16011 79948 16012 79988
rect 16052 79948 16053 79988
rect 16011 79939 16053 79948
rect 4107 79820 4149 79829
rect 4107 79780 4108 79820
rect 4148 79780 4149 79820
rect 4107 79771 4149 79780
rect 7275 79820 7317 79829
rect 7275 79780 7276 79820
rect 7316 79780 7317 79820
rect 7275 79771 7317 79780
rect 15811 79820 15869 79821
rect 15811 79780 15820 79820
rect 15860 79780 15869 79820
rect 15811 79779 15869 79780
rect 5211 79745 5253 79754
rect 1411 79736 1469 79737
rect 1411 79696 1420 79736
rect 1460 79696 1469 79736
rect 1411 79695 1469 79696
rect 2659 79736 2717 79737
rect 2659 79696 2668 79736
rect 2708 79696 2717 79736
rect 2659 79695 2717 79696
rect 3627 79736 3669 79745
rect 3627 79696 3628 79736
rect 3668 79696 3669 79736
rect 3627 79687 3669 79696
rect 3723 79736 3765 79745
rect 3723 79696 3724 79736
rect 3764 79696 3765 79736
rect 3723 79687 3765 79696
rect 4203 79736 4245 79745
rect 4203 79696 4204 79736
rect 4244 79696 4245 79736
rect 4203 79687 4245 79696
rect 4675 79736 4733 79737
rect 4675 79696 4684 79736
rect 4724 79696 4733 79736
rect 5211 79705 5212 79745
rect 5252 79705 5253 79745
rect 5211 79696 5253 79705
rect 5539 79736 5597 79737
rect 5539 79696 5548 79736
rect 5588 79696 5597 79736
rect 4675 79695 4733 79696
rect 5539 79695 5597 79696
rect 6787 79736 6845 79737
rect 6787 79696 6796 79736
rect 6836 79696 6845 79736
rect 6787 79695 6845 79696
rect 7179 79736 7221 79745
rect 7179 79696 7180 79736
rect 7220 79696 7221 79736
rect 7179 79687 7221 79696
rect 7371 79736 7413 79745
rect 7371 79696 7372 79736
rect 7412 79696 7413 79736
rect 7371 79687 7413 79696
rect 7939 79736 7997 79737
rect 7939 79696 7948 79736
rect 7988 79696 7997 79736
rect 7939 79695 7997 79696
rect 9187 79736 9245 79737
rect 9187 79696 9196 79736
rect 9236 79696 9245 79736
rect 9187 79695 9245 79696
rect 1227 79568 1269 79577
rect 1227 79528 1228 79568
rect 1268 79528 1269 79568
rect 1227 79519 1269 79528
rect 5355 79568 5397 79577
rect 5355 79528 5356 79568
rect 5396 79528 5397 79568
rect 5355 79519 5397 79528
rect 6987 79568 7029 79577
rect 6987 79528 6988 79568
rect 7028 79528 7029 79568
rect 6987 79519 7029 79528
rect 9387 79568 9429 79577
rect 9387 79528 9388 79568
rect 9428 79528 9429 79568
rect 9387 79519 9429 79528
rect 1152 79400 20452 79424
rect 1152 79360 4928 79400
rect 4968 79360 5010 79400
rect 5050 79360 5092 79400
rect 5132 79360 5174 79400
rect 5214 79360 5256 79400
rect 5296 79360 20048 79400
rect 20088 79360 20130 79400
rect 20170 79360 20212 79400
rect 20252 79360 20294 79400
rect 20334 79360 20376 79400
rect 20416 79360 20452 79400
rect 1152 79336 20452 79360
rect 5931 79232 5973 79241
rect 5931 79192 5932 79232
rect 5972 79192 5973 79232
rect 5931 79183 5973 79192
rect 7939 79232 7997 79233
rect 7939 79192 7948 79232
rect 7988 79192 7997 79232
rect 7939 79191 7997 79192
rect 16971 79232 17013 79241
rect 16971 79192 16972 79232
rect 17012 79192 17013 79232
rect 16971 79183 17013 79192
rect 1891 79064 1949 79065
rect 1891 79024 1900 79064
rect 1940 79024 1949 79064
rect 1891 79023 1949 79024
rect 3139 79064 3197 79065
rect 3139 79024 3148 79064
rect 3188 79024 3197 79064
rect 3139 79023 3197 79024
rect 4195 79064 4253 79065
rect 4195 79024 4204 79064
rect 4244 79024 4253 79064
rect 4195 79023 4253 79024
rect 5443 79064 5501 79065
rect 5443 79024 5452 79064
rect 5492 79024 5501 79064
rect 5443 79023 5501 79024
rect 5835 79064 5877 79073
rect 5835 79024 5836 79064
rect 5876 79024 5877 79064
rect 5835 79015 5877 79024
rect 6027 79064 6069 79073
rect 6027 79024 6028 79064
rect 6068 79024 6069 79064
rect 6027 79015 6069 79024
rect 6211 79064 6269 79065
rect 6211 79024 6220 79064
rect 6260 79024 6269 79064
rect 6211 79023 6269 79024
rect 7459 79064 7517 79065
rect 7459 79024 7468 79064
rect 7508 79024 7517 79064
rect 7459 79023 7517 79024
rect 7851 79064 7893 79073
rect 7851 79024 7852 79064
rect 7892 79024 7893 79064
rect 7851 79015 7893 79024
rect 8043 79064 8085 79073
rect 8043 79024 8044 79064
rect 8084 79024 8085 79064
rect 8043 79015 8085 79024
rect 8131 79064 8189 79065
rect 8131 79024 8140 79064
rect 8180 79024 8189 79064
rect 8131 79023 8189 79024
rect 8899 79064 8957 79065
rect 8899 79024 8908 79064
rect 8948 79024 8957 79064
rect 8899 79023 8957 79024
rect 10147 79064 10205 79065
rect 10147 79024 10156 79064
rect 10196 79024 10205 79064
rect 10147 79023 10205 79024
rect 16771 78980 16829 78981
rect 16771 78940 16780 78980
rect 16820 78940 16829 78980
rect 16771 78939 16829 78940
rect 3339 78812 3381 78821
rect 3339 78772 3340 78812
rect 3380 78772 3381 78812
rect 3339 78763 3381 78772
rect 5643 78812 5685 78821
rect 5643 78772 5644 78812
rect 5684 78772 5685 78812
rect 5643 78763 5685 78772
rect 7659 78812 7701 78821
rect 7659 78772 7660 78812
rect 7700 78772 7701 78812
rect 7659 78763 7701 78772
rect 10347 78812 10389 78821
rect 10347 78772 10348 78812
rect 10388 78772 10389 78812
rect 10347 78763 10389 78772
rect 1152 78644 20352 78668
rect 1152 78604 3688 78644
rect 3728 78604 3770 78644
rect 3810 78604 3852 78644
rect 3892 78604 3934 78644
rect 3974 78604 4016 78644
rect 4056 78604 18808 78644
rect 18848 78604 18890 78644
rect 18930 78604 18972 78644
rect 19012 78604 19054 78644
rect 19094 78604 19136 78644
rect 19176 78604 20352 78644
rect 1152 78580 20352 78604
rect 9003 78308 9045 78317
rect 9003 78268 9004 78308
rect 9044 78268 9045 78308
rect 9003 78259 9045 78268
rect 9963 78238 10005 78247
rect 1219 78224 1277 78225
rect 1219 78184 1228 78224
rect 1268 78184 1277 78224
rect 1219 78183 1277 78184
rect 2467 78224 2525 78225
rect 2467 78184 2476 78224
rect 2516 78184 2525 78224
rect 2467 78183 2525 78184
rect 3331 78224 3389 78225
rect 3331 78184 3340 78224
rect 3380 78184 3389 78224
rect 3331 78183 3389 78184
rect 4579 78224 4637 78225
rect 4579 78184 4588 78224
rect 4628 78184 4637 78224
rect 4579 78183 4637 78184
rect 5155 78224 5213 78225
rect 5155 78184 5164 78224
rect 5204 78184 5213 78224
rect 5155 78183 5213 78184
rect 6403 78224 6461 78225
rect 6403 78184 6412 78224
rect 6452 78184 6461 78224
rect 6403 78183 6461 78184
rect 6691 78224 6749 78225
rect 6691 78184 6700 78224
rect 6740 78184 6749 78224
rect 6691 78183 6749 78184
rect 7939 78224 7997 78225
rect 7939 78184 7948 78224
rect 7988 78184 7997 78224
rect 7939 78183 7997 78184
rect 8427 78224 8469 78233
rect 8427 78184 8428 78224
rect 8468 78184 8469 78224
rect 8427 78175 8469 78184
rect 8523 78224 8565 78233
rect 8523 78184 8524 78224
rect 8564 78184 8565 78224
rect 8523 78175 8565 78184
rect 8907 78224 8949 78233
rect 8907 78184 8908 78224
rect 8948 78184 8949 78224
rect 8907 78175 8949 78184
rect 9475 78224 9533 78225
rect 9475 78184 9484 78224
rect 9524 78184 9533 78224
rect 9963 78198 9964 78238
rect 10004 78198 10005 78238
rect 9963 78189 10005 78198
rect 9475 78183 9533 78184
rect 2667 78140 2709 78149
rect 2667 78100 2668 78140
rect 2708 78100 2709 78140
rect 2667 78091 2709 78100
rect 8139 78140 8181 78149
rect 8139 78100 8140 78140
rect 8180 78100 8181 78140
rect 8139 78091 8181 78100
rect 10155 78140 10197 78149
rect 10155 78100 10156 78140
rect 10196 78100 10197 78140
rect 10155 78091 10197 78100
rect 4779 78056 4821 78065
rect 4779 78016 4780 78056
rect 4820 78016 4821 78056
rect 4779 78007 4821 78016
rect 4971 78056 5013 78065
rect 4971 78016 4972 78056
rect 5012 78016 5013 78056
rect 4971 78007 5013 78016
rect 1152 77888 20452 77912
rect 1152 77848 4928 77888
rect 4968 77848 5010 77888
rect 5050 77848 5092 77888
rect 5132 77848 5174 77888
rect 5214 77848 5256 77888
rect 5296 77848 20048 77888
rect 20088 77848 20130 77888
rect 20170 77848 20212 77888
rect 20252 77848 20294 77888
rect 20334 77848 20376 77888
rect 20416 77848 20452 77888
rect 1152 77824 20452 77848
rect 4587 77636 4629 77645
rect 4587 77596 4588 77636
rect 4628 77596 4629 77636
rect 4587 77587 4629 77596
rect 9483 77636 9525 77645
rect 9483 77596 9484 77636
rect 9524 77596 9525 77636
rect 9483 77587 9525 77596
rect 2859 77552 2901 77561
rect 2859 77512 2860 77552
rect 2900 77512 2901 77552
rect 2859 77503 2901 77512
rect 2955 77552 2997 77561
rect 2955 77512 2956 77552
rect 2996 77512 2997 77552
rect 2955 77503 2997 77512
rect 3339 77552 3381 77561
rect 3339 77512 3340 77552
rect 3380 77512 3381 77552
rect 3339 77503 3381 77512
rect 3907 77552 3965 77553
rect 3907 77512 3916 77552
rect 3956 77512 3965 77552
rect 3907 77511 3965 77512
rect 4395 77547 4437 77556
rect 4395 77507 4396 77547
rect 4436 77507 4437 77547
rect 5155 77552 5213 77553
rect 5155 77512 5164 77552
rect 5204 77512 5213 77552
rect 5155 77511 5213 77512
rect 5451 77552 5493 77561
rect 5451 77512 5452 77552
rect 5492 77512 5493 77552
rect 4395 77498 4437 77507
rect 5451 77503 5493 77512
rect 5547 77552 5589 77561
rect 5547 77512 5548 77552
rect 5588 77512 5589 77552
rect 5547 77503 5589 77512
rect 6019 77552 6077 77553
rect 6019 77512 6028 77552
rect 6068 77512 6077 77552
rect 6019 77511 6077 77512
rect 7267 77552 7325 77553
rect 7267 77512 7276 77552
rect 7316 77512 7325 77552
rect 7267 77511 7325 77512
rect 7755 77552 7797 77561
rect 7755 77512 7756 77552
rect 7796 77512 7797 77552
rect 7755 77503 7797 77512
rect 7851 77552 7893 77561
rect 7851 77512 7852 77552
rect 7892 77512 7893 77552
rect 7851 77503 7893 77512
rect 8803 77552 8861 77553
rect 8803 77512 8812 77552
rect 8852 77512 8861 77552
rect 8803 77511 8861 77512
rect 9339 77542 9381 77551
rect 9339 77502 9340 77542
rect 9380 77502 9381 77542
rect 9339 77493 9381 77502
rect 3435 77468 3477 77477
rect 3435 77428 3436 77468
rect 3476 77428 3477 77468
rect 3435 77419 3477 77428
rect 8235 77468 8277 77477
rect 8235 77428 8236 77468
rect 8276 77428 8277 77468
rect 8235 77419 8277 77428
rect 8331 77468 8373 77477
rect 8331 77428 8332 77468
rect 8372 77428 8373 77468
rect 8331 77419 8373 77428
rect 5827 77384 5885 77385
rect 5827 77344 5836 77384
rect 5876 77344 5885 77384
rect 5827 77343 5885 77344
rect 7467 77300 7509 77309
rect 7467 77260 7468 77300
rect 7508 77260 7509 77300
rect 7467 77251 7509 77260
rect 1152 77132 20352 77156
rect 1152 77092 3688 77132
rect 3728 77092 3770 77132
rect 3810 77092 3852 77132
rect 3892 77092 3934 77132
rect 3974 77092 4016 77132
rect 4056 77092 18808 77132
rect 18848 77092 18890 77132
rect 18930 77092 18972 77132
rect 19012 77092 19054 77132
rect 19094 77092 19136 77132
rect 19176 77092 20352 77132
rect 1152 77068 20352 77092
rect 17163 76880 17205 76889
rect 17163 76840 17164 76880
rect 17204 76840 17205 76880
rect 17163 76831 17205 76840
rect 9003 76796 9045 76805
rect 9003 76756 9004 76796
rect 9044 76756 9045 76796
rect 9003 76747 9045 76756
rect 16963 76796 17021 76797
rect 16963 76756 16972 76796
rect 17012 76756 17021 76796
rect 16963 76755 17021 76756
rect 10011 76721 10053 76730
rect 2083 76712 2141 76713
rect 2083 76672 2092 76712
rect 2132 76672 2141 76712
rect 2083 76671 2141 76672
rect 3331 76712 3389 76713
rect 3331 76672 3340 76712
rect 3380 76672 3389 76712
rect 3331 76671 3389 76672
rect 4387 76712 4445 76713
rect 4387 76672 4396 76712
rect 4436 76672 4445 76712
rect 4387 76671 4445 76672
rect 5635 76712 5693 76713
rect 5635 76672 5644 76712
rect 5684 76672 5693 76712
rect 5635 76671 5693 76672
rect 6027 76712 6069 76721
rect 6027 76672 6028 76712
rect 6068 76672 6069 76712
rect 6027 76663 6069 76672
rect 6123 76712 6165 76721
rect 6123 76672 6124 76712
rect 6164 76672 6165 76712
rect 6123 76663 6165 76672
rect 6691 76712 6749 76713
rect 6691 76672 6700 76712
rect 6740 76672 6749 76712
rect 6691 76671 6749 76672
rect 7939 76712 7997 76713
rect 7939 76672 7948 76712
rect 7988 76672 7997 76712
rect 7939 76671 7997 76672
rect 8427 76712 8469 76721
rect 8427 76672 8428 76712
rect 8468 76672 8469 76712
rect 8427 76663 8469 76672
rect 8523 76712 8565 76721
rect 8523 76672 8524 76712
rect 8564 76672 8565 76712
rect 8523 76663 8565 76672
rect 8907 76712 8949 76721
rect 8907 76672 8908 76712
rect 8948 76672 8949 76712
rect 8907 76663 8949 76672
rect 9475 76712 9533 76713
rect 9475 76672 9484 76712
rect 9524 76672 9533 76712
rect 10011 76681 10012 76721
rect 10052 76681 10053 76721
rect 10011 76672 10053 76681
rect 10531 76712 10589 76713
rect 10531 76672 10540 76712
rect 10580 76672 10589 76712
rect 9475 76671 9533 76672
rect 10531 76671 10589 76672
rect 11779 76712 11837 76713
rect 11779 76672 11788 76712
rect 11828 76672 11837 76712
rect 11779 76671 11837 76672
rect 10347 76628 10389 76637
rect 10347 76588 10348 76628
rect 10388 76588 10389 76628
rect 10347 76579 10389 76588
rect 3531 76544 3573 76553
rect 3531 76504 3532 76544
rect 3572 76504 3573 76544
rect 3531 76495 3573 76504
rect 5835 76544 5877 76553
rect 5835 76504 5836 76544
rect 5876 76504 5877 76544
rect 5835 76495 5877 76504
rect 6307 76544 6365 76545
rect 6307 76504 6316 76544
rect 6356 76504 6365 76544
rect 6307 76503 6365 76504
rect 8139 76544 8181 76553
rect 8139 76504 8140 76544
rect 8180 76504 8181 76544
rect 8139 76495 8181 76504
rect 10155 76544 10197 76553
rect 10155 76504 10156 76544
rect 10196 76504 10197 76544
rect 10155 76495 10197 76504
rect 1152 76376 20452 76400
rect 1152 76336 4928 76376
rect 4968 76336 5010 76376
rect 5050 76336 5092 76376
rect 5132 76336 5174 76376
rect 5214 76336 5256 76376
rect 5296 76336 20048 76376
rect 20088 76336 20130 76376
rect 20170 76336 20212 76376
rect 20252 76336 20294 76376
rect 20334 76336 20376 76376
rect 20416 76336 20452 76376
rect 1152 76312 20452 76336
rect 3243 76208 3285 76217
rect 3243 76168 3244 76208
rect 3284 76168 3285 76208
rect 3243 76159 3285 76168
rect 6699 76208 6741 76217
rect 6699 76168 6700 76208
rect 6740 76168 6741 76208
rect 6699 76159 6741 76168
rect 7651 76208 7709 76209
rect 7651 76168 7660 76208
rect 7700 76168 7709 76208
rect 7651 76167 7709 76168
rect 9867 76208 9909 76217
rect 9867 76168 9868 76208
rect 9908 76168 9909 76208
rect 9867 76159 9909 76168
rect 10443 76208 10485 76217
rect 10443 76168 10444 76208
rect 10484 76168 10485 76208
rect 10443 76159 10485 76168
rect 11019 76124 11061 76133
rect 11019 76084 11020 76124
rect 11060 76084 11061 76124
rect 11019 76075 11061 76084
rect 1515 76040 1557 76049
rect 1515 76000 1516 76040
rect 1556 76000 1557 76040
rect 1515 75991 1557 76000
rect 1611 76040 1653 76049
rect 1611 76000 1612 76040
rect 1652 76000 1653 76040
rect 1611 75991 1653 76000
rect 2563 76040 2621 76041
rect 2563 76000 2572 76040
rect 2612 76000 2621 76040
rect 2563 75999 2621 76000
rect 3051 76035 3093 76044
rect 3051 75995 3052 76035
rect 3092 75995 3093 76035
rect 3051 75986 3093 75995
rect 4971 76040 5013 76049
rect 4971 76000 4972 76040
rect 5012 76000 5013 76040
rect 4971 75991 5013 76000
rect 5067 76040 5109 76049
rect 5067 76000 5068 76040
rect 5108 76000 5109 76040
rect 5067 75991 5109 76000
rect 6019 76040 6077 76041
rect 6019 76000 6028 76040
rect 6068 76000 6077 76040
rect 6019 75999 6077 76000
rect 6507 76035 6549 76044
rect 6507 75995 6508 76035
rect 6548 75995 6549 76035
rect 6507 75986 6549 75995
rect 6891 76040 6933 76049
rect 6891 76000 6892 76040
rect 6932 76000 6933 76040
rect 6891 75991 6933 76000
rect 6987 76040 7029 76049
rect 6987 76000 6988 76040
rect 7028 76000 7029 76040
rect 6987 75991 7029 76000
rect 7083 76040 7125 76049
rect 7083 76000 7084 76040
rect 7124 76000 7125 76040
rect 7083 75991 7125 76000
rect 7179 76040 7221 76049
rect 7179 76000 7180 76040
rect 7220 76000 7221 76040
rect 7179 75991 7221 76000
rect 7371 76040 7413 76049
rect 7371 76000 7372 76040
rect 7412 76000 7413 76040
rect 7371 75991 7413 76000
rect 7467 76040 7509 76049
rect 7467 76000 7468 76040
rect 7508 76000 7509 76040
rect 7467 75991 7509 76000
rect 7563 76040 7605 76049
rect 7563 76000 7564 76040
rect 7604 76000 7605 76040
rect 7563 75991 7605 76000
rect 8139 76040 8181 76049
rect 8139 76000 8140 76040
rect 8180 76000 8181 76040
rect 8139 75991 8181 76000
rect 8235 76040 8277 76049
rect 8235 76000 8236 76040
rect 8276 76000 8277 76040
rect 8235 75991 8277 76000
rect 8715 76040 8757 76049
rect 8715 76000 8716 76040
rect 8756 76000 8757 76040
rect 8715 75991 8757 76000
rect 9187 76040 9245 76041
rect 9187 76000 9196 76040
rect 9236 76000 9245 76040
rect 9187 75999 9245 76000
rect 9675 76035 9717 76044
rect 9675 75995 9676 76035
rect 9716 75995 9717 76035
rect 9675 75986 9717 75995
rect 10347 76040 10389 76049
rect 10347 76000 10348 76040
rect 10388 76000 10389 76040
rect 10347 75991 10389 76000
rect 10539 76040 10581 76049
rect 10539 76000 10540 76040
rect 10580 76000 10581 76040
rect 10539 75991 10581 76000
rect 11203 76040 11261 76041
rect 11203 76000 11212 76040
rect 11252 76000 11261 76040
rect 11203 75999 11261 76000
rect 12451 76040 12509 76041
rect 12451 76000 12460 76040
rect 12500 76000 12509 76040
rect 12451 75999 12509 76000
rect 1995 75956 2037 75965
rect 1995 75916 1996 75956
rect 2036 75916 2037 75956
rect 1995 75907 2037 75916
rect 2091 75956 2133 75965
rect 2091 75916 2092 75956
rect 2132 75916 2133 75956
rect 2091 75907 2133 75916
rect 5451 75956 5493 75965
rect 5451 75916 5452 75956
rect 5492 75916 5493 75956
rect 5451 75907 5493 75916
rect 5547 75956 5589 75965
rect 5547 75916 5548 75956
rect 5588 75916 5589 75956
rect 5547 75907 5589 75916
rect 8619 75956 8661 75965
rect 8619 75916 8620 75956
rect 8660 75916 8661 75956
rect 8619 75907 8661 75916
rect 10827 75872 10869 75881
rect 10827 75832 10828 75872
rect 10868 75832 10869 75872
rect 10827 75823 10869 75832
rect 1152 75620 20352 75644
rect 1152 75580 3688 75620
rect 3728 75580 3770 75620
rect 3810 75580 3852 75620
rect 3892 75580 3934 75620
rect 3974 75580 4016 75620
rect 4056 75580 18808 75620
rect 18848 75580 18890 75620
rect 18930 75580 18972 75620
rect 19012 75580 19054 75620
rect 19094 75580 19136 75620
rect 19176 75580 20352 75620
rect 1152 75556 20352 75580
rect 4779 75284 4821 75293
rect 4779 75244 4780 75284
rect 4820 75244 4821 75284
rect 4779 75235 4821 75244
rect 11307 75284 11349 75293
rect 11307 75244 11308 75284
rect 11348 75244 11349 75284
rect 11307 75235 11349 75244
rect 11403 75284 11445 75293
rect 11403 75244 11404 75284
rect 11444 75244 11445 75284
rect 11403 75235 11445 75244
rect 5835 75214 5877 75223
rect 1219 75200 1277 75201
rect 1219 75160 1228 75200
rect 1268 75160 1277 75200
rect 1219 75159 1277 75160
rect 2467 75200 2525 75201
rect 2467 75160 2476 75200
rect 2516 75160 2525 75200
rect 2467 75159 2525 75160
rect 4299 75200 4341 75209
rect 4299 75160 4300 75200
rect 4340 75160 4341 75200
rect 4299 75151 4341 75160
rect 4395 75200 4437 75209
rect 4395 75160 4396 75200
rect 4436 75160 4437 75200
rect 4395 75151 4437 75160
rect 4875 75200 4917 75209
rect 4875 75160 4876 75200
rect 4916 75160 4917 75200
rect 4875 75151 4917 75160
rect 5347 75200 5405 75201
rect 5347 75160 5356 75200
rect 5396 75160 5405 75200
rect 5835 75174 5836 75214
rect 5876 75174 5877 75214
rect 12411 75209 12453 75218
rect 5835 75165 5877 75174
rect 6211 75200 6269 75201
rect 5347 75159 5405 75160
rect 6211 75160 6220 75200
rect 6260 75160 6269 75200
rect 6211 75159 6269 75160
rect 7459 75200 7517 75201
rect 7459 75160 7468 75200
rect 7508 75160 7517 75200
rect 7459 75159 7517 75160
rect 9091 75200 9149 75201
rect 9091 75160 9100 75200
rect 9140 75160 9149 75200
rect 9091 75159 9149 75160
rect 10339 75200 10397 75201
rect 10339 75160 10348 75200
rect 10388 75160 10397 75200
rect 10339 75159 10397 75160
rect 10827 75200 10869 75209
rect 10827 75160 10828 75200
rect 10868 75160 10869 75200
rect 10827 75151 10869 75160
rect 10923 75200 10965 75209
rect 10923 75160 10924 75200
rect 10964 75160 10965 75200
rect 10923 75151 10965 75160
rect 11875 75200 11933 75201
rect 11875 75160 11884 75200
rect 11924 75160 11933 75200
rect 12411 75169 12412 75209
rect 12452 75169 12453 75209
rect 12411 75160 12453 75169
rect 11875 75159 11933 75160
rect 6027 75116 6069 75125
rect 6027 75076 6028 75116
rect 6068 75076 6069 75116
rect 6027 75067 6069 75076
rect 10539 75116 10581 75125
rect 10539 75076 10540 75116
rect 10580 75076 10581 75116
rect 10539 75067 10581 75076
rect 2667 75032 2709 75041
rect 2667 74992 2668 75032
rect 2708 74992 2709 75032
rect 2667 74983 2709 74992
rect 7659 75032 7701 75041
rect 7659 74992 7660 75032
rect 7700 74992 7701 75032
rect 7659 74983 7701 74992
rect 12555 75032 12597 75041
rect 12555 74992 12556 75032
rect 12596 74992 12597 75032
rect 12555 74983 12597 74992
rect 1152 74864 20452 74888
rect 1152 74824 4928 74864
rect 4968 74824 5010 74864
rect 5050 74824 5092 74864
rect 5132 74824 5174 74864
rect 5214 74824 5256 74864
rect 5296 74824 20048 74864
rect 20088 74824 20130 74864
rect 20170 74824 20212 74864
rect 20252 74824 20294 74864
rect 20334 74824 20376 74864
rect 20416 74824 20452 74864
rect 1152 74800 20452 74824
rect 8899 74738 8957 74739
rect 8899 74698 8908 74738
rect 8948 74698 8957 74738
rect 8899 74697 8957 74698
rect 7363 74696 7421 74697
rect 7363 74656 7372 74696
rect 7412 74656 7421 74696
rect 7363 74655 7421 74656
rect 9571 74696 9629 74697
rect 9571 74656 9580 74696
rect 9620 74656 9629 74696
rect 9571 74655 9629 74656
rect 12747 74696 12789 74705
rect 12747 74656 12748 74696
rect 12788 74656 12789 74696
rect 12747 74647 12789 74656
rect 9859 74612 9917 74613
rect 9859 74572 9868 74612
rect 9908 74572 9917 74612
rect 9859 74571 9917 74572
rect 1411 74528 1469 74529
rect 1411 74488 1420 74528
rect 1460 74488 1469 74528
rect 1411 74487 1469 74488
rect 2659 74528 2717 74529
rect 2659 74488 2668 74528
rect 2708 74488 2717 74528
rect 2659 74487 2717 74488
rect 2851 74528 2909 74529
rect 2851 74488 2860 74528
rect 2900 74488 2909 74528
rect 2851 74487 2909 74488
rect 4099 74528 4157 74529
rect 4099 74488 4108 74528
rect 4148 74488 4157 74528
rect 4099 74487 4157 74488
rect 5443 74528 5501 74529
rect 5443 74488 5452 74528
rect 5492 74488 5501 74528
rect 5443 74487 5501 74488
rect 5731 74528 5789 74529
rect 5731 74488 5740 74528
rect 5780 74488 5789 74528
rect 5731 74487 5789 74488
rect 6979 74528 7037 74529
rect 6979 74488 6988 74528
rect 7028 74488 7037 74528
rect 6979 74487 7037 74488
rect 7563 74528 7605 74537
rect 7563 74488 7564 74528
rect 7604 74488 7605 74528
rect 7563 74479 7605 74488
rect 7659 74528 7701 74537
rect 7659 74488 7660 74528
rect 7700 74488 7701 74528
rect 7659 74479 7701 74488
rect 8619 74528 8661 74537
rect 8619 74488 8620 74528
rect 8660 74488 8661 74528
rect 8619 74479 8661 74488
rect 8715 74528 8757 74537
rect 8715 74488 8716 74528
rect 8756 74488 8757 74528
rect 8715 74479 8757 74488
rect 9099 74528 9141 74537
rect 9099 74488 9100 74528
rect 9140 74488 9141 74528
rect 9099 74479 9141 74488
rect 9195 74528 9237 74537
rect 9195 74488 9196 74528
rect 9236 74488 9237 74528
rect 9195 74479 9237 74488
rect 9291 74528 9333 74537
rect 9291 74488 9292 74528
rect 9332 74488 9333 74528
rect 9291 74479 9333 74488
rect 9387 74528 9429 74537
rect 9387 74488 9388 74528
rect 9428 74488 9429 74528
rect 9387 74479 9429 74488
rect 9667 74528 9725 74529
rect 9667 74488 9676 74528
rect 9716 74488 9725 74528
rect 9667 74487 9725 74488
rect 10059 74528 10101 74537
rect 10059 74488 10060 74528
rect 10100 74488 10101 74528
rect 10059 74479 10101 74488
rect 10155 74528 10197 74537
rect 10155 74488 10156 74528
rect 10196 74488 10197 74528
rect 10155 74479 10197 74488
rect 10251 74528 10293 74537
rect 10251 74488 10252 74528
rect 10292 74488 10293 74528
rect 10251 74479 10293 74488
rect 10347 74528 10389 74537
rect 10347 74488 10348 74528
rect 10388 74488 10389 74528
rect 10347 74479 10389 74488
rect 11299 74528 11357 74529
rect 11299 74488 11308 74528
rect 11348 74488 11357 74528
rect 11299 74487 11357 74488
rect 12547 74528 12605 74529
rect 12547 74488 12556 74528
rect 12596 74488 12605 74528
rect 12547 74487 12605 74488
rect 5547 74360 5589 74369
rect 5547 74320 5548 74360
rect 5588 74320 5589 74360
rect 5547 74311 5589 74320
rect 10731 74360 10773 74369
rect 10731 74320 10732 74360
rect 10772 74320 10773 74360
rect 10731 74311 10773 74320
rect 1227 74276 1269 74285
rect 1227 74236 1228 74276
rect 1268 74236 1269 74276
rect 1227 74227 1269 74236
rect 4299 74276 4341 74285
rect 4299 74236 4300 74276
rect 4340 74236 4341 74276
rect 4299 74227 4341 74236
rect 7179 74276 7221 74285
rect 7179 74236 7180 74276
rect 7220 74236 7221 74276
rect 7179 74227 7221 74236
rect 1152 74108 20352 74132
rect 1152 74068 3688 74108
rect 3728 74068 3770 74108
rect 3810 74068 3852 74108
rect 3892 74068 3934 74108
rect 3974 74068 4016 74108
rect 4056 74068 18808 74108
rect 18848 74068 18890 74108
rect 18930 74068 18972 74108
rect 19012 74068 19054 74108
rect 19094 74068 19136 74108
rect 19176 74068 20352 74108
rect 1152 74044 20352 74068
rect 6795 73940 6837 73949
rect 6795 73900 6796 73940
rect 6836 73900 6837 73940
rect 6795 73891 6837 73900
rect 10827 73940 10869 73949
rect 10827 73900 10828 73940
rect 10868 73900 10869 73940
rect 10827 73891 10869 73900
rect 5259 73772 5301 73781
rect 5259 73732 5260 73772
rect 5300 73732 5301 73772
rect 5259 73723 5301 73732
rect 5355 73772 5397 73781
rect 5355 73732 5356 73772
rect 5396 73732 5397 73772
rect 5355 73723 5397 73732
rect 3339 73702 3381 73711
rect 1803 73688 1845 73697
rect 1803 73648 1804 73688
rect 1844 73648 1845 73688
rect 1803 73639 1845 73648
rect 1899 73688 1941 73697
rect 1899 73648 1900 73688
rect 1940 73648 1941 73688
rect 1899 73639 1941 73648
rect 2283 73688 2325 73697
rect 2283 73648 2284 73688
rect 2324 73648 2325 73688
rect 2283 73639 2325 73648
rect 2379 73688 2421 73697
rect 2379 73648 2380 73688
rect 2420 73648 2421 73688
rect 2379 73639 2421 73648
rect 2851 73688 2909 73689
rect 2851 73648 2860 73688
rect 2900 73648 2909 73688
rect 3339 73662 3340 73702
rect 3380 73662 3381 73702
rect 6315 73702 6357 73711
rect 3339 73653 3381 73662
rect 4779 73688 4821 73697
rect 2851 73647 2909 73648
rect 4779 73648 4780 73688
rect 4820 73648 4821 73688
rect 4779 73639 4821 73648
rect 4875 73688 4917 73697
rect 4875 73648 4876 73688
rect 4916 73648 4917 73688
rect 4875 73639 4917 73648
rect 5827 73688 5885 73689
rect 5827 73648 5836 73688
rect 5876 73648 5885 73688
rect 6315 73662 6316 73702
rect 6356 73662 6357 73702
rect 6315 73653 6357 73662
rect 6787 73688 6845 73689
rect 5827 73647 5885 73648
rect 6787 73648 6796 73688
rect 6836 73648 6845 73688
rect 6787 73647 6845 73648
rect 6883 73688 6941 73689
rect 6883 73648 6892 73688
rect 6932 73648 6941 73688
rect 6883 73647 6941 73648
rect 7083 73688 7125 73697
rect 7083 73648 7084 73688
rect 7124 73648 7125 73688
rect 7083 73639 7125 73648
rect 7179 73688 7221 73697
rect 7179 73648 7180 73688
rect 7220 73648 7221 73688
rect 7179 73639 7221 73648
rect 7272 73688 7330 73689
rect 7272 73648 7281 73688
rect 7321 73648 7330 73688
rect 7272 73647 7330 73648
rect 7755 73688 7797 73697
rect 7755 73648 7756 73688
rect 7796 73648 7797 73688
rect 7755 73639 7797 73648
rect 7851 73688 7893 73697
rect 7851 73648 7852 73688
rect 7892 73648 7893 73688
rect 7851 73639 7893 73648
rect 8227 73688 8285 73689
rect 8227 73648 8236 73688
rect 8276 73648 8285 73688
rect 8227 73647 8285 73648
rect 9475 73688 9533 73689
rect 9475 73648 9484 73688
rect 9524 73648 9533 73688
rect 9475 73647 9533 73648
rect 10059 73688 10101 73697
rect 10059 73648 10060 73688
rect 10100 73648 10101 73688
rect 10059 73639 10101 73648
rect 10155 73688 10197 73697
rect 10155 73648 10156 73688
rect 10196 73648 10197 73688
rect 10155 73639 10197 73648
rect 10251 73688 10293 73697
rect 10251 73648 10252 73688
rect 10292 73648 10293 73688
rect 10251 73639 10293 73648
rect 10347 73688 10389 73697
rect 10347 73648 10348 73688
rect 10388 73648 10389 73688
rect 10347 73639 10389 73648
rect 10531 73688 10589 73689
rect 10531 73648 10540 73688
rect 10580 73648 10589 73688
rect 10531 73647 10589 73648
rect 11011 73688 11069 73689
rect 11011 73648 11020 73688
rect 11060 73648 11069 73688
rect 11011 73647 11069 73648
rect 12259 73688 12317 73689
rect 12259 73648 12268 73688
rect 12308 73648 12317 73688
rect 12259 73647 12317 73648
rect 3531 73604 3573 73613
rect 3531 73564 3532 73604
rect 3572 73564 3573 73604
rect 3531 73555 3573 73564
rect 6507 73520 6549 73529
rect 6507 73480 6508 73520
rect 6548 73480 6549 73520
rect 6507 73471 6549 73480
rect 8035 73520 8093 73521
rect 8035 73480 8044 73520
rect 8084 73480 8093 73520
rect 8035 73479 8093 73480
rect 9675 73520 9717 73529
rect 9675 73480 9676 73520
rect 9716 73480 9717 73520
rect 9675 73471 9717 73480
rect 10635 73520 10677 73529
rect 10635 73480 10636 73520
rect 10676 73480 10677 73520
rect 10635 73471 10677 73480
rect 1152 73352 20452 73376
rect 1152 73312 4928 73352
rect 4968 73312 5010 73352
rect 5050 73312 5092 73352
rect 5132 73312 5174 73352
rect 5214 73312 5256 73352
rect 5296 73312 20048 73352
rect 20088 73312 20130 73352
rect 20170 73312 20212 73352
rect 20252 73312 20294 73352
rect 20334 73312 20376 73352
rect 20416 73312 20452 73352
rect 1152 73288 20452 73312
rect 8235 73100 8277 73109
rect 8235 73060 8236 73100
rect 8276 73060 8277 73100
rect 8235 73051 8277 73060
rect 10251 73100 10293 73109
rect 10251 73060 10252 73100
rect 10292 73060 10293 73100
rect 10251 73051 10293 73060
rect 10915 73058 10973 73059
rect 1219 73016 1277 73017
rect 1219 72976 1228 73016
rect 1268 72976 1277 73016
rect 1219 72975 1277 72976
rect 2467 73016 2525 73017
rect 2467 72976 2476 73016
rect 2516 72976 2525 73016
rect 2467 72975 2525 72976
rect 3043 73016 3101 73017
rect 3043 72976 3052 73016
rect 3092 72976 3101 73016
rect 3043 72975 3101 72976
rect 4291 73016 4349 73017
rect 4291 72976 4300 73016
rect 4340 72976 4349 73016
rect 4291 72975 4349 72976
rect 4483 73016 4541 73017
rect 4483 72976 4492 73016
rect 4532 72976 4541 73016
rect 4483 72975 4541 72976
rect 5731 73016 5789 73017
rect 5731 72976 5740 73016
rect 5780 72976 5789 73016
rect 5731 72975 5789 72976
rect 6315 73016 6357 73025
rect 6315 72976 6316 73016
rect 6356 72976 6357 73016
rect 6315 72967 6357 72976
rect 6507 73016 6549 73025
rect 6507 72976 6508 73016
rect 6548 72976 6549 73016
rect 6507 72967 6549 72976
rect 6603 73020 6645 73029
rect 6603 72980 6604 73020
rect 6644 72980 6645 73020
rect 6603 72971 6645 72980
rect 6787 73016 6845 73017
rect 6787 72976 6796 73016
rect 6836 72976 6845 73016
rect 6787 72975 6845 72976
rect 8035 73016 8093 73017
rect 8035 72976 8044 73016
rect 8084 72976 8093 73016
rect 8035 72975 8093 72976
rect 8523 73016 8565 73025
rect 8523 72976 8524 73016
rect 8564 72976 8565 73016
rect 8523 72967 8565 72976
rect 8619 73016 8661 73025
rect 8619 72976 8620 73016
rect 8660 72976 8661 73016
rect 8619 72967 8661 72976
rect 9571 73016 9629 73017
rect 9571 72976 9580 73016
rect 9620 72976 9629 73016
rect 9571 72975 9629 72976
rect 10059 73011 10101 73020
rect 10059 72971 10060 73011
rect 10100 72971 10101 73011
rect 10435 73016 10493 73017
rect 10435 72976 10444 73016
rect 10484 72976 10493 73016
rect 10435 72975 10493 72976
rect 10539 73016 10581 73025
rect 10539 72976 10540 73016
rect 10580 72976 10581 73016
rect 10059 72962 10101 72971
rect 10539 72967 10581 72976
rect 10731 73016 10773 73025
rect 10915 73018 10924 73058
rect 10964 73018 10973 73058
rect 10915 73017 10973 73018
rect 10731 72976 10732 73016
rect 10772 72976 10773 73016
rect 10731 72967 10773 72976
rect 12163 73016 12221 73017
rect 12163 72976 12172 73016
rect 12212 72976 12221 73016
rect 12163 72975 12221 72976
rect 9003 72932 9045 72941
rect 9003 72892 9004 72932
rect 9044 72892 9045 72932
rect 9003 72883 9045 72892
rect 9099 72932 9141 72941
rect 9099 72892 9100 72932
rect 9140 72892 9141 72932
rect 9099 72883 9141 72892
rect 16003 72932 16061 72933
rect 16003 72892 16012 72932
rect 16052 72892 16061 72932
rect 16003 72891 16061 72892
rect 6499 72848 6557 72849
rect 6499 72808 6508 72848
rect 6548 72808 6557 72848
rect 6499 72807 6557 72808
rect 16203 72848 16245 72857
rect 16203 72808 16204 72848
rect 16244 72808 16245 72848
rect 16203 72799 16245 72808
rect 2667 72764 2709 72773
rect 2667 72724 2668 72764
rect 2708 72724 2709 72764
rect 2667 72715 2709 72724
rect 2859 72764 2901 72773
rect 2859 72724 2860 72764
rect 2900 72724 2901 72764
rect 2859 72715 2901 72724
rect 5931 72764 5973 72773
rect 5931 72724 5932 72764
rect 5972 72724 5973 72764
rect 5931 72715 5973 72724
rect 10731 72764 10773 72773
rect 10731 72724 10732 72764
rect 10772 72724 10773 72764
rect 10731 72715 10773 72724
rect 12363 72764 12405 72773
rect 12363 72724 12364 72764
rect 12404 72724 12405 72764
rect 12363 72715 12405 72724
rect 1152 72596 20352 72620
rect 1152 72556 3688 72596
rect 3728 72556 3770 72596
rect 3810 72556 3852 72596
rect 3892 72556 3934 72596
rect 3974 72556 4016 72596
rect 4056 72556 18808 72596
rect 18848 72556 18890 72596
rect 18930 72556 18972 72596
rect 19012 72556 19054 72596
rect 19094 72556 19136 72596
rect 19176 72556 20352 72596
rect 1152 72532 20352 72556
rect 2571 72260 2613 72269
rect 2571 72220 2572 72260
rect 2612 72220 2613 72260
rect 2571 72211 2613 72220
rect 3531 72190 3573 72199
rect 1995 72176 2037 72185
rect 1995 72136 1996 72176
rect 2036 72136 2037 72176
rect 1995 72127 2037 72136
rect 2091 72176 2133 72185
rect 2091 72136 2092 72176
rect 2132 72136 2133 72176
rect 2091 72127 2133 72136
rect 2475 72176 2517 72185
rect 2475 72136 2476 72176
rect 2516 72136 2517 72176
rect 2475 72127 2517 72136
rect 3043 72176 3101 72177
rect 3043 72136 3052 72176
rect 3092 72136 3101 72176
rect 3531 72150 3532 72190
rect 3572 72150 3573 72190
rect 13467 72185 13509 72194
rect 17307 72185 17349 72194
rect 3531 72141 3573 72150
rect 4579 72176 4637 72177
rect 3043 72135 3101 72136
rect 4579 72136 4588 72176
rect 4628 72136 4637 72176
rect 4579 72135 4637 72136
rect 5827 72176 5885 72177
rect 5827 72136 5836 72176
rect 5876 72136 5885 72176
rect 5827 72135 5885 72136
rect 6219 72176 6261 72185
rect 6219 72136 6220 72176
rect 6260 72136 6261 72176
rect 6219 72127 6261 72136
rect 6315 72176 6357 72185
rect 6315 72136 6316 72176
rect 6356 72136 6357 72176
rect 6315 72127 6357 72136
rect 6411 72176 6453 72185
rect 6411 72136 6412 72176
rect 6452 72136 6453 72176
rect 6411 72127 6453 72136
rect 6787 72176 6845 72177
rect 6787 72136 6796 72176
rect 6836 72136 6845 72176
rect 6787 72135 6845 72136
rect 6979 72176 7037 72177
rect 6979 72136 6988 72176
rect 7028 72136 7037 72176
rect 6979 72135 7037 72136
rect 8227 72176 8285 72177
rect 8227 72136 8236 72176
rect 8276 72136 8285 72176
rect 8227 72135 8285 72136
rect 8619 72176 8661 72185
rect 8619 72136 8620 72176
rect 8660 72136 8661 72176
rect 8619 72127 8661 72136
rect 8811 72176 8853 72185
rect 8811 72136 8812 72176
rect 8852 72136 8853 72176
rect 8811 72127 8853 72136
rect 8907 72176 8949 72185
rect 8907 72136 8908 72176
rect 8948 72136 8949 72176
rect 8907 72127 8949 72136
rect 9099 72176 9141 72185
rect 9099 72136 9100 72176
rect 9140 72136 9141 72176
rect 9099 72127 9141 72136
rect 9195 72176 9237 72185
rect 9195 72136 9196 72176
rect 9236 72136 9237 72176
rect 9195 72127 9237 72136
rect 9291 72176 9333 72185
rect 9291 72136 9292 72176
rect 9332 72136 9333 72176
rect 9291 72127 9333 72136
rect 9387 72176 9429 72185
rect 9387 72136 9388 72176
rect 9428 72136 9429 72176
rect 9387 72127 9429 72136
rect 9579 72176 9621 72185
rect 9579 72136 9580 72176
rect 9620 72136 9621 72176
rect 9579 72127 9621 72136
rect 9771 72176 9813 72185
rect 9771 72136 9772 72176
rect 9812 72136 9813 72176
rect 9771 72127 9813 72136
rect 9867 72176 9909 72185
rect 9867 72136 9868 72176
rect 9908 72136 9909 72176
rect 9867 72127 9909 72136
rect 10059 72176 10101 72185
rect 10059 72136 10060 72176
rect 10100 72136 10101 72176
rect 10059 72127 10101 72136
rect 10347 72176 10389 72185
rect 10347 72136 10348 72176
rect 10388 72136 10389 72176
rect 10347 72127 10389 72136
rect 11883 72176 11925 72185
rect 11883 72136 11884 72176
rect 11924 72136 11925 72176
rect 11883 72127 11925 72136
rect 11979 72176 12021 72185
rect 11979 72136 11980 72176
rect 12020 72136 12021 72176
rect 11979 72127 12021 72136
rect 12363 72176 12405 72185
rect 12363 72136 12364 72176
rect 12404 72136 12405 72176
rect 12363 72127 12405 72136
rect 12459 72176 12501 72185
rect 12459 72136 12460 72176
rect 12500 72136 12501 72176
rect 12459 72127 12501 72136
rect 12931 72176 12989 72177
rect 12931 72136 12940 72176
rect 12980 72136 12989 72176
rect 13467 72145 13468 72185
rect 13508 72145 13509 72185
rect 13467 72136 13509 72145
rect 13987 72176 14045 72177
rect 13987 72136 13996 72176
rect 14036 72136 14045 72176
rect 12931 72135 12989 72136
rect 13987 72135 14045 72136
rect 15235 72176 15293 72177
rect 15235 72136 15244 72176
rect 15284 72136 15293 72176
rect 15235 72135 15293 72136
rect 15723 72176 15765 72185
rect 15723 72136 15724 72176
rect 15764 72136 15765 72176
rect 15723 72127 15765 72136
rect 15819 72176 15861 72185
rect 15819 72136 15820 72176
rect 15860 72136 15861 72176
rect 15819 72127 15861 72136
rect 16203 72176 16245 72185
rect 16203 72136 16204 72176
rect 16244 72136 16245 72176
rect 16203 72127 16245 72136
rect 16299 72176 16341 72185
rect 16299 72136 16300 72176
rect 16340 72136 16341 72176
rect 16299 72127 16341 72136
rect 16771 72176 16829 72177
rect 16771 72136 16780 72176
rect 16820 72136 16829 72176
rect 17307 72145 17308 72185
rect 17348 72145 17349 72185
rect 17307 72136 17349 72145
rect 16771 72135 16829 72136
rect 15435 72092 15477 72101
rect 15435 72052 15436 72092
rect 15476 72052 15477 72092
rect 15435 72043 15477 72052
rect 17451 72092 17493 72101
rect 17451 72052 17452 72092
rect 17492 72052 17493 72092
rect 17451 72043 17493 72052
rect 3723 72008 3765 72017
rect 3723 71968 3724 72008
rect 3764 71968 3765 72008
rect 3723 71959 3765 71968
rect 6027 72008 6069 72017
rect 6027 71968 6028 72008
rect 6068 71968 6069 72008
rect 6027 71959 6069 71968
rect 6499 72008 6557 72009
rect 6499 71968 6508 72008
rect 6548 71968 6557 72008
rect 6499 71967 6557 71968
rect 6699 72008 6741 72017
rect 6699 71968 6700 72008
rect 6740 71968 6741 72008
rect 6699 71959 6741 71968
rect 8427 72008 8469 72017
rect 8427 71968 8428 72008
rect 8468 71968 8469 72008
rect 8427 71959 8469 71968
rect 9675 72008 9717 72017
rect 9675 71968 9676 72008
rect 9716 71968 9717 72008
rect 9675 71959 9717 71968
rect 10251 72008 10293 72017
rect 10251 71968 10252 72008
rect 10292 71968 10293 72008
rect 10251 71959 10293 71968
rect 13611 72008 13653 72017
rect 13611 71968 13612 72008
rect 13652 71968 13653 72008
rect 13611 71959 13653 71968
rect 1152 71840 20452 71864
rect 1152 71800 4928 71840
rect 4968 71800 5010 71840
rect 5050 71800 5092 71840
rect 5132 71800 5174 71840
rect 5214 71800 5256 71840
rect 5296 71800 20048 71840
rect 20088 71800 20130 71840
rect 20170 71800 20212 71840
rect 20252 71800 20294 71840
rect 20334 71800 20376 71840
rect 20416 71800 20452 71840
rect 1152 71776 20452 71800
rect 5635 71672 5693 71673
rect 5635 71632 5644 71672
rect 5684 71632 5693 71672
rect 5635 71631 5693 71632
rect 9195 71672 9237 71681
rect 9195 71632 9196 71672
rect 9236 71632 9237 71672
rect 9195 71623 9237 71632
rect 13611 71672 13653 71681
rect 13611 71632 13612 71672
rect 13652 71632 13653 71672
rect 13611 71623 13653 71632
rect 17355 71672 17397 71681
rect 17355 71632 17356 71672
rect 17396 71632 17397 71672
rect 17355 71623 17397 71632
rect 15243 71588 15285 71597
rect 15243 71548 15244 71588
rect 15284 71548 15285 71588
rect 15243 71539 15285 71548
rect 1219 71504 1277 71505
rect 1219 71464 1228 71504
rect 1268 71464 1277 71504
rect 1219 71463 1277 71464
rect 2467 71504 2525 71505
rect 2467 71464 2476 71504
rect 2516 71464 2525 71504
rect 2467 71463 2525 71464
rect 2851 71504 2909 71505
rect 2851 71464 2860 71504
rect 2900 71464 2909 71504
rect 2851 71463 2909 71464
rect 4099 71504 4157 71505
rect 4099 71464 4108 71504
rect 4148 71464 4157 71504
rect 4099 71463 4157 71464
rect 5443 71504 5501 71505
rect 5443 71464 5452 71504
rect 5492 71464 5501 71504
rect 5443 71463 5501 71464
rect 5547 71504 5589 71513
rect 5547 71464 5548 71504
rect 5588 71464 5589 71504
rect 5547 71455 5589 71464
rect 5739 71504 5781 71513
rect 5739 71464 5740 71504
rect 5780 71464 5781 71504
rect 5739 71455 5781 71464
rect 5923 71504 5981 71505
rect 5923 71464 5932 71504
rect 5972 71464 5981 71504
rect 5923 71463 5981 71464
rect 7171 71504 7229 71505
rect 7171 71464 7180 71504
rect 7220 71464 7229 71504
rect 7171 71463 7229 71464
rect 7747 71504 7805 71505
rect 7747 71464 7756 71504
rect 7796 71464 7805 71504
rect 7747 71463 7805 71464
rect 8995 71504 9053 71505
rect 8995 71464 9004 71504
rect 9044 71464 9053 71504
rect 8995 71463 9053 71464
rect 9571 71504 9629 71505
rect 9571 71464 9580 71504
rect 9620 71464 9629 71504
rect 9571 71463 9629 71464
rect 10819 71504 10877 71505
rect 10819 71464 10828 71504
rect 10868 71464 10877 71504
rect 10819 71463 10877 71464
rect 12163 71504 12221 71505
rect 12163 71464 12172 71504
rect 12212 71464 12221 71504
rect 12163 71463 12221 71464
rect 13411 71504 13469 71505
rect 13411 71464 13420 71504
rect 13460 71464 13469 71504
rect 13411 71463 13469 71464
rect 13795 71504 13853 71505
rect 13795 71464 13804 71504
rect 13844 71464 13853 71504
rect 13795 71463 13853 71464
rect 15043 71504 15101 71505
rect 15043 71464 15052 71504
rect 15092 71464 15101 71504
rect 15043 71463 15101 71464
rect 15531 71504 15573 71513
rect 15531 71464 15532 71504
rect 15572 71464 15573 71504
rect 15531 71455 15573 71464
rect 15723 71504 15765 71513
rect 15723 71464 15724 71504
rect 15764 71464 15765 71504
rect 15723 71455 15765 71464
rect 15907 71504 15965 71505
rect 15907 71464 15916 71504
rect 15956 71464 15965 71504
rect 15907 71463 15965 71464
rect 17155 71504 17213 71505
rect 17155 71464 17164 71504
rect 17204 71464 17213 71504
rect 17155 71463 17213 71464
rect 17539 71504 17597 71505
rect 17539 71464 17548 71504
rect 17588 71464 17597 71504
rect 17539 71463 17597 71464
rect 18787 71504 18845 71505
rect 18787 71464 18796 71504
rect 18836 71464 18845 71504
rect 18787 71463 18845 71464
rect 19363 71504 19421 71505
rect 19363 71464 19372 71504
rect 19412 71464 19421 71504
rect 19363 71463 19421 71464
rect 7371 71336 7413 71345
rect 7371 71296 7372 71336
rect 7412 71296 7413 71336
rect 7371 71287 7413 71296
rect 9387 71336 9429 71345
rect 9387 71296 9388 71336
rect 9428 71296 9429 71336
rect 9387 71287 9429 71296
rect 2667 71252 2709 71261
rect 2667 71212 2668 71252
rect 2708 71212 2709 71252
rect 2667 71203 2709 71212
rect 4299 71252 4341 71261
rect 4299 71212 4300 71252
rect 4340 71212 4341 71252
rect 4299 71203 4341 71212
rect 15723 71252 15765 71261
rect 15723 71212 15724 71252
rect 15764 71212 15765 71252
rect 15723 71203 15765 71212
rect 18987 71252 19029 71261
rect 18987 71212 18988 71252
rect 19028 71212 19029 71252
rect 18987 71203 19029 71212
rect 19467 71252 19509 71261
rect 19467 71212 19468 71252
rect 19508 71212 19509 71252
rect 19467 71203 19509 71212
rect 1152 71084 20352 71108
rect 1152 71044 3688 71084
rect 3728 71044 3770 71084
rect 3810 71044 3852 71084
rect 3892 71044 3934 71084
rect 3974 71044 4016 71084
rect 4056 71044 18808 71084
rect 18848 71044 18890 71084
rect 18930 71044 18972 71084
rect 19012 71044 19054 71084
rect 19094 71044 19136 71084
rect 19176 71044 20352 71084
rect 1152 71020 20352 71044
rect 16395 70916 16437 70925
rect 16395 70876 16396 70916
rect 16436 70876 16437 70916
rect 16395 70867 16437 70876
rect 7467 70832 7509 70841
rect 7467 70792 7468 70832
rect 7508 70792 7509 70832
rect 7467 70783 7509 70792
rect 10347 70832 10389 70841
rect 10347 70792 10348 70832
rect 10388 70792 10389 70832
rect 10347 70783 10389 70792
rect 10539 70832 10581 70841
rect 10539 70792 10540 70832
rect 10580 70792 10581 70832
rect 10539 70783 10581 70792
rect 15051 70832 15093 70841
rect 15051 70792 15052 70832
rect 15092 70792 15093 70832
rect 15051 70783 15093 70792
rect 2955 70748 2997 70757
rect 2955 70708 2956 70748
rect 2996 70708 2997 70748
rect 2955 70699 2997 70708
rect 3051 70748 3093 70757
rect 3051 70708 3052 70748
rect 3092 70708 3093 70748
rect 3051 70699 3093 70708
rect 5643 70748 5685 70757
rect 5643 70708 5644 70748
rect 5684 70708 5685 70748
rect 5643 70699 5685 70708
rect 9627 70706 9669 70715
rect 4011 70678 4053 70687
rect 2475 70664 2517 70673
rect 2475 70624 2476 70664
rect 2516 70624 2517 70664
rect 2475 70615 2517 70624
rect 2571 70664 2613 70673
rect 2571 70624 2572 70664
rect 2612 70624 2613 70664
rect 2571 70615 2613 70624
rect 3523 70664 3581 70665
rect 3523 70624 3532 70664
rect 3572 70624 3581 70664
rect 4011 70638 4012 70678
rect 4052 70638 4053 70678
rect 6603 70678 6645 70687
rect 4011 70629 4053 70638
rect 5067 70664 5109 70673
rect 3523 70623 3581 70624
rect 5067 70624 5068 70664
rect 5108 70624 5109 70664
rect 5067 70615 5109 70624
rect 5163 70664 5205 70673
rect 5163 70624 5164 70664
rect 5204 70624 5205 70664
rect 5163 70615 5205 70624
rect 5547 70664 5589 70673
rect 5547 70624 5548 70664
rect 5588 70624 5589 70664
rect 5547 70615 5589 70624
rect 6115 70655 6173 70656
rect 6115 70615 6124 70655
rect 6164 70615 6173 70655
rect 6603 70638 6604 70678
rect 6644 70638 6645 70678
rect 9086 70677 9128 70686
rect 6603 70629 6645 70638
rect 6979 70664 7037 70665
rect 6979 70624 6988 70664
rect 7028 70624 7037 70664
rect 6979 70623 7037 70624
rect 7083 70664 7125 70673
rect 7083 70624 7084 70664
rect 7124 70624 7125 70664
rect 7083 70615 7125 70624
rect 7275 70664 7317 70673
rect 7275 70624 7276 70664
rect 7316 70624 7317 70664
rect 7275 70615 7317 70624
rect 7467 70664 7509 70673
rect 7467 70624 7468 70664
rect 7508 70624 7509 70664
rect 7467 70615 7509 70624
rect 7659 70664 7701 70673
rect 7659 70624 7660 70664
rect 7700 70624 7701 70664
rect 7659 70615 7701 70624
rect 8043 70664 8085 70673
rect 8043 70624 8044 70664
rect 8084 70624 8085 70664
rect 8043 70615 8085 70624
rect 8139 70664 8181 70673
rect 8139 70624 8140 70664
rect 8180 70624 8181 70664
rect 8139 70615 8181 70624
rect 8523 70664 8565 70673
rect 8523 70624 8524 70664
rect 8564 70624 8565 70664
rect 8523 70615 8565 70624
rect 8619 70664 8661 70673
rect 8619 70624 8620 70664
rect 8660 70624 8661 70664
rect 9086 70637 9087 70677
rect 9127 70637 9128 70677
rect 9627 70666 9628 70706
rect 9668 70666 9669 70706
rect 9627 70657 9669 70666
rect 10347 70664 10389 70673
rect 9086 70628 9128 70637
rect 8619 70615 8661 70624
rect 10347 70624 10348 70664
rect 10388 70624 10389 70664
rect 10347 70615 10389 70624
rect 10723 70664 10781 70665
rect 10723 70624 10732 70664
rect 10772 70624 10781 70664
rect 10723 70623 10781 70624
rect 11971 70664 12029 70665
rect 11971 70624 11980 70664
rect 12020 70624 12029 70664
rect 11971 70623 12029 70624
rect 13027 70664 13085 70665
rect 13027 70624 13036 70664
rect 13076 70624 13085 70664
rect 13027 70623 13085 70624
rect 14275 70664 14333 70665
rect 14275 70624 14284 70664
rect 14324 70624 14333 70664
rect 14275 70623 14333 70624
rect 14755 70664 14813 70665
rect 14755 70624 14764 70664
rect 14804 70624 14813 70664
rect 14755 70623 14813 70624
rect 14859 70664 14901 70673
rect 14859 70624 14860 70664
rect 14900 70624 14901 70664
rect 14859 70615 14901 70624
rect 15051 70664 15093 70673
rect 15051 70624 15052 70664
rect 15092 70624 15093 70664
rect 15051 70615 15093 70624
rect 15243 70664 15285 70673
rect 15243 70624 15244 70664
rect 15284 70624 15285 70664
rect 15243 70615 15285 70624
rect 15339 70664 15381 70673
rect 15339 70624 15340 70664
rect 15380 70624 15381 70664
rect 15339 70615 15381 70624
rect 15435 70664 15477 70673
rect 15435 70624 15436 70664
rect 15476 70624 15477 70664
rect 15435 70615 15477 70624
rect 15531 70664 15573 70673
rect 15531 70624 15532 70664
rect 15572 70624 15573 70664
rect 15531 70615 15573 70624
rect 15723 70664 15765 70673
rect 15723 70624 15724 70664
rect 15764 70624 15765 70664
rect 15723 70615 15765 70624
rect 15915 70664 15957 70673
rect 15915 70624 15916 70664
rect 15956 70624 15957 70664
rect 15915 70615 15957 70624
rect 16971 70664 17013 70673
rect 16971 70624 16972 70664
rect 17012 70624 17013 70664
rect 16971 70615 17013 70624
rect 17635 70664 17693 70665
rect 17635 70624 17644 70664
rect 17684 70624 17693 70664
rect 17635 70623 17693 70624
rect 18883 70664 18941 70665
rect 18883 70624 18892 70664
rect 18932 70624 18941 70664
rect 18883 70623 18941 70624
rect 19275 70664 19317 70673
rect 19275 70624 19276 70664
rect 19316 70624 19317 70664
rect 19275 70615 19317 70624
rect 19371 70664 19413 70673
rect 19371 70624 19372 70664
rect 19412 70624 19413 70664
rect 19371 70615 19413 70624
rect 19467 70664 19509 70673
rect 19467 70624 19468 70664
rect 19508 70624 19509 70664
rect 19467 70615 19509 70624
rect 19843 70664 19901 70665
rect 19843 70624 19852 70664
rect 19892 70624 19901 70664
rect 19843 70623 19901 70624
rect 6115 70614 6173 70615
rect 4203 70580 4245 70589
rect 4203 70540 4204 70580
rect 4244 70540 4245 70580
rect 4203 70531 4245 70540
rect 6795 70580 6837 70589
rect 6795 70540 6796 70580
rect 6836 70540 6837 70580
rect 6795 70531 6837 70540
rect 7179 70580 7221 70589
rect 7179 70540 7180 70580
rect 7220 70540 7221 70580
rect 7179 70531 7221 70540
rect 9771 70580 9813 70589
rect 9771 70540 9772 70580
rect 9812 70540 9813 70580
rect 9771 70531 9813 70540
rect 15819 70580 15861 70589
rect 15819 70540 15820 70580
rect 15860 70540 15861 70580
rect 15819 70531 15861 70540
rect 20035 70580 20093 70581
rect 20035 70540 20044 70580
rect 20084 70540 20093 70580
rect 20035 70539 20093 70540
rect 12171 70496 12213 70505
rect 12171 70456 12172 70496
rect 12212 70456 12213 70496
rect 12171 70447 12213 70456
rect 14475 70496 14517 70505
rect 14475 70456 14476 70496
rect 14516 70456 14517 70496
rect 14475 70447 14517 70456
rect 19083 70496 19125 70505
rect 19083 70456 19084 70496
rect 19124 70456 19125 70496
rect 19083 70447 19125 70456
rect 19555 70496 19613 70497
rect 19555 70456 19564 70496
rect 19604 70456 19613 70496
rect 19555 70455 19613 70456
rect 19747 70496 19805 70497
rect 19747 70456 19756 70496
rect 19796 70456 19805 70496
rect 19747 70455 19805 70456
rect 1152 70328 20452 70352
rect 1152 70288 4928 70328
rect 4968 70288 5010 70328
rect 5050 70288 5092 70328
rect 5132 70288 5174 70328
rect 5214 70288 5256 70328
rect 5296 70288 20048 70328
rect 20088 70288 20130 70328
rect 20170 70288 20212 70328
rect 20252 70288 20294 70328
rect 20334 70288 20376 70328
rect 20416 70288 20452 70328
rect 1152 70264 20452 70288
rect 16203 70160 16245 70169
rect 16203 70120 16204 70160
rect 16244 70120 16245 70160
rect 16203 70111 16245 70120
rect 16387 70160 16445 70161
rect 16387 70120 16396 70160
rect 16436 70120 16445 70160
rect 16387 70119 16445 70120
rect 16867 70160 16925 70161
rect 16867 70120 16876 70160
rect 16916 70120 16925 70160
rect 16867 70119 16925 70120
rect 13323 70076 13365 70085
rect 13323 70036 13324 70076
rect 13364 70036 13365 70076
rect 13323 70027 13365 70036
rect 19371 70076 19413 70085
rect 19371 70036 19372 70076
rect 19412 70036 19413 70076
rect 19371 70027 19413 70036
rect 1219 69992 1277 69993
rect 1219 69952 1228 69992
rect 1268 69952 1277 69992
rect 1219 69951 1277 69952
rect 2467 69992 2525 69993
rect 2467 69952 2476 69992
rect 2516 69952 2525 69992
rect 2467 69951 2525 69952
rect 3043 69992 3101 69993
rect 3043 69952 3052 69992
rect 3092 69952 3101 69992
rect 3043 69951 3101 69952
rect 4291 69992 4349 69993
rect 4291 69952 4300 69992
rect 4340 69952 4349 69992
rect 4291 69951 4349 69952
rect 4675 69992 4733 69993
rect 4675 69952 4684 69992
rect 4724 69952 4733 69992
rect 4675 69951 4733 69952
rect 5923 69992 5981 69993
rect 5923 69952 5932 69992
rect 5972 69952 5981 69992
rect 5923 69951 5981 69952
rect 6123 69992 6165 70001
rect 6123 69952 6124 69992
rect 6164 69952 6165 69992
rect 6123 69943 6165 69952
rect 6219 69992 6261 70001
rect 6219 69952 6220 69992
rect 6260 69952 6261 69992
rect 6219 69943 6261 69952
rect 6315 69992 6357 70001
rect 6315 69952 6316 69992
rect 6356 69952 6357 69992
rect 6315 69943 6357 69952
rect 6411 69992 6453 70001
rect 6411 69952 6412 69992
rect 6452 69952 6453 69992
rect 6411 69943 6453 69952
rect 6795 69992 6837 70001
rect 6795 69952 6796 69992
rect 6836 69952 6837 69992
rect 6795 69943 6837 69952
rect 6987 69992 7029 70001
rect 6987 69952 6988 69992
rect 7028 69952 7029 69992
rect 6987 69943 7029 69952
rect 8227 69992 8285 69993
rect 8227 69952 8236 69992
rect 8276 69952 8285 69992
rect 8227 69951 8285 69952
rect 9475 69992 9533 69993
rect 9475 69952 9484 69992
rect 9524 69952 9533 69992
rect 9475 69951 9533 69952
rect 9859 69992 9917 69993
rect 9859 69952 9868 69992
rect 9908 69952 9917 69992
rect 9859 69951 9917 69952
rect 11107 69992 11165 69993
rect 11107 69952 11116 69992
rect 11156 69952 11165 69992
rect 11107 69951 11165 69952
rect 11595 69992 11637 70001
rect 11595 69952 11596 69992
rect 11636 69952 11637 69992
rect 11595 69943 11637 69952
rect 11691 69992 11733 70001
rect 11691 69952 11692 69992
rect 11732 69952 11733 69992
rect 11691 69943 11733 69952
rect 12643 69992 12701 69993
rect 12643 69952 12652 69992
rect 12692 69952 12701 69992
rect 14475 69992 14517 70001
rect 12643 69951 12701 69952
rect 13179 69982 13221 69991
rect 13179 69942 13180 69982
rect 13220 69942 13221 69982
rect 14475 69952 14476 69992
rect 14516 69952 14517 69992
rect 14475 69943 14517 69952
rect 14571 69992 14613 70001
rect 14571 69952 14572 69992
rect 14612 69952 14613 69992
rect 14571 69943 14613 69952
rect 15523 69992 15581 69993
rect 15523 69952 15532 69992
rect 15572 69952 15581 69992
rect 16491 69992 16533 70001
rect 15523 69951 15581 69952
rect 16011 69978 16053 69987
rect 13179 69933 13221 69942
rect 16011 69938 16012 69978
rect 16052 69938 16053 69978
rect 16491 69952 16492 69992
rect 16532 69952 16533 69992
rect 16491 69943 16533 69952
rect 16587 69992 16629 70001
rect 16587 69952 16588 69992
rect 16628 69952 16629 69992
rect 16587 69943 16629 69952
rect 16683 69992 16725 70001
rect 16683 69952 16684 69992
rect 16724 69952 16725 69992
rect 16683 69943 16725 69952
rect 17067 69992 17109 70001
rect 17067 69952 17068 69992
rect 17108 69952 17109 69992
rect 17067 69943 17109 69952
rect 17163 69992 17205 70001
rect 17163 69952 17164 69992
rect 17204 69952 17205 69992
rect 17163 69943 17205 69952
rect 17643 69992 17685 70001
rect 17643 69952 17644 69992
rect 17684 69952 17685 69992
rect 17643 69943 17685 69952
rect 17739 69992 17781 70001
rect 17739 69952 17740 69992
rect 17780 69952 17781 69992
rect 17739 69943 17781 69952
rect 18123 69992 18165 70001
rect 18123 69952 18124 69992
rect 18164 69952 18165 69992
rect 18123 69943 18165 69952
rect 18691 69992 18749 69993
rect 18691 69952 18700 69992
rect 18740 69952 18749 69992
rect 18691 69951 18749 69952
rect 19179 69987 19221 69996
rect 19179 69947 19180 69987
rect 19220 69947 19221 69987
rect 19555 69992 19613 69993
rect 19555 69952 19564 69992
rect 19604 69952 19613 69992
rect 19555 69951 19613 69952
rect 19659 69992 19701 70001
rect 19659 69952 19660 69992
rect 19700 69952 19701 69992
rect 19179 69938 19221 69947
rect 19659 69943 19701 69952
rect 19851 69992 19893 70001
rect 19851 69952 19852 69992
rect 19892 69952 19893 69992
rect 19851 69943 19893 69952
rect 20043 69992 20085 70001
rect 20043 69952 20044 69992
rect 20084 69952 20085 69992
rect 20043 69943 20085 69952
rect 20235 69992 20277 70001
rect 20235 69952 20236 69992
rect 20276 69952 20277 69992
rect 20235 69943 20277 69952
rect 16011 69929 16053 69938
rect 6891 69908 6933 69917
rect 6891 69868 6892 69908
rect 6932 69868 6933 69908
rect 6891 69859 6933 69868
rect 12075 69908 12117 69917
rect 12075 69868 12076 69908
rect 12116 69868 12117 69908
rect 12075 69859 12117 69868
rect 12171 69908 12213 69917
rect 12171 69868 12172 69908
rect 12212 69868 12213 69908
rect 12171 69859 12213 69868
rect 14955 69908 14997 69917
rect 14955 69868 14956 69908
rect 14996 69868 14997 69908
rect 14955 69859 14997 69868
rect 15051 69908 15093 69917
rect 15051 69868 15052 69908
rect 15092 69868 15093 69908
rect 15051 69859 15093 69868
rect 18219 69908 18261 69917
rect 18219 69868 18220 69908
rect 18260 69868 18261 69908
rect 18219 69859 18261 69868
rect 20043 69824 20085 69833
rect 20043 69784 20044 69824
rect 20084 69784 20085 69824
rect 20043 69775 20085 69784
rect 2667 69740 2709 69749
rect 2667 69700 2668 69740
rect 2708 69700 2709 69740
rect 2667 69691 2709 69700
rect 2859 69740 2901 69749
rect 2859 69700 2860 69740
rect 2900 69700 2901 69740
rect 2859 69691 2901 69700
rect 4491 69740 4533 69749
rect 4491 69700 4492 69740
rect 4532 69700 4533 69740
rect 4491 69691 4533 69700
rect 9675 69740 9717 69749
rect 9675 69700 9676 69740
rect 9716 69700 9717 69740
rect 9675 69691 9717 69700
rect 11307 69740 11349 69749
rect 11307 69700 11308 69740
rect 11348 69700 11349 69740
rect 11307 69691 11349 69700
rect 19851 69740 19893 69749
rect 19851 69700 19852 69740
rect 19892 69700 19893 69740
rect 19851 69691 19893 69700
rect 1152 69572 20352 69596
rect 1152 69532 3688 69572
rect 3728 69532 3770 69572
rect 3810 69532 3852 69572
rect 3892 69532 3934 69572
rect 3974 69532 4016 69572
rect 4056 69532 18808 69572
rect 18848 69532 18890 69572
rect 18930 69532 18972 69572
rect 19012 69532 19054 69572
rect 19094 69532 19136 69572
rect 19176 69532 20352 69572
rect 1152 69508 20352 69532
rect 13419 69404 13461 69413
rect 13419 69364 13420 69404
rect 13460 69364 13461 69404
rect 13419 69355 13461 69364
rect 15147 69404 15189 69413
rect 15147 69364 15148 69404
rect 15188 69364 15189 69404
rect 15147 69355 15189 69364
rect 17835 69404 17877 69413
rect 17835 69364 17836 69404
rect 17876 69364 17877 69404
rect 17835 69355 17877 69364
rect 5451 69320 5493 69329
rect 5451 69280 5452 69320
rect 5492 69280 5493 69320
rect 5451 69271 5493 69280
rect 15331 69320 15389 69321
rect 15331 69280 15340 69320
rect 15380 69280 15389 69320
rect 15331 69279 15389 69280
rect 2475 69236 2517 69245
rect 2475 69196 2476 69236
rect 2516 69196 2517 69236
rect 2475 69187 2517 69196
rect 10443 69236 10485 69245
rect 10443 69196 10444 69236
rect 10484 69196 10485 69236
rect 10443 69187 10485 69196
rect 3435 69166 3477 69175
rect 1899 69152 1941 69161
rect 1899 69112 1900 69152
rect 1940 69112 1941 69152
rect 1899 69103 1941 69112
rect 1995 69152 2037 69161
rect 1995 69112 1996 69152
rect 2036 69112 2037 69152
rect 1995 69103 2037 69112
rect 2379 69152 2421 69161
rect 2379 69112 2380 69152
rect 2420 69112 2421 69152
rect 2379 69103 2421 69112
rect 2947 69152 3005 69153
rect 2947 69112 2956 69152
rect 2996 69112 3005 69152
rect 3435 69126 3436 69166
rect 3476 69126 3477 69166
rect 3435 69117 3477 69126
rect 4003 69152 4061 69153
rect 2947 69111 3005 69112
rect 4003 69112 4012 69152
rect 4052 69112 4061 69152
rect 4003 69111 4061 69112
rect 5251 69152 5309 69153
rect 5251 69112 5260 69152
rect 5300 69112 5309 69152
rect 5251 69111 5309 69112
rect 5635 69152 5693 69153
rect 5635 69112 5644 69152
rect 5684 69112 5693 69152
rect 5635 69111 5693 69112
rect 6883 69152 6941 69153
rect 6883 69112 6892 69152
rect 6932 69112 6941 69152
rect 6883 69111 6941 69112
rect 7075 69152 7133 69153
rect 7075 69112 7084 69152
rect 7124 69112 7133 69152
rect 7075 69111 7133 69112
rect 7179 69152 7221 69161
rect 7179 69112 7180 69152
rect 7220 69112 7221 69152
rect 7179 69103 7221 69112
rect 7371 69152 7413 69161
rect 7371 69112 7372 69152
rect 7412 69112 7413 69152
rect 7371 69103 7413 69112
rect 8227 69152 8285 69153
rect 8227 69112 8236 69152
rect 8276 69112 8285 69152
rect 8227 69111 8285 69112
rect 9475 69152 9533 69153
rect 9475 69112 9484 69152
rect 9524 69112 9533 69152
rect 9475 69111 9533 69112
rect 9963 69152 10005 69161
rect 9963 69112 9964 69152
rect 10004 69112 10005 69152
rect 9963 69103 10005 69112
rect 10059 69152 10101 69161
rect 10059 69112 10060 69152
rect 10100 69112 10101 69152
rect 10059 69103 10101 69112
rect 10539 69152 10581 69161
rect 11499 69157 11541 69166
rect 10539 69112 10540 69152
rect 10580 69112 10581 69152
rect 10539 69103 10581 69112
rect 11011 69152 11069 69153
rect 11011 69112 11020 69152
rect 11060 69112 11069 69152
rect 11011 69111 11069 69112
rect 11499 69117 11500 69157
rect 11540 69117 11541 69157
rect 11499 69108 11541 69117
rect 11971 69152 12029 69153
rect 11971 69112 11980 69152
rect 12020 69112 12029 69152
rect 11971 69111 12029 69112
rect 13219 69152 13277 69153
rect 13219 69112 13228 69152
rect 13268 69112 13277 69152
rect 13219 69111 13277 69112
rect 13699 69152 13757 69153
rect 13699 69112 13708 69152
rect 13748 69112 13757 69152
rect 13699 69111 13757 69112
rect 14947 69152 15005 69153
rect 14947 69112 14956 69152
rect 14996 69112 15005 69152
rect 14947 69111 15005 69112
rect 15723 69152 15765 69161
rect 15723 69112 15724 69152
rect 15764 69112 15765 69152
rect 15723 69103 15765 69112
rect 16003 69152 16061 69153
rect 16003 69112 16012 69152
rect 16052 69112 16061 69152
rect 16003 69111 16061 69112
rect 16387 69152 16445 69153
rect 16387 69112 16396 69152
rect 16436 69112 16445 69152
rect 16387 69111 16445 69112
rect 17635 69152 17693 69153
rect 17635 69112 17644 69152
rect 17684 69112 17693 69152
rect 17635 69111 17693 69112
rect 18219 69152 18261 69161
rect 18219 69112 18220 69152
rect 18260 69112 18261 69152
rect 18411 69152 18453 69161
rect 18219 69103 18261 69112
rect 18315 69131 18357 69140
rect 18315 69091 18316 69131
rect 18356 69091 18357 69131
rect 18411 69112 18412 69152
rect 18452 69112 18453 69152
rect 18411 69103 18453 69112
rect 18699 69152 18741 69161
rect 18699 69112 18700 69152
rect 18740 69112 18741 69152
rect 18699 69103 18741 69112
rect 18795 69152 18837 69161
rect 18795 69112 18796 69152
rect 18836 69112 18837 69152
rect 18795 69103 18837 69112
rect 18891 69152 18933 69161
rect 18891 69112 18892 69152
rect 18932 69112 18933 69152
rect 18891 69103 18933 69112
rect 18987 69152 19029 69161
rect 18987 69112 18988 69152
rect 19028 69112 19029 69152
rect 18987 69103 19029 69112
rect 19179 69152 19221 69161
rect 19179 69112 19180 69152
rect 19220 69112 19221 69152
rect 19179 69103 19221 69112
rect 19275 69152 19317 69161
rect 19275 69112 19276 69152
rect 19316 69112 19317 69152
rect 19275 69103 19317 69112
rect 19659 69152 19701 69161
rect 19659 69112 19660 69152
rect 19700 69112 19701 69152
rect 19659 69103 19701 69112
rect 19755 69152 19797 69161
rect 19755 69112 19756 69152
rect 19796 69112 19797 69152
rect 19755 69103 19797 69112
rect 18315 69082 18357 69091
rect 3627 69068 3669 69077
rect 3627 69028 3628 69068
rect 3668 69028 3669 69068
rect 3627 69019 3669 69028
rect 15627 69068 15669 69077
rect 15627 69028 15628 69068
rect 15668 69028 15669 69068
rect 15627 69019 15669 69028
rect 3819 68984 3861 68993
rect 3819 68944 3820 68984
rect 3860 68944 3861 68984
rect 3819 68935 3861 68944
rect 7267 68984 7325 68985
rect 7267 68944 7276 68984
rect 7316 68944 7325 68984
rect 7267 68943 7325 68944
rect 9675 68984 9717 68993
rect 9675 68944 9676 68984
rect 9716 68944 9717 68984
rect 9675 68935 9717 68944
rect 11691 68984 11733 68993
rect 11691 68944 11692 68984
rect 11732 68944 11733 68984
rect 11691 68935 11733 68944
rect 18499 68984 18557 68985
rect 18499 68944 18508 68984
rect 18548 68944 18557 68984
rect 18499 68943 18557 68944
rect 19459 68984 19517 68985
rect 19459 68944 19468 68984
rect 19508 68944 19517 68984
rect 19459 68943 19517 68944
rect 19939 68984 19997 68985
rect 19939 68944 19948 68984
rect 19988 68944 19997 68984
rect 19939 68943 19997 68944
rect 1152 68816 20452 68840
rect 1152 68776 4928 68816
rect 4968 68776 5010 68816
rect 5050 68776 5092 68816
rect 5132 68776 5174 68816
rect 5214 68776 5256 68816
rect 5296 68776 20048 68816
rect 20088 68776 20130 68816
rect 20170 68776 20212 68816
rect 20252 68776 20294 68816
rect 20334 68776 20376 68816
rect 20416 68776 20452 68816
rect 1152 68752 20452 68776
rect 6411 68648 6453 68657
rect 6411 68608 6412 68648
rect 6452 68608 6453 68648
rect 6411 68599 6453 68608
rect 10347 68648 10389 68657
rect 10347 68608 10348 68648
rect 10388 68608 10389 68648
rect 10347 68599 10389 68608
rect 8331 68564 8373 68573
rect 8331 68524 8332 68564
rect 8372 68524 8373 68564
rect 8331 68515 8373 68524
rect 6590 68491 6632 68500
rect 2371 68480 2429 68481
rect 2371 68440 2380 68480
rect 2420 68440 2429 68480
rect 2371 68439 2429 68440
rect 3619 68480 3677 68481
rect 3619 68440 3628 68480
rect 3668 68440 3677 68480
rect 3619 68439 3677 68440
rect 4099 68480 4157 68481
rect 4099 68440 4108 68480
rect 4148 68440 4157 68480
rect 4099 68439 4157 68440
rect 4203 68480 4245 68489
rect 4203 68440 4204 68480
rect 4244 68440 4245 68480
rect 4203 68431 4245 68440
rect 4395 68480 4437 68489
rect 4395 68440 4396 68480
rect 4436 68440 4437 68480
rect 4395 68431 4437 68440
rect 4683 68480 4725 68489
rect 4683 68440 4684 68480
rect 4724 68440 4725 68480
rect 4683 68431 4725 68440
rect 4779 68480 4821 68489
rect 4779 68440 4780 68480
rect 4820 68440 4821 68480
rect 4779 68431 4821 68440
rect 5163 68480 5205 68489
rect 5163 68440 5164 68480
rect 5204 68440 5205 68480
rect 5163 68431 5205 68440
rect 5731 68480 5789 68481
rect 5731 68440 5740 68480
rect 5780 68440 5789 68480
rect 5731 68439 5789 68440
rect 6219 68475 6261 68484
rect 6219 68435 6220 68475
rect 6260 68435 6261 68475
rect 6590 68451 6591 68491
rect 6631 68451 6632 68491
rect 6590 68442 6632 68451
rect 6883 68480 6941 68481
rect 6883 68440 6892 68480
rect 6932 68440 6941 68480
rect 6883 68439 6941 68440
rect 8131 68480 8189 68481
rect 8131 68440 8140 68480
rect 8180 68440 8189 68480
rect 8131 68439 8189 68440
rect 8619 68480 8661 68489
rect 8619 68440 8620 68480
rect 8660 68440 8661 68480
rect 6219 68426 6261 68435
rect 8619 68431 8661 68440
rect 8715 68480 8757 68489
rect 8715 68440 8716 68480
rect 8756 68440 8757 68480
rect 8715 68431 8757 68440
rect 9195 68480 9237 68489
rect 9195 68440 9196 68480
rect 9236 68440 9237 68480
rect 9195 68431 9237 68440
rect 9667 68480 9725 68481
rect 9667 68440 9676 68480
rect 9716 68440 9725 68480
rect 9667 68439 9725 68440
rect 10155 68475 10197 68484
rect 10155 68435 10156 68475
rect 10196 68435 10197 68475
rect 11491 68480 11549 68481
rect 11491 68440 11500 68480
rect 11540 68440 11549 68480
rect 11491 68439 11549 68440
rect 12739 68480 12797 68481
rect 12739 68440 12748 68480
rect 12788 68440 12797 68480
rect 12739 68439 12797 68440
rect 13699 68480 13757 68481
rect 13699 68440 13708 68480
rect 13748 68440 13757 68480
rect 13699 68439 13757 68440
rect 14947 68480 15005 68481
rect 14947 68440 14956 68480
rect 14996 68440 15005 68480
rect 14947 68439 15005 68440
rect 15331 68480 15389 68481
rect 15331 68440 15340 68480
rect 15380 68440 15389 68480
rect 15331 68439 15389 68440
rect 16579 68480 16637 68481
rect 16579 68440 16588 68480
rect 16628 68440 16637 68480
rect 16579 68439 16637 68440
rect 16963 68480 17021 68481
rect 16963 68440 16972 68480
rect 17012 68440 17021 68480
rect 16963 68439 17021 68440
rect 18211 68480 18269 68481
rect 18211 68440 18220 68480
rect 18260 68440 18269 68480
rect 18211 68439 18269 68440
rect 18603 68480 18645 68489
rect 18603 68440 18604 68480
rect 18644 68440 18645 68480
rect 10155 68426 10197 68435
rect 18603 68431 18645 68440
rect 18699 68480 18741 68489
rect 18699 68440 18700 68480
rect 18740 68440 18741 68480
rect 18699 68431 18741 68440
rect 18891 68480 18933 68489
rect 18891 68440 18892 68480
rect 18932 68440 18933 68480
rect 18891 68431 18933 68440
rect 19083 68480 19125 68489
rect 19083 68440 19084 68480
rect 19124 68440 19125 68480
rect 19083 68431 19125 68440
rect 19275 68480 19317 68489
rect 19275 68440 19276 68480
rect 19316 68440 19317 68480
rect 19275 68431 19317 68440
rect 19371 68480 19413 68489
rect 19371 68440 19372 68480
rect 19412 68440 19413 68480
rect 19371 68431 19413 68440
rect 5259 68396 5301 68405
rect 5259 68356 5260 68396
rect 5300 68356 5301 68396
rect 5259 68347 5301 68356
rect 9099 68396 9141 68405
rect 9099 68356 9100 68396
rect 9140 68356 9141 68396
rect 9099 68347 9141 68356
rect 19363 68312 19421 68313
rect 19363 68272 19372 68312
rect 19412 68272 19421 68312
rect 19363 68271 19421 68272
rect 3819 68228 3861 68237
rect 3819 68188 3820 68228
rect 3860 68188 3861 68228
rect 3819 68179 3861 68188
rect 4395 68228 4437 68237
rect 4395 68188 4396 68228
rect 4436 68188 4437 68228
rect 4395 68179 4437 68188
rect 6699 68228 6741 68237
rect 6699 68188 6700 68228
rect 6740 68188 6741 68228
rect 6699 68179 6741 68188
rect 12939 68228 12981 68237
rect 12939 68188 12940 68228
rect 12980 68188 12981 68228
rect 12939 68179 12981 68188
rect 15147 68228 15189 68237
rect 15147 68188 15148 68228
rect 15188 68188 15189 68228
rect 15147 68179 15189 68188
rect 16779 68228 16821 68237
rect 16779 68188 16780 68228
rect 16820 68188 16821 68228
rect 16779 68179 16821 68188
rect 18411 68228 18453 68237
rect 18411 68188 18412 68228
rect 18452 68188 18453 68228
rect 18411 68179 18453 68188
rect 1152 68060 20352 68084
rect 1152 68020 3688 68060
rect 3728 68020 3770 68060
rect 3810 68020 3852 68060
rect 3892 68020 3934 68060
rect 3974 68020 4016 68060
rect 4056 68020 18808 68060
rect 18848 68020 18890 68060
rect 18930 68020 18972 68060
rect 19012 68020 19054 68060
rect 19094 68020 19136 68060
rect 19176 68020 20352 68060
rect 1152 67996 20352 68020
rect 7371 67892 7413 67901
rect 7371 67852 7372 67892
rect 7412 67852 7413 67892
rect 7371 67843 7413 67852
rect 2859 67724 2901 67733
rect 2859 67684 2860 67724
rect 2900 67684 2901 67724
rect 2859 67675 2901 67684
rect 10155 67724 10197 67733
rect 10155 67684 10156 67724
rect 10196 67684 10197 67724
rect 10155 67675 10197 67684
rect 14187 67724 14229 67733
rect 14187 67684 14188 67724
rect 14228 67684 14229 67724
rect 14187 67675 14229 67684
rect 15339 67724 15381 67733
rect 15339 67684 15340 67724
rect 15380 67684 15381 67724
rect 15339 67675 15381 67684
rect 15435 67724 15477 67733
rect 15435 67684 15436 67724
rect 15476 67684 15477 67724
rect 15435 67675 15477 67684
rect 18027 67724 18069 67733
rect 18027 67684 18028 67724
rect 18068 67684 18069 67724
rect 18027 67675 18069 67684
rect 3963 67649 4005 67658
rect 2379 67640 2421 67649
rect 2379 67600 2380 67640
rect 2420 67600 2421 67640
rect 2379 67591 2421 67600
rect 2475 67640 2517 67649
rect 2475 67600 2476 67640
rect 2516 67600 2517 67640
rect 2475 67591 2517 67600
rect 2955 67640 2997 67649
rect 2955 67600 2956 67640
rect 2996 67600 2997 67640
rect 2955 67591 2997 67600
rect 3427 67640 3485 67641
rect 3427 67600 3436 67640
rect 3476 67600 3485 67640
rect 3963 67609 3964 67649
rect 4004 67609 4005 67649
rect 3963 67600 4005 67609
rect 4483 67640 4541 67641
rect 4483 67600 4492 67640
rect 4532 67600 4541 67640
rect 3427 67599 3485 67600
rect 4483 67599 4541 67600
rect 5731 67640 5789 67641
rect 5731 67600 5740 67640
rect 5780 67600 5789 67640
rect 5731 67599 5789 67600
rect 5923 67640 5981 67641
rect 5923 67600 5932 67640
rect 5972 67600 5981 67640
rect 5923 67599 5981 67600
rect 7171 67640 7229 67641
rect 7171 67600 7180 67640
rect 7220 67600 7229 67640
rect 7171 67599 7229 67600
rect 7843 67640 7901 67641
rect 7843 67600 7852 67640
rect 7892 67600 7901 67640
rect 7843 67599 7901 67600
rect 9091 67640 9149 67641
rect 9091 67600 9100 67640
rect 9140 67600 9149 67640
rect 9091 67599 9149 67600
rect 9579 67640 9621 67649
rect 9579 67600 9580 67640
rect 9620 67600 9621 67640
rect 9579 67591 9621 67600
rect 9675 67640 9717 67649
rect 9675 67600 9676 67640
rect 9716 67600 9717 67640
rect 9675 67591 9717 67600
rect 10059 67640 10101 67649
rect 11115 67645 11157 67654
rect 10059 67600 10060 67640
rect 10100 67600 10101 67640
rect 10059 67591 10101 67600
rect 10627 67640 10685 67641
rect 10627 67600 10636 67640
rect 10676 67600 10685 67640
rect 10627 67599 10685 67600
rect 11115 67605 11116 67645
rect 11156 67605 11157 67645
rect 11115 67596 11157 67605
rect 12067 67640 12125 67641
rect 12067 67600 12076 67640
rect 12116 67600 12125 67640
rect 12067 67599 12125 67600
rect 13315 67640 13373 67641
rect 13315 67600 13324 67640
rect 13364 67600 13373 67640
rect 13315 67599 13373 67600
rect 14091 67640 14133 67649
rect 14091 67600 14092 67640
rect 14132 67600 14133 67640
rect 14091 67591 14133 67600
rect 14283 67640 14325 67649
rect 14283 67600 14284 67640
rect 14324 67600 14325 67640
rect 14283 67591 14325 67600
rect 14859 67640 14901 67649
rect 14859 67600 14860 67640
rect 14900 67600 14901 67640
rect 14859 67591 14901 67600
rect 14955 67640 14997 67649
rect 16395 67645 16437 67654
rect 14955 67600 14956 67640
rect 14996 67600 14997 67640
rect 14955 67591 14997 67600
rect 15907 67640 15965 67641
rect 15907 67600 15916 67640
rect 15956 67600 15965 67640
rect 15907 67599 15965 67600
rect 16395 67605 16396 67645
rect 16436 67605 16437 67645
rect 16395 67596 16437 67605
rect 16779 67640 16821 67649
rect 16779 67600 16780 67640
rect 16820 67600 16821 67640
rect 16779 67591 16821 67600
rect 16971 67640 17013 67649
rect 16971 67600 16972 67640
rect 17012 67600 17013 67640
rect 16971 67591 17013 67600
rect 17059 67640 17117 67641
rect 17059 67600 17068 67640
rect 17108 67600 17117 67640
rect 17059 67599 17117 67600
rect 17547 67640 17589 67649
rect 17547 67600 17548 67640
rect 17588 67600 17589 67640
rect 17547 67591 17589 67600
rect 17643 67640 17685 67649
rect 17643 67600 17644 67640
rect 17684 67600 17685 67640
rect 17643 67591 17685 67600
rect 18123 67640 18165 67649
rect 19083 67645 19125 67654
rect 18123 67600 18124 67640
rect 18164 67600 18165 67640
rect 18123 67591 18165 67600
rect 18595 67640 18653 67641
rect 18595 67600 18604 67640
rect 18644 67600 18653 67640
rect 18595 67599 18653 67600
rect 19083 67605 19084 67645
rect 19124 67605 19125 67645
rect 19083 67596 19125 67605
rect 19467 67640 19509 67649
rect 19467 67600 19468 67640
rect 19508 67600 19509 67640
rect 19467 67591 19509 67600
rect 19563 67640 19605 67649
rect 19563 67600 19564 67640
rect 19604 67600 19605 67640
rect 19563 67591 19605 67600
rect 19659 67640 19701 67649
rect 19659 67600 19660 67640
rect 19700 67600 19701 67640
rect 19659 67591 19701 67600
rect 19947 67640 19989 67649
rect 19947 67600 19948 67640
rect 19988 67600 19989 67640
rect 19947 67591 19989 67600
rect 20235 67640 20277 67649
rect 20235 67600 20236 67640
rect 20276 67600 20277 67640
rect 20235 67591 20277 67600
rect 9291 67556 9333 67565
rect 9291 67516 9292 67556
rect 9332 67516 9333 67556
rect 9291 67507 9333 67516
rect 19275 67556 19317 67565
rect 19275 67516 19276 67556
rect 19316 67516 19317 67556
rect 19275 67507 19317 67516
rect 19755 67556 19797 67565
rect 19755 67516 19756 67556
rect 19796 67516 19797 67556
rect 19755 67507 19797 67516
rect 4107 67472 4149 67481
rect 4107 67432 4108 67472
rect 4148 67432 4149 67472
rect 4107 67423 4149 67432
rect 4299 67472 4341 67481
rect 4299 67432 4300 67472
rect 4340 67432 4341 67472
rect 4299 67423 4341 67432
rect 11307 67472 11349 67481
rect 11307 67432 11308 67472
rect 11348 67432 11349 67472
rect 11307 67423 11349 67432
rect 13515 67472 13557 67481
rect 13515 67432 13516 67472
rect 13556 67432 13557 67472
rect 13515 67423 13557 67432
rect 16587 67472 16629 67481
rect 16587 67432 16588 67472
rect 16628 67432 16629 67472
rect 16587 67423 16629 67432
rect 16867 67472 16925 67473
rect 16867 67432 16876 67472
rect 16916 67432 16925 67472
rect 16867 67431 16925 67432
rect 20043 67472 20085 67481
rect 20043 67432 20044 67472
rect 20084 67432 20085 67472
rect 20043 67423 20085 67432
rect 1152 67304 20452 67328
rect 1152 67264 4928 67304
rect 4968 67264 5010 67304
rect 5050 67264 5092 67304
rect 5132 67264 5174 67304
rect 5214 67264 5256 67304
rect 5296 67264 20048 67304
rect 20088 67264 20130 67304
rect 20170 67264 20212 67304
rect 20252 67264 20294 67304
rect 20334 67264 20376 67304
rect 20416 67264 20452 67304
rect 1152 67240 20452 67264
rect 9675 67136 9717 67145
rect 9675 67096 9676 67136
rect 9716 67096 9717 67136
rect 9675 67087 9717 67096
rect 11691 67136 11733 67145
rect 11691 67096 11692 67136
rect 11732 67096 11733 67136
rect 11691 67087 11733 67096
rect 13803 67136 13845 67145
rect 13803 67096 13804 67136
rect 13844 67096 13845 67136
rect 13803 67087 13845 67096
rect 19467 67136 19509 67145
rect 19467 67096 19468 67136
rect 19508 67096 19509 67136
rect 19467 67087 19509 67096
rect 8907 67052 8949 67061
rect 8907 67012 8908 67052
rect 8948 67012 8949 67052
rect 8907 67003 8949 67012
rect 1699 66968 1757 66969
rect 1699 66928 1708 66968
rect 1748 66928 1757 66968
rect 1699 66927 1757 66928
rect 2947 66968 3005 66969
rect 2947 66928 2956 66968
rect 2996 66928 3005 66968
rect 2947 66927 3005 66928
rect 3523 66968 3581 66969
rect 3523 66928 3532 66968
rect 3572 66928 3581 66968
rect 3523 66927 3581 66928
rect 4771 66968 4829 66969
rect 4771 66928 4780 66968
rect 4820 66928 4829 66968
rect 4771 66927 4829 66928
rect 5347 66968 5405 66969
rect 5347 66928 5356 66968
rect 5396 66928 5405 66968
rect 5347 66927 5405 66928
rect 6595 66968 6653 66969
rect 6595 66928 6604 66968
rect 6644 66928 6653 66968
rect 6595 66927 6653 66928
rect 6787 66968 6845 66969
rect 6787 66928 6796 66968
rect 6836 66928 6845 66968
rect 6787 66927 6845 66928
rect 8035 66968 8093 66969
rect 8035 66928 8044 66968
rect 8084 66928 8093 66968
rect 8035 66927 8093 66928
rect 8619 66968 8661 66977
rect 8619 66928 8620 66968
rect 8660 66928 8661 66968
rect 8619 66919 8661 66928
rect 8715 66968 8757 66977
rect 8715 66928 8716 66968
rect 8756 66928 8757 66968
rect 8715 66919 8757 66928
rect 8811 66968 8853 66977
rect 8811 66928 8812 66968
rect 8852 66928 8853 66968
rect 8811 66919 8853 66928
rect 9099 66968 9141 66977
rect 9099 66928 9100 66968
rect 9140 66928 9141 66968
rect 9099 66919 9141 66928
rect 9291 66968 9333 66977
rect 9291 66928 9292 66968
rect 9332 66928 9333 66968
rect 9291 66919 9333 66928
rect 9387 66968 9429 66977
rect 9387 66928 9388 66968
rect 9428 66928 9429 66968
rect 9387 66919 9429 66928
rect 9579 66968 9621 66977
rect 9579 66928 9580 66968
rect 9620 66928 9621 66968
rect 9579 66919 9621 66928
rect 9771 66968 9813 66977
rect 9771 66928 9772 66968
rect 9812 66928 9813 66968
rect 9771 66919 9813 66928
rect 10243 66968 10301 66969
rect 10243 66928 10252 66968
rect 10292 66928 10301 66968
rect 10243 66927 10301 66928
rect 11491 66968 11549 66969
rect 11491 66928 11500 66968
rect 11540 66928 11549 66968
rect 11491 66927 11549 66928
rect 12075 66968 12117 66977
rect 12075 66928 12076 66968
rect 12116 66928 12117 66968
rect 12075 66919 12117 66928
rect 12171 66968 12213 66977
rect 12171 66928 12172 66968
rect 12212 66928 12213 66968
rect 12171 66919 12213 66928
rect 13123 66968 13181 66969
rect 13123 66928 13132 66968
rect 13172 66928 13181 66968
rect 13123 66927 13181 66928
rect 13611 66963 13653 66972
rect 13611 66923 13612 66963
rect 13652 66923 13653 66963
rect 14179 66968 14237 66969
rect 14179 66928 14188 66968
rect 14228 66928 14237 66968
rect 14179 66927 14237 66928
rect 15427 66968 15485 66969
rect 15427 66928 15436 66968
rect 15476 66928 15485 66968
rect 15427 66927 15485 66928
rect 15619 66968 15677 66969
rect 15619 66928 15628 66968
rect 15668 66928 15677 66968
rect 15619 66927 15677 66928
rect 16867 66968 16925 66969
rect 16867 66928 16876 66968
rect 16916 66928 16925 66968
rect 16867 66927 16925 66928
rect 17251 66968 17309 66969
rect 17251 66928 17260 66968
rect 17300 66928 17309 66968
rect 17251 66927 17309 66928
rect 17355 66968 17397 66977
rect 17355 66928 17356 66968
rect 17396 66928 17397 66968
rect 13611 66914 13653 66923
rect 17355 66919 17397 66928
rect 17547 66968 17589 66977
rect 17547 66928 17548 66968
rect 17588 66928 17589 66968
rect 17547 66919 17589 66928
rect 18019 66968 18077 66969
rect 18019 66928 18028 66968
rect 18068 66928 18077 66968
rect 18019 66927 18077 66928
rect 19267 66968 19325 66969
rect 19267 66928 19276 66968
rect 19316 66928 19325 66968
rect 19267 66927 19325 66928
rect 19755 66968 19797 66977
rect 19755 66928 19756 66968
rect 19796 66928 19797 66968
rect 19755 66919 19797 66928
rect 12555 66884 12597 66893
rect 12555 66844 12556 66884
rect 12596 66844 12597 66884
rect 12555 66835 12597 66844
rect 12651 66884 12693 66893
rect 12651 66844 12652 66884
rect 12692 66844 12693 66884
rect 12651 66835 12693 66844
rect 8235 66800 8277 66809
rect 8235 66760 8236 66800
rect 8276 66760 8277 66800
rect 8235 66751 8277 66760
rect 9379 66800 9437 66801
rect 9379 66760 9388 66800
rect 9428 66760 9437 66800
rect 9379 66759 9437 66760
rect 13995 66800 14037 66809
rect 13995 66760 13996 66800
rect 14036 66760 14037 66800
rect 13995 66751 14037 66760
rect 17547 66800 17589 66809
rect 17547 66760 17548 66800
rect 17588 66760 17589 66800
rect 17547 66751 17589 66760
rect 19755 66800 19797 66809
rect 19755 66760 19756 66800
rect 19796 66760 19797 66800
rect 19755 66751 19797 66760
rect 19947 66800 19989 66809
rect 19947 66760 19948 66800
rect 19988 66760 19989 66800
rect 19947 66751 19989 66760
rect 3147 66716 3189 66725
rect 3147 66676 3148 66716
rect 3188 66676 3189 66716
rect 3147 66667 3189 66676
rect 4971 66716 5013 66725
rect 4971 66676 4972 66716
rect 5012 66676 5013 66716
rect 4971 66667 5013 66676
rect 5163 66716 5205 66725
rect 5163 66676 5164 66716
rect 5204 66676 5205 66716
rect 5163 66667 5205 66676
rect 17067 66716 17109 66725
rect 17067 66676 17068 66716
rect 17108 66676 17109 66716
rect 17067 66667 17109 66676
rect 1152 66548 20352 66572
rect 1152 66508 3688 66548
rect 3728 66508 3770 66548
rect 3810 66508 3852 66548
rect 3892 66508 3934 66548
rect 3974 66508 4016 66548
rect 4056 66508 18808 66548
rect 18848 66508 18890 66548
rect 18930 66508 18972 66548
rect 19012 66508 19054 66548
rect 19094 66508 19136 66548
rect 19176 66508 20352 66548
rect 1152 66484 20352 66508
rect 9099 66380 9141 66389
rect 9099 66340 9100 66380
rect 9140 66340 9141 66380
rect 9099 66331 9141 66340
rect 9675 66380 9717 66389
rect 9675 66340 9676 66380
rect 9716 66340 9717 66380
rect 9675 66331 9717 66340
rect 12363 66380 12405 66389
rect 12363 66340 12364 66380
rect 12404 66340 12405 66380
rect 12363 66331 12405 66340
rect 16107 66380 16149 66389
rect 16107 66340 16108 66380
rect 16148 66340 16149 66380
rect 16107 66331 16149 66340
rect 19851 66380 19893 66389
rect 19851 66340 19852 66380
rect 19892 66340 19893 66380
rect 19851 66331 19893 66340
rect 7171 66296 7229 66297
rect 7171 66256 7180 66296
rect 7220 66256 7229 66296
rect 7171 66255 7229 66256
rect 9963 66296 10005 66305
rect 9963 66256 9964 66296
rect 10004 66256 10005 66296
rect 9963 66247 10005 66256
rect 5067 66212 5109 66221
rect 5067 66172 5068 66212
rect 5108 66172 5109 66212
rect 5067 66163 5109 66172
rect 16875 66212 16917 66221
rect 16875 66172 16876 66212
rect 16916 66172 16917 66212
rect 16875 66163 16917 66172
rect 13507 66147 13565 66148
rect 1219 66128 1277 66129
rect 1219 66088 1228 66128
rect 1268 66088 1277 66128
rect 1219 66087 1277 66088
rect 2467 66128 2525 66129
rect 2467 66088 2476 66128
rect 2516 66088 2525 66128
rect 2467 66087 2525 66088
rect 3531 66128 3573 66137
rect 3531 66088 3532 66128
rect 3572 66088 3573 66128
rect 3531 66079 3573 66088
rect 3627 66128 3669 66137
rect 3627 66088 3628 66128
rect 3668 66088 3669 66128
rect 3627 66079 3669 66088
rect 3723 66128 3765 66137
rect 3723 66088 3724 66128
rect 3764 66088 3765 66128
rect 3723 66079 3765 66088
rect 3915 66128 3957 66137
rect 3915 66088 3916 66128
rect 3956 66088 3957 66128
rect 3915 66079 3957 66088
rect 4011 66128 4053 66137
rect 4011 66088 4012 66128
rect 4052 66088 4053 66128
rect 4011 66079 4053 66088
rect 4107 66128 4149 66137
rect 4107 66088 4108 66128
rect 4148 66088 4149 66128
rect 4107 66079 4149 66088
rect 4203 66128 4245 66137
rect 4203 66088 4204 66128
rect 4244 66088 4245 66128
rect 4203 66079 4245 66088
rect 4491 66128 4533 66137
rect 4491 66088 4492 66128
rect 4532 66088 4533 66128
rect 4491 66079 4533 66088
rect 4587 66128 4629 66137
rect 4587 66088 4588 66128
rect 4628 66088 4629 66128
rect 4587 66079 4629 66088
rect 4971 66128 5013 66137
rect 6027 66133 6069 66142
rect 4971 66088 4972 66128
rect 5012 66088 5013 66128
rect 4971 66079 5013 66088
rect 5539 66128 5597 66129
rect 5539 66088 5548 66128
rect 5588 66088 5597 66128
rect 5539 66087 5597 66088
rect 6027 66093 6028 66133
rect 6068 66093 6069 66133
rect 6027 66084 6069 66093
rect 6499 66128 6557 66129
rect 6499 66088 6508 66128
rect 6548 66088 6557 66128
rect 6499 66087 6557 66088
rect 6795 66128 6837 66137
rect 6795 66088 6796 66128
rect 6836 66088 6837 66128
rect 6795 66079 6837 66088
rect 6891 66128 6933 66137
rect 6891 66088 6892 66128
rect 6932 66088 6933 66128
rect 6891 66079 6933 66088
rect 7651 66128 7709 66129
rect 7651 66088 7660 66128
rect 7700 66088 7709 66128
rect 7651 66087 7709 66088
rect 8899 66128 8957 66129
rect 8899 66088 8908 66128
rect 8948 66088 8957 66128
rect 8899 66087 8957 66088
rect 9387 66128 9429 66137
rect 9387 66088 9388 66128
rect 9428 66088 9429 66128
rect 9387 66079 9429 66088
rect 9675 66121 9717 66130
rect 9675 66081 9676 66121
rect 9716 66081 9717 66121
rect 9675 66072 9717 66081
rect 9963 66128 10005 66137
rect 9963 66088 9964 66128
rect 10004 66088 10005 66128
rect 9963 66079 10005 66088
rect 12363 66128 12405 66137
rect 12363 66088 12364 66128
rect 12404 66088 12405 66128
rect 12363 66079 12405 66088
rect 12555 66128 12597 66137
rect 12555 66088 12556 66128
rect 12596 66088 12597 66128
rect 12555 66079 12597 66088
rect 12739 66128 12797 66129
rect 12739 66088 12748 66128
rect 12788 66088 12797 66128
rect 12739 66087 12797 66088
rect 12843 66128 12885 66137
rect 12843 66088 12844 66128
rect 12884 66088 12885 66128
rect 12843 66079 12885 66088
rect 13035 66128 13077 66137
rect 13035 66088 13036 66128
rect 13076 66088 13077 66128
rect 13035 66079 13077 66088
rect 13131 66128 13173 66137
rect 13131 66088 13132 66128
rect 13172 66088 13173 66128
rect 13131 66079 13173 66088
rect 13227 66128 13269 66137
rect 13227 66088 13228 66128
rect 13268 66088 13269 66128
rect 13507 66107 13516 66147
rect 13556 66107 13565 66147
rect 13507 66106 13565 66107
rect 13611 66128 13653 66137
rect 13227 66079 13269 66088
rect 13611 66088 13612 66128
rect 13652 66088 13653 66128
rect 13611 66079 13653 66088
rect 13803 66128 13845 66137
rect 13803 66088 13804 66128
rect 13844 66088 13845 66128
rect 13803 66079 13845 66088
rect 14179 66128 14237 66129
rect 14179 66088 14188 66128
rect 14228 66088 14237 66128
rect 14179 66087 14237 66088
rect 14283 66128 14325 66137
rect 14283 66088 14284 66128
rect 14324 66088 14325 66128
rect 14283 66079 14325 66088
rect 14475 66128 14517 66137
rect 14475 66088 14476 66128
rect 14516 66088 14517 66128
rect 14475 66079 14517 66088
rect 16003 66128 16061 66129
rect 16003 66088 16012 66128
rect 16052 66088 16061 66128
rect 16003 66087 16061 66088
rect 16299 66128 16341 66137
rect 16299 66088 16300 66128
rect 16340 66088 16341 66128
rect 16299 66079 16341 66088
rect 16395 66128 16437 66137
rect 16395 66088 16396 66128
rect 16436 66088 16437 66128
rect 16395 66079 16437 66088
rect 16491 66128 16533 66137
rect 16491 66088 16492 66128
rect 16532 66088 16533 66128
rect 16491 66079 16533 66088
rect 16587 66128 16629 66137
rect 16587 66088 16588 66128
rect 16628 66088 16629 66128
rect 16587 66079 16629 66088
rect 16779 66128 16821 66137
rect 16779 66088 16780 66128
rect 16820 66088 16821 66128
rect 16779 66079 16821 66088
rect 16971 66128 17013 66137
rect 16971 66088 16972 66128
rect 17012 66088 17013 66128
rect 16971 66079 17013 66088
rect 18403 66128 18461 66129
rect 18403 66088 18412 66128
rect 18452 66088 18461 66128
rect 18403 66087 18461 66088
rect 19651 66128 19709 66129
rect 19651 66088 19660 66128
rect 19700 66088 19709 66128
rect 19651 66087 19709 66088
rect 13707 66044 13749 66053
rect 13707 66004 13708 66044
rect 13748 66004 13749 66044
rect 13707 65995 13749 66004
rect 2667 65960 2709 65969
rect 2667 65920 2668 65960
rect 2708 65920 2709 65960
rect 2667 65911 2709 65920
rect 3427 65960 3485 65961
rect 3427 65920 3436 65960
rect 3476 65920 3485 65960
rect 3427 65919 3485 65920
rect 6219 65960 6261 65969
rect 6219 65920 6220 65960
rect 6260 65920 6261 65960
rect 6219 65911 6261 65920
rect 9099 65960 9141 65969
rect 9099 65920 9100 65960
rect 9140 65920 9141 65960
rect 9099 65911 9141 65920
rect 10155 65960 10197 65969
rect 10155 65920 10156 65960
rect 10196 65920 10197 65960
rect 10155 65911 10197 65920
rect 13315 65960 13373 65961
rect 13315 65920 13324 65960
rect 13364 65920 13373 65960
rect 13315 65919 13373 65920
rect 14371 65960 14429 65961
rect 14371 65920 14380 65960
rect 14420 65920 14429 65960
rect 14371 65919 14429 65920
rect 1152 65792 20452 65816
rect 1152 65752 4928 65792
rect 4968 65752 5010 65792
rect 5050 65752 5092 65792
rect 5132 65752 5174 65792
rect 5214 65752 5256 65792
rect 5296 65752 20048 65792
rect 20088 65752 20130 65792
rect 20170 65752 20212 65792
rect 20252 65752 20294 65792
rect 20334 65752 20376 65792
rect 20416 65752 20452 65792
rect 1152 65728 20452 65752
rect 5923 65624 5981 65625
rect 5923 65584 5932 65624
rect 5972 65584 5981 65624
rect 5923 65583 5981 65584
rect 9291 65624 9333 65633
rect 9291 65584 9292 65624
rect 9332 65584 9333 65624
rect 9291 65575 9333 65584
rect 9483 65624 9525 65633
rect 9483 65584 9484 65624
rect 9524 65584 9525 65624
rect 9483 65575 9525 65584
rect 13027 65624 13085 65625
rect 13027 65584 13036 65624
rect 13076 65584 13085 65624
rect 13027 65583 13085 65584
rect 3339 65540 3381 65549
rect 3339 65500 3340 65540
rect 3380 65500 3381 65540
rect 3339 65491 3381 65500
rect 6507 65540 6549 65549
rect 6507 65500 6508 65540
rect 6548 65500 6549 65540
rect 6507 65491 6549 65500
rect 13323 65540 13365 65549
rect 13323 65500 13324 65540
rect 13364 65500 13365 65540
rect 13323 65491 13365 65500
rect 15915 65540 15957 65549
rect 15915 65500 15916 65540
rect 15956 65500 15957 65540
rect 15915 65491 15957 65500
rect 17931 65540 17973 65549
rect 17931 65500 17932 65540
rect 17972 65500 17973 65540
rect 17931 65491 17973 65500
rect 12939 65477 12981 65486
rect 1611 65456 1653 65465
rect 1611 65416 1612 65456
rect 1652 65416 1653 65456
rect 1611 65407 1653 65416
rect 1707 65456 1749 65465
rect 1707 65416 1708 65456
rect 1748 65416 1749 65456
rect 1707 65407 1749 65416
rect 2091 65456 2133 65465
rect 2091 65416 2092 65456
rect 2132 65416 2133 65456
rect 2091 65407 2133 65416
rect 2187 65456 2229 65465
rect 2187 65416 2188 65456
rect 2228 65416 2229 65456
rect 2187 65407 2229 65416
rect 2659 65456 2717 65457
rect 2659 65416 2668 65456
rect 2708 65416 2717 65456
rect 2659 65415 2717 65416
rect 3147 65451 3189 65460
rect 3147 65411 3148 65451
rect 3188 65411 3189 65451
rect 4291 65456 4349 65457
rect 4291 65416 4300 65456
rect 4340 65416 4349 65456
rect 4291 65415 4349 65416
rect 5539 65456 5597 65457
rect 5539 65416 5548 65456
rect 5588 65416 5597 65456
rect 5539 65415 5597 65416
rect 6123 65456 6165 65465
rect 6123 65416 6124 65456
rect 6164 65416 6165 65456
rect 3147 65402 3189 65411
rect 6123 65407 6165 65416
rect 6219 65456 6261 65465
rect 6219 65416 6220 65456
rect 6260 65416 6261 65456
rect 6219 65407 6261 65416
rect 6411 65456 6453 65465
rect 6411 65416 6412 65456
rect 6452 65416 6453 65456
rect 6411 65407 6453 65416
rect 6603 65456 6645 65465
rect 6603 65416 6604 65456
rect 6644 65416 6645 65456
rect 6603 65407 6645 65416
rect 6691 65456 6749 65457
rect 6691 65416 6700 65456
rect 6740 65416 6749 65456
rect 6691 65415 6749 65416
rect 6987 65456 7029 65465
rect 6987 65416 6988 65456
rect 7028 65416 7029 65456
rect 6987 65407 7029 65416
rect 7275 65456 7317 65465
rect 7275 65416 7276 65456
rect 7316 65416 7317 65456
rect 7275 65407 7317 65416
rect 7563 65456 7605 65465
rect 7563 65416 7564 65456
rect 7604 65416 7605 65456
rect 7563 65407 7605 65416
rect 7659 65456 7701 65465
rect 7659 65416 7660 65456
rect 7700 65416 7701 65456
rect 7659 65407 7701 65416
rect 8043 65456 8085 65465
rect 8043 65416 8044 65456
rect 8084 65416 8085 65456
rect 8043 65407 8085 65416
rect 8139 65456 8181 65465
rect 8139 65416 8140 65456
rect 8180 65416 8181 65456
rect 8139 65407 8181 65416
rect 8611 65456 8669 65457
rect 8611 65416 8620 65456
rect 8660 65416 8669 65456
rect 8611 65415 8669 65416
rect 9099 65451 9141 65460
rect 9099 65411 9100 65451
rect 9140 65411 9141 65451
rect 9667 65456 9725 65457
rect 9667 65416 9676 65456
rect 9716 65416 9725 65456
rect 9667 65415 9725 65416
rect 10915 65456 10973 65457
rect 10915 65416 10924 65456
rect 10964 65416 10973 65456
rect 10915 65415 10973 65416
rect 11107 65456 11165 65457
rect 11107 65416 11116 65456
rect 11156 65416 11165 65456
rect 11107 65415 11165 65416
rect 12355 65456 12413 65457
rect 12355 65416 12364 65456
rect 12404 65416 12413 65456
rect 12355 65415 12413 65416
rect 12747 65456 12789 65465
rect 12747 65416 12748 65456
rect 12788 65416 12789 65456
rect 9099 65402 9141 65411
rect 12747 65407 12789 65416
rect 12843 65456 12885 65465
rect 12843 65416 12844 65456
rect 12884 65416 12885 65456
rect 12939 65437 12940 65477
rect 12980 65437 12981 65477
rect 12939 65428 12981 65437
rect 13227 65456 13269 65465
rect 12843 65407 12885 65416
rect 13227 65416 13228 65456
rect 13268 65416 13269 65456
rect 13227 65407 13269 65416
rect 13419 65456 13461 65465
rect 13419 65416 13420 65456
rect 13460 65416 13461 65456
rect 13419 65407 13461 65416
rect 13507 65456 13565 65457
rect 13507 65416 13516 65456
rect 13556 65416 13565 65456
rect 13507 65415 13565 65416
rect 14467 65456 14525 65457
rect 14467 65416 14476 65456
rect 14516 65416 14525 65456
rect 14467 65415 14525 65416
rect 15715 65456 15773 65457
rect 15715 65416 15724 65456
rect 15764 65416 15773 65456
rect 15715 65415 15773 65416
rect 16203 65456 16245 65465
rect 16203 65416 16204 65456
rect 16244 65416 16245 65456
rect 16203 65407 16245 65416
rect 16299 65456 16341 65465
rect 16299 65416 16300 65456
rect 16340 65416 16341 65456
rect 16299 65407 16341 65416
rect 16683 65456 16725 65465
rect 16683 65416 16684 65456
rect 16724 65416 16725 65456
rect 16683 65407 16725 65416
rect 17251 65456 17309 65457
rect 17251 65416 17260 65456
rect 17300 65416 17309 65456
rect 17251 65415 17309 65416
rect 17739 65442 17781 65451
rect 17739 65402 17740 65442
rect 17780 65402 17781 65442
rect 17739 65393 17781 65402
rect 16779 65372 16821 65381
rect 16779 65332 16780 65372
rect 16820 65332 16821 65372
rect 16779 65323 16821 65332
rect 6987 65288 7029 65297
rect 6987 65248 6988 65288
rect 7028 65248 7029 65288
rect 6987 65239 7029 65248
rect 12555 65288 12597 65297
rect 12555 65248 12556 65288
rect 12596 65248 12597 65288
rect 12555 65239 12597 65248
rect 5739 65204 5781 65213
rect 5739 65164 5740 65204
rect 5780 65164 5781 65204
rect 5739 65155 5781 65164
rect 1152 65036 20352 65060
rect 1152 64996 3688 65036
rect 3728 64996 3770 65036
rect 3810 64996 3852 65036
rect 3892 64996 3934 65036
rect 3974 64996 4016 65036
rect 4056 64996 18808 65036
rect 18848 64996 18890 65036
rect 18930 64996 18972 65036
rect 19012 64996 19054 65036
rect 19094 64996 19136 65036
rect 19176 64996 20352 65036
rect 1152 64972 20352 64996
rect 11019 64868 11061 64877
rect 11019 64828 11020 64868
rect 11060 64828 11061 64868
rect 11019 64819 11061 64828
rect 13707 64868 13749 64877
rect 13707 64828 13708 64868
rect 13748 64828 13749 64868
rect 13707 64819 13749 64828
rect 17643 64868 17685 64877
rect 17643 64828 17644 64868
rect 17684 64828 17685 64868
rect 17643 64819 17685 64828
rect 5259 64700 5301 64709
rect 5259 64660 5260 64700
rect 5300 64660 5301 64700
rect 5259 64651 5301 64660
rect 11787 64700 11829 64709
rect 11787 64660 11788 64700
rect 11828 64660 11829 64700
rect 11787 64651 11829 64660
rect 11883 64700 11925 64709
rect 11883 64660 11884 64700
rect 11924 64660 11925 64700
rect 11883 64651 11925 64660
rect 1219 64616 1277 64617
rect 1219 64576 1228 64616
rect 1268 64576 1277 64616
rect 1219 64575 1277 64576
rect 2467 64616 2525 64617
rect 2467 64576 2476 64616
rect 2516 64576 2525 64616
rect 2467 64575 2525 64576
rect 3523 64616 3581 64617
rect 3523 64576 3532 64616
rect 3572 64576 3581 64616
rect 3523 64575 3581 64576
rect 4771 64616 4829 64617
rect 4771 64576 4780 64616
rect 4820 64576 4829 64616
rect 4771 64575 4829 64576
rect 5163 64616 5205 64625
rect 5163 64576 5164 64616
rect 5204 64576 5205 64616
rect 5163 64567 5205 64576
rect 5355 64616 5397 64625
rect 5355 64576 5356 64616
rect 5396 64576 5397 64616
rect 5355 64567 5397 64576
rect 5539 64616 5597 64617
rect 5539 64576 5548 64616
rect 5588 64576 5597 64616
rect 5539 64575 5597 64576
rect 6787 64616 6845 64617
rect 6787 64576 6796 64616
rect 6836 64576 6845 64616
rect 6787 64575 6845 64576
rect 7363 64616 7421 64617
rect 7363 64576 7372 64616
rect 7412 64576 7421 64616
rect 7363 64575 7421 64576
rect 8611 64616 8669 64617
rect 8611 64576 8620 64616
rect 8660 64576 8669 64616
rect 8611 64575 8669 64576
rect 8907 64616 8949 64625
rect 8907 64576 8908 64616
rect 8948 64576 8949 64616
rect 8907 64567 8949 64576
rect 9003 64616 9045 64625
rect 9003 64576 9004 64616
rect 9044 64576 9045 64616
rect 9003 64567 9045 64576
rect 9571 64616 9629 64617
rect 9571 64576 9580 64616
rect 9620 64576 9629 64616
rect 9571 64575 9629 64576
rect 10819 64616 10877 64617
rect 10819 64576 10828 64616
rect 10868 64576 10877 64616
rect 10819 64575 10877 64576
rect 11307 64616 11349 64625
rect 11307 64576 11308 64616
rect 11348 64576 11349 64616
rect 11307 64567 11349 64576
rect 11403 64616 11445 64625
rect 12843 64621 12885 64630
rect 11403 64576 11404 64616
rect 11444 64576 11445 64616
rect 11403 64567 11445 64576
rect 12355 64616 12413 64617
rect 12355 64576 12364 64616
rect 12404 64576 12413 64616
rect 12355 64575 12413 64576
rect 12843 64581 12844 64621
rect 12884 64581 12885 64621
rect 12843 64572 12885 64581
rect 13227 64616 13269 64625
rect 13227 64576 13228 64616
rect 13268 64576 13269 64616
rect 13227 64567 13269 64576
rect 13323 64616 13365 64625
rect 13323 64576 13324 64616
rect 13364 64576 13365 64616
rect 13323 64567 13365 64576
rect 13419 64616 13461 64625
rect 13419 64576 13420 64616
rect 13460 64576 13461 64616
rect 13419 64567 13461 64576
rect 13515 64616 13557 64625
rect 13515 64576 13516 64616
rect 13556 64576 13557 64616
rect 13515 64567 13557 64576
rect 13707 64616 13749 64625
rect 13707 64576 13708 64616
rect 13748 64576 13749 64616
rect 13707 64567 13749 64576
rect 13899 64616 13941 64625
rect 13899 64576 13900 64616
rect 13940 64576 13941 64616
rect 13899 64567 13941 64576
rect 14083 64616 14141 64617
rect 14083 64576 14092 64616
rect 14132 64576 14141 64616
rect 14083 64575 14141 64576
rect 15331 64616 15389 64617
rect 15331 64576 15340 64616
rect 15380 64576 15389 64616
rect 15331 64575 15389 64576
rect 15723 64616 15765 64625
rect 15723 64576 15724 64616
rect 15764 64576 15765 64616
rect 15723 64567 15765 64576
rect 16011 64616 16053 64625
rect 16011 64576 16012 64616
rect 16052 64576 16053 64616
rect 16011 64567 16053 64576
rect 16195 64616 16253 64617
rect 16195 64576 16204 64616
rect 16244 64576 16253 64616
rect 16195 64575 16253 64576
rect 17443 64616 17501 64617
rect 17443 64576 17452 64616
rect 17492 64576 17501 64616
rect 17443 64575 17501 64576
rect 17827 64616 17885 64617
rect 17827 64576 17836 64616
rect 17876 64576 17885 64616
rect 17827 64575 17885 64576
rect 7179 64532 7221 64541
rect 7179 64492 7180 64532
rect 7220 64492 7221 64532
rect 7179 64483 7221 64492
rect 13035 64532 13077 64541
rect 13035 64492 13036 64532
rect 13076 64492 13077 64532
rect 13035 64483 13077 64492
rect 2667 64448 2709 64457
rect 2667 64408 2668 64448
rect 2708 64408 2709 64448
rect 2667 64399 2709 64408
rect 4971 64448 5013 64457
rect 4971 64408 4972 64448
rect 5012 64408 5013 64448
rect 4971 64399 5013 64408
rect 6987 64448 7029 64457
rect 6987 64408 6988 64448
rect 7028 64408 7029 64448
rect 6987 64399 7029 64408
rect 9187 64448 9245 64449
rect 9187 64408 9196 64448
rect 9236 64408 9245 64448
rect 9187 64407 9245 64408
rect 15531 64448 15573 64457
rect 15531 64408 15532 64448
rect 15572 64408 15573 64448
rect 15531 64399 15573 64408
rect 15915 64448 15957 64457
rect 15915 64408 15916 64448
rect 15956 64408 15957 64448
rect 15915 64399 15957 64408
rect 17931 64448 17973 64457
rect 17931 64408 17932 64448
rect 17972 64408 17973 64448
rect 17931 64399 17973 64408
rect 1152 64280 20452 64304
rect 1152 64240 4928 64280
rect 4968 64240 5010 64280
rect 5050 64240 5092 64280
rect 5132 64240 5174 64280
rect 5214 64240 5256 64280
rect 5296 64240 20048 64280
rect 20088 64240 20130 64280
rect 20170 64240 20212 64280
rect 20252 64240 20294 64280
rect 20334 64240 20376 64280
rect 20416 64240 20452 64280
rect 1152 64216 20452 64240
rect 4011 64112 4053 64121
rect 4011 64072 4012 64112
rect 4052 64072 4053 64112
rect 4011 64063 4053 64072
rect 7179 64112 7221 64121
rect 7179 64072 7180 64112
rect 7220 64072 7221 64112
rect 7179 64063 7221 64072
rect 8323 64112 8381 64113
rect 8323 64072 8332 64112
rect 8372 64072 8381 64112
rect 8323 64071 8381 64072
rect 12267 64112 12309 64121
rect 12267 64072 12268 64112
rect 12308 64072 12309 64112
rect 17347 64112 17405 64113
rect 8131 64070 8189 64071
rect 8131 64030 8140 64070
rect 8180 64030 8189 64070
rect 12267 64063 12309 64072
rect 15531 64070 15573 64079
rect 17347 64072 17356 64112
rect 17396 64072 17405 64112
rect 17347 64071 17405 64072
rect 18019 64112 18077 64113
rect 18019 64072 18028 64112
rect 18068 64072 18077 64112
rect 18019 64071 18077 64072
rect 8131 64029 8189 64030
rect 12939 64028 12981 64037
rect 12939 63988 12940 64028
rect 12980 63988 12981 64028
rect 15531 64030 15532 64070
rect 15572 64030 15573 64070
rect 15531 64021 15573 64030
rect 12939 63979 12981 63988
rect 2283 63944 2325 63953
rect 2283 63904 2284 63944
rect 2324 63904 2325 63944
rect 2283 63895 2325 63904
rect 2379 63944 2421 63953
rect 2379 63904 2380 63944
rect 2420 63904 2421 63944
rect 2379 63895 2421 63904
rect 2763 63944 2805 63953
rect 2763 63904 2764 63944
rect 2804 63904 2805 63944
rect 2763 63895 2805 63904
rect 2859 63944 2901 63953
rect 2859 63904 2860 63944
rect 2900 63904 2901 63944
rect 2859 63895 2901 63904
rect 3331 63944 3389 63945
rect 3331 63904 3340 63944
rect 3380 63904 3389 63944
rect 3331 63903 3389 63904
rect 3819 63939 3861 63948
rect 3819 63899 3820 63939
rect 3860 63899 3861 63939
rect 3819 63890 3861 63899
rect 5451 63944 5493 63953
rect 5451 63904 5452 63944
rect 5492 63904 5493 63944
rect 5451 63895 5493 63904
rect 5547 63944 5589 63953
rect 5547 63904 5548 63944
rect 5588 63904 5589 63944
rect 5547 63895 5589 63904
rect 6027 63944 6069 63953
rect 6027 63904 6028 63944
rect 6068 63904 6069 63944
rect 6027 63895 6069 63904
rect 6499 63944 6557 63945
rect 6499 63904 6508 63944
rect 6548 63904 6557 63944
rect 6499 63903 6557 63904
rect 6987 63939 7029 63948
rect 6987 63899 6988 63939
rect 7028 63899 7029 63939
rect 6987 63890 7029 63899
rect 7851 63944 7893 63953
rect 7851 63904 7852 63944
rect 7892 63904 7893 63944
rect 7851 63895 7893 63904
rect 7947 63944 7989 63953
rect 7947 63904 7948 63944
rect 7988 63904 7989 63944
rect 7947 63895 7989 63904
rect 8419 63944 8477 63945
rect 8419 63904 8428 63944
rect 8468 63904 8477 63944
rect 8419 63903 8477 63904
rect 8803 63944 8861 63945
rect 8803 63904 8812 63944
rect 8852 63904 8861 63944
rect 8803 63903 8861 63904
rect 10051 63944 10109 63945
rect 10051 63904 10060 63944
rect 10100 63904 10109 63944
rect 10051 63903 10109 63904
rect 10819 63944 10877 63945
rect 10819 63904 10828 63944
rect 10868 63904 10877 63944
rect 10819 63903 10877 63904
rect 12067 63944 12125 63945
rect 12067 63904 12076 63944
rect 12116 63904 12125 63944
rect 12067 63903 12125 63904
rect 12547 63944 12605 63945
rect 12547 63904 12556 63944
rect 12596 63904 12605 63944
rect 12547 63903 12605 63904
rect 12843 63944 12885 63953
rect 12843 63904 12844 63944
rect 12884 63904 12885 63944
rect 12843 63895 12885 63904
rect 13803 63944 13845 63953
rect 13803 63904 13804 63944
rect 13844 63904 13845 63944
rect 13803 63895 13845 63904
rect 13899 63944 13941 63953
rect 13899 63904 13900 63944
rect 13940 63904 13941 63944
rect 13899 63895 13941 63904
rect 14379 63944 14421 63953
rect 14379 63904 14380 63944
rect 14420 63904 14421 63944
rect 14379 63895 14421 63904
rect 14851 63944 14909 63945
rect 14851 63904 14860 63944
rect 14900 63904 14909 63944
rect 15723 63944 15765 63953
rect 14851 63903 14909 63904
rect 15339 63930 15381 63939
rect 15339 63890 15340 63930
rect 15380 63890 15381 63930
rect 15723 63904 15724 63944
rect 15764 63904 15765 63944
rect 15723 63895 15765 63904
rect 15915 63944 15957 63953
rect 15915 63904 15916 63944
rect 15956 63904 15957 63944
rect 15915 63895 15957 63904
rect 16011 63944 16053 63953
rect 16011 63904 16012 63944
rect 16052 63904 16053 63944
rect 16011 63895 16053 63904
rect 16203 63944 16245 63953
rect 16203 63904 16204 63944
rect 16244 63904 16245 63944
rect 16203 63895 16245 63904
rect 16395 63944 16437 63953
rect 16395 63904 16396 63944
rect 16436 63904 16437 63944
rect 16395 63895 16437 63904
rect 16491 63944 16533 63953
rect 16491 63904 16492 63944
rect 16532 63904 16533 63944
rect 16491 63895 16533 63904
rect 16779 63944 16821 63953
rect 16779 63904 16780 63944
rect 16820 63904 16821 63944
rect 16779 63895 16821 63904
rect 17342 63944 17400 63945
rect 17342 63904 17351 63944
rect 17391 63904 17400 63944
rect 17342 63903 17400 63904
rect 17451 63944 17493 63953
rect 17451 63904 17452 63944
rect 17492 63904 17493 63944
rect 17451 63895 17493 63904
rect 17547 63944 17589 63953
rect 17547 63904 17548 63944
rect 17588 63904 17589 63944
rect 17547 63895 17589 63904
rect 17731 63944 17789 63945
rect 17731 63904 17740 63944
rect 17780 63904 17789 63944
rect 17731 63903 17789 63904
rect 17827 63944 17885 63945
rect 17827 63904 17836 63944
rect 17876 63904 17885 63944
rect 17827 63903 17885 63904
rect 18219 63944 18261 63953
rect 18219 63904 18220 63944
rect 18260 63904 18261 63944
rect 18219 63895 18261 63904
rect 18315 63944 18357 63953
rect 18315 63904 18316 63944
rect 18356 63904 18357 63944
rect 18315 63895 18357 63904
rect 15339 63881 15381 63890
rect 5931 63860 5973 63869
rect 5931 63820 5932 63860
rect 5972 63820 5973 63860
rect 5931 63811 5973 63820
rect 14283 63860 14325 63869
rect 14283 63820 14284 63860
rect 14324 63820 14325 63860
rect 14283 63811 14325 63820
rect 13219 63776 13277 63777
rect 13219 63736 13228 63776
rect 13268 63736 13277 63776
rect 13219 63735 13277 63736
rect 16483 63776 16541 63777
rect 16483 63736 16492 63776
rect 16532 63736 16541 63776
rect 16483 63735 16541 63736
rect 16779 63776 16821 63785
rect 16779 63736 16780 63776
rect 16820 63736 16821 63776
rect 16779 63727 16821 63736
rect 8611 63692 8669 63693
rect 8611 63652 8620 63692
rect 8660 63652 8669 63692
rect 8611 63651 8669 63652
rect 10251 63692 10293 63701
rect 10251 63652 10252 63692
rect 10292 63652 10293 63692
rect 10251 63643 10293 63652
rect 16971 63692 17013 63701
rect 16971 63652 16972 63692
rect 17012 63652 17013 63692
rect 16971 63643 17013 63652
rect 1152 63524 20352 63548
rect 1152 63484 3688 63524
rect 3728 63484 3770 63524
rect 3810 63484 3852 63524
rect 3892 63484 3934 63524
rect 3974 63484 4016 63524
rect 4056 63484 18808 63524
rect 18848 63484 18890 63524
rect 18930 63484 18972 63524
rect 19012 63484 19054 63524
rect 19094 63484 19136 63524
rect 19176 63484 20352 63524
rect 1152 63460 20352 63484
rect 14667 63356 14709 63365
rect 14667 63316 14668 63356
rect 14708 63316 14709 63356
rect 14667 63307 14709 63316
rect 14859 63356 14901 63365
rect 14859 63316 14860 63356
rect 14900 63316 14901 63356
rect 14859 63307 14901 63316
rect 17931 63356 17973 63365
rect 17931 63316 17932 63356
rect 17972 63316 17973 63356
rect 17931 63307 17973 63316
rect 18115 63272 18173 63273
rect 18115 63232 18124 63272
rect 18164 63232 18173 63272
rect 18115 63231 18173 63232
rect 3243 63188 3285 63197
rect 3243 63148 3244 63188
rect 3284 63148 3285 63188
rect 3243 63139 3285 63148
rect 3339 63188 3381 63197
rect 3339 63148 3340 63188
rect 3380 63148 3381 63188
rect 3339 63139 3381 63148
rect 8139 63188 8181 63197
rect 8139 63148 8140 63188
rect 8180 63148 8181 63188
rect 8139 63139 8181 63148
rect 8235 63188 8277 63197
rect 8235 63148 8236 63188
rect 8276 63148 8277 63188
rect 11211 63188 11253 63197
rect 8235 63139 8277 63148
rect 10251 63146 10293 63155
rect 2763 63123 2805 63132
rect 2763 63083 2764 63123
rect 2804 63083 2805 63123
rect 4299 63118 4341 63127
rect 2763 63074 2805 63083
rect 2859 63104 2901 63113
rect 2859 63064 2860 63104
rect 2900 63064 2901 63104
rect 2859 63055 2901 63064
rect 3811 63104 3869 63105
rect 3811 63064 3820 63104
rect 3860 63064 3869 63104
rect 4299 63078 4300 63118
rect 4340 63078 4341 63118
rect 9195 63118 9237 63127
rect 4299 63069 4341 63078
rect 5923 63104 5981 63105
rect 3811 63063 3869 63064
rect 5923 63064 5932 63104
rect 5972 63064 5981 63104
rect 5923 63063 5981 63064
rect 7171 63104 7229 63105
rect 7171 63064 7180 63104
rect 7220 63064 7229 63104
rect 7171 63063 7229 63064
rect 7659 63104 7701 63113
rect 7659 63064 7660 63104
rect 7700 63064 7701 63104
rect 7659 63055 7701 63064
rect 7755 63104 7797 63113
rect 7755 63064 7756 63104
rect 7796 63064 7797 63104
rect 7755 63055 7797 63064
rect 8707 63104 8765 63105
rect 8707 63064 8716 63104
rect 8756 63064 8765 63104
rect 9195 63078 9196 63118
rect 9236 63078 9237 63118
rect 9195 63069 9237 63078
rect 9763 63104 9821 63105
rect 8707 63063 8765 63064
rect 9763 63064 9772 63104
rect 9812 63064 9821 63104
rect 9763 63063 9821 63064
rect 9867 63104 9909 63113
rect 9867 63064 9868 63104
rect 9908 63064 9909 63104
rect 9867 63055 9909 63064
rect 10059 63104 10101 63113
rect 10059 63064 10060 63104
rect 10100 63064 10101 63104
rect 10251 63106 10252 63146
rect 10292 63106 10293 63146
rect 11211 63148 11212 63188
rect 11252 63148 11253 63188
rect 11211 63139 11253 63148
rect 10251 63097 10293 63106
rect 10347 63104 10389 63113
rect 10059 63055 10101 63064
rect 10347 63064 10348 63104
rect 10388 63064 10389 63104
rect 10347 63055 10389 63064
rect 10443 63104 10485 63113
rect 10443 63064 10444 63104
rect 10484 63064 10485 63104
rect 10443 63055 10485 63064
rect 10539 63104 10581 63113
rect 10539 63064 10540 63104
rect 10580 63064 10581 63104
rect 10539 63055 10581 63064
rect 10731 63104 10773 63113
rect 10731 63064 10732 63104
rect 10772 63064 10773 63104
rect 10731 63055 10773 63064
rect 10923 63104 10965 63113
rect 10923 63064 10924 63104
rect 10964 63064 10965 63104
rect 10923 63055 10965 63064
rect 11107 63104 11165 63105
rect 11107 63064 11116 63104
rect 11156 63064 11165 63104
rect 11107 63063 11165 63064
rect 12555 63104 12597 63113
rect 12555 63064 12556 63104
rect 12596 63064 12597 63104
rect 12555 63055 12597 63064
rect 12651 63104 12693 63113
rect 12651 63064 12652 63104
rect 12692 63064 12693 63104
rect 12651 63055 12693 63064
rect 13219 63104 13277 63105
rect 13219 63064 13228 63104
rect 13268 63064 13277 63104
rect 13219 63063 13277 63064
rect 14467 63104 14525 63105
rect 14467 63064 14476 63104
rect 14516 63064 14525 63104
rect 14467 63063 14525 63064
rect 15043 63104 15101 63105
rect 15043 63064 15052 63104
rect 15092 63064 15101 63104
rect 15043 63063 15101 63064
rect 16291 63104 16349 63105
rect 16291 63064 16300 63104
rect 16340 63064 16349 63104
rect 16291 63063 16349 63064
rect 16483 63104 16541 63105
rect 16483 63064 16492 63104
rect 16532 63064 16541 63104
rect 16483 63063 16541 63064
rect 17731 63104 17789 63105
rect 17731 63064 17740 63104
rect 17780 63064 17789 63104
rect 17731 63063 17789 63064
rect 18123 63104 18165 63113
rect 18123 63064 18124 63104
rect 18164 63064 18165 63104
rect 18123 63055 18165 63064
rect 18219 63104 18261 63113
rect 18219 63064 18220 63104
rect 18260 63064 18261 63104
rect 18219 63055 18261 63064
rect 18411 63104 18453 63113
rect 18411 63064 18412 63104
rect 18452 63064 18453 63104
rect 18411 63055 18453 63064
rect 4491 63020 4533 63029
rect 4491 62980 4492 63020
rect 4532 62980 4533 63020
rect 4491 62971 4533 62980
rect 7371 63020 7413 63029
rect 7371 62980 7372 63020
rect 7412 62980 7413 63020
rect 7371 62971 7413 62980
rect 9387 63020 9429 63029
rect 9387 62980 9388 63020
rect 9428 62980 9429 63020
rect 9387 62971 9429 62980
rect 9963 63020 10005 63029
rect 9963 62980 9964 63020
rect 10004 62980 10005 63020
rect 9963 62971 10005 62980
rect 10827 63020 10869 63029
rect 10827 62980 10828 63020
rect 10868 62980 10869 63020
rect 10827 62971 10869 62980
rect 12835 62936 12893 62937
rect 12835 62896 12844 62936
rect 12884 62896 12893 62936
rect 12835 62895 12893 62896
rect 14667 62936 14709 62945
rect 14667 62896 14668 62936
rect 14708 62896 14709 62936
rect 14667 62887 14709 62896
rect 14859 62936 14901 62945
rect 14859 62896 14860 62936
rect 14900 62896 14901 62936
rect 14859 62887 14901 62896
rect 1152 62768 20452 62792
rect 1152 62728 4928 62768
rect 4968 62728 5010 62768
rect 5050 62728 5092 62768
rect 5132 62728 5174 62768
rect 5214 62728 5256 62768
rect 5296 62728 20048 62768
rect 20088 62728 20130 62768
rect 20170 62728 20212 62768
rect 20252 62728 20294 62768
rect 20334 62728 20376 62768
rect 20416 62728 20452 62768
rect 1152 62704 20452 62728
rect 9379 62600 9437 62601
rect 9379 62560 9388 62600
rect 9428 62560 9437 62600
rect 9379 62559 9437 62560
rect 9859 62600 9917 62601
rect 9859 62560 9868 62600
rect 9908 62560 9917 62600
rect 9859 62559 9917 62560
rect 13707 62600 13749 62609
rect 13707 62560 13708 62600
rect 13748 62560 13749 62600
rect 13707 62551 13749 62560
rect 15043 62600 15101 62601
rect 15043 62560 15052 62600
rect 15092 62560 15101 62600
rect 15043 62559 15101 62560
rect 15715 62600 15773 62601
rect 15715 62560 15724 62600
rect 15764 62560 15773 62600
rect 15715 62559 15773 62560
rect 17931 62600 17973 62609
rect 17931 62560 17932 62600
rect 17972 62560 17973 62600
rect 17931 62551 17973 62560
rect 1699 62432 1757 62433
rect 1699 62392 1708 62432
rect 1748 62392 1757 62432
rect 1699 62391 1757 62392
rect 2947 62432 3005 62433
rect 2947 62392 2956 62432
rect 2996 62392 3005 62432
rect 2947 62391 3005 62392
rect 4195 62432 4253 62433
rect 4195 62392 4204 62432
rect 4244 62392 4253 62432
rect 4195 62391 4253 62392
rect 5443 62432 5501 62433
rect 5443 62392 5452 62432
rect 5492 62392 5501 62432
rect 5443 62391 5501 62392
rect 5827 62432 5885 62433
rect 5827 62392 5836 62432
rect 5876 62392 5885 62432
rect 5827 62391 5885 62392
rect 7075 62432 7133 62433
rect 7075 62392 7084 62432
rect 7124 62392 7133 62432
rect 7075 62391 7133 62392
rect 7459 62432 7517 62433
rect 7459 62392 7468 62432
rect 7508 62392 7517 62432
rect 7459 62391 7517 62392
rect 8707 62432 8765 62433
rect 8707 62392 8716 62432
rect 8756 62392 8765 62432
rect 8707 62391 8765 62392
rect 9099 62432 9141 62441
rect 9099 62392 9100 62432
rect 9140 62392 9141 62432
rect 9099 62383 9141 62392
rect 9195 62432 9237 62441
rect 9195 62392 9196 62432
rect 9236 62392 9237 62432
rect 9195 62383 9237 62392
rect 9291 62432 9333 62441
rect 9291 62392 9292 62432
rect 9332 62392 9333 62432
rect 9291 62383 9333 62392
rect 9579 62432 9621 62441
rect 9579 62392 9580 62432
rect 9620 62392 9621 62432
rect 9579 62383 9621 62392
rect 9675 62432 9717 62441
rect 9675 62392 9676 62432
rect 9716 62392 9717 62432
rect 9675 62383 9717 62392
rect 9771 62432 9813 62441
rect 9771 62392 9772 62432
rect 9812 62392 9813 62432
rect 9771 62383 9813 62392
rect 10243 62432 10301 62433
rect 10243 62392 10252 62432
rect 10292 62392 10301 62432
rect 10243 62391 10301 62392
rect 11491 62432 11549 62433
rect 11491 62392 11500 62432
rect 11540 62392 11549 62432
rect 11491 62391 11549 62392
rect 11979 62432 12021 62441
rect 11979 62392 11980 62432
rect 12020 62392 12021 62432
rect 11979 62383 12021 62392
rect 12075 62432 12117 62441
rect 12075 62392 12076 62432
rect 12116 62392 12117 62432
rect 12075 62383 12117 62392
rect 12459 62432 12501 62441
rect 12459 62392 12460 62432
rect 12500 62392 12501 62432
rect 12459 62383 12501 62392
rect 13027 62432 13085 62433
rect 13027 62392 13036 62432
rect 13076 62392 13085 62432
rect 14763 62432 14805 62441
rect 13027 62391 13085 62392
rect 13515 62418 13557 62427
rect 13515 62378 13516 62418
rect 13556 62378 13557 62418
rect 14763 62392 14764 62432
rect 14804 62392 14805 62432
rect 14763 62383 14805 62392
rect 14859 62432 14901 62441
rect 14859 62392 14860 62432
rect 14900 62392 14901 62432
rect 14859 62383 14901 62392
rect 14955 62432 14997 62441
rect 14955 62392 14956 62432
rect 14996 62392 14997 62432
rect 14955 62383 14997 62392
rect 15243 62432 15285 62441
rect 15243 62392 15244 62432
rect 15284 62392 15285 62432
rect 15243 62383 15285 62392
rect 15339 62432 15381 62441
rect 15339 62392 15340 62432
rect 15380 62392 15381 62432
rect 15339 62383 15381 62392
rect 15435 62432 15477 62441
rect 15435 62392 15436 62432
rect 15476 62392 15477 62432
rect 15435 62383 15477 62392
rect 15531 62432 15573 62441
rect 15531 62392 15532 62432
rect 15572 62392 15573 62432
rect 15531 62383 15573 62392
rect 15811 62432 15869 62433
rect 15811 62392 15820 62432
rect 15860 62392 15869 62432
rect 15811 62391 15869 62392
rect 16483 62432 16541 62433
rect 16483 62392 16492 62432
rect 16532 62392 16541 62432
rect 16483 62391 16541 62392
rect 17731 62432 17789 62433
rect 17731 62392 17740 62432
rect 17780 62392 17789 62432
rect 17731 62391 17789 62392
rect 13515 62369 13557 62378
rect 12555 62348 12597 62357
rect 12555 62308 12556 62348
rect 12596 62308 12597 62348
rect 12555 62299 12597 62308
rect 11691 62264 11733 62273
rect 11691 62224 11692 62264
rect 11732 62224 11733 62264
rect 11691 62215 11733 62224
rect 3147 62180 3189 62189
rect 3147 62140 3148 62180
rect 3188 62140 3189 62180
rect 3147 62131 3189 62140
rect 5643 62180 5685 62189
rect 5643 62140 5644 62180
rect 5684 62140 5685 62180
rect 5643 62131 5685 62140
rect 7275 62180 7317 62189
rect 7275 62140 7276 62180
rect 7316 62140 7317 62180
rect 7275 62131 7317 62140
rect 8907 62180 8949 62189
rect 8907 62140 8908 62180
rect 8948 62140 8949 62180
rect 8907 62131 8949 62140
rect 16003 62180 16061 62181
rect 16003 62140 16012 62180
rect 16052 62140 16061 62180
rect 16003 62139 16061 62140
rect 1152 62012 20352 62036
rect 1152 61972 3688 62012
rect 3728 61972 3770 62012
rect 3810 61972 3852 62012
rect 3892 61972 3934 62012
rect 3974 61972 4016 62012
rect 4056 61972 18808 62012
rect 18848 61972 18890 62012
rect 18930 61972 18972 62012
rect 19012 61972 19054 62012
rect 19094 61972 19136 62012
rect 19176 61972 20352 62012
rect 1152 61948 20352 61972
rect 13611 61844 13653 61853
rect 13611 61804 13612 61844
rect 13652 61804 13653 61844
rect 13611 61795 13653 61804
rect 2667 61676 2709 61685
rect 2667 61636 2668 61676
rect 2708 61636 2709 61676
rect 2667 61627 2709 61636
rect 6219 61676 6261 61685
rect 6219 61636 6220 61676
rect 6260 61636 6261 61676
rect 6219 61627 6261 61636
rect 3723 61606 3765 61615
rect 2187 61592 2229 61601
rect 2187 61552 2188 61592
rect 2228 61552 2229 61592
rect 2187 61543 2229 61552
rect 2283 61592 2325 61601
rect 2283 61552 2284 61592
rect 2324 61552 2325 61592
rect 2283 61543 2325 61552
rect 2763 61592 2805 61601
rect 2763 61552 2764 61592
rect 2804 61552 2805 61592
rect 2763 61543 2805 61552
rect 3235 61592 3293 61593
rect 3235 61552 3244 61592
rect 3284 61552 3293 61592
rect 3723 61566 3724 61606
rect 3764 61566 3765 61606
rect 7179 61606 7221 61615
rect 3723 61557 3765 61566
rect 5643 61592 5685 61601
rect 3235 61551 3293 61552
rect 5643 61552 5644 61592
rect 5684 61552 5685 61592
rect 5643 61543 5685 61552
rect 5739 61592 5781 61601
rect 5739 61552 5740 61592
rect 5780 61552 5781 61592
rect 5739 61543 5781 61552
rect 6123 61592 6165 61601
rect 6123 61552 6124 61592
rect 6164 61552 6165 61592
rect 6123 61543 6165 61552
rect 6691 61592 6749 61593
rect 6691 61552 6700 61592
rect 6740 61552 6749 61592
rect 7179 61566 7180 61606
rect 7220 61566 7221 61606
rect 7179 61557 7221 61566
rect 7747 61592 7805 61593
rect 6691 61551 6749 61552
rect 7747 61552 7756 61592
rect 7796 61552 7805 61592
rect 7747 61551 7805 61552
rect 8995 61592 9053 61593
rect 8995 61552 9004 61592
rect 9044 61552 9053 61592
rect 8995 61551 9053 61552
rect 9667 61592 9725 61593
rect 9667 61552 9676 61592
rect 9716 61552 9725 61592
rect 9667 61551 9725 61552
rect 10915 61592 10973 61593
rect 10915 61552 10924 61592
rect 10964 61552 10973 61592
rect 10915 61551 10973 61552
rect 12163 61592 12221 61593
rect 12163 61552 12172 61592
rect 12212 61552 12221 61592
rect 12163 61551 12221 61552
rect 13411 61592 13469 61593
rect 13411 61552 13420 61592
rect 13460 61552 13469 61592
rect 13411 61551 13469 61552
rect 14379 61592 14421 61601
rect 14379 61552 14380 61592
rect 14420 61552 14421 61592
rect 14379 61543 14421 61552
rect 14571 61592 14613 61601
rect 14571 61552 14572 61592
rect 14612 61552 14613 61592
rect 14571 61543 14613 61552
rect 14763 61592 14805 61601
rect 14763 61552 14764 61592
rect 14804 61552 14805 61592
rect 14763 61543 14805 61552
rect 14859 61592 14901 61601
rect 14859 61552 14860 61592
rect 14900 61552 14901 61592
rect 15907 61592 15965 61593
rect 14859 61543 14901 61552
rect 15243 61571 15285 61580
rect 15243 61531 15244 61571
rect 15284 61531 15285 61571
rect 15243 61522 15285 61531
rect 15339 61571 15381 61580
rect 15339 61531 15340 61571
rect 15380 61531 15381 61571
rect 15339 61522 15381 61531
rect 15435 61571 15477 61580
rect 15435 61531 15436 61571
rect 15476 61531 15477 61571
rect 15907 61552 15916 61592
rect 15956 61552 15965 61592
rect 15907 61551 15965 61552
rect 17155 61592 17213 61593
rect 17155 61552 17164 61592
rect 17204 61552 17213 61592
rect 17155 61551 17213 61552
rect 15435 61522 15477 61531
rect 3915 61508 3957 61517
rect 3915 61468 3916 61508
rect 3956 61468 3957 61508
rect 3915 61459 3957 61468
rect 7563 61508 7605 61517
rect 7563 61468 7564 61508
rect 7604 61468 7605 61508
rect 7563 61459 7605 61468
rect 7371 61424 7413 61433
rect 7371 61384 7372 61424
rect 7412 61384 7413 61424
rect 7371 61375 7413 61384
rect 11115 61424 11157 61433
rect 11115 61384 11116 61424
rect 11156 61384 11157 61424
rect 11115 61375 11157 61384
rect 14475 61424 14517 61433
rect 14475 61384 14476 61424
rect 14516 61384 14517 61424
rect 14475 61375 14517 61384
rect 15043 61424 15101 61425
rect 15043 61384 15052 61424
rect 15092 61384 15101 61424
rect 15043 61383 15101 61384
rect 15523 61424 15581 61425
rect 15523 61384 15532 61424
rect 15572 61384 15581 61424
rect 15523 61383 15581 61384
rect 15723 61424 15765 61433
rect 15723 61384 15724 61424
rect 15764 61384 15765 61424
rect 15723 61375 15765 61384
rect 1152 61256 20452 61280
rect 1152 61216 4928 61256
rect 4968 61216 5010 61256
rect 5050 61216 5092 61256
rect 5132 61216 5174 61256
rect 5214 61216 5256 61256
rect 5296 61216 20048 61256
rect 20088 61216 20130 61256
rect 20170 61216 20212 61256
rect 20252 61216 20294 61256
rect 20334 61216 20376 61256
rect 20416 61216 20452 61256
rect 1152 61192 20452 61216
rect 10923 61088 10965 61097
rect 10923 61048 10924 61088
rect 10964 61048 10965 61088
rect 10923 61039 10965 61048
rect 15627 61088 15669 61097
rect 15627 61048 15628 61088
rect 15668 61048 15669 61088
rect 15627 61039 15669 61048
rect 4587 61004 4629 61013
rect 4587 60964 4588 61004
rect 4628 60964 4629 61004
rect 4587 60955 4629 60964
rect 6795 61004 6837 61013
rect 6795 60964 6796 61004
rect 6836 60964 6837 61004
rect 6795 60955 6837 60964
rect 8907 61004 8949 61013
rect 8907 60964 8908 61004
rect 8948 60964 8949 61004
rect 8907 60955 8949 60964
rect 2859 60920 2901 60929
rect 2859 60880 2860 60920
rect 2900 60880 2901 60920
rect 2859 60871 2901 60880
rect 2955 60920 2997 60929
rect 2955 60880 2956 60920
rect 2996 60880 2997 60920
rect 2955 60871 2997 60880
rect 3435 60920 3477 60929
rect 3435 60880 3436 60920
rect 3476 60880 3477 60920
rect 3435 60871 3477 60880
rect 3907 60920 3965 60921
rect 3907 60880 3916 60920
rect 3956 60880 3965 60920
rect 5059 60920 5117 60921
rect 3907 60879 3965 60880
rect 4443 60910 4485 60919
rect 4443 60870 4444 60910
rect 4484 60870 4485 60910
rect 5059 60880 5068 60920
rect 5108 60880 5117 60920
rect 5059 60879 5117 60880
rect 5347 60920 5405 60921
rect 5347 60880 5356 60920
rect 5396 60880 5405 60920
rect 5347 60879 5405 60880
rect 6595 60920 6653 60921
rect 6595 60880 6604 60920
rect 6644 60880 6653 60920
rect 6595 60879 6653 60880
rect 6987 60920 7029 60929
rect 6987 60880 6988 60920
rect 7028 60880 7029 60920
rect 6987 60871 7029 60880
rect 7179 60920 7221 60929
rect 7179 60880 7180 60920
rect 7220 60880 7221 60920
rect 7179 60871 7221 60880
rect 7275 60920 7317 60929
rect 7275 60880 7276 60920
rect 7316 60880 7317 60920
rect 7275 60871 7317 60880
rect 7459 60920 7517 60921
rect 7459 60880 7468 60920
rect 7508 60880 7517 60920
rect 7459 60879 7517 60880
rect 8707 60920 8765 60921
rect 8707 60880 8716 60920
rect 8756 60880 8765 60920
rect 8707 60879 8765 60880
rect 9195 60920 9237 60929
rect 9195 60880 9196 60920
rect 9236 60880 9237 60920
rect 9195 60871 9237 60880
rect 9291 60920 9333 60929
rect 9291 60880 9292 60920
rect 9332 60880 9333 60920
rect 9291 60871 9333 60880
rect 9675 60920 9717 60929
rect 9675 60880 9676 60920
rect 9716 60880 9717 60920
rect 9675 60871 9717 60880
rect 10243 60920 10301 60921
rect 10243 60880 10252 60920
rect 10292 60880 10301 60920
rect 11107 60920 11165 60921
rect 10243 60879 10301 60880
rect 10779 60910 10821 60919
rect 4443 60861 4485 60870
rect 10779 60870 10780 60910
rect 10820 60870 10821 60910
rect 11107 60880 11116 60920
rect 11156 60880 11165 60920
rect 12747 60920 12789 60929
rect 11107 60879 11165 60880
rect 12355 60899 12413 60900
rect 10779 60861 10821 60870
rect 12355 60859 12364 60899
rect 12404 60859 12413 60899
rect 12747 60880 12748 60920
rect 12788 60880 12789 60920
rect 12747 60871 12789 60880
rect 12843 60920 12885 60929
rect 12843 60880 12844 60920
rect 12884 60880 12885 60920
rect 12843 60871 12885 60880
rect 13035 60920 13077 60929
rect 13035 60880 13036 60920
rect 13076 60880 13077 60920
rect 13035 60871 13077 60880
rect 13899 60920 13941 60929
rect 13899 60880 13900 60920
rect 13940 60880 13941 60920
rect 13899 60871 13941 60880
rect 13995 60920 14037 60929
rect 13995 60880 13996 60920
rect 14036 60880 14037 60920
rect 13995 60871 14037 60880
rect 14379 60920 14421 60929
rect 14379 60880 14380 60920
rect 14420 60880 14421 60920
rect 14379 60871 14421 60880
rect 14947 60920 15005 60921
rect 14947 60880 14956 60920
rect 14996 60880 15005 60920
rect 15819 60920 15861 60929
rect 14947 60879 15005 60880
rect 15435 60906 15477 60915
rect 12355 60858 12413 60859
rect 15435 60866 15436 60906
rect 15476 60866 15477 60906
rect 15819 60880 15820 60920
rect 15860 60880 15861 60920
rect 15819 60871 15861 60880
rect 16011 60920 16053 60929
rect 16011 60880 16012 60920
rect 16052 60880 16053 60920
rect 16011 60871 16053 60880
rect 16099 60920 16157 60921
rect 16099 60880 16108 60920
rect 16148 60880 16157 60920
rect 16099 60879 16157 60880
rect 16387 60920 16445 60921
rect 16387 60880 16396 60920
rect 16436 60880 16445 60920
rect 16387 60879 16445 60880
rect 17635 60920 17693 60921
rect 17635 60880 17644 60920
rect 17684 60880 17693 60920
rect 17635 60879 17693 60880
rect 18211 60920 18269 60921
rect 18211 60880 18220 60920
rect 18260 60880 18269 60920
rect 18211 60879 18269 60880
rect 19459 60920 19517 60921
rect 19459 60880 19468 60920
rect 19508 60880 19517 60920
rect 19459 60879 19517 60880
rect 15435 60857 15477 60866
rect 3339 60836 3381 60845
rect 3339 60796 3340 60836
rect 3380 60796 3381 60836
rect 3339 60787 3381 60796
rect 9771 60836 9813 60845
rect 9771 60796 9772 60836
rect 9812 60796 9813 60836
rect 9771 60787 9813 60796
rect 14475 60836 14517 60845
rect 14475 60796 14476 60836
rect 14516 60796 14517 60836
rect 14475 60787 14517 60796
rect 7267 60752 7325 60753
rect 7267 60712 7276 60752
rect 7316 60712 7325 60752
rect 7267 60711 7325 60712
rect 12939 60752 12981 60761
rect 12939 60712 12940 60752
rect 12980 60712 12981 60752
rect 12939 60703 12981 60712
rect 5163 60668 5205 60677
rect 5163 60628 5164 60668
rect 5204 60628 5205 60668
rect 5163 60619 5205 60628
rect 12555 60668 12597 60677
rect 12555 60628 12556 60668
rect 12596 60628 12597 60668
rect 12555 60619 12597 60628
rect 15819 60668 15861 60677
rect 15819 60628 15820 60668
rect 15860 60628 15861 60668
rect 15819 60619 15861 60628
rect 17835 60668 17877 60677
rect 17835 60628 17836 60668
rect 17876 60628 17877 60668
rect 17835 60619 17877 60628
rect 19659 60668 19701 60677
rect 19659 60628 19660 60668
rect 19700 60628 19701 60668
rect 19659 60619 19701 60628
rect 1152 60500 20352 60524
rect 1152 60460 3688 60500
rect 3728 60460 3770 60500
rect 3810 60460 3852 60500
rect 3892 60460 3934 60500
rect 3974 60460 4016 60500
rect 4056 60460 18808 60500
rect 18848 60460 18890 60500
rect 18930 60460 18972 60500
rect 19012 60460 19054 60500
rect 19094 60460 19136 60500
rect 19176 60460 20352 60500
rect 1152 60436 20352 60460
rect 14187 60332 14229 60341
rect 14187 60292 14188 60332
rect 14228 60292 14229 60332
rect 14187 60283 14229 60292
rect 9675 60164 9717 60173
rect 9675 60124 9676 60164
rect 9716 60124 9717 60164
rect 9675 60115 9717 60124
rect 9771 60164 9813 60173
rect 9771 60124 9772 60164
rect 9812 60124 9813 60164
rect 9771 60115 9813 60124
rect 10731 60089 10773 60098
rect 19083 60094 19125 60103
rect 1411 60080 1469 60081
rect 1411 60040 1420 60080
rect 1460 60040 1469 60080
rect 1411 60039 1469 60040
rect 2659 60080 2717 60081
rect 2659 60040 2668 60080
rect 2708 60040 2717 60080
rect 2659 60039 2717 60040
rect 4291 60080 4349 60081
rect 4291 60040 4300 60080
rect 4340 60040 4349 60080
rect 4291 60039 4349 60040
rect 5347 60080 5405 60081
rect 5347 60040 5356 60080
rect 5396 60040 5405 60080
rect 5347 60039 5405 60040
rect 6595 60080 6653 60081
rect 6595 60040 6604 60080
rect 6644 60040 6653 60080
rect 6595 60039 6653 60040
rect 6987 60080 7029 60089
rect 6987 60040 6988 60080
rect 7028 60040 7029 60080
rect 3043 60038 3101 60039
rect 3043 59998 3052 60038
rect 3092 59998 3101 60038
rect 6987 60031 7029 60040
rect 7083 60080 7125 60089
rect 7083 60040 7084 60080
rect 7124 60040 7125 60080
rect 7083 60031 7125 60040
rect 7459 60080 7517 60081
rect 7459 60040 7468 60080
rect 7508 60040 7517 60080
rect 7459 60039 7517 60040
rect 8707 60080 8765 60081
rect 8707 60040 8716 60080
rect 8756 60040 8765 60080
rect 8707 60039 8765 60040
rect 9195 60080 9237 60089
rect 9195 60040 9196 60080
rect 9236 60040 9237 60080
rect 9195 60031 9237 60040
rect 9291 60080 9333 60089
rect 9291 60040 9292 60080
rect 9332 60040 9333 60080
rect 9291 60031 9333 60040
rect 10243 60080 10301 60081
rect 10243 60040 10252 60080
rect 10292 60040 10301 60080
rect 10731 60049 10732 60089
rect 10772 60049 10773 60089
rect 10731 60040 10773 60049
rect 11875 60080 11933 60081
rect 11875 60040 11884 60080
rect 11924 60040 11933 60080
rect 10243 60039 10301 60040
rect 11875 60039 11933 60040
rect 12267 60080 12309 60089
rect 12267 60040 12268 60080
rect 12308 60040 12309 60080
rect 12267 60031 12309 60040
rect 12363 60080 12405 60089
rect 12363 60040 12364 60080
rect 12404 60040 12405 60080
rect 12363 60031 12405 60040
rect 12747 60080 12789 60089
rect 12747 60040 12748 60080
rect 12788 60040 12789 60080
rect 12747 60031 12789 60040
rect 12843 60080 12885 60089
rect 13803 60085 13845 60094
rect 12843 60040 12844 60080
rect 12884 60040 12885 60080
rect 12843 60031 12885 60040
rect 13315 60080 13373 60081
rect 13315 60040 13324 60080
rect 13364 60040 13373 60080
rect 13315 60039 13373 60040
rect 13803 60045 13804 60085
rect 13844 60045 13845 60085
rect 13803 60036 13845 60045
rect 14371 60080 14429 60081
rect 14371 60040 14380 60080
rect 14420 60040 14429 60080
rect 14371 60039 14429 60040
rect 15619 60080 15677 60081
rect 15619 60040 15628 60080
rect 15668 60040 15677 60080
rect 15619 60039 15677 60040
rect 15811 60080 15869 60081
rect 15811 60040 15820 60080
rect 15860 60040 15869 60080
rect 15811 60039 15869 60040
rect 17059 60080 17117 60081
rect 17059 60040 17068 60080
rect 17108 60040 17117 60080
rect 17059 60039 17117 60040
rect 17547 60080 17589 60089
rect 17547 60040 17548 60080
rect 17588 60040 17589 60080
rect 17547 60031 17589 60040
rect 17643 60080 17685 60089
rect 17643 60040 17644 60080
rect 17684 60040 17685 60080
rect 17643 60031 17685 60040
rect 18027 60080 18069 60089
rect 18027 60040 18028 60080
rect 18068 60040 18069 60080
rect 18027 60031 18069 60040
rect 18123 60080 18165 60089
rect 18123 60040 18124 60080
rect 18164 60040 18165 60080
rect 18123 60031 18165 60040
rect 18595 60080 18653 60081
rect 18595 60040 18604 60080
rect 18644 60040 18653 60080
rect 19083 60054 19084 60094
rect 19124 60054 19125 60094
rect 19083 60045 19125 60054
rect 18595 60039 18653 60040
rect 3043 59997 3101 59998
rect 6795 59996 6837 60005
rect 6795 59956 6796 59996
rect 6836 59956 6837 59996
rect 6795 59947 6837 59956
rect 8907 59996 8949 60005
rect 8907 59956 8908 59996
rect 8948 59956 8949 59996
rect 8907 59947 8949 59956
rect 2859 59912 2901 59921
rect 2859 59872 2860 59912
rect 2900 59872 2901 59912
rect 2859 59863 2901 59872
rect 4491 59912 4533 59921
rect 4491 59872 4492 59912
rect 4532 59872 4533 59912
rect 4491 59863 4533 59872
rect 7267 59912 7325 59913
rect 7267 59872 7276 59912
rect 7316 59872 7325 59912
rect 7267 59871 7325 59872
rect 10923 59912 10965 59921
rect 10923 59872 10924 59912
rect 10964 59872 10965 59912
rect 10923 59863 10965 59872
rect 11979 59912 12021 59921
rect 11979 59872 11980 59912
rect 12020 59872 12021 59912
rect 11979 59863 12021 59872
rect 13995 59912 14037 59921
rect 13995 59872 13996 59912
rect 14036 59872 14037 59912
rect 13995 59863 14037 59872
rect 17259 59912 17301 59921
rect 17259 59872 17260 59912
rect 17300 59872 17301 59912
rect 17259 59863 17301 59872
rect 19275 59912 19317 59921
rect 19275 59872 19276 59912
rect 19316 59872 19317 59912
rect 19275 59863 19317 59872
rect 1152 59744 20452 59768
rect 1152 59704 4928 59744
rect 4968 59704 5010 59744
rect 5050 59704 5092 59744
rect 5132 59704 5174 59744
rect 5214 59704 5256 59744
rect 5296 59704 20048 59744
rect 20088 59704 20130 59744
rect 20170 59704 20212 59744
rect 20252 59704 20294 59744
rect 20334 59704 20376 59744
rect 20416 59704 20452 59744
rect 1152 59680 20452 59704
rect 10923 59576 10965 59585
rect 10923 59536 10924 59576
rect 10964 59536 10965 59576
rect 10923 59527 10965 59536
rect 12747 59576 12789 59585
rect 12747 59536 12748 59576
rect 12788 59536 12789 59576
rect 12747 59527 12789 59536
rect 14379 59576 14421 59585
rect 14379 59536 14380 59576
rect 14420 59536 14421 59576
rect 14379 59527 14421 59536
rect 14571 59576 14613 59585
rect 14571 59536 14572 59576
rect 14612 59536 14613 59576
rect 14571 59527 14613 59536
rect 4299 59492 4341 59501
rect 4299 59452 4300 59492
rect 4340 59452 4341 59492
rect 4299 59443 4341 59452
rect 17155 59492 17213 59493
rect 17155 59452 17164 59492
rect 17204 59452 17213 59492
rect 17155 59451 17213 59452
rect 19275 59492 19317 59501
rect 19275 59452 19276 59492
rect 19316 59452 19317 59492
rect 19275 59443 19317 59452
rect 2571 59408 2613 59417
rect 2571 59368 2572 59408
rect 2612 59368 2613 59408
rect 2571 59359 2613 59368
rect 2667 59408 2709 59417
rect 2667 59368 2668 59408
rect 2708 59368 2709 59408
rect 2667 59359 2709 59368
rect 3051 59408 3093 59417
rect 3051 59368 3052 59408
rect 3092 59368 3093 59408
rect 3051 59359 3093 59368
rect 3147 59408 3189 59417
rect 3147 59368 3148 59408
rect 3188 59368 3189 59408
rect 3147 59359 3189 59368
rect 3619 59408 3677 59409
rect 3619 59368 3628 59408
rect 3668 59368 3677 59408
rect 5155 59408 5213 59409
rect 3619 59367 3677 59368
rect 4155 59398 4197 59407
rect 4155 59358 4156 59398
rect 4196 59358 4197 59398
rect 5155 59368 5164 59408
rect 5204 59368 5213 59408
rect 5155 59367 5213 59368
rect 6403 59408 6461 59409
rect 6403 59368 6412 59408
rect 6452 59368 6461 59408
rect 6403 59367 6461 59368
rect 6787 59408 6845 59409
rect 6787 59368 6796 59408
rect 6836 59368 6845 59408
rect 6787 59367 6845 59368
rect 8035 59408 8093 59409
rect 8035 59368 8044 59408
rect 8084 59368 8093 59408
rect 8035 59367 8093 59368
rect 8419 59408 8477 59409
rect 8419 59368 8428 59408
rect 8468 59368 8477 59408
rect 8419 59367 8477 59368
rect 8515 59408 8573 59409
rect 8515 59368 8524 59408
rect 8564 59368 8573 59408
rect 8515 59367 8573 59368
rect 8715 59408 8757 59417
rect 8715 59368 8716 59408
rect 8756 59368 8757 59408
rect 8715 59359 8757 59368
rect 8811 59408 8853 59417
rect 8811 59368 8812 59408
rect 8852 59368 8853 59408
rect 8811 59359 8853 59368
rect 8904 59408 8962 59409
rect 8904 59368 8913 59408
rect 8953 59368 8962 59408
rect 8904 59367 8962 59368
rect 9475 59408 9533 59409
rect 9475 59368 9484 59408
rect 9524 59368 9533 59408
rect 9475 59367 9533 59368
rect 10723 59408 10781 59409
rect 10723 59368 10732 59408
rect 10772 59368 10781 59408
rect 10723 59367 10781 59368
rect 11299 59408 11357 59409
rect 11299 59368 11308 59408
rect 11348 59368 11357 59408
rect 11299 59367 11357 59368
rect 12547 59408 12605 59409
rect 12547 59368 12556 59408
rect 12596 59368 12605 59408
rect 12547 59367 12605 59368
rect 12931 59408 12989 59409
rect 12931 59368 12940 59408
rect 12980 59368 12989 59408
rect 12931 59367 12989 59368
rect 14179 59408 14237 59409
rect 14179 59368 14188 59408
rect 14228 59368 14237 59408
rect 14179 59367 14237 59368
rect 14755 59408 14813 59409
rect 14755 59368 14764 59408
rect 14804 59368 14813 59408
rect 14755 59367 14813 59368
rect 16003 59408 16061 59409
rect 16003 59368 16012 59408
rect 16052 59368 16061 59408
rect 16003 59367 16061 59368
rect 16291 59408 16349 59409
rect 16291 59368 16300 59408
rect 16340 59368 16349 59408
rect 16291 59367 16349 59368
rect 17547 59408 17589 59417
rect 17547 59368 17548 59408
rect 17588 59368 17589 59408
rect 17547 59359 17589 59368
rect 17643 59408 17685 59417
rect 17643 59368 17644 59408
rect 17684 59368 17685 59408
rect 17643 59359 17685 59368
rect 18595 59408 18653 59409
rect 18595 59368 18604 59408
rect 18644 59368 18653 59408
rect 18595 59367 18653 59368
rect 19083 59394 19125 59403
rect 4155 59349 4197 59358
rect 19083 59354 19084 59394
rect 19124 59354 19125 59394
rect 19083 59345 19125 59354
rect 2083 59324 2141 59325
rect 2083 59284 2092 59324
rect 2132 59284 2141 59324
rect 2083 59283 2141 59284
rect 18027 59324 18069 59333
rect 18027 59284 18028 59324
rect 18068 59284 18069 59324
rect 18027 59275 18069 59284
rect 18123 59324 18165 59333
rect 18123 59284 18124 59324
rect 18164 59284 18165 59324
rect 18123 59275 18165 59284
rect 1899 59156 1941 59165
rect 1899 59116 1900 59156
rect 1940 59116 1941 59156
rect 1899 59107 1941 59116
rect 6603 59156 6645 59165
rect 6603 59116 6604 59156
rect 6644 59116 6645 59156
rect 6603 59107 6645 59116
rect 8235 59156 8277 59165
rect 8235 59116 8236 59156
rect 8276 59116 8277 59156
rect 8235 59107 8277 59116
rect 8427 59156 8469 59165
rect 8427 59116 8428 59156
rect 8468 59116 8469 59156
rect 8427 59107 8469 59116
rect 12747 59156 12789 59165
rect 12747 59116 12748 59156
rect 12788 59116 12789 59156
rect 12747 59107 12789 59116
rect 16971 59156 17013 59165
rect 16971 59116 16972 59156
rect 17012 59116 17013 59156
rect 16971 59107 17013 59116
rect 1152 58988 20352 59012
rect 1152 58948 3688 58988
rect 3728 58948 3770 58988
rect 3810 58948 3852 58988
rect 3892 58948 3934 58988
rect 3974 58948 4016 58988
rect 4056 58948 18808 58988
rect 18848 58948 18890 58988
rect 18930 58948 18972 58988
rect 19012 58948 19054 58988
rect 19094 58948 19136 58988
rect 19176 58948 20352 58988
rect 1152 58924 20352 58948
rect 19851 58820 19893 58829
rect 19851 58780 19852 58820
rect 19892 58780 19893 58820
rect 19851 58771 19893 58780
rect 12555 58736 12597 58745
rect 12555 58696 12556 58736
rect 12596 58696 12597 58736
rect 12555 58687 12597 58696
rect 15531 58736 15573 58745
rect 15531 58696 15532 58736
rect 15572 58696 15573 58736
rect 15531 58687 15573 58696
rect 1219 58568 1277 58569
rect 1219 58528 1228 58568
rect 1268 58528 1277 58568
rect 1219 58527 1277 58528
rect 2467 58568 2525 58569
rect 2467 58528 2476 58568
rect 2516 58528 2525 58568
rect 2467 58527 2525 58528
rect 3715 58568 3773 58569
rect 3715 58528 3724 58568
rect 3764 58528 3773 58568
rect 3715 58527 3773 58528
rect 4963 58568 5021 58569
rect 4963 58528 4972 58568
rect 5012 58528 5021 58568
rect 4963 58527 5021 58528
rect 5347 58568 5405 58569
rect 5347 58528 5356 58568
rect 5396 58528 5405 58568
rect 5347 58527 5405 58528
rect 6595 58568 6653 58569
rect 6595 58528 6604 58568
rect 6644 58528 6653 58568
rect 6595 58527 6653 58528
rect 7363 58568 7421 58569
rect 7363 58528 7372 58568
rect 7412 58528 7421 58568
rect 7363 58527 7421 58528
rect 8611 58568 8669 58569
rect 8611 58528 8620 58568
rect 8660 58528 8669 58568
rect 8611 58527 8669 58528
rect 8995 58568 9053 58569
rect 8995 58528 9004 58568
rect 9044 58528 9053 58568
rect 8995 58527 9053 58528
rect 10243 58568 10301 58569
rect 10243 58528 10252 58568
rect 10292 58528 10301 58568
rect 10243 58527 10301 58528
rect 11107 58568 11165 58569
rect 11107 58528 11116 58568
rect 11156 58528 11165 58568
rect 11107 58527 11165 58528
rect 12355 58568 12413 58569
rect 12355 58528 12364 58568
rect 12404 58528 12413 58568
rect 12355 58527 12413 58528
rect 12830 58568 12888 58569
rect 12830 58528 12839 58568
rect 12879 58528 12888 58568
rect 12830 58527 12888 58528
rect 12939 58568 12981 58577
rect 12939 58528 12940 58568
rect 12980 58528 12981 58568
rect 12939 58519 12981 58528
rect 13035 58568 13077 58577
rect 13035 58528 13036 58568
rect 13076 58528 13077 58568
rect 13035 58519 13077 58528
rect 13219 58568 13277 58569
rect 13219 58528 13228 58568
rect 13268 58528 13277 58568
rect 13219 58527 13277 58528
rect 13315 58568 13373 58569
rect 13315 58528 13324 58568
rect 13364 58528 13373 58568
rect 13315 58527 13373 58528
rect 13515 58568 13557 58577
rect 13515 58528 13516 58568
rect 13556 58528 13557 58568
rect 13515 58519 13557 58528
rect 13611 58568 13653 58577
rect 13611 58528 13612 58568
rect 13652 58528 13653 58568
rect 13611 58519 13653 58528
rect 14083 58568 14141 58569
rect 14083 58528 14092 58568
rect 14132 58528 14141 58568
rect 14083 58527 14141 58528
rect 15331 58568 15389 58569
rect 15331 58528 15340 58568
rect 15380 58528 15389 58568
rect 15331 58527 15389 58528
rect 16011 58568 16053 58577
rect 16011 58528 16012 58568
rect 16052 58528 16053 58568
rect 16011 58519 16053 58528
rect 16107 58568 16149 58577
rect 16107 58528 16108 58568
rect 16148 58528 16149 58568
rect 16107 58519 16149 58528
rect 16299 58568 16341 58577
rect 16299 58528 16300 58568
rect 16340 58528 16341 58568
rect 16299 58519 16341 58528
rect 16395 58568 16437 58577
rect 16395 58528 16396 58568
rect 16436 58528 16437 58568
rect 16395 58519 16437 58528
rect 16491 58568 16533 58577
rect 16491 58528 16492 58568
rect 16532 58528 16533 58568
rect 16491 58519 16533 58528
rect 16587 58568 16629 58577
rect 16587 58528 16588 58568
rect 16628 58528 16629 58568
rect 16587 58519 16629 58528
rect 16771 58568 16829 58569
rect 16771 58528 16780 58568
rect 16820 58528 16829 58568
rect 16771 58527 16829 58528
rect 18019 58568 18077 58569
rect 18019 58528 18028 58568
rect 18068 58528 18077 58568
rect 18019 58527 18077 58528
rect 18403 58568 18461 58569
rect 18403 58528 18412 58568
rect 18452 58528 18461 58568
rect 18403 58527 18461 58528
rect 19651 58568 19709 58569
rect 19651 58528 19660 58568
rect 19700 58528 19709 58568
rect 19651 58527 19709 58528
rect 2667 58400 2709 58409
rect 2667 58360 2668 58400
rect 2708 58360 2709 58400
rect 2667 58351 2709 58360
rect 5163 58400 5205 58409
rect 5163 58360 5164 58400
rect 5204 58360 5205 58400
rect 5163 58351 5205 58360
rect 6795 58400 6837 58409
rect 6795 58360 6796 58400
rect 6836 58360 6837 58400
rect 6795 58351 6837 58360
rect 8811 58400 8853 58409
rect 8811 58360 8812 58400
rect 8852 58360 8853 58400
rect 8811 58351 8853 58360
rect 10443 58400 10485 58409
rect 10443 58360 10444 58400
rect 10484 58360 10485 58400
rect 10443 58351 10485 58360
rect 13123 58400 13181 58401
rect 13123 58360 13132 58400
rect 13172 58360 13181 58400
rect 13123 58359 13181 58360
rect 13795 58400 13853 58401
rect 13795 58360 13804 58400
rect 13844 58360 13853 58400
rect 13795 58359 13853 58360
rect 15811 58400 15869 58401
rect 15811 58360 15820 58400
rect 15860 58360 15869 58400
rect 15811 58359 15869 58360
rect 18219 58400 18261 58409
rect 18219 58360 18220 58400
rect 18260 58360 18261 58400
rect 18219 58351 18261 58360
rect 1152 58232 20452 58256
rect 1152 58192 4928 58232
rect 4968 58192 5010 58232
rect 5050 58192 5092 58232
rect 5132 58192 5174 58232
rect 5214 58192 5256 58232
rect 5296 58192 20048 58232
rect 20088 58192 20130 58232
rect 20170 58192 20212 58232
rect 20252 58192 20294 58232
rect 20334 58192 20376 58232
rect 20416 58192 20452 58232
rect 1152 58168 20452 58192
rect 5355 57980 5397 57989
rect 5355 57940 5356 57980
rect 5396 57940 5397 57980
rect 5355 57931 5397 57940
rect 10155 57980 10197 57989
rect 10155 57940 10156 57980
rect 10196 57940 10197 57980
rect 10155 57931 10197 57940
rect 2083 57896 2141 57897
rect 2083 57856 2092 57896
rect 2132 57856 2141 57896
rect 2083 57855 2141 57856
rect 3331 57896 3389 57897
rect 3331 57856 3340 57896
rect 3380 57856 3389 57896
rect 3331 57855 3389 57856
rect 3627 57896 3669 57905
rect 3627 57856 3628 57896
rect 3668 57856 3669 57896
rect 3627 57847 3669 57856
rect 3723 57896 3765 57905
rect 3723 57856 3724 57896
rect 3764 57856 3765 57896
rect 3723 57847 3765 57856
rect 4675 57896 4733 57897
rect 4675 57856 4684 57896
rect 4724 57856 4733 57896
rect 6307 57896 6365 57897
rect 4675 57855 4733 57856
rect 5211 57886 5253 57895
rect 5211 57846 5212 57886
rect 5252 57846 5253 57886
rect 6307 57856 6316 57896
rect 6356 57856 6365 57896
rect 6307 57855 6365 57856
rect 7555 57896 7613 57897
rect 7555 57856 7564 57896
rect 7604 57856 7613 57896
rect 7555 57855 7613 57856
rect 8427 57896 8469 57905
rect 8427 57856 8428 57896
rect 8468 57856 8469 57896
rect 8427 57847 8469 57856
rect 8523 57896 8565 57905
rect 8523 57856 8524 57896
rect 8564 57856 8565 57896
rect 8523 57847 8565 57856
rect 8907 57896 8949 57905
rect 8907 57856 8908 57896
rect 8948 57856 8949 57896
rect 8907 57847 8949 57856
rect 9475 57896 9533 57897
rect 9475 57856 9484 57896
rect 9524 57856 9533 57896
rect 9475 57855 9533 57856
rect 9963 57891 10005 57900
rect 9963 57851 9964 57891
rect 10004 57851 10005 57891
rect 11683 57896 11741 57897
rect 11683 57856 11692 57896
rect 11732 57856 11741 57896
rect 11683 57855 11741 57856
rect 12931 57896 12989 57897
rect 12931 57856 12940 57896
rect 12980 57856 12989 57896
rect 12931 57855 12989 57856
rect 13507 57896 13565 57897
rect 13507 57856 13516 57896
rect 13556 57856 13565 57896
rect 13507 57855 13565 57856
rect 14755 57896 14813 57897
rect 14755 57856 14764 57896
rect 14804 57856 14813 57896
rect 14755 57855 14813 57856
rect 15907 57896 15965 57897
rect 15907 57856 15916 57896
rect 15956 57856 15965 57896
rect 15907 57855 15965 57856
rect 17155 57896 17213 57897
rect 17155 57856 17164 57896
rect 17204 57856 17213 57896
rect 17155 57855 17213 57856
rect 17539 57896 17597 57897
rect 17539 57856 17548 57896
rect 17588 57856 17597 57896
rect 17539 57855 17597 57856
rect 17643 57896 17685 57905
rect 17643 57856 17644 57896
rect 17684 57856 17685 57896
rect 5211 57837 5253 57846
rect 9963 57842 10005 57851
rect 17643 57847 17685 57856
rect 4107 57812 4149 57821
rect 4107 57772 4108 57812
rect 4148 57772 4149 57812
rect 4107 57763 4149 57772
rect 4203 57812 4245 57821
rect 4203 57772 4204 57812
rect 4244 57772 4245 57812
rect 4203 57763 4245 57772
rect 9003 57812 9045 57821
rect 9003 57772 9004 57812
rect 9044 57772 9045 57812
rect 9003 57763 9045 57772
rect 11491 57812 11549 57813
rect 11491 57772 11500 57812
rect 11540 57772 11549 57812
rect 11491 57771 11549 57772
rect 11307 57728 11349 57737
rect 11307 57688 11308 57728
rect 11348 57688 11349 57728
rect 11307 57679 11349 57688
rect 13323 57728 13365 57737
rect 13323 57688 13324 57728
rect 13364 57688 13365 57728
rect 13323 57679 13365 57688
rect 1899 57644 1941 57653
rect 1899 57604 1900 57644
rect 1940 57604 1941 57644
rect 1899 57595 1941 57604
rect 7755 57644 7797 57653
rect 7755 57604 7756 57644
rect 7796 57604 7797 57644
rect 7755 57595 7797 57604
rect 13131 57644 13173 57653
rect 13131 57604 13132 57644
rect 13172 57604 13173 57644
rect 13131 57595 13173 57604
rect 17355 57644 17397 57653
rect 17355 57604 17356 57644
rect 17396 57604 17397 57644
rect 17355 57595 17397 57604
rect 1152 57476 20352 57500
rect 1152 57436 3688 57476
rect 3728 57436 3770 57476
rect 3810 57436 3852 57476
rect 3892 57436 3934 57476
rect 3974 57436 4016 57476
rect 4056 57436 18808 57476
rect 18848 57436 18890 57476
rect 18930 57436 18972 57476
rect 19012 57436 19054 57476
rect 19094 57436 19136 57476
rect 19176 57436 20352 57476
rect 1152 57412 20352 57436
rect 1803 57308 1845 57317
rect 1803 57268 1804 57308
rect 1844 57268 1845 57308
rect 1803 57259 1845 57268
rect 16299 57308 16341 57317
rect 16299 57268 16300 57308
rect 16340 57268 16341 57308
rect 16299 57259 16341 57268
rect 1987 57140 2045 57141
rect 1987 57100 1996 57140
rect 2036 57100 2045 57140
rect 1987 57099 2045 57100
rect 7755 57140 7797 57149
rect 7755 57100 7756 57140
rect 7796 57100 7797 57140
rect 7755 57091 7797 57100
rect 9667 57140 9725 57141
rect 9667 57100 9676 57140
rect 9716 57100 9725 57140
rect 9667 57099 9725 57100
rect 12171 57140 12213 57149
rect 12171 57100 12172 57140
rect 12212 57100 12213 57140
rect 12171 57091 12213 57100
rect 14283 57140 14325 57149
rect 14283 57100 14284 57140
rect 14324 57100 14325 57140
rect 14283 57091 14325 57100
rect 14379 57140 14421 57149
rect 14379 57100 14380 57140
rect 14420 57100 14421 57140
rect 14379 57091 14421 57100
rect 16003 57140 16061 57141
rect 16003 57100 16012 57140
rect 16052 57100 16061 57140
rect 16003 57099 16061 57100
rect 16483 57140 16541 57141
rect 16483 57100 16492 57140
rect 16532 57100 16541 57140
rect 16483 57099 16541 57100
rect 20131 57098 20189 57099
rect 8715 57070 8757 57079
rect 2179 57056 2237 57057
rect 2179 57016 2188 57056
rect 2228 57016 2237 57056
rect 2179 57015 2237 57016
rect 3427 57056 3485 57057
rect 3427 57016 3436 57056
rect 3476 57016 3485 57056
rect 3427 57015 3485 57016
rect 3811 57056 3869 57057
rect 3811 57016 3820 57056
rect 3860 57016 3869 57056
rect 3811 57015 3869 57016
rect 5059 57056 5117 57057
rect 5059 57016 5068 57056
rect 5108 57016 5117 57056
rect 5059 57015 5117 57016
rect 5443 57056 5501 57057
rect 5443 57016 5452 57056
rect 5492 57016 5501 57056
rect 5443 57015 5501 57016
rect 6691 57056 6749 57057
rect 6691 57016 6700 57056
rect 6740 57016 6749 57056
rect 6691 57015 6749 57016
rect 7179 57056 7221 57065
rect 7179 57016 7180 57056
rect 7220 57016 7221 57056
rect 7179 57007 7221 57016
rect 7275 57056 7317 57065
rect 7275 57016 7276 57056
rect 7316 57016 7317 57056
rect 7275 57007 7317 57016
rect 7659 57056 7701 57065
rect 7659 57016 7660 57056
rect 7700 57016 7701 57056
rect 7659 57007 7701 57016
rect 8227 57056 8285 57057
rect 8227 57016 8236 57056
rect 8276 57016 8285 57056
rect 8715 57030 8716 57070
rect 8756 57030 8757 57070
rect 13131 57070 13173 57079
rect 8715 57021 8757 57030
rect 9859 57056 9917 57057
rect 8227 57015 8285 57016
rect 9859 57016 9868 57056
rect 9908 57016 9917 57056
rect 9859 57015 9917 57016
rect 11107 57056 11165 57057
rect 11107 57016 11116 57056
rect 11156 57016 11165 57056
rect 11107 57015 11165 57016
rect 11595 57056 11637 57065
rect 11595 57016 11596 57056
rect 11636 57016 11637 57056
rect 11595 57007 11637 57016
rect 11691 57056 11733 57065
rect 11691 57016 11692 57056
rect 11732 57016 11733 57056
rect 11691 57007 11733 57016
rect 12075 57056 12117 57065
rect 12075 57016 12076 57056
rect 12116 57016 12117 57056
rect 12075 57007 12117 57016
rect 12643 57056 12701 57057
rect 12643 57016 12652 57056
rect 12692 57016 12701 57056
rect 13131 57030 13132 57070
rect 13172 57030 13173 57070
rect 15339 57070 15381 57079
rect 13131 57021 13173 57030
rect 13803 57056 13845 57065
rect 12643 57015 12701 57016
rect 13803 57016 13804 57056
rect 13844 57016 13845 57056
rect 13803 57007 13845 57016
rect 13899 57056 13941 57065
rect 13899 57016 13900 57056
rect 13940 57016 13941 57056
rect 13899 57007 13941 57016
rect 14851 57056 14909 57057
rect 14851 57016 14860 57056
rect 14900 57016 14909 57056
rect 15339 57030 15340 57070
rect 15380 57030 15381 57070
rect 18315 57070 18357 57079
rect 15339 57021 15381 57030
rect 16779 57056 16821 57065
rect 14851 57015 14909 57016
rect 16779 57016 16780 57056
rect 16820 57016 16821 57056
rect 16779 57007 16821 57016
rect 16875 57056 16917 57065
rect 16875 57016 16876 57056
rect 16916 57016 16917 57056
rect 16875 57007 16917 57016
rect 17259 57056 17301 57065
rect 17259 57016 17260 57056
rect 17300 57016 17301 57056
rect 17259 57007 17301 57016
rect 17355 57056 17397 57065
rect 17355 57016 17356 57056
rect 17396 57016 17397 57056
rect 17355 57007 17397 57016
rect 17827 57056 17885 57057
rect 17827 57016 17836 57056
rect 17876 57016 17885 57056
rect 18315 57030 18316 57070
rect 18356 57030 18357 57070
rect 20131 57058 20140 57098
rect 20180 57058 20189 57098
rect 20131 57057 20189 57058
rect 18315 57021 18357 57030
rect 18883 57056 18941 57057
rect 17827 57015 17885 57016
rect 18883 57016 18892 57056
rect 18932 57016 18941 57056
rect 18883 57015 18941 57016
rect 8907 56972 8949 56981
rect 8907 56932 8908 56972
rect 8948 56932 8949 56972
rect 8907 56923 8949 56932
rect 11307 56972 11349 56981
rect 11307 56932 11308 56972
rect 11348 56932 11349 56972
rect 11307 56923 11349 56932
rect 13323 56972 13365 56981
rect 13323 56932 13324 56972
rect 13364 56932 13365 56972
rect 13323 56923 13365 56932
rect 18507 56972 18549 56981
rect 18507 56932 18508 56972
rect 18548 56932 18549 56972
rect 18507 56923 18549 56932
rect 3627 56888 3669 56897
rect 3627 56848 3628 56888
rect 3668 56848 3669 56888
rect 3627 56839 3669 56848
rect 5259 56888 5301 56897
rect 5259 56848 5260 56888
rect 5300 56848 5301 56888
rect 5259 56839 5301 56848
rect 6891 56888 6933 56897
rect 6891 56848 6892 56888
rect 6932 56848 6933 56888
rect 6891 56839 6933 56848
rect 9483 56888 9525 56897
rect 9483 56848 9484 56888
rect 9524 56848 9525 56888
rect 9483 56839 9525 56848
rect 15531 56888 15573 56897
rect 15531 56848 15532 56888
rect 15572 56848 15573 56888
rect 15531 56839 15573 56848
rect 15819 56888 15861 56897
rect 15819 56848 15820 56888
rect 15860 56848 15861 56888
rect 15819 56839 15861 56848
rect 18699 56888 18741 56897
rect 18699 56848 18700 56888
rect 18740 56848 18741 56888
rect 18699 56839 18741 56848
rect 1152 56720 20452 56744
rect 1152 56680 4928 56720
rect 4968 56680 5010 56720
rect 5050 56680 5092 56720
rect 5132 56680 5174 56720
rect 5214 56680 5256 56720
rect 5296 56680 20048 56720
rect 20088 56680 20130 56720
rect 20170 56680 20212 56720
rect 20252 56680 20294 56720
rect 20334 56680 20376 56720
rect 20416 56680 20452 56720
rect 1152 56656 20452 56680
rect 12363 56552 12405 56561
rect 12363 56512 12364 56552
rect 12404 56512 12405 56552
rect 12363 56503 12405 56512
rect 16683 56552 16725 56561
rect 16683 56512 16684 56552
rect 16724 56512 16725 56552
rect 16683 56503 16725 56512
rect 16875 56552 16917 56561
rect 16875 56512 16876 56552
rect 16916 56512 16917 56552
rect 16875 56503 16917 56512
rect 19563 56552 19605 56561
rect 19563 56512 19564 56552
rect 19604 56512 19605 56552
rect 19563 56503 19605 56512
rect 3051 56468 3093 56477
rect 3051 56428 3052 56468
rect 3092 56428 3093 56468
rect 3051 56419 3093 56428
rect 7179 56468 7221 56477
rect 7179 56428 7180 56468
rect 7220 56428 7221 56468
rect 7179 56419 7221 56428
rect 9195 56468 9237 56477
rect 9195 56428 9196 56468
rect 9236 56428 9237 56468
rect 9195 56419 9237 56428
rect 19179 56468 19221 56477
rect 19179 56428 19180 56468
rect 19220 56428 19221 56468
rect 19179 56419 19221 56428
rect 1411 56384 1469 56385
rect 1411 56344 1420 56384
rect 1460 56344 1469 56384
rect 1411 56343 1469 56344
rect 2659 56384 2717 56385
rect 2659 56344 2668 56384
rect 2708 56344 2717 56384
rect 2659 56343 2717 56344
rect 3243 56379 3285 56388
rect 3243 56339 3244 56379
rect 3284 56339 3285 56379
rect 3715 56384 3773 56385
rect 3715 56344 3724 56384
rect 3764 56344 3773 56384
rect 3715 56343 3773 56344
rect 4203 56384 4245 56393
rect 4203 56344 4204 56384
rect 4244 56344 4245 56384
rect 3243 56330 3285 56339
rect 4203 56335 4245 56344
rect 4683 56384 4725 56393
rect 4683 56344 4684 56384
rect 4724 56344 4725 56384
rect 4683 56335 4725 56344
rect 4779 56384 4821 56393
rect 4779 56344 4780 56384
rect 4820 56344 4821 56384
rect 4779 56335 4821 56344
rect 5731 56384 5789 56385
rect 5731 56344 5740 56384
rect 5780 56344 5789 56384
rect 5731 56343 5789 56344
rect 6979 56384 7037 56385
rect 6979 56344 6988 56384
rect 7028 56344 7037 56384
rect 6979 56343 7037 56344
rect 7467 56384 7509 56393
rect 7467 56344 7468 56384
rect 7508 56344 7509 56384
rect 7467 56335 7509 56344
rect 7563 56384 7605 56393
rect 7563 56344 7564 56384
rect 7604 56344 7605 56384
rect 7563 56335 7605 56344
rect 7947 56384 7989 56393
rect 7947 56344 7948 56384
rect 7988 56344 7989 56384
rect 7947 56335 7989 56344
rect 8043 56384 8085 56393
rect 8043 56344 8044 56384
rect 8084 56344 8085 56384
rect 8043 56335 8085 56344
rect 8515 56384 8573 56385
rect 8515 56344 8524 56384
rect 8564 56344 8573 56384
rect 8515 56343 8573 56344
rect 9003 56379 9045 56388
rect 9003 56339 9004 56379
rect 9044 56339 9045 56379
rect 10723 56384 10781 56385
rect 10723 56344 10732 56384
rect 10772 56344 10781 56384
rect 10723 56343 10781 56344
rect 13219 56384 13277 56385
rect 13219 56344 13228 56384
rect 13268 56344 13277 56384
rect 13219 56343 13277 56344
rect 14467 56384 14525 56385
rect 14467 56344 14476 56384
rect 14516 56344 14525 56384
rect 14467 56343 14525 56344
rect 15235 56384 15293 56385
rect 15235 56344 15244 56384
rect 15284 56344 15293 56384
rect 15235 56343 15293 56344
rect 16483 56384 16541 56385
rect 16483 56344 16492 56384
rect 16532 56344 16541 56384
rect 16483 56343 16541 56344
rect 17451 56384 17493 56393
rect 17451 56344 17452 56384
rect 17492 56344 17493 56384
rect 9003 56330 9045 56339
rect 11971 56342 12029 56343
rect 4299 56300 4341 56309
rect 11971 56302 11980 56342
rect 12020 56302 12029 56342
rect 17451 56335 17493 56344
rect 17547 56384 17589 56393
rect 17547 56344 17548 56384
rect 17588 56344 17589 56384
rect 17547 56335 17589 56344
rect 17931 56384 17973 56393
rect 17931 56344 17932 56384
rect 17972 56344 17973 56384
rect 17931 56335 17973 56344
rect 18499 56384 18557 56385
rect 18499 56344 18508 56384
rect 18548 56344 18557 56384
rect 18499 56343 18557 56344
rect 18987 56379 19029 56388
rect 18987 56339 18988 56379
rect 19028 56339 19029 56379
rect 18987 56330 19029 56339
rect 11971 56301 12029 56302
rect 4299 56260 4300 56300
rect 4340 56260 4341 56300
rect 4299 56251 4341 56260
rect 10339 56300 10397 56301
rect 10339 56260 10348 56300
rect 10388 56260 10397 56300
rect 10339 56259 10397 56260
rect 12547 56300 12605 56301
rect 12547 56260 12556 56300
rect 12596 56260 12605 56300
rect 12547 56259 12605 56260
rect 15043 56300 15101 56301
rect 15043 56260 15052 56300
rect 15092 56260 15101 56300
rect 15043 56259 15101 56260
rect 17059 56300 17117 56301
rect 17059 56260 17068 56300
rect 17108 56260 17117 56300
rect 17059 56259 17117 56260
rect 18027 56300 18069 56309
rect 18027 56260 18028 56300
rect 18068 56260 18069 56300
rect 18027 56251 18069 56260
rect 19363 56300 19421 56301
rect 19363 56260 19372 56300
rect 19412 56260 19421 56300
rect 19363 56259 19421 56260
rect 2859 56216 2901 56225
rect 2859 56176 2860 56216
rect 2900 56176 2901 56216
rect 2859 56167 2901 56176
rect 10539 56132 10581 56141
rect 10539 56092 10540 56132
rect 10580 56092 10581 56132
rect 10539 56083 10581 56092
rect 12171 56132 12213 56141
rect 12171 56092 12172 56132
rect 12212 56092 12213 56132
rect 12171 56083 12213 56092
rect 14667 56132 14709 56141
rect 14667 56092 14668 56132
rect 14708 56092 14709 56132
rect 14667 56083 14709 56092
rect 14859 56132 14901 56141
rect 14859 56092 14860 56132
rect 14900 56092 14901 56132
rect 14859 56083 14901 56092
rect 1152 55964 20352 55988
rect 1152 55924 3688 55964
rect 3728 55924 3770 55964
rect 3810 55924 3852 55964
rect 3892 55924 3934 55964
rect 3974 55924 4016 55964
rect 4056 55924 18808 55964
rect 18848 55924 18890 55964
rect 18930 55924 18972 55964
rect 19012 55924 19054 55964
rect 19094 55924 19136 55964
rect 19176 55924 20352 55964
rect 1152 55900 20352 55924
rect 2859 55712 2901 55721
rect 2859 55672 2860 55712
rect 2900 55672 2901 55712
rect 2859 55663 2901 55672
rect 19563 55712 19605 55721
rect 19563 55672 19564 55712
rect 19604 55672 19605 55712
rect 19563 55663 19605 55672
rect 10051 55639 10109 55640
rect 3235 55628 3293 55629
rect 3235 55588 3244 55628
rect 3284 55588 3293 55628
rect 3235 55587 3293 55588
rect 5643 55628 5685 55637
rect 5643 55588 5644 55628
rect 5684 55588 5685 55628
rect 5643 55579 5685 55588
rect 5739 55628 5781 55637
rect 5739 55588 5740 55628
rect 5780 55588 5781 55628
rect 5739 55579 5781 55588
rect 8427 55628 8469 55637
rect 8427 55588 8428 55628
rect 8468 55588 8469 55628
rect 8427 55579 8469 55588
rect 8523 55628 8565 55637
rect 8523 55588 8524 55628
rect 8564 55588 8565 55628
rect 10051 55599 10060 55639
rect 10100 55599 10109 55639
rect 10051 55598 10109 55599
rect 11211 55628 11253 55637
rect 8523 55579 8565 55588
rect 11211 55588 11212 55628
rect 11252 55588 11253 55628
rect 11211 55579 11253 55588
rect 11307 55628 11349 55637
rect 11307 55588 11308 55628
rect 11348 55588 11349 55628
rect 11307 55579 11349 55588
rect 19363 55628 19421 55629
rect 19363 55588 19372 55628
rect 19412 55588 19421 55628
rect 19363 55587 19421 55588
rect 6699 55558 6741 55567
rect 12267 55558 12309 55567
rect 1411 55544 1469 55545
rect 1411 55504 1420 55544
rect 1460 55504 1469 55544
rect 1411 55503 1469 55504
rect 2659 55544 2717 55545
rect 2659 55504 2668 55544
rect 2708 55504 2717 55544
rect 2659 55503 2717 55504
rect 3427 55544 3485 55545
rect 3427 55504 3436 55544
rect 3476 55504 3485 55544
rect 3427 55503 3485 55504
rect 4675 55544 4733 55545
rect 4675 55504 4684 55544
rect 4724 55504 4733 55544
rect 4675 55503 4733 55504
rect 5163 55544 5205 55553
rect 5163 55504 5164 55544
rect 5204 55504 5205 55544
rect 5163 55495 5205 55504
rect 5259 55544 5301 55553
rect 5259 55504 5260 55544
rect 5300 55504 5301 55544
rect 5259 55495 5301 55504
rect 6211 55544 6269 55545
rect 6211 55504 6220 55544
rect 6260 55504 6269 55544
rect 6699 55518 6700 55558
rect 6740 55518 6741 55558
rect 6699 55509 6741 55518
rect 7947 55544 7989 55553
rect 6211 55503 6269 55504
rect 7947 55504 7948 55544
rect 7988 55504 7989 55544
rect 7947 55495 7989 55504
rect 8043 55544 8085 55553
rect 9483 55549 9525 55558
rect 8043 55504 8044 55544
rect 8084 55504 8085 55544
rect 8043 55495 8085 55504
rect 8995 55544 9053 55545
rect 8995 55504 9004 55544
rect 9044 55504 9053 55544
rect 8995 55503 9053 55504
rect 9483 55509 9484 55549
rect 9524 55509 9525 55549
rect 9483 55500 9525 55509
rect 10731 55544 10773 55553
rect 10731 55504 10732 55544
rect 10772 55504 10773 55544
rect 10731 55495 10773 55504
rect 10827 55544 10869 55553
rect 10827 55504 10828 55544
rect 10868 55504 10869 55544
rect 10827 55495 10869 55504
rect 11779 55544 11837 55545
rect 11779 55504 11788 55544
rect 11828 55504 11837 55544
rect 12267 55518 12268 55558
rect 12308 55518 12309 55558
rect 12267 55509 12309 55518
rect 13123 55544 13181 55545
rect 11779 55503 11837 55504
rect 13123 55504 13132 55544
rect 13172 55504 13181 55544
rect 13123 55503 13181 55504
rect 14371 55544 14429 55545
rect 14371 55504 14380 55544
rect 14420 55504 14429 55544
rect 14371 55503 14429 55504
rect 15043 55544 15101 55545
rect 15043 55504 15052 55544
rect 15092 55504 15101 55544
rect 15043 55503 15101 55504
rect 16291 55544 16349 55545
rect 16291 55504 16300 55544
rect 16340 55504 16349 55544
rect 16291 55503 16349 55504
rect 16867 55544 16925 55545
rect 16867 55504 16876 55544
rect 16916 55504 16925 55544
rect 16867 55503 16925 55504
rect 18115 55544 18173 55545
rect 18115 55504 18124 55544
rect 18164 55504 18173 55544
rect 18115 55503 18173 55504
rect 6891 55460 6933 55469
rect 6891 55420 6892 55460
rect 6932 55420 6933 55460
rect 6891 55411 6933 55420
rect 9675 55460 9717 55469
rect 9675 55420 9676 55460
rect 9716 55420 9717 55460
rect 9675 55411 9717 55420
rect 12459 55460 12501 55469
rect 12459 55420 12460 55460
rect 12500 55420 12501 55460
rect 12459 55411 12501 55420
rect 3051 55376 3093 55385
rect 3051 55336 3052 55376
rect 3092 55336 3093 55376
rect 3051 55327 3093 55336
rect 4875 55376 4917 55385
rect 4875 55336 4876 55376
rect 4916 55336 4917 55376
rect 4875 55327 4917 55336
rect 9867 55376 9909 55385
rect 9867 55336 9868 55376
rect 9908 55336 9909 55376
rect 9867 55327 9909 55336
rect 14571 55376 14613 55385
rect 14571 55336 14572 55376
rect 14612 55336 14613 55376
rect 14571 55327 14613 55336
rect 16491 55376 16533 55385
rect 16491 55336 16492 55376
rect 16532 55336 16533 55376
rect 16491 55327 16533 55336
rect 16683 55376 16725 55385
rect 16683 55336 16684 55376
rect 16724 55336 16725 55376
rect 16683 55327 16725 55336
rect 1152 55208 20452 55232
rect 1152 55168 4928 55208
rect 4968 55168 5010 55208
rect 5050 55168 5092 55208
rect 5132 55168 5174 55208
rect 5214 55168 5256 55208
rect 5296 55168 20048 55208
rect 20088 55168 20130 55208
rect 20170 55168 20212 55208
rect 20252 55168 20294 55208
rect 20334 55168 20376 55208
rect 20416 55168 20452 55208
rect 1152 55144 20452 55168
rect 9387 55040 9429 55049
rect 9387 55000 9388 55040
rect 9428 55000 9429 55040
rect 9387 54991 9429 55000
rect 11019 55040 11061 55049
rect 11019 55000 11020 55040
rect 11060 55000 11061 55040
rect 11019 54991 11061 55000
rect 16779 55040 16821 55049
rect 16779 55000 16780 55040
rect 16820 55000 16821 55040
rect 16779 54991 16821 55000
rect 20235 55040 20277 55049
rect 20235 55000 20236 55040
rect 20276 55000 20277 55040
rect 20235 54991 20277 55000
rect 2187 54956 2229 54965
rect 2187 54916 2188 54956
rect 2228 54916 2229 54956
rect 2187 54907 2229 54916
rect 12747 54956 12789 54965
rect 12747 54916 12748 54956
rect 12788 54916 12789 54956
rect 12747 54907 12789 54916
rect 14763 54956 14805 54965
rect 14763 54916 14764 54956
rect 14804 54916 14805 54956
rect 14763 54907 14805 54916
rect 19083 54956 19125 54965
rect 19083 54916 19084 54956
rect 19124 54916 19125 54956
rect 19083 54907 19125 54916
rect 2851 54872 2909 54873
rect 2331 54862 2373 54871
rect 2331 54822 2332 54862
rect 2372 54822 2373 54862
rect 2851 54832 2860 54872
rect 2900 54832 2909 54872
rect 2851 54831 2909 54832
rect 3339 54872 3381 54881
rect 3339 54832 3340 54872
rect 3380 54832 3381 54872
rect 3339 54823 3381 54832
rect 3819 54872 3861 54881
rect 3819 54832 3820 54872
rect 3860 54832 3861 54872
rect 3819 54823 3861 54832
rect 3915 54872 3957 54881
rect 3915 54832 3916 54872
rect 3956 54832 3957 54872
rect 3915 54823 3957 54832
rect 5443 54872 5501 54873
rect 5443 54832 5452 54872
rect 5492 54832 5501 54872
rect 5443 54831 5501 54832
rect 6691 54872 6749 54873
rect 6691 54832 6700 54872
rect 6740 54832 6749 54872
rect 6691 54831 6749 54832
rect 7939 54872 7997 54873
rect 7939 54832 7948 54872
rect 7988 54832 7997 54872
rect 7939 54831 7997 54832
rect 9187 54872 9245 54873
rect 9187 54832 9196 54872
rect 9236 54832 9245 54872
rect 9187 54831 9245 54832
rect 9571 54872 9629 54873
rect 9571 54832 9580 54872
rect 9620 54832 9629 54872
rect 9571 54831 9629 54832
rect 10819 54872 10877 54873
rect 10819 54832 10828 54872
rect 10868 54832 10877 54872
rect 10819 54831 10877 54832
rect 11299 54872 11357 54873
rect 11299 54832 11308 54872
rect 11348 54832 11357 54872
rect 13035 54872 13077 54881
rect 11299 54831 11357 54832
rect 12547 54851 12605 54852
rect 2331 54813 2373 54822
rect 12547 54811 12556 54851
rect 12596 54811 12605 54851
rect 13035 54832 13036 54872
rect 13076 54832 13077 54872
rect 13035 54823 13077 54832
rect 13131 54872 13173 54881
rect 13131 54832 13132 54872
rect 13172 54832 13173 54872
rect 13131 54823 13173 54832
rect 13611 54872 13653 54881
rect 13611 54832 13612 54872
rect 13652 54832 13653 54872
rect 13611 54823 13653 54832
rect 14083 54872 14141 54873
rect 14083 54832 14092 54872
rect 14132 54832 14141 54872
rect 14083 54831 14141 54832
rect 14571 54867 14613 54876
rect 14571 54827 14572 54867
rect 14612 54827 14613 54867
rect 14571 54818 14613 54827
rect 15051 54872 15093 54881
rect 15051 54832 15052 54872
rect 15092 54832 15093 54872
rect 15051 54823 15093 54832
rect 15147 54872 15189 54881
rect 15147 54832 15148 54872
rect 15188 54832 15189 54872
rect 15147 54823 15189 54832
rect 15531 54872 15573 54881
rect 15531 54832 15532 54872
rect 15572 54832 15573 54872
rect 15531 54823 15573 54832
rect 15627 54872 15669 54881
rect 15627 54832 15628 54872
rect 15668 54832 15669 54872
rect 15627 54823 15669 54832
rect 16099 54872 16157 54873
rect 16099 54832 16108 54872
rect 16148 54832 16157 54872
rect 16099 54831 16157 54832
rect 16587 54867 16629 54876
rect 16587 54827 16588 54867
rect 16628 54827 16629 54867
rect 16587 54818 16629 54827
rect 17355 54872 17397 54881
rect 17355 54832 17356 54872
rect 17396 54832 17397 54872
rect 17355 54823 17397 54832
rect 17451 54872 17493 54881
rect 17451 54832 17452 54872
rect 17492 54832 17493 54872
rect 17451 54823 17493 54832
rect 17931 54872 17973 54881
rect 17931 54832 17932 54872
rect 17972 54832 17973 54872
rect 17931 54823 17973 54832
rect 18403 54872 18461 54873
rect 18403 54832 18412 54872
rect 18452 54832 18461 54872
rect 18403 54831 18461 54832
rect 18939 54830 18981 54839
rect 12547 54810 12605 54811
rect 1987 54788 2045 54789
rect 1987 54748 1996 54788
rect 2036 54748 2045 54788
rect 1987 54747 2045 54748
rect 3435 54788 3477 54797
rect 3435 54748 3436 54788
rect 3476 54748 3477 54788
rect 3435 54739 3477 54748
rect 13515 54788 13557 54797
rect 13515 54748 13516 54788
rect 13556 54748 13557 54788
rect 13515 54739 13557 54748
rect 17835 54788 17877 54797
rect 17835 54748 17836 54788
rect 17876 54748 17877 54788
rect 18939 54790 18940 54830
rect 18980 54790 18981 54830
rect 18939 54781 18981 54790
rect 19459 54788 19517 54789
rect 17835 54739 17877 54748
rect 19459 54748 19468 54788
rect 19508 54748 19517 54788
rect 19459 54747 19517 54748
rect 19651 54788 19709 54789
rect 19651 54748 19660 54788
rect 19700 54748 19709 54788
rect 19651 54747 19709 54748
rect 20035 54788 20093 54789
rect 20035 54748 20044 54788
rect 20084 54748 20093 54788
rect 20035 54747 20093 54748
rect 1803 54620 1845 54629
rect 1803 54580 1804 54620
rect 1844 54580 1845 54620
rect 1803 54571 1845 54580
rect 6891 54620 6933 54629
rect 6891 54580 6892 54620
rect 6932 54580 6933 54620
rect 6891 54571 6933 54580
rect 19275 54620 19317 54629
rect 19275 54580 19276 54620
rect 19316 54580 19317 54620
rect 19275 54571 19317 54580
rect 19851 54620 19893 54629
rect 19851 54580 19852 54620
rect 19892 54580 19893 54620
rect 19851 54571 19893 54580
rect 1152 54452 20352 54476
rect 1152 54412 3688 54452
rect 3728 54412 3770 54452
rect 3810 54412 3852 54452
rect 3892 54412 3934 54452
rect 3974 54412 4016 54452
rect 4056 54412 18808 54452
rect 18848 54412 18890 54452
rect 18930 54412 18972 54452
rect 19012 54412 19054 54452
rect 19094 54412 19136 54452
rect 19176 54412 20352 54452
rect 1152 54388 20352 54412
rect 19275 54284 19317 54293
rect 19275 54244 19276 54284
rect 19316 54244 19317 54284
rect 19275 54235 19317 54244
rect 17163 54200 17205 54209
rect 17163 54160 17164 54200
rect 17204 54160 17205 54200
rect 17163 54151 17205 54160
rect 9955 54116 10013 54117
rect 9955 54076 9964 54116
rect 10004 54076 10013 54116
rect 9955 54075 10013 54076
rect 12163 54116 12221 54117
rect 12163 54076 12172 54116
rect 12212 54076 12221 54116
rect 12163 54075 12221 54076
rect 17347 54116 17405 54117
rect 17347 54076 17356 54116
rect 17396 54076 17405 54116
rect 17347 54075 17405 54076
rect 19459 54116 19517 54117
rect 19459 54076 19468 54116
rect 19508 54076 19517 54116
rect 19459 54075 19517 54076
rect 19843 54116 19901 54117
rect 19843 54076 19852 54116
rect 19892 54076 19901 54116
rect 19843 54075 19901 54076
rect 4875 54046 4917 54055
rect 1219 54032 1277 54033
rect 1219 53992 1228 54032
rect 1268 53992 1277 54032
rect 1219 53991 1277 53992
rect 2467 54032 2525 54033
rect 2467 53992 2476 54032
rect 2516 53992 2525 54032
rect 2467 53991 2525 53992
rect 3339 54032 3381 54041
rect 3339 53992 3340 54032
rect 3380 53992 3381 54032
rect 3339 53983 3381 53992
rect 3435 54032 3477 54041
rect 3435 53992 3436 54032
rect 3476 53992 3477 54032
rect 3435 53983 3477 53992
rect 3819 54032 3861 54041
rect 3819 53992 3820 54032
rect 3860 53992 3861 54032
rect 3819 53983 3861 53992
rect 3915 54032 3957 54041
rect 3915 53992 3916 54032
rect 3956 53992 3957 54032
rect 3915 53983 3957 53992
rect 4387 54032 4445 54033
rect 4387 53992 4396 54032
rect 4436 53992 4445 54032
rect 4875 54006 4876 54046
rect 4916 54006 4917 54046
rect 4875 53997 4917 54006
rect 6691 54032 6749 54033
rect 4387 53991 4445 53992
rect 6691 53992 6700 54032
rect 6740 53992 6749 54032
rect 6691 53991 6749 53992
rect 7939 54032 7997 54033
rect 7939 53992 7948 54032
rect 7988 53992 7997 54032
rect 7939 53991 7997 53992
rect 8323 54032 8381 54033
rect 8323 53992 8332 54032
rect 8372 53992 8381 54032
rect 8323 53991 8381 53992
rect 9571 54032 9629 54033
rect 9571 53992 9580 54032
rect 9620 53992 9629 54032
rect 9571 53991 9629 53992
rect 10339 54032 10397 54033
rect 10339 53992 10348 54032
rect 10388 53992 10397 54032
rect 10339 53991 10397 53992
rect 11587 54032 11645 54033
rect 11587 53992 11596 54032
rect 11636 53992 11645 54032
rect 11587 53991 11645 53992
rect 13795 54032 13853 54033
rect 13795 53992 13804 54032
rect 13844 53992 13853 54032
rect 13795 53991 13853 53992
rect 15043 54032 15101 54033
rect 15043 53992 15052 54032
rect 15092 53992 15101 54032
rect 15043 53991 15101 53992
rect 15523 54032 15581 54033
rect 15523 53992 15532 54032
rect 15572 53992 15581 54032
rect 15523 53991 15581 53992
rect 16771 54032 16829 54033
rect 16771 53992 16780 54032
rect 16820 53992 16829 54032
rect 16771 53991 16829 53992
rect 17827 54032 17885 54033
rect 17827 53992 17836 54032
rect 17876 53992 17885 54032
rect 17827 53991 17885 53992
rect 19075 54032 19133 54033
rect 19075 53992 19084 54032
rect 19124 53992 19133 54032
rect 19075 53991 19133 53992
rect 5067 53948 5109 53957
rect 5067 53908 5068 53948
rect 5108 53908 5109 53948
rect 5067 53899 5109 53908
rect 2667 53864 2709 53873
rect 2667 53824 2668 53864
rect 2708 53824 2709 53864
rect 2667 53815 2709 53824
rect 8139 53864 8181 53873
rect 8139 53824 8140 53864
rect 8180 53824 8181 53864
rect 8139 53815 8181 53824
rect 9771 53864 9813 53873
rect 9771 53824 9772 53864
rect 9812 53824 9813 53864
rect 9771 53815 9813 53824
rect 10155 53864 10197 53873
rect 10155 53824 10156 53864
rect 10196 53824 10197 53864
rect 10155 53815 10197 53824
rect 11787 53864 11829 53873
rect 11787 53824 11788 53864
rect 11828 53824 11829 53864
rect 11787 53815 11829 53824
rect 11979 53864 12021 53873
rect 11979 53824 11980 53864
rect 12020 53824 12021 53864
rect 11979 53815 12021 53824
rect 15243 53864 15285 53873
rect 15243 53824 15244 53864
rect 15284 53824 15285 53864
rect 15243 53815 15285 53824
rect 16971 53864 17013 53873
rect 16971 53824 16972 53864
rect 17012 53824 17013 53864
rect 16971 53815 17013 53824
rect 19659 53864 19701 53873
rect 19659 53824 19660 53864
rect 19700 53824 19701 53864
rect 19659 53815 19701 53824
rect 20043 53864 20085 53873
rect 20043 53824 20044 53864
rect 20084 53824 20085 53864
rect 20043 53815 20085 53824
rect 1152 53696 20452 53720
rect 1152 53656 4928 53696
rect 4968 53656 5010 53696
rect 5050 53656 5092 53696
rect 5132 53656 5174 53696
rect 5214 53656 5256 53696
rect 5296 53656 20048 53696
rect 20088 53656 20130 53696
rect 20170 53656 20212 53696
rect 20252 53656 20294 53696
rect 20334 53656 20376 53696
rect 20416 53656 20452 53696
rect 1152 53632 20452 53656
rect 3147 53528 3189 53537
rect 3147 53488 3148 53528
rect 3188 53488 3189 53528
rect 3147 53479 3189 53488
rect 9291 53528 9333 53537
rect 9291 53488 9292 53528
rect 9332 53488 9333 53528
rect 9291 53479 9333 53488
rect 16875 53528 16917 53537
rect 16875 53488 16876 53528
rect 16916 53488 16917 53528
rect 16875 53479 16917 53488
rect 2955 53444 2997 53453
rect 2955 53404 2956 53444
rect 2996 53404 2997 53444
rect 2955 53395 2997 53404
rect 7275 53444 7317 53453
rect 7275 53404 7276 53444
rect 7316 53404 7317 53444
rect 7275 53395 7317 53404
rect 1507 53360 1565 53361
rect 1507 53320 1516 53360
rect 1556 53320 1565 53360
rect 1507 53319 1565 53320
rect 2755 53360 2813 53361
rect 2755 53320 2764 53360
rect 2804 53320 2813 53360
rect 3811 53360 3869 53361
rect 2755 53319 2813 53320
rect 3291 53350 3333 53359
rect 3291 53310 3292 53350
rect 3332 53310 3333 53350
rect 3811 53320 3820 53360
rect 3860 53320 3869 53360
rect 3811 53319 3869 53320
rect 4779 53360 4821 53369
rect 4779 53320 4780 53360
rect 4820 53320 4821 53360
rect 4779 53311 4821 53320
rect 4875 53360 4917 53369
rect 4875 53320 4876 53360
rect 4916 53320 4917 53360
rect 4875 53311 4917 53320
rect 5827 53360 5885 53361
rect 5827 53320 5836 53360
rect 5876 53320 5885 53360
rect 5827 53319 5885 53320
rect 7075 53360 7133 53361
rect 7075 53320 7084 53360
rect 7124 53320 7133 53360
rect 7075 53319 7133 53320
rect 7563 53360 7605 53369
rect 7563 53320 7564 53360
rect 7604 53320 7605 53360
rect 7563 53311 7605 53320
rect 7659 53360 7701 53369
rect 7659 53320 7660 53360
rect 7700 53320 7701 53360
rect 7659 53311 7701 53320
rect 8611 53360 8669 53361
rect 8611 53320 8620 53360
rect 8660 53320 8669 53360
rect 8611 53319 8669 53320
rect 9099 53355 9141 53364
rect 9099 53315 9100 53355
rect 9140 53315 9141 53355
rect 9475 53360 9533 53361
rect 9475 53320 9484 53360
rect 9524 53320 9533 53360
rect 9475 53319 9533 53320
rect 10723 53360 10781 53361
rect 10723 53320 10732 53360
rect 10772 53320 10781 53360
rect 10723 53319 10781 53320
rect 11107 53360 11165 53361
rect 11107 53320 11116 53360
rect 11156 53320 11165 53360
rect 11107 53319 11165 53320
rect 12355 53360 12413 53361
rect 12355 53320 12364 53360
rect 12404 53320 12413 53360
rect 12355 53319 12413 53320
rect 12739 53360 12797 53361
rect 12739 53320 12748 53360
rect 12788 53320 12797 53360
rect 12739 53319 12797 53320
rect 13987 53360 14045 53361
rect 13987 53320 13996 53360
rect 14036 53320 14045 53360
rect 13987 53319 14045 53320
rect 15147 53360 15189 53369
rect 15147 53320 15148 53360
rect 15188 53320 15189 53360
rect 3291 53301 3333 53310
rect 9099 53306 9141 53315
rect 15147 53311 15189 53320
rect 15243 53360 15285 53369
rect 15243 53320 15244 53360
rect 15284 53320 15285 53360
rect 15243 53311 15285 53320
rect 15723 53360 15765 53369
rect 15723 53320 15724 53360
rect 15764 53320 15765 53360
rect 15723 53311 15765 53320
rect 16195 53360 16253 53361
rect 16195 53320 16204 53360
rect 16244 53320 16253 53360
rect 16195 53319 16253 53320
rect 16683 53355 16725 53364
rect 16683 53315 16684 53355
rect 16724 53315 16725 53355
rect 18499 53360 18557 53361
rect 18499 53320 18508 53360
rect 18548 53320 18557 53360
rect 18499 53319 18557 53320
rect 19747 53360 19805 53361
rect 19747 53320 19756 53360
rect 19796 53320 19805 53360
rect 19747 53319 19805 53320
rect 16683 53306 16725 53315
rect 4299 53276 4341 53285
rect 4299 53236 4300 53276
rect 4340 53236 4341 53276
rect 4299 53227 4341 53236
rect 4395 53276 4437 53285
rect 4395 53236 4396 53276
rect 4436 53236 4437 53276
rect 4395 53227 4437 53236
rect 8043 53276 8085 53285
rect 8043 53236 8044 53276
rect 8084 53236 8085 53276
rect 8043 53227 8085 53236
rect 8139 53276 8181 53285
rect 8139 53236 8140 53276
rect 8180 53236 8181 53276
rect 8139 53227 8181 53236
rect 15627 53276 15669 53285
rect 15627 53236 15628 53276
rect 15668 53236 15669 53276
rect 15627 53227 15669 53236
rect 17251 53276 17309 53277
rect 17251 53236 17260 53276
rect 17300 53236 17309 53276
rect 17251 53235 17309 53236
rect 14187 53192 14229 53201
rect 14187 53152 14188 53192
rect 14228 53152 14229 53192
rect 14187 53143 14229 53152
rect 10923 53108 10965 53117
rect 10923 53068 10924 53108
rect 10964 53068 10965 53108
rect 10923 53059 10965 53068
rect 12555 53108 12597 53117
rect 12555 53068 12556 53108
rect 12596 53068 12597 53108
rect 12555 53059 12597 53068
rect 17067 53108 17109 53117
rect 17067 53068 17068 53108
rect 17108 53068 17109 53108
rect 17067 53059 17109 53068
rect 19947 53108 19989 53117
rect 19947 53068 19948 53108
rect 19988 53068 19989 53108
rect 19947 53059 19989 53068
rect 1152 52940 20352 52964
rect 1152 52900 3688 52940
rect 3728 52900 3770 52940
rect 3810 52900 3852 52940
rect 3892 52900 3934 52940
rect 3974 52900 4016 52940
rect 4056 52900 18808 52940
rect 18848 52900 18890 52940
rect 18930 52900 18972 52940
rect 19012 52900 19054 52940
rect 19094 52900 19136 52940
rect 19176 52900 20352 52940
rect 1152 52876 20352 52900
rect 1803 52772 1845 52781
rect 1803 52732 1804 52772
rect 1844 52732 1845 52772
rect 1803 52723 1845 52732
rect 1603 52604 1661 52605
rect 1603 52564 1612 52604
rect 1652 52564 1661 52604
rect 1603 52563 1661 52564
rect 1987 52604 2045 52605
rect 1987 52564 1996 52604
rect 2036 52564 2045 52604
rect 1987 52563 2045 52564
rect 10923 52604 10965 52613
rect 10923 52564 10924 52604
rect 10964 52564 10965 52604
rect 10923 52555 10965 52564
rect 19555 52604 19613 52605
rect 19555 52564 19564 52604
rect 19604 52564 19613 52604
rect 19555 52563 19613 52564
rect 19747 52604 19805 52605
rect 19747 52564 19756 52604
rect 19796 52564 19805 52604
rect 19747 52563 19805 52564
rect 8427 52534 8469 52543
rect 2371 52520 2429 52521
rect 2371 52480 2380 52520
rect 2420 52480 2429 52520
rect 2371 52479 2429 52480
rect 3619 52520 3677 52521
rect 3619 52480 3628 52520
rect 3668 52480 3677 52520
rect 3619 52479 3677 52480
rect 3811 52520 3869 52521
rect 3811 52480 3820 52520
rect 3860 52480 3869 52520
rect 3811 52479 3869 52480
rect 5059 52520 5117 52521
rect 5059 52480 5068 52520
rect 5108 52480 5117 52520
rect 5059 52479 5117 52480
rect 6891 52520 6933 52529
rect 6891 52480 6892 52520
rect 6932 52480 6933 52520
rect 6891 52471 6933 52480
rect 6987 52520 7029 52529
rect 6987 52480 6988 52520
rect 7028 52480 7029 52520
rect 6987 52471 7029 52480
rect 7371 52520 7413 52529
rect 7371 52480 7372 52520
rect 7412 52480 7413 52520
rect 7371 52471 7413 52480
rect 7467 52520 7509 52529
rect 7467 52480 7468 52520
rect 7508 52480 7509 52520
rect 7467 52471 7509 52480
rect 7939 52520 7997 52521
rect 7939 52480 7948 52520
rect 7988 52480 7997 52520
rect 8427 52494 8428 52534
rect 8468 52494 8469 52534
rect 11883 52534 11925 52543
rect 8427 52485 8469 52494
rect 10347 52520 10389 52529
rect 7939 52479 7997 52480
rect 10347 52480 10348 52520
rect 10388 52480 10389 52520
rect 10347 52471 10389 52480
rect 10443 52520 10485 52529
rect 10443 52480 10444 52520
rect 10484 52480 10485 52520
rect 10443 52471 10485 52480
rect 10827 52520 10869 52529
rect 10827 52480 10828 52520
rect 10868 52480 10869 52520
rect 10827 52471 10869 52480
rect 11395 52520 11453 52521
rect 11395 52480 11404 52520
rect 11444 52480 11453 52520
rect 11883 52494 11884 52534
rect 11924 52494 11925 52534
rect 14187 52534 14229 52543
rect 11883 52485 11925 52494
rect 12651 52520 12693 52529
rect 11395 52479 11453 52480
rect 12651 52480 12652 52520
rect 12692 52480 12693 52520
rect 12651 52471 12693 52480
rect 12747 52520 12789 52529
rect 12747 52480 12748 52520
rect 12788 52480 12789 52520
rect 12747 52471 12789 52480
rect 13131 52520 13173 52529
rect 13131 52480 13132 52520
rect 13172 52480 13173 52520
rect 13131 52471 13173 52480
rect 13227 52520 13269 52529
rect 13227 52480 13228 52520
rect 13268 52480 13269 52520
rect 13227 52471 13269 52480
rect 13718 52519 13760 52528
rect 13718 52479 13719 52519
rect 13759 52479 13760 52519
rect 14187 52494 14188 52534
rect 14228 52494 14229 52534
rect 14187 52485 14229 52494
rect 14563 52520 14621 52521
rect 14563 52480 14572 52520
rect 14612 52480 14621 52520
rect 14563 52479 14621 52480
rect 15811 52520 15869 52521
rect 15811 52480 15820 52520
rect 15860 52480 15869 52520
rect 15811 52479 15869 52480
rect 17443 52520 17501 52521
rect 17443 52480 17452 52520
rect 17492 52480 17501 52520
rect 17443 52479 17501 52480
rect 18691 52520 18749 52521
rect 18691 52480 18700 52520
rect 18740 52480 18749 52520
rect 18691 52479 18749 52480
rect 13718 52470 13760 52479
rect 8619 52436 8661 52445
rect 8619 52396 8620 52436
rect 8660 52396 8661 52436
rect 8619 52387 8661 52396
rect 12075 52436 12117 52445
rect 12075 52396 12076 52436
rect 12116 52396 12117 52436
rect 12075 52387 12117 52396
rect 14379 52436 14421 52445
rect 14379 52396 14380 52436
rect 14420 52396 14421 52436
rect 14379 52387 14421 52396
rect 1419 52352 1461 52361
rect 1419 52312 1420 52352
rect 1460 52312 1461 52352
rect 1419 52303 1461 52312
rect 2187 52352 2229 52361
rect 2187 52312 2188 52352
rect 2228 52312 2229 52352
rect 2187 52303 2229 52312
rect 5259 52352 5301 52361
rect 5259 52312 5260 52352
rect 5300 52312 5301 52352
rect 5259 52303 5301 52312
rect 16011 52352 16053 52361
rect 16011 52312 16012 52352
rect 16052 52312 16053 52352
rect 16011 52303 16053 52312
rect 18891 52352 18933 52361
rect 18891 52312 18892 52352
rect 18932 52312 18933 52352
rect 18891 52303 18933 52312
rect 19371 52352 19413 52361
rect 19371 52312 19372 52352
rect 19412 52312 19413 52352
rect 19371 52303 19413 52312
rect 19947 52352 19989 52361
rect 19947 52312 19948 52352
rect 19988 52312 19989 52352
rect 19947 52303 19989 52312
rect 1152 52184 20452 52208
rect 1152 52144 4928 52184
rect 4968 52144 5010 52184
rect 5050 52144 5092 52184
rect 5132 52144 5174 52184
rect 5214 52144 5256 52184
rect 5296 52144 20048 52184
rect 20088 52144 20130 52184
rect 20170 52144 20212 52184
rect 20252 52144 20294 52184
rect 20334 52144 20376 52184
rect 20416 52144 20452 52184
rect 1152 52120 20452 52144
rect 17451 52016 17493 52025
rect 17451 51976 17452 52016
rect 17492 51976 17493 52016
rect 17451 51967 17493 51976
rect 20043 52016 20085 52025
rect 20043 51976 20044 52016
rect 20084 51976 20085 52016
rect 20043 51967 20085 51976
rect 2379 51932 2421 51941
rect 2379 51892 2380 51932
rect 2420 51892 2421 51932
rect 2379 51883 2421 51892
rect 2571 51843 2613 51852
rect 2571 51803 2572 51843
rect 2612 51803 2613 51843
rect 3043 51848 3101 51849
rect 3043 51808 3052 51848
rect 3092 51808 3101 51848
rect 3043 51807 3101 51808
rect 3531 51848 3573 51857
rect 3531 51808 3532 51848
rect 3572 51808 3573 51848
rect 2571 51794 2613 51803
rect 3531 51799 3573 51808
rect 4011 51848 4053 51857
rect 4011 51808 4012 51848
rect 4052 51808 4053 51848
rect 4011 51799 4053 51808
rect 4107 51848 4149 51857
rect 4107 51808 4108 51848
rect 4148 51808 4149 51848
rect 4107 51799 4149 51808
rect 5923 51848 5981 51849
rect 5923 51808 5932 51848
rect 5972 51808 5981 51848
rect 5923 51807 5981 51808
rect 7171 51848 7229 51849
rect 7171 51808 7180 51848
rect 7220 51808 7229 51848
rect 7171 51807 7229 51808
rect 8611 51848 8669 51849
rect 8611 51808 8620 51848
rect 8660 51808 8669 51848
rect 8611 51807 8669 51808
rect 9859 51848 9917 51849
rect 9859 51808 9868 51848
rect 9908 51808 9917 51848
rect 9859 51807 9917 51808
rect 10243 51848 10301 51849
rect 10243 51808 10252 51848
rect 10292 51808 10301 51848
rect 10243 51807 10301 51808
rect 11491 51848 11549 51849
rect 11491 51808 11500 51848
rect 11540 51808 11549 51848
rect 11491 51807 11549 51808
rect 11875 51848 11933 51849
rect 11875 51808 11884 51848
rect 11924 51808 11933 51848
rect 11875 51807 11933 51808
rect 13123 51848 13181 51849
rect 13123 51808 13132 51848
rect 13172 51808 13181 51848
rect 13123 51807 13181 51808
rect 13507 51848 13565 51849
rect 13507 51808 13516 51848
rect 13556 51808 13565 51848
rect 13507 51807 13565 51808
rect 14755 51848 14813 51849
rect 14755 51808 14764 51848
rect 14804 51808 14813 51848
rect 14755 51807 14813 51808
rect 15723 51848 15765 51857
rect 15723 51808 15724 51848
rect 15764 51808 15765 51848
rect 15723 51799 15765 51808
rect 15819 51848 15861 51857
rect 15819 51808 15820 51848
rect 15860 51808 15861 51848
rect 15819 51799 15861 51808
rect 16299 51848 16341 51857
rect 16299 51808 16300 51848
rect 16340 51808 16341 51848
rect 16299 51799 16341 51808
rect 16771 51848 16829 51849
rect 16771 51808 16780 51848
rect 16820 51808 16829 51848
rect 18315 51848 18357 51857
rect 16771 51807 16829 51808
rect 17259 51834 17301 51843
rect 17259 51794 17260 51834
rect 17300 51794 17301 51834
rect 18315 51808 18316 51848
rect 18356 51808 18357 51848
rect 18315 51799 18357 51808
rect 18411 51848 18453 51857
rect 18411 51808 18412 51848
rect 18452 51808 18453 51848
rect 18411 51799 18453 51808
rect 18891 51848 18933 51857
rect 18891 51808 18892 51848
rect 18932 51808 18933 51848
rect 18891 51799 18933 51808
rect 19363 51848 19421 51849
rect 19363 51808 19372 51848
rect 19412 51808 19421 51848
rect 19363 51807 19421 51808
rect 19851 51843 19893 51852
rect 19851 51803 19852 51843
rect 19892 51803 19893 51843
rect 19851 51794 19893 51803
rect 17259 51785 17301 51794
rect 1699 51764 1757 51765
rect 1699 51724 1708 51764
rect 1748 51724 1757 51764
rect 1699 51723 1757 51724
rect 2083 51764 2141 51765
rect 2083 51724 2092 51764
rect 2132 51724 2141 51764
rect 2083 51723 2141 51724
rect 3627 51764 3669 51773
rect 3627 51724 3628 51764
rect 3668 51724 3669 51764
rect 3627 51715 3669 51724
rect 16203 51764 16245 51773
rect 16203 51724 16204 51764
rect 16244 51724 16245 51764
rect 16203 51715 16245 51724
rect 18795 51764 18837 51773
rect 18795 51724 18796 51764
rect 18836 51724 18837 51764
rect 18795 51715 18837 51724
rect 1515 51596 1557 51605
rect 1515 51556 1516 51596
rect 1556 51556 1557 51596
rect 1515 51547 1557 51556
rect 1899 51596 1941 51605
rect 1899 51556 1900 51596
rect 1940 51556 1941 51596
rect 1899 51547 1941 51556
rect 7371 51596 7413 51605
rect 7371 51556 7372 51596
rect 7412 51556 7413 51596
rect 7371 51547 7413 51556
rect 10059 51596 10101 51605
rect 10059 51556 10060 51596
rect 10100 51556 10101 51596
rect 10059 51547 10101 51556
rect 11691 51596 11733 51605
rect 11691 51556 11692 51596
rect 11732 51556 11733 51596
rect 11691 51547 11733 51556
rect 13323 51596 13365 51605
rect 13323 51556 13324 51596
rect 13364 51556 13365 51596
rect 13323 51547 13365 51556
rect 14955 51596 14997 51605
rect 14955 51556 14956 51596
rect 14996 51556 14997 51596
rect 14955 51547 14997 51556
rect 1152 51428 20352 51452
rect 1152 51388 3688 51428
rect 3728 51388 3770 51428
rect 3810 51388 3852 51428
rect 3892 51388 3934 51428
rect 3974 51388 4016 51428
rect 4056 51388 18808 51428
rect 18848 51388 18890 51428
rect 18930 51388 18972 51428
rect 19012 51388 19054 51428
rect 19094 51388 19136 51428
rect 19176 51388 20352 51428
rect 1152 51364 20352 51388
rect 2859 51260 2901 51269
rect 2859 51220 2860 51260
rect 2900 51220 2901 51260
rect 2859 51211 2901 51220
rect 12363 51260 12405 51269
rect 12363 51220 12364 51260
rect 12404 51220 12405 51260
rect 12363 51211 12405 51220
rect 17643 51260 17685 51269
rect 17643 51220 17644 51260
rect 17684 51220 17685 51260
rect 17643 51211 17685 51220
rect 3043 51092 3101 51093
rect 3043 51052 3052 51092
rect 3092 51052 3101 51092
rect 3043 51051 3101 51052
rect 5931 51092 5973 51101
rect 5931 51052 5932 51092
rect 5972 51052 5973 51092
rect 5931 51043 5973 51052
rect 8043 51092 8085 51101
rect 8043 51052 8044 51092
rect 8084 51052 8085 51092
rect 8043 51043 8085 51052
rect 12547 51092 12605 51093
rect 12547 51052 12556 51092
rect 12596 51052 12605 51092
rect 19747 51092 19805 51093
rect 12547 51051 12605 51052
rect 14811 51050 14853 51059
rect 19747 51052 19756 51092
rect 19796 51052 19805 51092
rect 19747 51051 19805 51052
rect 19939 51092 19997 51093
rect 19939 51052 19948 51092
rect 19988 51052 19997 51092
rect 19939 51051 19997 51052
rect 6891 51022 6933 51031
rect 11979 51022 12021 51031
rect 1219 51008 1277 51009
rect 1219 50968 1228 51008
rect 1268 50968 1277 51008
rect 1219 50967 1277 50968
rect 2467 51008 2525 51009
rect 2467 50968 2476 51008
rect 2516 50968 2525 51008
rect 2467 50967 2525 50968
rect 3331 51008 3389 51009
rect 3331 50968 3340 51008
rect 3380 50968 3389 51008
rect 3331 50967 3389 50968
rect 4579 51008 4637 51009
rect 4579 50968 4588 51008
rect 4628 50968 4637 51008
rect 4579 50967 4637 50968
rect 5355 51008 5397 51017
rect 5355 50968 5356 51008
rect 5396 50968 5397 51008
rect 5355 50959 5397 50968
rect 5451 51008 5493 51017
rect 5451 50968 5452 51008
rect 5492 50968 5493 51008
rect 5451 50959 5493 50968
rect 5835 51008 5877 51017
rect 5835 50968 5836 51008
rect 5876 50968 5877 51008
rect 5835 50959 5877 50968
rect 6403 51008 6461 51009
rect 6403 50968 6412 51008
rect 6452 50968 6461 51008
rect 6891 50982 6892 51022
rect 6932 50982 6933 51022
rect 6891 50973 6933 50982
rect 7563 51008 7605 51017
rect 6403 50967 6461 50968
rect 7563 50968 7564 51008
rect 7604 50968 7605 51008
rect 7563 50959 7605 50968
rect 7659 51008 7701 51017
rect 7659 50968 7660 51008
rect 7700 50968 7701 51008
rect 7659 50959 7701 50968
rect 8139 51008 8181 51017
rect 9099 51013 9141 51022
rect 8139 50968 8140 51008
rect 8180 50968 8181 51008
rect 8139 50959 8181 50968
rect 8611 51008 8669 51009
rect 8611 50968 8620 51008
rect 8660 50968 8669 51008
rect 8611 50967 8669 50968
rect 9099 50973 9100 51013
rect 9140 50973 9141 51013
rect 9099 50964 9141 50973
rect 10443 51008 10485 51017
rect 10443 50968 10444 51008
rect 10484 50968 10485 51008
rect 10443 50959 10485 50968
rect 10539 51008 10581 51017
rect 10539 50968 10540 51008
rect 10580 50968 10581 51008
rect 10539 50959 10581 50968
rect 10923 51008 10965 51017
rect 10923 50968 10924 51008
rect 10964 50968 10965 51008
rect 10923 50959 10965 50968
rect 11019 51008 11061 51017
rect 11019 50968 11020 51008
rect 11060 50968 11061 51008
rect 11019 50959 11061 50968
rect 11491 51008 11549 51009
rect 11491 50968 11500 51008
rect 11540 50968 11549 51008
rect 11979 50982 11980 51022
rect 12020 50982 12021 51022
rect 11979 50973 12021 50982
rect 13227 51008 13269 51017
rect 11491 50967 11549 50968
rect 13227 50968 13228 51008
rect 13268 50968 13269 51008
rect 13227 50959 13269 50968
rect 13323 51008 13365 51017
rect 13323 50968 13324 51008
rect 13364 50968 13365 51008
rect 13323 50959 13365 50968
rect 13707 51008 13749 51017
rect 13707 50968 13708 51008
rect 13748 50968 13749 51008
rect 13707 50959 13749 50968
rect 13803 51008 13845 51017
rect 14811 51010 14812 51050
rect 14852 51010 14853 51050
rect 13803 50968 13804 51008
rect 13844 50968 13845 51008
rect 13803 50959 13845 50968
rect 14275 51008 14333 51009
rect 14275 50968 14284 51008
rect 14324 50968 14333 51008
rect 14811 51001 14853 51010
rect 16195 51008 16253 51009
rect 14275 50967 14333 50968
rect 16195 50968 16204 51008
rect 16244 50968 16253 51008
rect 16195 50967 16253 50968
rect 17443 51008 17501 51009
rect 17443 50968 17452 51008
rect 17492 50968 17501 51008
rect 17443 50967 17501 50968
rect 17923 51008 17981 51009
rect 17923 50968 17932 51008
rect 17972 50968 17981 51008
rect 17923 50967 17981 50968
rect 19171 51008 19229 51009
rect 19171 50968 19180 51008
rect 19220 50968 19229 51008
rect 19171 50967 19229 50968
rect 9291 50924 9333 50933
rect 9291 50884 9292 50924
rect 9332 50884 9333 50924
rect 9291 50875 9333 50884
rect 12171 50924 12213 50933
rect 12171 50884 12172 50924
rect 12212 50884 12213 50924
rect 12171 50875 12213 50884
rect 2667 50840 2709 50849
rect 2667 50800 2668 50840
rect 2708 50800 2709 50840
rect 2667 50791 2709 50800
rect 4779 50840 4821 50849
rect 4779 50800 4780 50840
rect 4820 50800 4821 50840
rect 4779 50791 4821 50800
rect 7083 50840 7125 50849
rect 7083 50800 7084 50840
rect 7124 50800 7125 50840
rect 7083 50791 7125 50800
rect 14955 50840 14997 50849
rect 14955 50800 14956 50840
rect 14996 50800 14997 50840
rect 14955 50791 14997 50800
rect 19371 50840 19413 50849
rect 19371 50800 19372 50840
rect 19412 50800 19413 50840
rect 19371 50791 19413 50800
rect 19563 50840 19605 50849
rect 19563 50800 19564 50840
rect 19604 50800 19605 50840
rect 19563 50791 19605 50800
rect 20139 50840 20181 50849
rect 20139 50800 20140 50840
rect 20180 50800 20181 50840
rect 20139 50791 20181 50800
rect 1152 50672 20452 50696
rect 1152 50632 4928 50672
rect 4968 50632 5010 50672
rect 5050 50632 5092 50672
rect 5132 50632 5174 50672
rect 5214 50632 5256 50672
rect 5296 50632 20048 50672
rect 20088 50632 20130 50672
rect 20170 50632 20212 50672
rect 20252 50632 20294 50672
rect 20334 50632 20376 50672
rect 20416 50632 20452 50672
rect 1152 50608 20452 50632
rect 9003 50504 9045 50513
rect 9003 50464 9004 50504
rect 9044 50464 9045 50504
rect 9003 50455 9045 50464
rect 19275 50504 19317 50513
rect 19275 50464 19276 50504
rect 19316 50464 19317 50504
rect 19275 50455 19317 50464
rect 4683 50420 4725 50429
rect 4683 50380 4684 50420
rect 4724 50380 4725 50420
rect 4683 50371 4725 50380
rect 1411 50336 1469 50337
rect 1411 50296 1420 50336
rect 1460 50296 1469 50336
rect 1411 50295 1469 50296
rect 2659 50336 2717 50337
rect 2659 50296 2668 50336
rect 2708 50296 2717 50336
rect 2659 50295 2717 50296
rect 3043 50336 3101 50337
rect 3043 50296 3052 50336
rect 3092 50296 3101 50336
rect 3043 50295 3101 50296
rect 4291 50336 4349 50337
rect 4291 50296 4300 50336
rect 4340 50296 4349 50336
rect 5347 50336 5405 50337
rect 4291 50295 4349 50296
rect 4875 50322 4917 50331
rect 4875 50282 4876 50322
rect 4916 50282 4917 50322
rect 5347 50296 5356 50336
rect 5396 50296 5405 50336
rect 5347 50295 5405 50296
rect 6315 50336 6357 50345
rect 6315 50296 6316 50336
rect 6356 50296 6357 50336
rect 6315 50287 6357 50296
rect 6411 50336 6453 50345
rect 6411 50296 6412 50336
rect 6452 50296 6453 50336
rect 6411 50287 6453 50296
rect 7555 50336 7613 50337
rect 7555 50296 7564 50336
rect 7604 50296 7613 50336
rect 7555 50295 7613 50296
rect 8803 50336 8861 50337
rect 8803 50296 8812 50336
rect 8852 50296 8861 50336
rect 8803 50295 8861 50296
rect 9187 50336 9245 50337
rect 9187 50296 9196 50336
rect 9236 50296 9245 50336
rect 9187 50295 9245 50296
rect 10435 50336 10493 50337
rect 10435 50296 10444 50336
rect 10484 50296 10493 50336
rect 10435 50295 10493 50296
rect 11587 50336 11645 50337
rect 11587 50296 11596 50336
rect 11636 50296 11645 50336
rect 11587 50295 11645 50296
rect 12835 50336 12893 50337
rect 12835 50296 12844 50336
rect 12884 50296 12893 50336
rect 12835 50295 12893 50296
rect 13987 50336 14045 50337
rect 13987 50296 13996 50336
rect 14036 50296 14045 50336
rect 13987 50295 14045 50296
rect 15235 50336 15293 50337
rect 15235 50296 15244 50336
rect 15284 50296 15293 50336
rect 15235 50295 15293 50296
rect 17155 50336 17213 50337
rect 17155 50296 17164 50336
rect 17204 50296 17213 50336
rect 17155 50295 17213 50296
rect 17547 50336 17589 50345
rect 17547 50296 17548 50336
rect 17588 50296 17589 50336
rect 17547 50287 17589 50296
rect 17643 50336 17685 50345
rect 17643 50296 17644 50336
rect 17684 50296 17685 50336
rect 17643 50287 17685 50296
rect 18123 50336 18165 50345
rect 18123 50296 18124 50336
rect 18164 50296 18165 50336
rect 18123 50287 18165 50296
rect 18595 50336 18653 50337
rect 18595 50296 18604 50336
rect 18644 50296 18653 50336
rect 18595 50295 18653 50296
rect 19131 50326 19173 50335
rect 4875 50273 4917 50282
rect 19131 50286 19132 50326
rect 19172 50286 19173 50326
rect 19131 50277 19173 50286
rect 5835 50252 5877 50261
rect 5835 50212 5836 50252
rect 5876 50212 5877 50252
rect 5835 50203 5877 50212
rect 5931 50252 5973 50261
rect 5931 50212 5932 50252
rect 5972 50212 5973 50252
rect 5931 50203 5973 50212
rect 13411 50252 13469 50253
rect 13411 50212 13420 50252
rect 13460 50212 13469 50252
rect 13411 50211 13469 50212
rect 16003 50252 16061 50253
rect 16003 50212 16012 50252
rect 16052 50212 16061 50252
rect 16003 50211 16061 50212
rect 18027 50252 18069 50261
rect 18027 50212 18028 50252
rect 18068 50212 18069 50252
rect 18027 50203 18069 50212
rect 19459 50252 19517 50253
rect 19459 50212 19468 50252
rect 19508 50212 19517 50252
rect 19459 50211 19517 50212
rect 19843 50252 19901 50253
rect 19843 50212 19852 50252
rect 19892 50212 19901 50252
rect 19843 50211 19901 50212
rect 13227 50168 13269 50177
rect 13227 50128 13228 50168
rect 13268 50128 13269 50168
rect 13227 50119 13269 50128
rect 20043 50168 20085 50177
rect 20043 50128 20044 50168
rect 20084 50128 20085 50168
rect 20043 50119 20085 50128
rect 2859 50084 2901 50093
rect 2859 50044 2860 50084
rect 2900 50044 2901 50084
rect 2859 50035 2901 50044
rect 4491 50084 4533 50093
rect 4491 50044 4492 50084
rect 4532 50044 4533 50084
rect 4491 50035 4533 50044
rect 10635 50084 10677 50093
rect 10635 50044 10636 50084
rect 10676 50044 10677 50084
rect 10635 50035 10677 50044
rect 13035 50084 13077 50093
rect 13035 50044 13036 50084
rect 13076 50044 13077 50084
rect 13035 50035 13077 50044
rect 15435 50084 15477 50093
rect 15435 50044 15436 50084
rect 15476 50044 15477 50084
rect 15435 50035 15477 50044
rect 15819 50084 15861 50093
rect 15819 50044 15820 50084
rect 15860 50044 15861 50084
rect 15819 50035 15861 50044
rect 16491 50084 16533 50093
rect 16491 50044 16492 50084
rect 16532 50044 16533 50084
rect 16491 50035 16533 50044
rect 19659 50084 19701 50093
rect 19659 50044 19660 50084
rect 19700 50044 19701 50084
rect 19659 50035 19701 50044
rect 1152 49916 20352 49940
rect 1152 49876 3688 49916
rect 3728 49876 3770 49916
rect 3810 49876 3852 49916
rect 3892 49876 3934 49916
rect 3974 49876 4016 49916
rect 4056 49876 18808 49916
rect 18848 49876 18890 49916
rect 18930 49876 18972 49916
rect 19012 49876 19054 49916
rect 19094 49876 19136 49916
rect 19176 49876 20352 49916
rect 1152 49852 20352 49876
rect 1899 49748 1941 49757
rect 1899 49708 1900 49748
rect 1940 49708 1941 49748
rect 1899 49699 1941 49708
rect 7275 49748 7317 49757
rect 7275 49708 7276 49748
rect 7316 49708 7317 49748
rect 7275 49699 7317 49708
rect 17259 49748 17301 49757
rect 17259 49708 17260 49748
rect 17300 49708 17301 49748
rect 17259 49699 17301 49708
rect 18987 49748 19029 49757
rect 18987 49708 18988 49748
rect 19028 49708 19029 49748
rect 18987 49699 19029 49708
rect 11307 49664 11349 49673
rect 11307 49624 11308 49664
rect 11348 49624 11349 49664
rect 11307 49615 11349 49624
rect 1699 49580 1757 49581
rect 1699 49540 1708 49580
rect 1748 49540 1757 49580
rect 1699 49539 1757 49540
rect 2083 49580 2141 49581
rect 2083 49540 2092 49580
rect 2132 49540 2141 49580
rect 2083 49539 2141 49540
rect 3435 49580 3477 49589
rect 3435 49540 3436 49580
rect 3476 49540 3477 49580
rect 3435 49531 3477 49540
rect 3531 49580 3573 49589
rect 3531 49540 3532 49580
rect 3572 49540 3573 49580
rect 3531 49531 3573 49540
rect 12075 49580 12117 49589
rect 12075 49540 12076 49580
rect 12116 49540 12117 49580
rect 12075 49531 12117 49540
rect 12171 49580 12213 49589
rect 12171 49540 12172 49580
rect 12212 49540 12213 49580
rect 12171 49531 12213 49540
rect 15915 49580 15957 49589
rect 15915 49540 15916 49580
rect 15956 49540 15957 49580
rect 15915 49531 15957 49540
rect 19171 49580 19229 49581
rect 19171 49540 19180 49580
rect 19220 49540 19229 49580
rect 19171 49539 19229 49540
rect 19363 49580 19421 49581
rect 19363 49540 19372 49580
rect 19412 49540 19421 49580
rect 19363 49539 19421 49540
rect 19747 49580 19805 49581
rect 19747 49540 19756 49580
rect 19796 49540 19805 49580
rect 19747 49539 19805 49540
rect 2475 49510 2517 49519
rect 2475 49470 2476 49510
rect 2516 49470 2517 49510
rect 13131 49510 13173 49519
rect 2475 49461 2517 49470
rect 2947 49496 3005 49497
rect 2947 49456 2956 49496
rect 2996 49456 3005 49496
rect 2947 49455 3005 49456
rect 3915 49496 3957 49505
rect 3915 49456 3916 49496
rect 3956 49456 3957 49496
rect 3915 49447 3957 49456
rect 4011 49496 4053 49505
rect 4011 49456 4012 49496
rect 4052 49456 4053 49496
rect 4011 49447 4053 49456
rect 5827 49496 5885 49497
rect 5827 49456 5836 49496
rect 5876 49456 5885 49496
rect 5827 49455 5885 49456
rect 7075 49496 7133 49497
rect 7075 49456 7084 49496
rect 7124 49456 7133 49496
rect 7075 49455 7133 49456
rect 7459 49496 7517 49497
rect 7459 49456 7468 49496
rect 7508 49456 7517 49496
rect 7459 49455 7517 49456
rect 8707 49496 8765 49497
rect 8707 49456 8716 49496
rect 8756 49456 8765 49496
rect 8707 49455 8765 49456
rect 9859 49496 9917 49497
rect 9859 49456 9868 49496
rect 9908 49456 9917 49496
rect 9859 49455 9917 49456
rect 11107 49496 11165 49497
rect 11107 49456 11116 49496
rect 11156 49456 11165 49496
rect 11107 49455 11165 49456
rect 11595 49496 11637 49505
rect 11595 49456 11596 49496
rect 11636 49456 11637 49496
rect 11595 49447 11637 49456
rect 11691 49496 11733 49505
rect 11691 49456 11692 49496
rect 11732 49456 11733 49496
rect 11691 49447 11733 49456
rect 12643 49496 12701 49497
rect 12643 49456 12652 49496
rect 12692 49456 12701 49496
rect 13131 49470 13132 49510
rect 13172 49470 13173 49510
rect 16923 49505 16965 49514
rect 13131 49461 13173 49470
rect 13507 49496 13565 49497
rect 12643 49455 12701 49456
rect 13507 49456 13516 49496
rect 13556 49456 13565 49496
rect 13507 49455 13565 49456
rect 14755 49496 14813 49497
rect 14755 49456 14764 49496
rect 14804 49456 14813 49496
rect 14755 49455 14813 49456
rect 15339 49496 15381 49505
rect 15339 49456 15340 49496
rect 15380 49456 15381 49496
rect 15819 49496 15861 49505
rect 15339 49447 15381 49456
rect 15435 49476 15477 49485
rect 15435 49436 15436 49476
rect 15476 49436 15477 49476
rect 15819 49456 15820 49496
rect 15860 49456 15861 49496
rect 15819 49447 15861 49456
rect 16387 49496 16445 49497
rect 16387 49456 16396 49496
rect 16436 49456 16445 49496
rect 16923 49465 16924 49505
rect 16964 49465 16965 49505
rect 16923 49456 16965 49465
rect 17443 49496 17501 49497
rect 17443 49456 17452 49496
rect 17492 49456 17501 49496
rect 16387 49455 16445 49456
rect 17443 49455 17501 49456
rect 18691 49496 18749 49497
rect 18691 49456 18700 49496
rect 18740 49456 18749 49496
rect 18691 49455 18749 49456
rect 15435 49427 15477 49436
rect 2283 49412 2325 49421
rect 2283 49372 2284 49412
rect 2324 49372 2325 49412
rect 2283 49363 2325 49372
rect 13323 49412 13365 49421
rect 13323 49372 13324 49412
rect 13364 49372 13365 49412
rect 13323 49363 13365 49372
rect 17067 49412 17109 49421
rect 17067 49372 17068 49412
rect 17108 49372 17109 49412
rect 17067 49363 17109 49372
rect 1515 49328 1557 49337
rect 1515 49288 1516 49328
rect 1556 49288 1557 49328
rect 1515 49279 1557 49288
rect 8907 49328 8949 49337
rect 8907 49288 8908 49328
rect 8948 49288 8949 49328
rect 8907 49279 8949 49288
rect 14955 49328 14997 49337
rect 14955 49288 14956 49328
rect 14996 49288 14997 49328
rect 14955 49279 14997 49288
rect 19563 49328 19605 49337
rect 19563 49288 19564 49328
rect 19604 49288 19605 49328
rect 19563 49279 19605 49288
rect 19947 49328 19989 49337
rect 19947 49288 19948 49328
rect 19988 49288 19989 49328
rect 19947 49279 19989 49288
rect 1152 49160 20452 49184
rect 1152 49120 4928 49160
rect 4968 49120 5010 49160
rect 5050 49120 5092 49160
rect 5132 49120 5174 49160
rect 5214 49120 5256 49160
rect 5296 49120 20048 49160
rect 20088 49120 20130 49160
rect 20170 49120 20212 49160
rect 20252 49120 20294 49160
rect 20334 49120 20376 49160
rect 20416 49120 20452 49160
rect 1152 49096 20452 49120
rect 2859 48992 2901 49001
rect 2859 48952 2860 48992
rect 2900 48952 2901 48992
rect 2859 48943 2901 48952
rect 14955 48992 14997 49001
rect 14955 48952 14956 48992
rect 14996 48952 14997 48992
rect 14955 48943 14997 48952
rect 17067 48992 17109 49001
rect 17067 48952 17068 48992
rect 17108 48952 17109 48992
rect 17067 48943 17109 48952
rect 19755 48992 19797 49001
rect 19755 48952 19756 48992
rect 19796 48952 19797 48992
rect 19755 48943 19797 48952
rect 10539 48908 10581 48917
rect 10539 48868 10540 48908
rect 10580 48868 10581 48908
rect 10539 48859 10581 48868
rect 12939 48908 12981 48917
rect 12939 48868 12940 48908
rect 12980 48868 12981 48908
rect 12939 48859 12981 48868
rect 1219 48824 1277 48825
rect 1219 48784 1228 48824
rect 1268 48784 1277 48824
rect 1219 48783 1277 48784
rect 2467 48824 2525 48825
rect 2467 48784 2476 48824
rect 2516 48784 2525 48824
rect 2467 48783 2525 48784
rect 3427 48824 3485 48825
rect 3427 48784 3436 48824
rect 3476 48784 3485 48824
rect 3427 48783 3485 48784
rect 4675 48824 4733 48825
rect 4675 48784 4684 48824
rect 4724 48784 4733 48824
rect 4675 48783 4733 48784
rect 5059 48824 5117 48825
rect 5059 48784 5068 48824
rect 5108 48784 5117 48824
rect 5059 48783 5117 48784
rect 6307 48824 6365 48825
rect 6307 48784 6316 48824
rect 6356 48784 6365 48824
rect 6307 48783 6365 48784
rect 6787 48824 6845 48825
rect 6787 48784 6796 48824
rect 6836 48784 6845 48824
rect 6787 48783 6845 48784
rect 8035 48824 8093 48825
rect 8035 48784 8044 48824
rect 8084 48784 8093 48824
rect 8035 48783 8093 48784
rect 8811 48824 8853 48833
rect 8811 48784 8812 48824
rect 8852 48784 8853 48824
rect 8811 48775 8853 48784
rect 8907 48824 8949 48833
rect 8907 48784 8908 48824
rect 8948 48784 8949 48824
rect 8907 48775 8949 48784
rect 9291 48824 9333 48833
rect 9291 48784 9292 48824
rect 9332 48784 9333 48824
rect 9291 48775 9333 48784
rect 9387 48824 9429 48833
rect 9387 48784 9388 48824
rect 9428 48784 9429 48824
rect 9387 48775 9429 48784
rect 9859 48824 9917 48825
rect 9859 48784 9868 48824
rect 9908 48784 9917 48824
rect 11491 48824 11549 48825
rect 9859 48783 9917 48784
rect 10395 48814 10437 48823
rect 10395 48774 10396 48814
rect 10436 48774 10437 48814
rect 11491 48784 11500 48824
rect 11540 48784 11549 48824
rect 11491 48783 11549 48784
rect 12739 48824 12797 48825
rect 12739 48784 12748 48824
rect 12788 48784 12797 48824
rect 12739 48783 12797 48784
rect 13227 48824 13269 48833
rect 13227 48784 13228 48824
rect 13268 48784 13269 48824
rect 13227 48775 13269 48784
rect 13323 48824 13365 48833
rect 13323 48784 13324 48824
rect 13364 48784 13365 48824
rect 13323 48775 13365 48784
rect 14275 48824 14333 48825
rect 14275 48784 14284 48824
rect 14324 48784 14333 48824
rect 15619 48824 15677 48825
rect 14275 48783 14333 48784
rect 14811 48814 14853 48823
rect 10395 48765 10437 48774
rect 14811 48774 14812 48814
rect 14852 48774 14853 48814
rect 15619 48784 15628 48824
rect 15668 48784 15677 48824
rect 15619 48783 15677 48784
rect 16867 48824 16925 48825
rect 16867 48784 16876 48824
rect 16916 48784 16925 48824
rect 16867 48783 16925 48784
rect 18027 48824 18069 48833
rect 18027 48784 18028 48824
rect 18068 48784 18069 48824
rect 18027 48775 18069 48784
rect 18123 48824 18165 48833
rect 18123 48784 18124 48824
rect 18164 48784 18165 48824
rect 18123 48775 18165 48784
rect 18603 48824 18645 48833
rect 18603 48784 18604 48824
rect 18644 48784 18645 48824
rect 18603 48775 18645 48784
rect 19075 48824 19133 48825
rect 19075 48784 19084 48824
rect 19124 48784 19133 48824
rect 19075 48783 19133 48784
rect 19611 48782 19653 48791
rect 14811 48765 14853 48774
rect 3043 48740 3101 48741
rect 3043 48700 3052 48740
rect 3092 48700 3101 48740
rect 3043 48699 3101 48700
rect 13707 48740 13749 48749
rect 13707 48700 13708 48740
rect 13748 48700 13749 48740
rect 13707 48691 13749 48700
rect 13803 48740 13845 48749
rect 13803 48700 13804 48740
rect 13844 48700 13845 48740
rect 13803 48691 13845 48700
rect 18507 48740 18549 48749
rect 18507 48700 18508 48740
rect 18548 48700 18549 48740
rect 19611 48742 19612 48782
rect 19652 48742 19653 48782
rect 19611 48733 19653 48742
rect 19939 48740 19997 48741
rect 18507 48691 18549 48700
rect 19939 48700 19948 48740
rect 19988 48700 19997 48740
rect 19939 48699 19997 48700
rect 2667 48572 2709 48581
rect 2667 48532 2668 48572
rect 2708 48532 2709 48572
rect 2667 48523 2709 48532
rect 4875 48572 4917 48581
rect 4875 48532 4876 48572
rect 4916 48532 4917 48572
rect 4875 48523 4917 48532
rect 6507 48572 6549 48581
rect 6507 48532 6508 48572
rect 6548 48532 6549 48572
rect 6507 48523 6549 48532
rect 8235 48572 8277 48581
rect 8235 48532 8236 48572
rect 8276 48532 8277 48572
rect 8235 48523 8277 48532
rect 20139 48572 20181 48581
rect 20139 48532 20140 48572
rect 20180 48532 20181 48572
rect 20139 48523 20181 48532
rect 1152 48404 20352 48428
rect 1152 48364 3688 48404
rect 3728 48364 3770 48404
rect 3810 48364 3852 48404
rect 3892 48364 3934 48404
rect 3974 48364 4016 48404
rect 4056 48364 18808 48404
rect 18848 48364 18890 48404
rect 18930 48364 18972 48404
rect 19012 48364 19054 48404
rect 19094 48364 19136 48404
rect 19176 48364 20352 48404
rect 1152 48340 20352 48364
rect 1611 48236 1653 48245
rect 1611 48196 1612 48236
rect 1652 48196 1653 48236
rect 1611 48187 1653 48196
rect 16203 48236 16245 48245
rect 16203 48196 16204 48236
rect 16244 48196 16245 48236
rect 16203 48187 16245 48196
rect 18027 48236 18069 48245
rect 18027 48196 18028 48236
rect 18068 48196 18069 48236
rect 18027 48187 18069 48196
rect 19659 48236 19701 48245
rect 19659 48196 19660 48236
rect 19700 48196 19701 48236
rect 19659 48187 19701 48196
rect 1795 48068 1853 48069
rect 1795 48028 1804 48068
rect 1844 48028 1853 48068
rect 1795 48027 1853 48028
rect 6411 48068 6453 48077
rect 6411 48028 6412 48068
rect 6452 48028 6453 48068
rect 6411 48019 6453 48028
rect 6507 48068 6549 48077
rect 6507 48028 6508 48068
rect 6548 48028 6549 48068
rect 6507 48019 6549 48028
rect 8907 48068 8949 48077
rect 8907 48028 8908 48068
rect 8948 48028 8949 48068
rect 8907 48019 8949 48028
rect 9003 48068 9045 48077
rect 9003 48028 9004 48068
rect 9044 48028 9045 48068
rect 9003 48019 9045 48028
rect 16387 48068 16445 48069
rect 16387 48028 16396 48068
rect 16436 48028 16445 48068
rect 16387 48027 16445 48028
rect 19843 48068 19901 48069
rect 19843 48028 19852 48068
rect 19892 48028 19901 48068
rect 19843 48027 19901 48028
rect 5451 47989 5493 47998
rect 1987 47984 2045 47985
rect 1987 47944 1996 47984
rect 2036 47944 2045 47984
rect 1987 47943 2045 47944
rect 3235 47984 3293 47985
rect 3235 47944 3244 47984
rect 3284 47944 3293 47984
rect 3235 47943 3293 47944
rect 3619 47984 3677 47985
rect 3619 47944 3628 47984
rect 3668 47944 3677 47984
rect 3619 47943 3677 47944
rect 4867 47984 4925 47985
rect 4867 47944 4876 47984
rect 4916 47944 4925 47984
rect 4867 47943 4925 47944
rect 5451 47949 5452 47989
rect 5492 47949 5493 47989
rect 5451 47940 5493 47949
rect 5923 47984 5981 47985
rect 5923 47944 5932 47984
rect 5972 47944 5981 47984
rect 5923 47943 5981 47944
rect 6891 47984 6933 47993
rect 6891 47944 6892 47984
rect 6932 47944 6933 47984
rect 6891 47935 6933 47944
rect 6987 47984 7029 47993
rect 6987 47944 6988 47984
rect 7028 47944 7029 47984
rect 6987 47935 7029 47944
rect 7947 47989 7989 47998
rect 7947 47949 7948 47989
rect 7988 47949 7989 47989
rect 7947 47940 7989 47949
rect 8419 47984 8477 47985
rect 8419 47944 8428 47984
rect 8468 47944 8477 47984
rect 8419 47943 8477 47944
rect 9387 47984 9429 47993
rect 9387 47944 9388 47984
rect 9428 47944 9429 47984
rect 9387 47935 9429 47944
rect 9483 47984 9525 47993
rect 9483 47944 9484 47984
rect 9524 47944 9525 47984
rect 9483 47935 9525 47944
rect 10243 47984 10301 47985
rect 10243 47944 10252 47984
rect 10292 47944 10301 47984
rect 10243 47943 10301 47944
rect 11491 47984 11549 47985
rect 11491 47944 11500 47984
rect 11540 47944 11549 47984
rect 11491 47943 11549 47944
rect 13603 47984 13661 47985
rect 13603 47944 13612 47984
rect 13652 47944 13661 47984
rect 13603 47943 13661 47944
rect 14851 47984 14909 47985
rect 14851 47944 14860 47984
rect 14900 47944 14909 47984
rect 14851 47943 14909 47944
rect 16579 47984 16637 47985
rect 16579 47944 16588 47984
rect 16628 47944 16637 47984
rect 16579 47943 16637 47944
rect 17827 47984 17885 47985
rect 17827 47944 17836 47984
rect 17876 47944 17885 47984
rect 17827 47943 17885 47944
rect 18211 47984 18269 47985
rect 18211 47944 18220 47984
rect 18260 47944 18269 47984
rect 18211 47943 18269 47944
rect 19459 47984 19517 47985
rect 19459 47944 19468 47984
rect 19508 47944 19517 47984
rect 19459 47943 19517 47944
rect 5067 47900 5109 47909
rect 5067 47860 5068 47900
rect 5108 47860 5109 47900
rect 5067 47851 5109 47860
rect 5259 47900 5301 47909
rect 5259 47860 5260 47900
rect 5300 47860 5301 47900
rect 5259 47851 5301 47860
rect 7755 47900 7797 47909
rect 7755 47860 7756 47900
rect 7796 47860 7797 47900
rect 7755 47851 7797 47860
rect 3435 47816 3477 47825
rect 3435 47776 3436 47816
rect 3476 47776 3477 47816
rect 3435 47767 3477 47776
rect 11691 47816 11733 47825
rect 11691 47776 11692 47816
rect 11732 47776 11733 47816
rect 11691 47767 11733 47776
rect 15051 47816 15093 47825
rect 15051 47776 15052 47816
rect 15092 47776 15093 47816
rect 15051 47767 15093 47776
rect 20043 47816 20085 47825
rect 20043 47776 20044 47816
rect 20084 47776 20085 47816
rect 20043 47767 20085 47776
rect 1152 47648 20452 47672
rect 1152 47608 4928 47648
rect 4968 47608 5010 47648
rect 5050 47608 5092 47648
rect 5132 47608 5174 47648
rect 5214 47608 5256 47648
rect 5296 47608 20048 47648
rect 20088 47608 20130 47648
rect 20170 47608 20212 47648
rect 20252 47608 20294 47648
rect 20334 47608 20376 47648
rect 20416 47608 20452 47648
rect 1152 47584 20452 47608
rect 1803 47480 1845 47489
rect 1803 47440 1804 47480
rect 1844 47440 1845 47480
rect 1803 47431 1845 47440
rect 6699 47480 6741 47489
rect 6699 47440 6700 47480
rect 6740 47440 6741 47480
rect 6699 47431 6741 47440
rect 8043 47480 8085 47489
rect 8043 47440 8044 47480
rect 8084 47440 8085 47480
rect 8043 47431 8085 47440
rect 10635 47480 10677 47489
rect 10635 47440 10636 47480
rect 10676 47440 10677 47480
rect 10635 47431 10677 47440
rect 16779 47480 16821 47489
rect 16779 47440 16780 47480
rect 16820 47440 16821 47480
rect 16779 47431 16821 47440
rect 4011 47396 4053 47405
rect 4011 47356 4012 47396
rect 4052 47356 4053 47396
rect 4011 47347 4053 47356
rect 2283 47312 2325 47321
rect 2283 47272 2284 47312
rect 2324 47272 2325 47312
rect 2283 47263 2325 47272
rect 2379 47312 2421 47321
rect 2379 47272 2380 47312
rect 2420 47272 2421 47312
rect 2379 47263 2421 47272
rect 2859 47312 2901 47321
rect 2859 47272 2860 47312
rect 2900 47272 2901 47312
rect 2859 47263 2901 47272
rect 3331 47312 3389 47313
rect 3331 47272 3340 47312
rect 3380 47272 3389 47312
rect 3331 47271 3389 47272
rect 3819 47307 3861 47316
rect 3819 47267 3820 47307
rect 3860 47267 3861 47307
rect 3819 47258 3861 47267
rect 4971 47312 5013 47321
rect 4971 47272 4972 47312
rect 5012 47272 5013 47312
rect 4971 47263 5013 47272
rect 5067 47312 5109 47321
rect 5067 47272 5068 47312
rect 5108 47272 5109 47312
rect 5067 47263 5109 47272
rect 5451 47312 5493 47321
rect 5451 47272 5452 47312
rect 5492 47272 5493 47312
rect 5451 47263 5493 47272
rect 5547 47312 5589 47321
rect 5547 47272 5548 47312
rect 5588 47272 5589 47312
rect 5547 47263 5589 47272
rect 6019 47312 6077 47313
rect 6019 47272 6028 47312
rect 6068 47272 6077 47312
rect 8227 47312 8285 47313
rect 6019 47271 6077 47272
rect 6555 47302 6597 47311
rect 6555 47262 6556 47302
rect 6596 47262 6597 47302
rect 8227 47272 8236 47312
rect 8276 47272 8285 47312
rect 8227 47271 8285 47272
rect 9475 47312 9533 47313
rect 9475 47272 9484 47312
rect 9524 47272 9533 47312
rect 9475 47271 9533 47272
rect 11107 47312 11165 47313
rect 11107 47272 11116 47312
rect 11156 47272 11165 47312
rect 11107 47271 11165 47272
rect 12355 47312 12413 47313
rect 12355 47272 12364 47312
rect 12404 47272 12413 47312
rect 12355 47271 12413 47272
rect 12739 47312 12797 47313
rect 12739 47272 12748 47312
rect 12788 47272 12797 47312
rect 12739 47271 12797 47272
rect 13987 47312 14045 47313
rect 13987 47272 13996 47312
rect 14036 47272 14045 47312
rect 13987 47271 14045 47272
rect 15051 47312 15093 47321
rect 15051 47272 15052 47312
rect 15092 47272 15093 47312
rect 15051 47263 15093 47272
rect 15147 47312 15189 47321
rect 15147 47272 15148 47312
rect 15188 47272 15189 47312
rect 15147 47263 15189 47272
rect 15531 47312 15573 47321
rect 15531 47272 15532 47312
rect 15572 47272 15573 47312
rect 15531 47263 15573 47272
rect 15627 47312 15669 47321
rect 15627 47272 15628 47312
rect 15668 47272 15669 47312
rect 15627 47263 15669 47272
rect 16099 47312 16157 47313
rect 16099 47272 16108 47312
rect 16148 47272 16157 47312
rect 16963 47312 17021 47313
rect 16099 47271 16157 47272
rect 16635 47270 16677 47279
rect 16963 47272 16972 47312
rect 17012 47272 17021 47312
rect 16963 47271 17021 47272
rect 18211 47312 18269 47313
rect 18211 47272 18220 47312
rect 18260 47272 18269 47312
rect 18211 47271 18269 47272
rect 18595 47312 18653 47313
rect 18595 47272 18604 47312
rect 18644 47272 18653 47312
rect 18595 47271 18653 47272
rect 19843 47312 19901 47313
rect 19843 47272 19852 47312
rect 19892 47272 19901 47312
rect 19843 47271 19901 47272
rect 6555 47253 6597 47262
rect 1987 47228 2045 47229
rect 1987 47188 1996 47228
rect 2036 47188 2045 47228
rect 1987 47187 2045 47188
rect 2763 47228 2805 47237
rect 16635 47230 16636 47270
rect 16676 47230 16677 47270
rect 2763 47188 2764 47228
rect 2804 47188 2805 47228
rect 2763 47179 2805 47188
rect 10819 47228 10877 47229
rect 10819 47188 10828 47228
rect 10868 47188 10877 47228
rect 16635 47221 16677 47230
rect 10819 47187 10877 47188
rect 12555 47060 12597 47069
rect 12555 47020 12556 47060
rect 12596 47020 12597 47060
rect 12555 47011 12597 47020
rect 14187 47060 14229 47069
rect 14187 47020 14188 47060
rect 14228 47020 14229 47060
rect 14187 47011 14229 47020
rect 18411 47060 18453 47069
rect 18411 47020 18412 47060
rect 18452 47020 18453 47060
rect 18411 47011 18453 47020
rect 20043 47060 20085 47069
rect 20043 47020 20044 47060
rect 20084 47020 20085 47060
rect 20043 47011 20085 47020
rect 1152 46892 20352 46916
rect 1152 46852 3688 46892
rect 3728 46852 3770 46892
rect 3810 46852 3852 46892
rect 3892 46852 3934 46892
rect 3974 46852 4016 46892
rect 4056 46852 18808 46892
rect 18848 46852 18890 46892
rect 18930 46852 18972 46892
rect 19012 46852 19054 46892
rect 19094 46852 19136 46892
rect 19176 46852 20352 46892
rect 1152 46828 20352 46852
rect 16683 46724 16725 46733
rect 16683 46684 16684 46724
rect 16724 46684 16725 46724
rect 16683 46675 16725 46684
rect 5931 46640 5973 46649
rect 5931 46600 5932 46640
rect 5972 46600 5973 46640
rect 5931 46591 5973 46600
rect 11875 46556 11933 46557
rect 11875 46516 11884 46556
rect 11924 46516 11933 46556
rect 11875 46515 11933 46516
rect 13131 46556 13173 46565
rect 13131 46516 13132 46556
rect 13172 46516 13173 46556
rect 18411 46556 18453 46565
rect 13131 46507 13173 46516
rect 14139 46514 14181 46523
rect 11451 46481 11493 46490
rect 1219 46472 1277 46473
rect 1219 46432 1228 46472
rect 1268 46432 1277 46472
rect 1219 46431 1277 46432
rect 2467 46472 2525 46473
rect 2467 46432 2476 46472
rect 2516 46432 2525 46472
rect 2467 46431 2525 46432
rect 4483 46472 4541 46473
rect 4483 46432 4492 46472
rect 4532 46432 4541 46472
rect 4483 46431 4541 46432
rect 5731 46472 5789 46473
rect 5731 46432 5740 46472
rect 5780 46432 5789 46472
rect 5731 46431 5789 46432
rect 6115 46472 6173 46473
rect 6115 46432 6124 46472
rect 6164 46432 6173 46472
rect 6115 46431 6173 46432
rect 7363 46472 7421 46473
rect 7363 46432 7372 46472
rect 7412 46432 7421 46472
rect 7363 46431 7421 46432
rect 8131 46472 8189 46473
rect 8131 46432 8140 46472
rect 8180 46432 8189 46472
rect 8131 46431 8189 46432
rect 9379 46472 9437 46473
rect 9379 46432 9388 46472
rect 9428 46432 9437 46472
rect 9379 46431 9437 46432
rect 9867 46472 9909 46481
rect 9867 46432 9868 46472
rect 9908 46432 9909 46472
rect 9867 46423 9909 46432
rect 9963 46472 10005 46481
rect 9963 46432 9964 46472
rect 10004 46432 10005 46472
rect 9963 46423 10005 46432
rect 10347 46472 10389 46481
rect 10347 46432 10348 46472
rect 10388 46432 10389 46472
rect 10347 46423 10389 46432
rect 10443 46472 10485 46481
rect 10443 46432 10444 46472
rect 10484 46432 10485 46472
rect 10443 46423 10485 46432
rect 10915 46472 10973 46473
rect 10915 46432 10924 46472
rect 10964 46432 10973 46472
rect 11451 46441 11452 46481
rect 11492 46441 11493 46481
rect 11451 46432 11493 46441
rect 12555 46472 12597 46481
rect 12555 46432 12556 46472
rect 12596 46432 12597 46472
rect 10915 46431 10973 46432
rect 12555 46423 12597 46432
rect 12651 46472 12693 46481
rect 12651 46432 12652 46472
rect 12692 46432 12693 46472
rect 12651 46423 12693 46432
rect 13035 46472 13077 46481
rect 14139 46474 14140 46514
rect 14180 46474 14181 46514
rect 18411 46516 18412 46556
rect 18452 46516 18453 46556
rect 19843 46556 19901 46557
rect 18411 46507 18453 46516
rect 19515 46514 19557 46523
rect 19843 46516 19852 46556
rect 19892 46516 19901 46556
rect 19843 46515 19901 46516
rect 13035 46432 13036 46472
rect 13076 46432 13077 46472
rect 13035 46423 13077 46432
rect 13603 46472 13661 46473
rect 13603 46432 13612 46472
rect 13652 46432 13661 46472
rect 14139 46465 14181 46474
rect 15235 46472 15293 46473
rect 13603 46431 13661 46432
rect 15235 46432 15244 46472
rect 15284 46432 15293 46472
rect 15235 46431 15293 46432
rect 16483 46472 16541 46473
rect 16483 46432 16492 46472
rect 16532 46432 16541 46472
rect 16483 46431 16541 46432
rect 17931 46472 17973 46481
rect 17931 46432 17932 46472
rect 17972 46432 17973 46472
rect 17931 46423 17973 46432
rect 18027 46472 18069 46481
rect 18027 46432 18028 46472
rect 18068 46432 18069 46472
rect 18027 46423 18069 46432
rect 18507 46472 18549 46481
rect 19515 46474 19516 46514
rect 19556 46474 19557 46514
rect 18507 46432 18508 46472
rect 18548 46432 18549 46472
rect 18507 46423 18549 46432
rect 18979 46472 19037 46473
rect 18979 46432 18988 46472
rect 19028 46432 19037 46472
rect 19515 46465 19557 46474
rect 18979 46431 19037 46432
rect 2667 46304 2709 46313
rect 2667 46264 2668 46304
rect 2708 46264 2709 46304
rect 2667 46255 2709 46264
rect 7563 46304 7605 46313
rect 7563 46264 7564 46304
rect 7604 46264 7605 46304
rect 7563 46255 7605 46264
rect 9579 46304 9621 46313
rect 9579 46264 9580 46304
rect 9620 46264 9621 46304
rect 9579 46255 9621 46264
rect 11595 46304 11637 46313
rect 11595 46264 11596 46304
rect 11636 46264 11637 46304
rect 11595 46255 11637 46264
rect 12075 46304 12117 46313
rect 12075 46264 12076 46304
rect 12116 46264 12117 46304
rect 12075 46255 12117 46264
rect 14283 46304 14325 46313
rect 14283 46264 14284 46304
rect 14324 46264 14325 46304
rect 14283 46255 14325 46264
rect 19659 46304 19701 46313
rect 19659 46264 19660 46304
rect 19700 46264 19701 46304
rect 19659 46255 19701 46264
rect 20043 46304 20085 46313
rect 20043 46264 20044 46304
rect 20084 46264 20085 46304
rect 20043 46255 20085 46264
rect 1152 46136 20452 46160
rect 1152 46096 4928 46136
rect 4968 46096 5010 46136
rect 5050 46096 5092 46136
rect 5132 46096 5174 46136
rect 5214 46096 5256 46136
rect 5296 46096 20048 46136
rect 20088 46096 20130 46136
rect 20170 46096 20212 46136
rect 20252 46096 20294 46136
rect 20334 46096 20376 46136
rect 20416 46096 20452 46136
rect 1152 46072 20452 46096
rect 1515 45968 1557 45977
rect 1515 45928 1516 45968
rect 1556 45928 1557 45968
rect 1515 45919 1557 45928
rect 1899 45968 1941 45977
rect 1899 45928 1900 45968
rect 1940 45928 1941 45968
rect 1899 45919 1941 45928
rect 11211 45968 11253 45977
rect 11211 45928 11212 45968
rect 11252 45928 11253 45968
rect 11211 45919 11253 45928
rect 12939 45968 12981 45977
rect 12939 45928 12940 45968
rect 12980 45928 12981 45968
rect 12939 45919 12981 45928
rect 19179 45968 19221 45977
rect 19179 45928 19180 45968
rect 19220 45928 19221 45968
rect 19179 45919 19221 45928
rect 14859 45884 14901 45893
rect 14859 45844 14860 45884
rect 14900 45844 14901 45884
rect 14859 45835 14901 45844
rect 16875 45884 16917 45893
rect 16875 45844 16876 45884
rect 16916 45844 16917 45884
rect 16875 45835 16917 45844
rect 2659 45800 2717 45801
rect 2659 45760 2668 45800
rect 2708 45760 2717 45800
rect 2659 45759 2717 45760
rect 3907 45800 3965 45801
rect 3907 45760 3916 45800
rect 3956 45760 3965 45800
rect 3907 45759 3965 45760
rect 4099 45800 4157 45801
rect 4099 45760 4108 45800
rect 4148 45760 4157 45800
rect 4099 45759 4157 45760
rect 5347 45800 5405 45801
rect 5347 45760 5356 45800
rect 5396 45760 5405 45800
rect 5347 45759 5405 45760
rect 6307 45800 6365 45801
rect 6307 45760 6316 45800
rect 6356 45760 6365 45800
rect 6307 45759 6365 45760
rect 7555 45800 7613 45801
rect 7555 45760 7564 45800
rect 7604 45760 7613 45800
rect 7555 45759 7613 45760
rect 9483 45800 9525 45809
rect 9483 45760 9484 45800
rect 9524 45760 9525 45800
rect 9483 45751 9525 45760
rect 9579 45800 9621 45809
rect 9579 45760 9580 45800
rect 9620 45760 9621 45800
rect 9579 45751 9621 45760
rect 10059 45800 10101 45809
rect 10059 45760 10060 45800
rect 10100 45760 10101 45800
rect 10059 45751 10101 45760
rect 10531 45800 10589 45801
rect 10531 45760 10540 45800
rect 10580 45760 10589 45800
rect 13411 45800 13469 45801
rect 10531 45759 10589 45760
rect 11019 45786 11061 45795
rect 11019 45746 11020 45786
rect 11060 45746 11061 45786
rect 13411 45760 13420 45800
rect 13460 45760 13469 45800
rect 13411 45759 13469 45760
rect 14659 45800 14717 45801
rect 14659 45760 14668 45800
rect 14708 45760 14717 45800
rect 14659 45759 14717 45760
rect 15147 45800 15189 45809
rect 15147 45760 15148 45800
rect 15188 45760 15189 45800
rect 15147 45751 15189 45760
rect 15243 45800 15285 45809
rect 15243 45760 15244 45800
rect 15284 45760 15285 45800
rect 15243 45751 15285 45760
rect 15723 45800 15765 45809
rect 15723 45760 15724 45800
rect 15764 45760 15765 45800
rect 15723 45751 15765 45760
rect 16195 45800 16253 45801
rect 16195 45760 16204 45800
rect 16244 45760 16253 45800
rect 17059 45800 17117 45801
rect 16195 45759 16253 45760
rect 16683 45786 16725 45795
rect 11019 45737 11061 45746
rect 16683 45746 16684 45786
rect 16724 45746 16725 45786
rect 17059 45760 17068 45800
rect 17108 45760 17117 45800
rect 17059 45759 17117 45760
rect 18307 45800 18365 45801
rect 18307 45760 18316 45800
rect 18356 45760 18365 45800
rect 18307 45759 18365 45760
rect 16683 45737 16725 45746
rect 1699 45716 1757 45717
rect 1699 45676 1708 45716
rect 1748 45676 1757 45716
rect 1699 45675 1757 45676
rect 2083 45716 2141 45717
rect 2083 45676 2092 45716
rect 2132 45676 2141 45716
rect 2083 45675 2141 45676
rect 9963 45716 10005 45725
rect 9963 45676 9964 45716
rect 10004 45676 10005 45716
rect 9963 45667 10005 45676
rect 11587 45716 11645 45717
rect 11587 45676 11596 45716
rect 11636 45676 11645 45716
rect 11587 45675 11645 45676
rect 13123 45716 13181 45717
rect 13123 45676 13132 45716
rect 13172 45676 13181 45716
rect 13123 45675 13181 45676
rect 15627 45716 15669 45725
rect 15627 45676 15628 45716
rect 15668 45676 15669 45716
rect 15627 45667 15669 45676
rect 18979 45716 19037 45717
rect 18979 45676 18988 45716
rect 19028 45676 19037 45716
rect 18979 45675 19037 45676
rect 19363 45716 19421 45717
rect 19363 45676 19372 45716
rect 19412 45676 19421 45716
rect 19363 45675 19421 45676
rect 19555 45716 19613 45717
rect 19555 45676 19564 45716
rect 19604 45676 19613 45716
rect 19555 45675 19613 45676
rect 2475 45548 2517 45557
rect 2475 45508 2476 45548
rect 2516 45508 2517 45548
rect 2475 45499 2517 45508
rect 5547 45548 5589 45557
rect 5547 45508 5548 45548
rect 5588 45508 5589 45548
rect 5547 45499 5589 45508
rect 7755 45548 7797 45557
rect 7755 45508 7756 45548
rect 7796 45508 7797 45548
rect 7755 45499 7797 45508
rect 11403 45548 11445 45557
rect 11403 45508 11404 45548
rect 11444 45508 11445 45548
rect 11403 45499 11445 45508
rect 18507 45548 18549 45557
rect 18507 45508 18508 45548
rect 18548 45508 18549 45548
rect 18507 45499 18549 45508
rect 18795 45548 18837 45557
rect 18795 45508 18796 45548
rect 18836 45508 18837 45548
rect 18795 45499 18837 45508
rect 19755 45548 19797 45557
rect 19755 45508 19756 45548
rect 19796 45508 19797 45548
rect 19755 45499 19797 45508
rect 1152 45380 20352 45404
rect 1152 45340 3688 45380
rect 3728 45340 3770 45380
rect 3810 45340 3852 45380
rect 3892 45340 3934 45380
rect 3974 45340 4016 45380
rect 4056 45340 18808 45380
rect 18848 45340 18890 45380
rect 18930 45340 18972 45380
rect 19012 45340 19054 45380
rect 19094 45340 19136 45380
rect 19176 45340 20352 45380
rect 1152 45316 20352 45340
rect 1515 45212 1557 45221
rect 1515 45172 1516 45212
rect 1556 45172 1557 45212
rect 1515 45163 1557 45172
rect 9387 45212 9429 45221
rect 9387 45172 9388 45212
rect 9428 45172 9429 45212
rect 9387 45163 9429 45172
rect 11019 45212 11061 45221
rect 11019 45172 11020 45212
rect 11060 45172 11061 45212
rect 11019 45163 11061 45172
rect 13707 45212 13749 45221
rect 13707 45172 13708 45212
rect 13748 45172 13749 45212
rect 13707 45163 13749 45172
rect 16683 45212 16725 45221
rect 16683 45172 16684 45212
rect 16724 45172 16725 45212
rect 16683 45163 16725 45172
rect 16875 45212 16917 45221
rect 16875 45172 16876 45212
rect 16916 45172 16917 45212
rect 16875 45163 16917 45172
rect 1699 45044 1757 45045
rect 1699 45004 1708 45044
rect 1748 45004 1757 45044
rect 1699 45003 1757 45004
rect 2083 45044 2141 45045
rect 2083 45004 2092 45044
rect 2132 45004 2141 45044
rect 6123 45044 6165 45053
rect 2083 45003 2141 45004
rect 2523 45002 2565 45011
rect 2523 44962 2524 45002
rect 2564 44962 2565 45002
rect 6123 45004 6124 45044
rect 6164 45004 6165 45044
rect 6123 44995 6165 45004
rect 13891 45044 13949 45045
rect 13891 45004 13900 45044
rect 13940 45004 13949 45044
rect 13891 45003 13949 45004
rect 17059 45044 17117 45045
rect 17059 45004 17068 45044
rect 17108 45004 17117 45044
rect 17059 45003 17117 45004
rect 18411 45044 18453 45053
rect 18411 45004 18412 45044
rect 18452 45004 18453 45044
rect 18411 44995 18453 45004
rect 18507 45044 18549 45053
rect 18507 45004 18508 45044
rect 18548 45004 18549 45044
rect 18507 44995 18549 45004
rect 19843 45044 19901 45045
rect 19843 45004 19852 45044
rect 19892 45004 19901 45044
rect 19843 45003 19901 45004
rect 7179 44974 7221 44983
rect 2523 44953 2565 44962
rect 3043 44960 3101 44961
rect 3043 44920 3052 44960
rect 3092 44920 3101 44960
rect 3043 44919 3101 44920
rect 3531 44960 3573 44969
rect 3531 44920 3532 44960
rect 3572 44920 3573 44960
rect 3531 44911 3573 44920
rect 3627 44960 3669 44969
rect 3627 44920 3628 44960
rect 3668 44920 3669 44960
rect 3627 44911 3669 44920
rect 4011 44960 4053 44969
rect 4011 44920 4012 44960
rect 4052 44920 4053 44960
rect 4011 44911 4053 44920
rect 4107 44960 4149 44969
rect 4107 44920 4108 44960
rect 4148 44920 4149 44960
rect 4107 44911 4149 44920
rect 5643 44960 5685 44969
rect 5643 44920 5644 44960
rect 5684 44920 5685 44960
rect 5643 44911 5685 44920
rect 5739 44960 5781 44969
rect 5739 44920 5740 44960
rect 5780 44920 5781 44960
rect 5739 44911 5781 44920
rect 6219 44960 6261 44969
rect 6219 44920 6220 44960
rect 6260 44920 6261 44960
rect 6219 44911 6261 44920
rect 6691 44960 6749 44961
rect 6691 44920 6700 44960
rect 6740 44920 6749 44960
rect 7179 44934 7180 44974
rect 7220 44934 7221 44974
rect 19515 44969 19557 44978
rect 7179 44925 7221 44934
rect 7939 44960 7997 44961
rect 6691 44919 6749 44920
rect 7939 44920 7948 44960
rect 7988 44920 7997 44960
rect 7939 44919 7997 44920
rect 9187 44960 9245 44961
rect 9187 44920 9196 44960
rect 9236 44920 9245 44960
rect 9187 44919 9245 44920
rect 9571 44960 9629 44961
rect 9571 44920 9580 44960
rect 9620 44920 9629 44960
rect 9571 44919 9629 44920
rect 10819 44960 10877 44961
rect 10819 44920 10828 44960
rect 10868 44920 10877 44960
rect 10819 44919 10877 44920
rect 12067 44960 12125 44961
rect 12067 44920 12076 44960
rect 12116 44920 12125 44960
rect 12067 44919 12125 44920
rect 13315 44960 13373 44961
rect 13315 44920 13324 44960
rect 13364 44920 13373 44960
rect 13315 44919 13373 44920
rect 15235 44960 15293 44961
rect 15235 44920 15244 44960
rect 15284 44920 15293 44960
rect 15235 44919 15293 44920
rect 16483 44960 16541 44961
rect 16483 44920 16492 44960
rect 16532 44920 16541 44960
rect 16483 44919 16541 44920
rect 17931 44960 17973 44969
rect 17931 44920 17932 44960
rect 17972 44920 17973 44960
rect 17931 44911 17973 44920
rect 18027 44960 18069 44969
rect 18027 44920 18028 44960
rect 18068 44920 18069 44960
rect 18027 44911 18069 44920
rect 18979 44960 19037 44961
rect 18979 44920 18988 44960
rect 19028 44920 19037 44960
rect 19515 44929 19516 44969
rect 19556 44929 19557 44969
rect 19515 44920 19557 44929
rect 18979 44919 19037 44920
rect 2379 44876 2421 44885
rect 2379 44836 2380 44876
rect 2420 44836 2421 44876
rect 2379 44827 2421 44836
rect 7371 44876 7413 44885
rect 7371 44836 7372 44876
rect 7412 44836 7413 44876
rect 7371 44827 7413 44836
rect 19659 44876 19701 44885
rect 19659 44836 19660 44876
rect 19700 44836 19701 44876
rect 19659 44827 19701 44836
rect 1899 44792 1941 44801
rect 1899 44752 1900 44792
rect 1940 44752 1941 44792
rect 1899 44743 1941 44752
rect 13515 44792 13557 44801
rect 13515 44752 13516 44792
rect 13556 44752 13557 44792
rect 13515 44743 13557 44752
rect 20043 44792 20085 44801
rect 20043 44752 20044 44792
rect 20084 44752 20085 44792
rect 20043 44743 20085 44752
rect 1152 44624 20452 44648
rect 1152 44584 4928 44624
rect 4968 44584 5010 44624
rect 5050 44584 5092 44624
rect 5132 44584 5174 44624
rect 5214 44584 5256 44624
rect 5296 44584 20048 44624
rect 20088 44584 20130 44624
rect 20170 44584 20212 44624
rect 20252 44584 20294 44624
rect 20334 44584 20376 44624
rect 20416 44584 20452 44624
rect 1152 44560 20452 44584
rect 1803 44456 1845 44465
rect 1803 44416 1804 44456
rect 1844 44416 1845 44456
rect 1803 44407 1845 44416
rect 7275 44456 7317 44465
rect 7275 44416 7276 44456
rect 7316 44416 7317 44456
rect 7275 44407 7317 44416
rect 9675 44456 9717 44465
rect 9675 44416 9676 44456
rect 9716 44416 9717 44456
rect 9675 44407 9717 44416
rect 13515 44456 13557 44465
rect 13515 44416 13516 44456
rect 13556 44416 13557 44456
rect 13515 44407 13557 44416
rect 15435 44456 15477 44465
rect 15435 44416 15436 44456
rect 15476 44416 15477 44456
rect 15435 44407 15477 44416
rect 19563 44456 19605 44465
rect 19563 44416 19564 44456
rect 19604 44416 19605 44456
rect 19563 44407 19605 44416
rect 17451 44372 17493 44381
rect 17451 44332 17452 44372
rect 17492 44332 17493 44372
rect 13987 44330 14045 44331
rect 2371 44288 2429 44289
rect 2371 44248 2380 44288
rect 2420 44248 2429 44288
rect 2371 44247 2429 44248
rect 3619 44288 3677 44289
rect 3619 44248 3628 44288
rect 3668 44248 3677 44288
rect 3619 44247 3677 44248
rect 3811 44288 3869 44289
rect 3811 44248 3820 44288
rect 3860 44248 3869 44288
rect 3811 44247 3869 44248
rect 5059 44288 5117 44289
rect 5059 44248 5068 44288
rect 5108 44248 5117 44288
rect 5059 44247 5117 44248
rect 5547 44288 5589 44297
rect 5547 44248 5548 44288
rect 5588 44248 5589 44288
rect 5547 44239 5589 44248
rect 5643 44288 5685 44297
rect 5643 44248 5644 44288
rect 5684 44248 5685 44288
rect 5643 44239 5685 44248
rect 6027 44288 6069 44297
rect 6027 44248 6028 44288
rect 6068 44248 6069 44288
rect 6027 44239 6069 44248
rect 6123 44288 6165 44297
rect 6123 44248 6124 44288
rect 6164 44248 6165 44288
rect 6123 44239 6165 44248
rect 6595 44288 6653 44289
rect 6595 44248 6604 44288
rect 6644 44248 6653 44288
rect 6595 44247 6653 44248
rect 7083 44283 7125 44292
rect 7083 44243 7084 44283
rect 7124 44243 7125 44283
rect 10051 44288 10109 44289
rect 10051 44248 10060 44288
rect 10100 44248 10109 44288
rect 10051 44247 10109 44248
rect 11299 44288 11357 44289
rect 11299 44248 11308 44288
rect 11348 44248 11357 44288
rect 11299 44247 11357 44248
rect 11787 44288 11829 44297
rect 11787 44248 11788 44288
rect 11828 44248 11829 44288
rect 7083 44234 7125 44243
rect 11787 44239 11829 44248
rect 11883 44288 11925 44297
rect 11883 44248 11884 44288
rect 11924 44248 11925 44288
rect 11883 44239 11925 44248
rect 12363 44288 12405 44297
rect 13987 44290 13996 44330
rect 14036 44290 14045 44330
rect 17451 44323 17493 44332
rect 13987 44289 14045 44290
rect 12363 44248 12364 44288
rect 12404 44248 12405 44288
rect 12363 44239 12405 44248
rect 12835 44288 12893 44289
rect 12835 44248 12844 44288
rect 12884 44248 12893 44288
rect 15235 44288 15293 44289
rect 12835 44247 12893 44248
rect 13323 44274 13365 44283
rect 13323 44234 13324 44274
rect 13364 44234 13365 44274
rect 15235 44248 15244 44288
rect 15284 44248 15293 44288
rect 15235 44247 15293 44248
rect 15723 44288 15765 44297
rect 15723 44248 15724 44288
rect 15764 44248 15765 44288
rect 15723 44239 15765 44248
rect 15819 44288 15861 44297
rect 15819 44248 15820 44288
rect 15860 44248 15861 44288
rect 15819 44239 15861 44248
rect 16203 44288 16245 44297
rect 16203 44248 16204 44288
rect 16244 44248 16245 44288
rect 16203 44239 16245 44248
rect 16299 44288 16341 44297
rect 16299 44248 16300 44288
rect 16340 44248 16341 44288
rect 16299 44239 16341 44248
rect 16771 44288 16829 44289
rect 16771 44248 16780 44288
rect 16820 44248 16829 44288
rect 18115 44288 18173 44289
rect 16771 44247 16829 44248
rect 17259 44274 17301 44283
rect 13323 44225 13365 44234
rect 17259 44234 17260 44274
rect 17300 44234 17301 44274
rect 18115 44248 18124 44288
rect 18164 44248 18173 44288
rect 18115 44247 18173 44248
rect 19363 44288 19421 44289
rect 19363 44248 19372 44288
rect 19412 44248 19421 44288
rect 19363 44247 19421 44248
rect 17259 44225 17301 44234
rect 1987 44204 2045 44205
rect 1987 44164 1996 44204
rect 2036 44164 2045 44204
rect 1987 44163 2045 44164
rect 9187 44204 9245 44205
rect 9187 44164 9196 44204
rect 9236 44164 9245 44204
rect 9187 44163 9245 44164
rect 9859 44204 9917 44205
rect 9859 44164 9868 44204
rect 9908 44164 9917 44204
rect 9859 44163 9917 44164
rect 12267 44204 12309 44213
rect 12267 44164 12268 44204
rect 12308 44164 12309 44204
rect 12267 44155 12309 44164
rect 19747 44204 19805 44205
rect 19747 44164 19756 44204
rect 19796 44164 19805 44204
rect 19747 44163 19805 44164
rect 5259 44120 5301 44129
rect 5259 44080 5260 44120
rect 5300 44080 5301 44120
rect 5259 44071 5301 44080
rect 2187 44036 2229 44045
rect 2187 43996 2188 44036
rect 2228 43996 2229 44036
rect 2187 43987 2229 43996
rect 9003 44036 9045 44045
rect 9003 43996 9004 44036
rect 9044 43996 9045 44036
rect 9003 43987 9045 43996
rect 11499 44036 11541 44045
rect 11499 43996 11500 44036
rect 11540 43996 11541 44036
rect 11499 43987 11541 43996
rect 19947 44036 19989 44045
rect 19947 43996 19948 44036
rect 19988 43996 19989 44036
rect 19947 43987 19989 43996
rect 1152 43868 20352 43892
rect 1152 43828 3688 43868
rect 3728 43828 3770 43868
rect 3810 43828 3852 43868
rect 3892 43828 3934 43868
rect 3974 43828 4016 43868
rect 4056 43828 18808 43868
rect 18848 43828 18890 43868
rect 18930 43828 18972 43868
rect 19012 43828 19054 43868
rect 19094 43828 19136 43868
rect 19176 43828 20352 43868
rect 1152 43804 20352 43828
rect 11403 43700 11445 43709
rect 11403 43660 11404 43700
rect 11444 43660 11445 43700
rect 11403 43651 11445 43660
rect 15051 43700 15093 43709
rect 15051 43660 15052 43700
rect 15092 43660 15093 43700
rect 15051 43651 15093 43660
rect 17259 43700 17301 43709
rect 17259 43660 17260 43700
rect 17300 43660 17301 43700
rect 17259 43651 17301 43660
rect 17451 43700 17493 43709
rect 17451 43660 17452 43700
rect 17492 43660 17493 43700
rect 17451 43651 17493 43660
rect 19179 43700 19221 43709
rect 19179 43660 19180 43700
rect 19220 43660 19221 43700
rect 19179 43651 19221 43660
rect 3627 43532 3669 43541
rect 3627 43492 3628 43532
rect 3668 43492 3669 43532
rect 3627 43483 3669 43492
rect 8523 43532 8565 43541
rect 8523 43492 8524 43532
rect 8564 43492 8565 43532
rect 8523 43483 8565 43492
rect 12267 43532 12309 43541
rect 12267 43492 12268 43532
rect 12308 43492 12309 43532
rect 12267 43483 12309 43492
rect 14083 43532 14141 43533
rect 14083 43492 14092 43532
rect 14132 43492 14141 43532
rect 14083 43491 14141 43492
rect 14851 43532 14909 43533
rect 14851 43492 14860 43532
rect 14900 43492 14909 43532
rect 14851 43491 14909 43492
rect 17635 43532 17693 43533
rect 17635 43492 17644 43532
rect 17684 43492 17693 43532
rect 17635 43491 17693 43492
rect 17827 43532 17885 43533
rect 17827 43492 17836 43532
rect 17876 43492 17885 43532
rect 17827 43491 17885 43492
rect 18979 43532 19037 43533
rect 18979 43492 18988 43532
rect 19028 43492 19037 43532
rect 18979 43491 19037 43492
rect 19363 43532 19421 43533
rect 19363 43492 19372 43532
rect 19412 43492 19421 43532
rect 19363 43491 19421 43492
rect 2667 43462 2709 43471
rect 2667 43422 2668 43462
rect 2708 43422 2709 43462
rect 9531 43457 9573 43466
rect 13275 43457 13317 43466
rect 2667 43413 2709 43422
rect 3139 43448 3197 43449
rect 3139 43408 3148 43448
rect 3188 43408 3197 43448
rect 3139 43407 3197 43408
rect 3723 43448 3765 43457
rect 3723 43408 3724 43448
rect 3764 43408 3765 43448
rect 3723 43399 3765 43408
rect 4107 43448 4149 43457
rect 4107 43408 4108 43448
rect 4148 43408 4149 43448
rect 4107 43399 4149 43408
rect 4203 43448 4245 43457
rect 4203 43408 4204 43448
rect 4244 43408 4245 43448
rect 4203 43399 4245 43408
rect 6211 43448 6269 43449
rect 6211 43408 6220 43448
rect 6260 43408 6269 43448
rect 6211 43407 6269 43408
rect 7459 43448 7517 43449
rect 7459 43408 7468 43448
rect 7508 43408 7517 43448
rect 7459 43407 7517 43408
rect 7947 43448 7989 43457
rect 7947 43408 7948 43448
rect 7988 43408 7989 43448
rect 7947 43399 7989 43408
rect 8043 43448 8085 43457
rect 8043 43408 8044 43448
rect 8084 43408 8085 43448
rect 8043 43399 8085 43408
rect 8427 43448 8469 43457
rect 8427 43408 8428 43448
rect 8468 43408 8469 43448
rect 8427 43399 8469 43408
rect 8995 43448 9053 43449
rect 8995 43408 9004 43448
rect 9044 43408 9053 43448
rect 9531 43417 9532 43457
rect 9572 43417 9573 43457
rect 9531 43408 9573 43417
rect 9955 43448 10013 43449
rect 9955 43408 9964 43448
rect 10004 43408 10013 43448
rect 8995 43407 9053 43408
rect 9955 43407 10013 43408
rect 11203 43448 11261 43449
rect 11203 43408 11212 43448
rect 11252 43408 11261 43448
rect 11203 43407 11261 43408
rect 11691 43448 11733 43457
rect 11691 43408 11692 43448
rect 11732 43408 11733 43448
rect 11691 43399 11733 43408
rect 11787 43448 11829 43457
rect 11787 43408 11788 43448
rect 11828 43408 11829 43448
rect 11787 43399 11829 43408
rect 12171 43448 12213 43457
rect 12171 43408 12172 43448
rect 12212 43408 12213 43448
rect 12171 43399 12213 43408
rect 12739 43448 12797 43449
rect 12739 43408 12748 43448
rect 12788 43408 12797 43448
rect 13275 43417 13276 43457
rect 13316 43417 13317 43457
rect 13275 43408 13317 43417
rect 15811 43448 15869 43449
rect 15811 43408 15820 43448
rect 15860 43408 15869 43448
rect 12739 43407 12797 43408
rect 15811 43407 15869 43408
rect 17059 43448 17117 43449
rect 17059 43408 17068 43448
rect 17108 43408 17117 43448
rect 17059 43407 17117 43408
rect 2475 43364 2517 43373
rect 2475 43324 2476 43364
rect 2516 43324 2517 43364
rect 2475 43315 2517 43324
rect 7659 43364 7701 43373
rect 7659 43324 7660 43364
rect 7700 43324 7701 43364
rect 7659 43315 7701 43324
rect 9675 43364 9717 43373
rect 9675 43324 9676 43364
rect 9716 43324 9717 43364
rect 9675 43315 9717 43324
rect 13419 43280 13461 43289
rect 13419 43240 13420 43280
rect 13460 43240 13461 43280
rect 13419 43231 13461 43240
rect 13899 43280 13941 43289
rect 13899 43240 13900 43280
rect 13940 43240 13941 43280
rect 13899 43231 13941 43240
rect 18027 43280 18069 43289
rect 18027 43240 18028 43280
rect 18068 43240 18069 43280
rect 18027 43231 18069 43240
rect 19563 43280 19605 43289
rect 19563 43240 19564 43280
rect 19604 43240 19605 43280
rect 19563 43231 19605 43240
rect 1152 43112 20452 43136
rect 1152 43072 4928 43112
rect 4968 43072 5010 43112
rect 5050 43072 5092 43112
rect 5132 43072 5174 43112
rect 5214 43072 5256 43112
rect 5296 43072 20048 43112
rect 20088 43072 20130 43112
rect 20170 43072 20212 43112
rect 20252 43072 20294 43112
rect 20334 43072 20376 43112
rect 20416 43072 20452 43112
rect 1152 43048 20452 43072
rect 9579 42944 9621 42953
rect 9579 42904 9580 42944
rect 9620 42904 9621 42944
rect 9579 42895 9621 42904
rect 2667 42860 2709 42869
rect 2667 42820 2668 42860
rect 2708 42820 2709 42860
rect 2667 42811 2709 42820
rect 4683 42860 4725 42869
rect 4683 42820 4684 42860
rect 4724 42820 4725 42860
rect 4683 42811 4725 42820
rect 6699 42860 6741 42869
rect 6699 42820 6700 42860
rect 6740 42820 6741 42860
rect 6699 42811 6741 42820
rect 13803 42860 13845 42869
rect 13803 42820 13804 42860
rect 13844 42820 13845 42860
rect 13803 42811 13845 42820
rect 1219 42776 1277 42777
rect 1219 42736 1228 42776
rect 1268 42736 1277 42776
rect 1219 42735 1277 42736
rect 2467 42776 2525 42777
rect 2467 42736 2476 42776
rect 2516 42736 2525 42776
rect 2467 42735 2525 42736
rect 3235 42776 3293 42777
rect 3235 42736 3244 42776
rect 3284 42736 3293 42776
rect 3235 42735 3293 42736
rect 4483 42776 4541 42777
rect 4483 42736 4492 42776
rect 4532 42736 4541 42776
rect 4483 42735 4541 42736
rect 4971 42776 5013 42785
rect 4971 42736 4972 42776
rect 5012 42736 5013 42776
rect 4971 42727 5013 42736
rect 5067 42776 5109 42785
rect 5067 42736 5068 42776
rect 5108 42736 5109 42776
rect 5067 42727 5109 42736
rect 6019 42776 6077 42777
rect 6019 42736 6028 42776
rect 6068 42736 6077 42776
rect 8131 42776 8189 42777
rect 6019 42735 6077 42736
rect 6555 42734 6597 42743
rect 8131 42736 8140 42776
rect 8180 42736 8189 42776
rect 8131 42735 8189 42736
rect 9379 42776 9437 42777
rect 9379 42736 9388 42776
rect 9428 42736 9437 42776
rect 9379 42735 9437 42736
rect 12355 42776 12413 42777
rect 12355 42736 12364 42776
rect 12404 42736 12413 42776
rect 12355 42735 12413 42736
rect 13603 42776 13661 42777
rect 13603 42736 13612 42776
rect 13652 42736 13661 42776
rect 13603 42735 13661 42736
rect 5451 42692 5493 42701
rect 5451 42652 5452 42692
rect 5492 42652 5493 42692
rect 5451 42643 5493 42652
rect 5547 42692 5589 42701
rect 5547 42652 5548 42692
rect 5588 42652 5589 42692
rect 6555 42694 6556 42734
rect 6596 42694 6597 42734
rect 6555 42685 6597 42694
rect 18595 42692 18653 42693
rect 5547 42643 5589 42652
rect 18595 42652 18604 42692
rect 18644 42652 18653 42692
rect 18595 42651 18653 42652
rect 18979 42692 19037 42693
rect 18979 42652 18988 42692
rect 19028 42652 19037 42692
rect 18979 42651 19037 42652
rect 19363 42692 19421 42693
rect 19363 42652 19372 42692
rect 19412 42652 19421 42692
rect 19363 42651 19421 42652
rect 19747 42692 19805 42693
rect 19747 42652 19756 42692
rect 19796 42652 19805 42692
rect 19747 42651 19805 42652
rect 19179 42608 19221 42617
rect 19179 42568 19180 42608
rect 19220 42568 19221 42608
rect 19179 42559 19221 42568
rect 19563 42608 19605 42617
rect 19563 42568 19564 42608
rect 19604 42568 19605 42608
rect 19563 42559 19605 42568
rect 18795 42524 18837 42533
rect 18795 42484 18796 42524
rect 18836 42484 18837 42524
rect 18795 42475 18837 42484
rect 19947 42524 19989 42533
rect 19947 42484 19948 42524
rect 19988 42484 19989 42524
rect 19947 42475 19989 42484
rect 1152 42356 20352 42380
rect 1152 42316 3688 42356
rect 3728 42316 3770 42356
rect 3810 42316 3852 42356
rect 3892 42316 3934 42356
rect 3974 42316 4016 42356
rect 4056 42316 18808 42356
rect 18848 42316 18890 42356
rect 18930 42316 18972 42356
rect 19012 42316 19054 42356
rect 19094 42316 19136 42356
rect 19176 42316 20352 42356
rect 1152 42292 20352 42316
rect 1899 42188 1941 42197
rect 1899 42148 1900 42188
rect 1940 42148 1941 42188
rect 1899 42139 1941 42148
rect 6699 42188 6741 42197
rect 6699 42148 6700 42188
rect 6740 42148 6741 42188
rect 6699 42139 6741 42148
rect 17163 42188 17205 42197
rect 17163 42148 17164 42188
rect 17204 42148 17205 42188
rect 17163 42139 17205 42148
rect 19275 42188 19317 42197
rect 19275 42148 19276 42188
rect 19316 42148 19317 42188
rect 19275 42139 19317 42148
rect 20043 42188 20085 42197
rect 20043 42148 20044 42188
rect 20084 42148 20085 42188
rect 20043 42139 20085 42148
rect 4875 42104 4917 42113
rect 4875 42064 4876 42104
rect 4916 42064 4917 42104
rect 4875 42055 4917 42064
rect 18891 42104 18933 42113
rect 18891 42064 18892 42104
rect 18932 42064 18933 42104
rect 18891 42055 18933 42064
rect 2083 42020 2141 42021
rect 2083 41980 2092 42020
rect 2132 41980 2141 42020
rect 2083 41979 2141 41980
rect 3435 42020 3477 42029
rect 3435 41980 3436 42020
rect 3476 41980 3477 42020
rect 3435 41971 3477 41980
rect 16963 42020 17021 42021
rect 16963 41980 16972 42020
rect 17012 41980 17021 42020
rect 16963 41979 17021 41980
rect 18307 42020 18365 42021
rect 18307 41980 18316 42020
rect 18356 41980 18365 42020
rect 18307 41979 18365 41980
rect 18691 42020 18749 42021
rect 18691 41980 18700 42020
rect 18740 41980 18749 42020
rect 18691 41979 18749 41980
rect 19075 42020 19133 42021
rect 19075 41980 19084 42020
rect 19124 41980 19133 42020
rect 19075 41979 19133 41980
rect 19459 42020 19517 42021
rect 19459 41980 19468 42020
rect 19508 41980 19517 42020
rect 19459 41979 19517 41980
rect 19843 42020 19901 42021
rect 19843 41980 19852 42020
rect 19892 41980 19901 42020
rect 19843 41979 19901 41980
rect 2475 41941 2517 41950
rect 2475 41901 2476 41941
rect 2516 41901 2517 41941
rect 2475 41892 2517 41901
rect 2947 41936 3005 41937
rect 2947 41896 2956 41936
rect 2996 41896 3005 41936
rect 2947 41895 3005 41896
rect 3531 41936 3573 41945
rect 3531 41896 3532 41936
rect 3572 41896 3573 41936
rect 3531 41887 3573 41896
rect 3915 41936 3957 41945
rect 3915 41896 3916 41936
rect 3956 41896 3957 41936
rect 3915 41887 3957 41896
rect 4011 41936 4053 41945
rect 4011 41896 4012 41936
rect 4052 41896 4053 41936
rect 4011 41887 4053 41896
rect 5251 41936 5309 41937
rect 5251 41896 5260 41936
rect 5300 41896 5309 41936
rect 5251 41895 5309 41896
rect 6499 41936 6557 41937
rect 6499 41896 6508 41936
rect 6548 41896 6557 41936
rect 6499 41895 6557 41896
rect 7555 41936 7613 41937
rect 7555 41896 7564 41936
rect 7604 41896 7613 41936
rect 7555 41895 7613 41896
rect 8803 41936 8861 41937
rect 8803 41896 8812 41936
rect 8852 41896 8861 41936
rect 8803 41895 8861 41896
rect 9187 41936 9245 41937
rect 9187 41896 9196 41936
rect 9236 41896 9245 41936
rect 9187 41895 9245 41896
rect 10435 41936 10493 41937
rect 10435 41896 10444 41936
rect 10484 41896 10493 41936
rect 10435 41895 10493 41896
rect 10819 41936 10877 41937
rect 10819 41896 10828 41936
rect 10868 41896 10877 41936
rect 10819 41895 10877 41896
rect 12067 41936 12125 41937
rect 12067 41896 12076 41936
rect 12116 41896 12125 41936
rect 12067 41895 12125 41896
rect 2283 41852 2325 41861
rect 2283 41812 2284 41852
rect 2324 41812 2325 41852
rect 2283 41803 2325 41812
rect 9003 41768 9045 41777
rect 9003 41728 9004 41768
rect 9044 41728 9045 41768
rect 9003 41719 9045 41728
rect 10635 41768 10677 41777
rect 10635 41728 10636 41768
rect 10676 41728 10677 41768
rect 10635 41719 10677 41728
rect 12267 41768 12309 41777
rect 12267 41728 12268 41768
rect 12308 41728 12309 41768
rect 12267 41719 12309 41728
rect 18507 41768 18549 41777
rect 18507 41728 18508 41768
rect 18548 41728 18549 41768
rect 18507 41719 18549 41728
rect 19659 41768 19701 41777
rect 19659 41728 19660 41768
rect 19700 41728 19701 41768
rect 19659 41719 19701 41728
rect 1152 41600 20452 41624
rect 1152 41560 4928 41600
rect 4968 41560 5010 41600
rect 5050 41560 5092 41600
rect 5132 41560 5174 41600
rect 5214 41560 5256 41600
rect 5296 41560 20048 41600
rect 20088 41560 20130 41600
rect 20170 41560 20212 41600
rect 20252 41560 20294 41600
rect 20334 41560 20376 41600
rect 20416 41560 20452 41600
rect 1152 41536 20452 41560
rect 3339 41432 3381 41441
rect 3339 41392 3340 41432
rect 3380 41392 3381 41432
rect 3339 41383 3381 41392
rect 9283 41432 9341 41433
rect 9283 41392 9292 41432
rect 9332 41392 9341 41432
rect 9283 41391 9341 41392
rect 12939 41432 12981 41441
rect 12939 41392 12940 41432
rect 12980 41392 12981 41432
rect 12939 41383 12981 41392
rect 19083 41432 19125 41441
rect 19083 41392 19084 41432
rect 19124 41392 19125 41432
rect 19083 41383 19125 41392
rect 5067 41348 5109 41357
rect 5067 41308 5068 41348
rect 5108 41308 5109 41348
rect 5067 41299 5109 41308
rect 7083 41348 7125 41357
rect 7083 41308 7084 41348
rect 7124 41308 7125 41348
rect 7083 41299 7125 41308
rect 9099 41348 9141 41357
rect 9099 41308 9100 41348
rect 9140 41308 9141 41348
rect 9099 41299 9141 41308
rect 12171 41348 12213 41357
rect 12171 41308 12172 41348
rect 12212 41308 12213 41348
rect 12171 41299 12213 41308
rect 1891 41264 1949 41265
rect 1891 41224 1900 41264
rect 1940 41224 1949 41264
rect 1891 41223 1949 41224
rect 3139 41264 3197 41265
rect 3139 41224 3148 41264
rect 3188 41224 3197 41264
rect 3139 41223 3197 41224
rect 3619 41264 3677 41265
rect 3619 41224 3628 41264
rect 3668 41224 3677 41264
rect 3619 41223 3677 41224
rect 4867 41264 4925 41265
rect 4867 41224 4876 41264
rect 4916 41224 4925 41264
rect 4867 41223 4925 41224
rect 5355 41264 5397 41273
rect 5355 41224 5356 41264
rect 5396 41224 5397 41264
rect 5355 41215 5397 41224
rect 5451 41264 5493 41273
rect 5451 41224 5452 41264
rect 5492 41224 5493 41264
rect 5451 41215 5493 41224
rect 6403 41264 6461 41265
rect 6403 41224 6412 41264
rect 6452 41224 6461 41264
rect 7651 41264 7709 41265
rect 6403 41223 6461 41224
rect 6939 41254 6981 41263
rect 6939 41214 6940 41254
rect 6980 41214 6981 41254
rect 7651 41224 7660 41264
rect 7700 41224 7709 41264
rect 7651 41223 7709 41224
rect 8899 41264 8957 41265
rect 8899 41224 8908 41264
rect 8948 41224 8957 41264
rect 8899 41223 8957 41224
rect 10443 41264 10485 41273
rect 10443 41224 10444 41264
rect 10484 41224 10485 41264
rect 10443 41215 10485 41224
rect 10539 41264 10581 41273
rect 10539 41224 10540 41264
rect 10580 41224 10581 41264
rect 10539 41215 10581 41224
rect 11019 41264 11061 41273
rect 11019 41224 11020 41264
rect 11060 41224 11061 41264
rect 11019 41215 11061 41224
rect 11491 41264 11549 41265
rect 11491 41224 11500 41264
rect 11540 41224 11549 41264
rect 11491 41223 11549 41224
rect 12027 41254 12069 41263
rect 6939 41205 6981 41214
rect 12027 41214 12028 41254
rect 12068 41214 12069 41254
rect 12027 41205 12069 41214
rect 5835 41180 5877 41189
rect 5835 41140 5836 41180
rect 5876 41140 5877 41180
rect 5835 41131 5877 41140
rect 5931 41180 5973 41189
rect 5931 41140 5932 41180
rect 5972 41140 5973 41180
rect 5931 41131 5973 41140
rect 10923 41180 10965 41189
rect 10923 41140 10924 41180
rect 10964 41140 10965 41180
rect 10923 41131 10965 41140
rect 12739 41180 12797 41181
rect 12739 41140 12748 41180
rect 12788 41140 12797 41180
rect 12739 41139 12797 41140
rect 18883 41180 18941 41181
rect 18883 41140 18892 41180
rect 18932 41140 18941 41180
rect 18883 41139 18941 41140
rect 19267 41180 19325 41181
rect 19267 41140 19276 41180
rect 19316 41140 19325 41180
rect 19267 41139 19325 41140
rect 19651 41180 19709 41181
rect 19651 41140 19660 41180
rect 19700 41140 19709 41180
rect 19651 41139 19709 41140
rect 19467 41012 19509 41021
rect 19467 40972 19468 41012
rect 19508 40972 19509 41012
rect 19467 40963 19509 40972
rect 19851 41012 19893 41021
rect 19851 40972 19852 41012
rect 19892 40972 19893 41012
rect 19851 40963 19893 40972
rect 1152 40844 20352 40868
rect 1152 40804 3688 40844
rect 3728 40804 3770 40844
rect 3810 40804 3852 40844
rect 3892 40804 3934 40844
rect 3974 40804 4016 40844
rect 4056 40804 18808 40844
rect 18848 40804 18890 40844
rect 18930 40804 18972 40844
rect 19012 40804 19054 40844
rect 19094 40804 19136 40844
rect 19176 40804 20352 40844
rect 1152 40780 20352 40804
rect 2667 40676 2709 40685
rect 2667 40636 2668 40676
rect 2708 40636 2709 40676
rect 2667 40627 2709 40636
rect 7371 40676 7413 40685
rect 7371 40636 7372 40676
rect 7412 40636 7413 40676
rect 7371 40627 7413 40636
rect 13227 40676 13269 40685
rect 13227 40636 13228 40676
rect 13268 40636 13269 40676
rect 13227 40627 13269 40636
rect 19083 40676 19125 40685
rect 19083 40636 19084 40676
rect 19124 40636 19125 40676
rect 19083 40627 19125 40636
rect 19467 40676 19509 40685
rect 19467 40636 19468 40676
rect 19508 40636 19509 40676
rect 19467 40627 19509 40636
rect 9963 40508 10005 40517
rect 9963 40468 9964 40508
rect 10004 40468 10005 40508
rect 2467 40466 2525 40467
rect 2467 40426 2476 40466
rect 2516 40426 2525 40466
rect 9963 40459 10005 40468
rect 13027 40508 13085 40509
rect 13027 40468 13036 40508
rect 13076 40468 13085 40508
rect 13027 40467 13085 40468
rect 18883 40508 18941 40509
rect 18883 40468 18892 40508
rect 18932 40468 18941 40508
rect 18883 40467 18941 40468
rect 19267 40508 19325 40509
rect 19267 40468 19276 40508
rect 19316 40468 19325 40508
rect 19267 40467 19325 40468
rect 19651 40508 19709 40509
rect 19651 40468 19660 40508
rect 19700 40468 19709 40508
rect 19651 40467 19709 40468
rect 20035 40508 20093 40509
rect 20035 40468 20044 40508
rect 20084 40468 20093 40508
rect 20035 40467 20093 40468
rect 10923 40438 10965 40447
rect 2467 40425 2525 40426
rect 1219 40424 1277 40425
rect 1219 40384 1228 40424
rect 1268 40384 1277 40424
rect 1219 40383 1277 40384
rect 3907 40424 3965 40425
rect 3907 40384 3916 40424
rect 3956 40384 3965 40424
rect 3907 40383 3965 40384
rect 5155 40424 5213 40425
rect 5155 40384 5164 40424
rect 5204 40384 5213 40424
rect 5155 40383 5213 40384
rect 5923 40424 5981 40425
rect 5923 40384 5932 40424
rect 5972 40384 5981 40424
rect 5923 40383 5981 40384
rect 7171 40424 7229 40425
rect 7171 40384 7180 40424
rect 7220 40384 7229 40424
rect 7171 40383 7229 40384
rect 7747 40424 7805 40425
rect 7747 40384 7756 40424
rect 7796 40384 7805 40424
rect 7747 40383 7805 40384
rect 8995 40424 9053 40425
rect 8995 40384 9004 40424
rect 9044 40384 9053 40424
rect 8995 40383 9053 40384
rect 9387 40424 9429 40433
rect 9387 40384 9388 40424
rect 9428 40384 9429 40424
rect 9387 40375 9429 40384
rect 9483 40424 9525 40433
rect 9483 40384 9484 40424
rect 9524 40384 9525 40424
rect 9483 40375 9525 40384
rect 9867 40424 9909 40433
rect 9867 40384 9868 40424
rect 9908 40384 9909 40424
rect 9867 40375 9909 40384
rect 10435 40424 10493 40425
rect 10435 40384 10444 40424
rect 10484 40384 10493 40424
rect 10923 40398 10924 40438
rect 10964 40398 10965 40438
rect 10923 40389 10965 40398
rect 10435 40383 10493 40384
rect 7563 40340 7605 40349
rect 7563 40300 7564 40340
rect 7604 40300 7605 40340
rect 7563 40291 7605 40300
rect 5355 40256 5397 40265
rect 5355 40216 5356 40256
rect 5396 40216 5397 40256
rect 5355 40207 5397 40216
rect 11115 40256 11157 40265
rect 11115 40216 11116 40256
rect 11156 40216 11157 40256
rect 11115 40207 11157 40216
rect 19851 40256 19893 40265
rect 19851 40216 19852 40256
rect 19892 40216 19893 40256
rect 19851 40207 19893 40216
rect 20235 40256 20277 40265
rect 20235 40216 20236 40256
rect 20276 40216 20277 40256
rect 20235 40207 20277 40216
rect 1152 40088 20452 40112
rect 1152 40048 4928 40088
rect 4968 40048 5010 40088
rect 5050 40048 5092 40088
rect 5132 40048 5174 40088
rect 5214 40048 5256 40088
rect 5296 40048 20048 40088
rect 20088 40048 20130 40088
rect 20170 40048 20212 40088
rect 20252 40048 20294 40088
rect 20334 40048 20376 40088
rect 20416 40048 20452 40088
rect 1152 40024 20452 40048
rect 3723 39920 3765 39929
rect 3723 39880 3724 39920
rect 3764 39880 3765 39920
rect 3723 39871 3765 39880
rect 5739 39920 5781 39929
rect 5739 39880 5740 39920
rect 5780 39880 5781 39920
rect 5739 39871 5781 39880
rect 9387 39920 9429 39929
rect 9387 39880 9388 39920
rect 9428 39880 9429 39920
rect 9387 39871 9429 39880
rect 19563 39920 19605 39929
rect 19563 39880 19564 39920
rect 19604 39880 19605 39920
rect 19563 39871 19605 39880
rect 19947 39920 19989 39929
rect 19947 39880 19948 39920
rect 19988 39880 19989 39920
rect 19947 39871 19989 39880
rect 1995 39752 2037 39761
rect 1995 39712 1996 39752
rect 2036 39712 2037 39752
rect 1995 39703 2037 39712
rect 2091 39752 2133 39761
rect 2091 39712 2092 39752
rect 2132 39712 2133 39752
rect 2091 39703 2133 39712
rect 3043 39752 3101 39753
rect 3043 39712 3052 39752
rect 3092 39712 3101 39752
rect 3043 39711 3101 39712
rect 3531 39747 3573 39756
rect 3531 39707 3532 39747
rect 3572 39707 3573 39747
rect 3531 39698 3573 39707
rect 4011 39752 4053 39761
rect 4011 39712 4012 39752
rect 4052 39712 4053 39752
rect 4011 39703 4053 39712
rect 4107 39752 4149 39761
rect 4107 39712 4108 39752
rect 4148 39712 4149 39752
rect 4107 39703 4149 39712
rect 5059 39752 5117 39753
rect 5059 39712 5068 39752
rect 5108 39712 5117 39752
rect 5059 39711 5117 39712
rect 5547 39747 5589 39756
rect 5547 39707 5548 39747
rect 5588 39707 5589 39747
rect 5547 39698 5589 39707
rect 5931 39752 5973 39761
rect 5931 39712 5932 39752
rect 5972 39712 5973 39752
rect 5931 39703 5973 39712
rect 6123 39752 6165 39761
rect 6123 39712 6124 39752
rect 6164 39712 6165 39752
rect 6123 39703 6165 39712
rect 6219 39752 6261 39761
rect 6219 39712 6220 39752
rect 6260 39712 6261 39752
rect 6219 39703 6261 39712
rect 6403 39752 6461 39753
rect 6403 39712 6412 39752
rect 6452 39712 6461 39752
rect 6403 39711 6461 39712
rect 6499 39752 6557 39753
rect 6499 39712 6508 39752
rect 6548 39712 6557 39752
rect 6499 39711 6557 39712
rect 6699 39752 6741 39761
rect 6699 39712 6700 39752
rect 6740 39712 6741 39752
rect 6699 39703 6741 39712
rect 6795 39752 6837 39761
rect 6795 39712 6796 39752
rect 6836 39712 6837 39752
rect 6795 39703 6837 39712
rect 6888 39752 6946 39753
rect 6888 39712 6897 39752
rect 6937 39712 6946 39752
rect 6888 39711 6946 39712
rect 7651 39752 7709 39753
rect 7651 39712 7660 39752
rect 7700 39712 7709 39752
rect 7651 39711 7709 39712
rect 8899 39752 8957 39753
rect 8899 39712 8908 39752
rect 8948 39712 8957 39752
rect 8899 39711 8957 39712
rect 10627 39752 10685 39753
rect 10627 39712 10636 39752
rect 10676 39712 10685 39752
rect 10627 39711 10685 39712
rect 11875 39752 11933 39753
rect 11875 39712 11884 39752
rect 11924 39712 11933 39752
rect 11875 39711 11933 39712
rect 12651 39752 12693 39761
rect 12651 39712 12652 39752
rect 12692 39712 12693 39752
rect 12651 39703 12693 39712
rect 12843 39752 12885 39761
rect 12843 39712 12844 39752
rect 12884 39712 12885 39752
rect 12843 39703 12885 39712
rect 12939 39752 12981 39761
rect 12939 39712 12940 39752
rect 12980 39712 12981 39752
rect 12939 39703 12981 39712
rect 2475 39668 2517 39677
rect 2475 39628 2476 39668
rect 2516 39628 2517 39668
rect 2475 39619 2517 39628
rect 2571 39668 2613 39677
rect 2571 39628 2572 39668
rect 2612 39628 2613 39668
rect 2571 39619 2613 39628
rect 4491 39668 4533 39677
rect 4491 39628 4492 39668
rect 4532 39628 4533 39668
rect 4491 39619 4533 39628
rect 4587 39668 4629 39677
rect 4587 39628 4588 39668
rect 4628 39628 4629 39668
rect 4587 39619 4629 39628
rect 18979 39668 19037 39669
rect 18979 39628 18988 39668
rect 19028 39628 19037 39668
rect 18979 39627 19037 39628
rect 19363 39668 19421 39669
rect 19363 39628 19372 39668
rect 19412 39628 19421 39668
rect 19363 39627 19421 39628
rect 19747 39668 19805 39669
rect 19747 39628 19756 39668
rect 19796 39628 19805 39668
rect 19747 39627 19805 39628
rect 6211 39584 6269 39585
rect 6211 39544 6220 39584
rect 6260 39544 6269 39584
rect 6211 39543 6269 39544
rect 9291 39584 9333 39593
rect 9291 39544 9292 39584
rect 9332 39544 9333 39584
rect 9291 39535 9333 39544
rect 12835 39584 12893 39585
rect 12835 39544 12844 39584
rect 12884 39544 12893 39584
rect 12835 39543 12893 39544
rect 6411 39500 6453 39509
rect 6411 39460 6412 39500
rect 6452 39460 6453 39500
rect 6411 39451 6453 39460
rect 9099 39500 9141 39509
rect 9099 39460 9100 39500
rect 9140 39460 9141 39500
rect 9099 39451 9141 39460
rect 10443 39500 10485 39509
rect 10443 39460 10444 39500
rect 10484 39460 10485 39500
rect 10443 39451 10485 39460
rect 19179 39500 19221 39509
rect 19179 39460 19180 39500
rect 19220 39460 19221 39500
rect 19179 39451 19221 39460
rect 1152 39332 20352 39356
rect 1152 39292 3688 39332
rect 3728 39292 3770 39332
rect 3810 39292 3852 39332
rect 3892 39292 3934 39332
rect 3974 39292 4016 39332
rect 4056 39292 18808 39332
rect 18848 39292 18890 39332
rect 18930 39292 18972 39332
rect 19012 39292 19054 39332
rect 19094 39292 19136 39332
rect 19176 39292 20352 39332
rect 1152 39268 20352 39292
rect 3435 39164 3477 39173
rect 3435 39124 3436 39164
rect 3476 39124 3477 39164
rect 3435 39115 3477 39124
rect 6699 39164 6741 39173
rect 6699 39124 6700 39164
rect 6740 39124 6741 39164
rect 6699 39115 6741 39124
rect 12939 39164 12981 39173
rect 12939 39124 12940 39164
rect 12980 39124 12981 39164
rect 12939 39115 12981 39124
rect 9195 38996 9237 39005
rect 9195 38956 9196 38996
rect 9236 38956 9237 38996
rect 9195 38947 9237 38956
rect 14467 38996 14525 38997
rect 14467 38956 14476 38996
rect 14516 38956 14525 38996
rect 14467 38955 14525 38956
rect 19363 38996 19421 38997
rect 19363 38956 19372 38996
rect 19412 38956 19421 38996
rect 19363 38955 19421 38956
rect 12739 38954 12797 38955
rect 10155 38926 10197 38935
rect 1987 38912 2045 38913
rect 1987 38872 1996 38912
rect 2036 38872 2045 38912
rect 1987 38871 2045 38872
rect 3235 38912 3293 38913
rect 3235 38872 3244 38912
rect 3284 38872 3293 38912
rect 3235 38871 3293 38872
rect 3619 38912 3677 38913
rect 3619 38872 3628 38912
rect 3668 38872 3677 38912
rect 3619 38871 3677 38872
rect 4867 38912 4925 38913
rect 4867 38872 4876 38912
rect 4916 38872 4925 38912
rect 4867 38871 4925 38872
rect 5251 38912 5309 38913
rect 5251 38872 5260 38912
rect 5300 38872 5309 38912
rect 5251 38871 5309 38872
rect 6499 38912 6557 38913
rect 6499 38872 6508 38912
rect 6548 38872 6557 38912
rect 6499 38871 6557 38872
rect 6883 38912 6941 38913
rect 6883 38872 6892 38912
rect 6932 38872 6941 38912
rect 6883 38871 6941 38872
rect 8131 38912 8189 38913
rect 8131 38872 8140 38912
rect 8180 38872 8189 38912
rect 8131 38871 8189 38872
rect 8619 38912 8661 38921
rect 8619 38872 8620 38912
rect 8660 38872 8661 38912
rect 8619 38863 8661 38872
rect 8715 38912 8757 38921
rect 8715 38872 8716 38912
rect 8756 38872 8757 38912
rect 8715 38863 8757 38872
rect 9099 38912 9141 38921
rect 9099 38872 9100 38912
rect 9140 38872 9141 38912
rect 9099 38863 9141 38872
rect 9667 38912 9725 38913
rect 9667 38872 9676 38912
rect 9716 38872 9725 38912
rect 10155 38886 10156 38926
rect 10196 38886 10197 38926
rect 12739 38914 12748 38954
rect 12788 38914 12797 38954
rect 12739 38913 12797 38914
rect 10155 38877 10197 38886
rect 11491 38912 11549 38913
rect 9667 38871 9725 38872
rect 11491 38872 11500 38912
rect 11540 38872 11549 38912
rect 11491 38871 11549 38872
rect 13131 38912 13173 38921
rect 13131 38872 13132 38912
rect 13172 38872 13173 38912
rect 13131 38863 13173 38872
rect 13419 38912 13461 38921
rect 13419 38872 13420 38912
rect 13460 38872 13461 38912
rect 13419 38863 13461 38872
rect 8331 38828 8373 38837
rect 8331 38788 8332 38828
rect 8372 38788 8373 38828
rect 8331 38779 8373 38788
rect 5067 38744 5109 38753
rect 5067 38704 5068 38744
rect 5108 38704 5109 38744
rect 5067 38695 5109 38704
rect 10347 38744 10389 38753
rect 10347 38704 10348 38744
rect 10388 38704 10389 38744
rect 10347 38695 10389 38704
rect 13323 38744 13365 38753
rect 13323 38704 13324 38744
rect 13364 38704 13365 38744
rect 13323 38695 13365 38704
rect 14667 38744 14709 38753
rect 14667 38704 14668 38744
rect 14708 38704 14709 38744
rect 14667 38695 14709 38704
rect 19563 38744 19605 38753
rect 19563 38704 19564 38744
rect 19604 38704 19605 38744
rect 19563 38695 19605 38704
rect 1152 38576 20452 38600
rect 1152 38536 4928 38576
rect 4968 38536 5010 38576
rect 5050 38536 5092 38576
rect 5132 38536 5174 38576
rect 5214 38536 5256 38576
rect 5296 38536 20048 38576
rect 20088 38536 20130 38576
rect 20170 38536 20212 38576
rect 20252 38536 20294 38576
rect 20334 38536 20376 38576
rect 20416 38536 20452 38576
rect 1152 38512 20452 38536
rect 3051 38408 3093 38417
rect 3051 38368 3052 38408
rect 3092 38368 3093 38408
rect 3051 38359 3093 38368
rect 7179 38408 7221 38417
rect 7179 38368 7180 38408
rect 7220 38368 7221 38408
rect 7179 38359 7221 38368
rect 7459 38408 7517 38409
rect 7459 38368 7468 38408
rect 7508 38368 7517 38408
rect 7459 38367 7517 38368
rect 8043 38408 8085 38417
rect 8043 38368 8044 38408
rect 8084 38368 8085 38408
rect 8043 38359 8085 38368
rect 12939 38408 12981 38417
rect 12939 38368 12940 38408
rect 12980 38368 12981 38408
rect 12939 38359 12981 38368
rect 14571 38408 14613 38417
rect 14571 38368 14572 38408
rect 14612 38368 14613 38408
rect 14571 38359 14613 38368
rect 5163 38324 5205 38333
rect 5163 38284 5164 38324
rect 5204 38284 5205 38324
rect 5163 38275 5205 38284
rect 10251 38324 10293 38333
rect 10251 38284 10252 38324
rect 10292 38284 10293 38324
rect 10251 38275 10293 38284
rect 13803 38324 13845 38333
rect 13803 38284 13804 38324
rect 13844 38284 13845 38324
rect 13803 38275 13845 38284
rect 1603 38240 1661 38241
rect 1603 38200 1612 38240
rect 1652 38200 1661 38240
rect 1603 38199 1661 38200
rect 2851 38240 2909 38241
rect 2851 38200 2860 38240
rect 2900 38200 2909 38240
rect 2851 38199 2909 38200
rect 3715 38240 3773 38241
rect 3715 38200 3724 38240
rect 3764 38200 3773 38240
rect 3715 38199 3773 38200
rect 4963 38240 5021 38241
rect 4963 38200 4972 38240
rect 5012 38200 5021 38240
rect 4963 38199 5021 38200
rect 5451 38240 5493 38249
rect 5451 38200 5452 38240
rect 5492 38200 5493 38240
rect 5451 38191 5493 38200
rect 5547 38240 5589 38249
rect 5547 38200 5548 38240
rect 5588 38200 5589 38240
rect 5547 38191 5589 38200
rect 6499 38240 6557 38241
rect 6499 38200 6508 38240
rect 6548 38200 6557 38240
rect 6499 38199 6557 38200
rect 6987 38235 7029 38244
rect 6987 38195 6988 38235
rect 7028 38195 7029 38235
rect 6987 38186 7029 38195
rect 7659 38240 7701 38249
rect 7659 38200 7660 38240
rect 7700 38200 7701 38240
rect 7659 38191 7701 38200
rect 7755 38240 7797 38249
rect 7755 38200 7756 38240
rect 7796 38200 7797 38240
rect 7755 38191 7797 38200
rect 7939 38240 7997 38241
rect 7939 38200 7948 38240
rect 7988 38200 7997 38240
rect 7939 38199 7997 38200
rect 8523 38240 8565 38249
rect 8523 38200 8524 38240
rect 8564 38200 8565 38240
rect 8523 38191 8565 38200
rect 8619 38240 8661 38249
rect 8619 38200 8620 38240
rect 8660 38200 8661 38240
rect 8619 38191 8661 38200
rect 9003 38240 9045 38249
rect 9003 38200 9004 38240
rect 9044 38200 9045 38240
rect 9003 38191 9045 38200
rect 9099 38240 9141 38249
rect 9099 38200 9100 38240
rect 9140 38200 9141 38240
rect 9099 38191 9141 38200
rect 9571 38240 9629 38241
rect 9571 38200 9580 38240
rect 9620 38200 9629 38240
rect 11491 38240 11549 38241
rect 9571 38199 9629 38200
rect 10059 38226 10101 38235
rect 10059 38186 10060 38226
rect 10100 38186 10101 38226
rect 11491 38200 11500 38240
rect 11540 38200 11549 38240
rect 11491 38199 11549 38200
rect 12739 38240 12797 38241
rect 12739 38200 12748 38240
rect 12788 38200 12797 38240
rect 12739 38199 12797 38200
rect 13131 38240 13173 38249
rect 13131 38200 13132 38240
rect 13172 38200 13173 38240
rect 13131 38191 13173 38200
rect 13323 38240 13365 38249
rect 13323 38200 13324 38240
rect 13364 38200 13365 38240
rect 13323 38191 13365 38200
rect 13419 38240 13461 38249
rect 13419 38200 13420 38240
rect 13460 38200 13461 38240
rect 13419 38191 13461 38200
rect 13603 38240 13661 38241
rect 13603 38200 13612 38240
rect 13652 38200 13661 38240
rect 13603 38199 13661 38200
rect 13707 38240 13749 38249
rect 13707 38200 13708 38240
rect 13748 38200 13749 38240
rect 13707 38191 13749 38200
rect 13899 38240 13941 38249
rect 13899 38200 13900 38240
rect 13940 38200 13941 38240
rect 13899 38191 13941 38200
rect 14091 38240 14133 38249
rect 14091 38200 14092 38240
rect 14132 38200 14133 38240
rect 14091 38191 14133 38200
rect 14179 38240 14237 38241
rect 14179 38200 14188 38240
rect 14228 38200 14237 38240
rect 14179 38199 14237 38200
rect 10059 38177 10101 38186
rect 5931 38156 5973 38165
rect 5931 38116 5932 38156
rect 5972 38116 5973 38156
rect 5931 38107 5973 38116
rect 6027 38156 6069 38165
rect 6027 38116 6028 38156
rect 6068 38116 6069 38156
rect 6027 38107 6069 38116
rect 14371 38156 14429 38157
rect 14371 38116 14380 38156
rect 14420 38116 14429 38156
rect 18595 38156 18653 38157
rect 14371 38115 14429 38116
rect 15331 38145 15389 38146
rect 15331 38105 15340 38145
rect 15380 38105 15389 38145
rect 18595 38116 18604 38156
rect 18644 38116 18653 38156
rect 18595 38115 18653 38116
rect 19363 38156 19421 38157
rect 19363 38116 19372 38156
rect 19412 38116 19421 38156
rect 19363 38115 19421 38116
rect 15331 38104 15389 38105
rect 13411 38072 13469 38073
rect 13411 38032 13420 38072
rect 13460 38032 13469 38072
rect 13411 38031 13469 38032
rect 15531 38072 15573 38081
rect 15531 38032 15532 38072
rect 15572 38032 15573 38072
rect 15531 38023 15573 38032
rect 19563 38072 19605 38081
rect 19563 38032 19564 38072
rect 19604 38032 19605 38072
rect 19563 38023 19605 38032
rect 12939 37988 12981 37997
rect 12939 37948 12940 37988
rect 12980 37948 12981 37988
rect 12939 37939 12981 37948
rect 18795 37988 18837 37997
rect 18795 37948 18796 37988
rect 18836 37948 18837 37988
rect 18795 37939 18837 37948
rect 1152 37820 20352 37844
rect 1152 37780 3688 37820
rect 3728 37780 3770 37820
rect 3810 37780 3852 37820
rect 3892 37780 3934 37820
rect 3974 37780 4016 37820
rect 4056 37780 18808 37820
rect 18848 37780 18890 37820
rect 18930 37780 18972 37820
rect 19012 37780 19054 37820
rect 19094 37780 19136 37820
rect 19176 37780 20352 37820
rect 1152 37756 20352 37780
rect 15051 37652 15093 37661
rect 15051 37612 15052 37652
rect 15092 37612 15093 37652
rect 15051 37603 15093 37612
rect 19947 37652 19989 37661
rect 19947 37612 19948 37652
rect 19988 37612 19989 37652
rect 19947 37603 19989 37612
rect 10443 37568 10485 37577
rect 10443 37528 10444 37568
rect 10484 37528 10485 37568
rect 10443 37519 10485 37528
rect 11875 37568 11933 37569
rect 11875 37528 11884 37568
rect 11924 37528 11933 37568
rect 11875 37527 11933 37528
rect 12555 37568 12597 37577
rect 12555 37528 12556 37568
rect 12596 37528 12597 37568
rect 12555 37519 12597 37528
rect 19563 37568 19605 37577
rect 19563 37528 19564 37568
rect 19604 37528 19605 37568
rect 19563 37519 19605 37528
rect 18979 37484 19037 37485
rect 18979 37444 18988 37484
rect 19028 37444 19037 37484
rect 18979 37443 19037 37444
rect 19363 37484 19421 37485
rect 19363 37444 19372 37484
rect 19412 37444 19421 37484
rect 19363 37443 19421 37444
rect 19747 37484 19805 37485
rect 19747 37444 19756 37484
rect 19796 37444 19805 37484
rect 19747 37443 19805 37444
rect 3963 37409 4005 37418
rect 2379 37400 2421 37409
rect 2379 37360 2380 37400
rect 2420 37360 2421 37400
rect 2379 37351 2421 37360
rect 2475 37400 2517 37409
rect 2475 37360 2476 37400
rect 2516 37360 2517 37400
rect 2475 37351 2517 37360
rect 2859 37400 2901 37409
rect 2859 37360 2860 37400
rect 2900 37360 2901 37400
rect 2859 37351 2901 37360
rect 2955 37400 2997 37409
rect 2955 37360 2956 37400
rect 2996 37360 2997 37400
rect 2955 37351 2997 37360
rect 3427 37400 3485 37401
rect 3427 37360 3436 37400
rect 3476 37360 3485 37400
rect 3963 37369 3964 37409
rect 4004 37369 4005 37409
rect 3963 37360 4005 37369
rect 4291 37400 4349 37401
rect 4291 37360 4300 37400
rect 4340 37360 4349 37400
rect 3427 37359 3485 37360
rect 4291 37359 4349 37360
rect 5539 37400 5597 37401
rect 5539 37360 5548 37400
rect 5588 37360 5597 37400
rect 5539 37359 5597 37360
rect 6027 37400 6069 37409
rect 6027 37360 6028 37400
rect 6068 37360 6069 37400
rect 6027 37351 6069 37360
rect 6123 37400 6165 37409
rect 6123 37360 6124 37400
rect 6164 37360 6165 37400
rect 6123 37351 6165 37360
rect 6507 37400 6549 37409
rect 6507 37360 6508 37400
rect 6548 37360 6549 37400
rect 6507 37351 6549 37360
rect 6603 37400 6645 37409
rect 7563 37405 7605 37414
rect 6603 37360 6604 37400
rect 6644 37360 6645 37400
rect 6603 37351 6645 37360
rect 7075 37400 7133 37401
rect 7075 37360 7084 37400
rect 7124 37360 7133 37400
rect 7075 37359 7133 37360
rect 7563 37365 7564 37405
rect 7604 37365 7605 37405
rect 7563 37356 7605 37365
rect 8995 37400 9053 37401
rect 8995 37360 9004 37400
rect 9044 37360 9053 37400
rect 8995 37359 9053 37360
rect 10243 37400 10301 37401
rect 10243 37360 10252 37400
rect 10292 37360 10301 37400
rect 10243 37359 10301 37360
rect 11115 37400 11157 37409
rect 11115 37360 11116 37400
rect 11156 37360 11157 37400
rect 11115 37351 11157 37360
rect 11307 37400 11349 37409
rect 11307 37360 11308 37400
rect 11348 37360 11349 37400
rect 11307 37351 11349 37360
rect 11395 37400 11453 37401
rect 11395 37360 11404 37400
rect 11444 37360 11453 37400
rect 11395 37359 11453 37360
rect 11595 37400 11637 37409
rect 11595 37360 11596 37400
rect 11636 37360 11637 37400
rect 11595 37351 11637 37360
rect 11787 37400 11829 37409
rect 11787 37360 11788 37400
rect 11828 37360 11829 37400
rect 11787 37351 11829 37360
rect 11883 37400 11925 37409
rect 11883 37360 11884 37400
rect 11924 37360 11925 37400
rect 11883 37351 11925 37360
rect 12075 37400 12117 37409
rect 12075 37360 12076 37400
rect 12116 37360 12117 37400
rect 12075 37351 12117 37360
rect 12267 37400 12309 37409
rect 12267 37360 12268 37400
rect 12308 37360 12309 37400
rect 12267 37351 12309 37360
rect 12355 37400 12413 37401
rect 12355 37360 12364 37400
rect 12404 37360 12413 37400
rect 12355 37359 12413 37360
rect 12555 37400 12597 37409
rect 12555 37360 12556 37400
rect 12596 37360 12597 37400
rect 12555 37351 12597 37360
rect 12843 37400 12885 37409
rect 12843 37360 12844 37400
rect 12884 37360 12885 37400
rect 12843 37351 12885 37360
rect 13027 37400 13085 37401
rect 13027 37360 13036 37400
rect 13076 37360 13085 37400
rect 13027 37359 13085 37360
rect 13131 37400 13173 37409
rect 13131 37360 13132 37400
rect 13172 37360 13173 37400
rect 13131 37351 13173 37360
rect 13315 37400 13373 37401
rect 13315 37360 13324 37400
rect 13364 37360 13373 37400
rect 13315 37359 13373 37360
rect 13603 37400 13661 37401
rect 13603 37360 13612 37400
rect 13652 37360 13661 37400
rect 13603 37359 13661 37360
rect 14851 37400 14909 37401
rect 14851 37360 14860 37400
rect 14900 37360 14909 37400
rect 14851 37359 14909 37360
rect 5739 37316 5781 37325
rect 5739 37276 5740 37316
rect 5780 37276 5781 37316
rect 5739 37267 5781 37276
rect 12171 37316 12213 37325
rect 12171 37276 12172 37316
rect 12212 37276 12213 37316
rect 12171 37267 12213 37276
rect 4107 37232 4149 37241
rect 4107 37192 4108 37232
rect 4148 37192 4149 37232
rect 4107 37183 4149 37192
rect 7755 37232 7797 37241
rect 7755 37192 7756 37232
rect 7796 37192 7797 37232
rect 7755 37183 7797 37192
rect 11203 37232 11261 37233
rect 11203 37192 11212 37232
rect 11252 37192 11261 37232
rect 11203 37191 11261 37192
rect 13323 37232 13365 37241
rect 13323 37192 13324 37232
rect 13364 37192 13365 37232
rect 13323 37183 13365 37192
rect 19179 37232 19221 37241
rect 19179 37192 19180 37232
rect 19220 37192 19221 37232
rect 19179 37183 19221 37192
rect 1152 37064 20452 37088
rect 1152 37024 4928 37064
rect 4968 37024 5010 37064
rect 5050 37024 5092 37064
rect 5132 37024 5174 37064
rect 5214 37024 5256 37064
rect 5296 37024 20048 37064
rect 20088 37024 20130 37064
rect 20170 37024 20212 37064
rect 20252 37024 20294 37064
rect 20334 37024 20376 37064
rect 20416 37024 20452 37064
rect 1152 37000 20452 37024
rect 2667 36896 2709 36905
rect 2667 36856 2668 36896
rect 2708 36856 2709 36896
rect 2667 36847 2709 36856
rect 4299 36896 4341 36905
rect 4299 36856 4300 36896
rect 4340 36856 4341 36896
rect 4299 36847 4341 36856
rect 8907 36896 8949 36905
rect 8907 36856 8908 36896
rect 8948 36856 8949 36896
rect 8907 36847 8949 36856
rect 10827 36896 10869 36905
rect 10827 36856 10828 36896
rect 10868 36856 10869 36896
rect 10827 36847 10869 36856
rect 12355 36896 12413 36897
rect 12355 36856 12364 36896
rect 12404 36856 12413 36896
rect 12355 36855 12413 36856
rect 13035 36896 13077 36905
rect 13035 36856 13036 36896
rect 13076 36856 13077 36896
rect 13035 36847 13077 36856
rect 13795 36896 13853 36897
rect 13795 36856 13804 36896
rect 13844 36856 13853 36896
rect 13795 36855 13853 36856
rect 19563 36896 19605 36905
rect 19563 36856 19564 36896
rect 19604 36856 19605 36896
rect 19563 36847 19605 36856
rect 11299 36743 11357 36744
rect 1219 36728 1277 36729
rect 1219 36688 1228 36728
rect 1268 36688 1277 36728
rect 1219 36687 1277 36688
rect 2467 36728 2525 36729
rect 2467 36688 2476 36728
rect 2516 36688 2525 36728
rect 2467 36687 2525 36688
rect 2851 36728 2909 36729
rect 2851 36688 2860 36728
rect 2900 36688 2909 36728
rect 2851 36687 2909 36688
rect 4099 36728 4157 36729
rect 4099 36688 4108 36728
rect 4148 36688 4157 36728
rect 4099 36687 4157 36688
rect 4483 36728 4541 36729
rect 4483 36688 4492 36728
rect 4532 36688 4541 36728
rect 4483 36687 4541 36688
rect 4683 36728 4725 36737
rect 4683 36688 4684 36728
rect 4724 36688 4725 36728
rect 4683 36679 4725 36688
rect 4771 36728 4829 36729
rect 4771 36688 4780 36728
rect 4820 36688 4829 36728
rect 4771 36687 4829 36688
rect 4963 36728 5021 36729
rect 4963 36688 4972 36728
rect 5012 36688 5021 36728
rect 4963 36687 5021 36688
rect 5163 36728 5205 36737
rect 5163 36688 5164 36728
rect 5204 36688 5205 36728
rect 5163 36679 5205 36688
rect 5827 36728 5885 36729
rect 5827 36688 5836 36728
rect 5876 36688 5885 36728
rect 5827 36687 5885 36688
rect 7075 36728 7133 36729
rect 7075 36688 7084 36728
rect 7124 36688 7133 36728
rect 7075 36687 7133 36688
rect 7459 36728 7517 36729
rect 7459 36688 7468 36728
rect 7508 36688 7517 36728
rect 7459 36687 7517 36688
rect 8707 36728 8765 36729
rect 8707 36688 8716 36728
rect 8756 36688 8765 36728
rect 8707 36687 8765 36688
rect 10243 36728 10301 36729
rect 10243 36688 10252 36728
rect 10292 36688 10301 36728
rect 10243 36687 10301 36688
rect 10347 36728 10389 36737
rect 10347 36688 10348 36728
rect 10388 36688 10389 36728
rect 10347 36679 10389 36688
rect 10539 36728 10581 36737
rect 10539 36688 10540 36728
rect 10580 36688 10581 36728
rect 10539 36679 10581 36688
rect 10731 36728 10773 36737
rect 10731 36688 10732 36728
rect 10772 36688 10773 36728
rect 10731 36679 10773 36688
rect 10923 36728 10965 36737
rect 10923 36688 10924 36728
rect 10964 36688 10965 36728
rect 10923 36679 10965 36688
rect 11019 36728 11061 36737
rect 11019 36688 11020 36728
rect 11060 36688 11061 36728
rect 11299 36703 11308 36743
rect 11348 36703 11357 36743
rect 11299 36702 11357 36703
rect 11595 36728 11637 36737
rect 11019 36679 11061 36688
rect 11595 36688 11596 36728
rect 11636 36688 11637 36728
rect 11595 36679 11637 36688
rect 11691 36728 11733 36737
rect 11691 36688 11692 36728
rect 11732 36688 11733 36728
rect 11691 36679 11733 36688
rect 12163 36728 12221 36729
rect 12163 36688 12172 36728
rect 12212 36688 12221 36728
rect 12163 36687 12221 36688
rect 12259 36728 12317 36729
rect 12259 36688 12268 36728
rect 12308 36688 12317 36728
rect 12259 36687 12317 36688
rect 12459 36728 12501 36737
rect 12459 36688 12460 36728
rect 12500 36688 12501 36728
rect 12459 36679 12501 36688
rect 12555 36728 12597 36737
rect 12555 36688 12556 36728
rect 12596 36688 12597 36728
rect 12555 36679 12597 36688
rect 12648 36728 12706 36729
rect 12648 36688 12657 36728
rect 12697 36688 12706 36728
rect 12648 36687 12706 36688
rect 12931 36728 12989 36729
rect 12931 36688 12940 36728
rect 12980 36688 12989 36728
rect 12931 36687 12989 36688
rect 13227 36728 13269 36737
rect 13227 36688 13228 36728
rect 13268 36688 13269 36728
rect 13227 36679 13269 36688
rect 13603 36728 13661 36729
rect 13603 36688 13612 36728
rect 13652 36688 13661 36728
rect 13603 36687 13661 36688
rect 13899 36728 13941 36737
rect 13899 36688 13900 36728
rect 13940 36688 13941 36728
rect 13899 36679 13941 36688
rect 13995 36728 14037 36737
rect 13995 36688 13996 36728
rect 14036 36688 14037 36728
rect 13995 36679 14037 36688
rect 14091 36728 14133 36737
rect 14091 36688 14092 36728
rect 14132 36688 14133 36728
rect 14091 36679 14133 36688
rect 14275 36728 14333 36729
rect 14275 36688 14284 36728
rect 14324 36688 14333 36728
rect 14275 36687 14333 36688
rect 13323 36644 13365 36653
rect 13323 36604 13324 36644
rect 13364 36604 13365 36644
rect 13323 36595 13365 36604
rect 13515 36644 13557 36653
rect 13515 36604 13516 36644
rect 13556 36604 13557 36644
rect 13515 36595 13557 36604
rect 18979 36644 19037 36645
rect 18979 36604 18988 36644
rect 19028 36604 19037 36644
rect 18979 36603 19037 36604
rect 19363 36644 19421 36645
rect 19363 36604 19372 36644
rect 19412 36604 19421 36644
rect 19363 36603 19421 36604
rect 5067 36560 5109 36569
rect 5067 36520 5068 36560
rect 5108 36520 5109 36560
rect 5067 36511 5109 36520
rect 7275 36560 7317 36569
rect 7275 36520 7276 36560
rect 7316 36520 7317 36560
rect 7275 36511 7317 36520
rect 10539 36560 10581 36569
rect 10539 36520 10540 36560
rect 10580 36520 10581 36560
rect 10539 36511 10581 36520
rect 11971 36560 12029 36561
rect 11971 36520 11980 36560
rect 12020 36520 12029 36560
rect 11971 36519 12029 36520
rect 13419 36560 13461 36569
rect 13419 36520 13420 36560
rect 13460 36520 13461 36560
rect 13419 36511 13461 36520
rect 14379 36560 14421 36569
rect 14379 36520 14380 36560
rect 14420 36520 14421 36560
rect 14379 36511 14421 36520
rect 4491 36476 4533 36485
rect 4491 36436 4492 36476
rect 4532 36436 4533 36476
rect 4491 36427 4533 36436
rect 19179 36476 19221 36485
rect 19179 36436 19180 36476
rect 19220 36436 19221 36476
rect 19179 36427 19221 36436
rect 1152 36308 20352 36332
rect 1152 36268 3688 36308
rect 3728 36268 3770 36308
rect 3810 36268 3852 36308
rect 3892 36268 3934 36308
rect 3974 36268 4016 36308
rect 4056 36268 18808 36308
rect 18848 36268 18890 36308
rect 18930 36268 18972 36308
rect 19012 36268 19054 36308
rect 19094 36268 19136 36308
rect 19176 36268 20352 36308
rect 1152 36244 20352 36268
rect 2667 36140 2709 36149
rect 2667 36100 2668 36140
rect 2708 36100 2709 36140
rect 2667 36091 2709 36100
rect 4299 36140 4341 36149
rect 4299 36100 4300 36140
rect 4340 36100 4341 36140
rect 4299 36091 4341 36100
rect 11019 36140 11061 36149
rect 11019 36100 11020 36140
rect 11060 36100 11061 36140
rect 11019 36091 11061 36100
rect 12267 36140 12309 36149
rect 12267 36100 12268 36140
rect 12308 36100 12309 36140
rect 12267 36091 12309 36100
rect 19563 36140 19605 36149
rect 19563 36100 19564 36140
rect 19604 36100 19605 36140
rect 19563 36091 19605 36100
rect 13315 36056 13373 36057
rect 13315 36016 13324 36056
rect 13364 36016 13373 36056
rect 13315 36015 13373 36016
rect 19179 36056 19221 36065
rect 19179 36016 19180 36056
rect 19220 36016 19221 36056
rect 19179 36007 19221 36016
rect 10443 35972 10485 35981
rect 10443 35932 10444 35972
rect 10484 35932 10485 35972
rect 10443 35923 10485 35932
rect 18979 35972 19037 35973
rect 18979 35932 18988 35972
rect 19028 35932 19037 35972
rect 18979 35931 19037 35932
rect 19363 35972 19421 35973
rect 19363 35932 19372 35972
rect 19412 35932 19421 35972
rect 19363 35931 19421 35932
rect 19747 35972 19805 35973
rect 19747 35932 19756 35972
rect 19796 35932 19805 35972
rect 19747 35931 19805 35932
rect 9915 35897 9957 35906
rect 1219 35888 1277 35889
rect 1219 35848 1228 35888
rect 1268 35848 1277 35888
rect 1219 35847 1277 35848
rect 2467 35888 2525 35889
rect 2467 35848 2476 35888
rect 2516 35848 2525 35888
rect 2467 35847 2525 35848
rect 2851 35888 2909 35889
rect 2851 35848 2860 35888
rect 2900 35848 2909 35888
rect 2851 35847 2909 35848
rect 4099 35888 4157 35889
rect 4099 35848 4108 35888
rect 4148 35848 4157 35888
rect 4099 35847 4157 35848
rect 4491 35888 4533 35897
rect 4491 35848 4492 35888
rect 4532 35848 4533 35888
rect 4491 35839 4533 35848
rect 4587 35888 4629 35897
rect 4587 35848 4588 35888
rect 4628 35848 4629 35888
rect 4587 35839 4629 35848
rect 4963 35888 5021 35889
rect 4963 35848 4972 35888
rect 5012 35848 5021 35888
rect 4963 35847 5021 35848
rect 6211 35888 6269 35889
rect 6211 35848 6220 35888
rect 6260 35848 6269 35888
rect 6211 35847 6269 35848
rect 6595 35888 6653 35889
rect 6595 35848 6604 35888
rect 6644 35848 6653 35888
rect 6595 35847 6653 35848
rect 7843 35888 7901 35889
rect 7843 35848 7852 35888
rect 7892 35848 7901 35888
rect 7843 35847 7901 35848
rect 8331 35888 8373 35897
rect 8331 35848 8332 35888
rect 8372 35848 8373 35888
rect 8331 35839 8373 35848
rect 8427 35888 8469 35897
rect 8427 35848 8428 35888
rect 8468 35848 8469 35888
rect 8427 35839 8469 35848
rect 8811 35888 8853 35897
rect 8811 35848 8812 35888
rect 8852 35848 8853 35888
rect 8811 35839 8853 35848
rect 8907 35888 8949 35897
rect 8907 35848 8908 35888
rect 8948 35848 8949 35888
rect 8907 35839 8949 35848
rect 9379 35888 9437 35889
rect 9379 35848 9388 35888
rect 9428 35848 9437 35888
rect 9915 35857 9916 35897
rect 9956 35857 9957 35897
rect 9915 35848 9957 35857
rect 10251 35888 10293 35897
rect 10251 35848 10252 35888
rect 10292 35848 10293 35888
rect 9379 35847 9437 35848
rect 10251 35839 10293 35848
rect 10539 35888 10581 35897
rect 10539 35848 10540 35888
rect 10580 35848 10581 35888
rect 10539 35839 10581 35848
rect 10731 35888 10773 35897
rect 10731 35848 10732 35888
rect 10772 35848 10773 35888
rect 10731 35839 10773 35848
rect 11019 35888 11061 35897
rect 11019 35848 11020 35888
rect 11060 35848 11061 35888
rect 11019 35839 11061 35848
rect 11307 35888 11349 35897
rect 11307 35848 11308 35888
rect 11348 35848 11349 35888
rect 11307 35839 11349 35848
rect 11595 35888 11637 35897
rect 11595 35848 11596 35888
rect 11636 35848 11637 35888
rect 11595 35839 11637 35848
rect 11779 35888 11837 35889
rect 11779 35848 11788 35888
rect 11828 35848 11837 35888
rect 11779 35847 11837 35848
rect 11883 35888 11925 35897
rect 11883 35848 11884 35888
rect 11924 35848 11925 35888
rect 11883 35839 11925 35848
rect 12067 35888 12125 35889
rect 12067 35848 12076 35888
rect 12116 35848 12125 35888
rect 12067 35847 12125 35848
rect 12267 35888 12309 35897
rect 12267 35848 12268 35888
rect 12308 35848 12309 35888
rect 12267 35839 12309 35848
rect 12555 35888 12597 35897
rect 12555 35848 12556 35888
rect 12596 35848 12597 35888
rect 12555 35839 12597 35848
rect 12747 35888 12789 35897
rect 12747 35848 12748 35888
rect 12788 35848 12789 35888
rect 12747 35839 12789 35848
rect 12843 35888 12885 35897
rect 12843 35848 12844 35888
rect 12884 35848 12885 35888
rect 12843 35839 12885 35848
rect 13227 35888 13269 35897
rect 13227 35848 13228 35888
rect 13268 35848 13269 35888
rect 13227 35839 13269 35848
rect 13323 35888 13365 35897
rect 13323 35848 13324 35888
rect 13364 35848 13365 35888
rect 13323 35839 13365 35848
rect 13515 35888 13557 35897
rect 13515 35848 13516 35888
rect 13556 35848 13557 35888
rect 13515 35839 13557 35848
rect 13707 35888 13749 35897
rect 13707 35848 13708 35888
rect 13748 35848 13749 35888
rect 13707 35839 13749 35848
rect 13803 35888 13845 35897
rect 13803 35848 13804 35888
rect 13844 35848 13845 35888
rect 13803 35839 13845 35848
rect 13899 35888 13941 35897
rect 13899 35848 13900 35888
rect 13940 35848 13941 35888
rect 13899 35839 13941 35848
rect 13995 35888 14037 35897
rect 13995 35848 13996 35888
rect 14036 35848 14037 35888
rect 13995 35839 14037 35848
rect 14187 35888 14229 35897
rect 14187 35848 14188 35888
rect 14228 35848 14229 35888
rect 14187 35839 14229 35848
rect 14283 35888 14325 35897
rect 14283 35848 14284 35888
rect 14324 35848 14325 35888
rect 14283 35839 14325 35848
rect 14379 35888 14421 35897
rect 14379 35848 14380 35888
rect 14420 35848 14421 35888
rect 14379 35839 14421 35848
rect 8043 35804 8085 35813
rect 8043 35764 8044 35804
rect 8084 35764 8085 35804
rect 8043 35755 8085 35764
rect 4299 35720 4341 35729
rect 4299 35680 4300 35720
rect 4340 35680 4341 35720
rect 4299 35671 4341 35680
rect 4771 35720 4829 35721
rect 4771 35680 4780 35720
rect 4820 35680 4829 35720
rect 4771 35679 4829 35680
rect 6411 35720 6453 35729
rect 6411 35680 6412 35720
rect 6452 35680 6453 35720
rect 6411 35671 6453 35680
rect 10059 35720 10101 35729
rect 10059 35680 10060 35720
rect 10100 35680 10101 35720
rect 10059 35671 10101 35680
rect 11499 35720 11541 35729
rect 11499 35680 11500 35720
rect 11540 35680 11541 35720
rect 11499 35671 11541 35680
rect 12075 35720 12117 35729
rect 12075 35680 12076 35720
rect 12116 35680 12117 35720
rect 12075 35671 12117 35680
rect 13027 35720 13085 35721
rect 13027 35680 13036 35720
rect 13076 35680 13085 35720
rect 13027 35679 13085 35680
rect 14467 35720 14525 35721
rect 14467 35680 14476 35720
rect 14516 35680 14525 35720
rect 14467 35679 14525 35680
rect 19947 35720 19989 35729
rect 19947 35680 19948 35720
rect 19988 35680 19989 35720
rect 19947 35671 19989 35680
rect 1152 35552 20452 35576
rect 1152 35512 4928 35552
rect 4968 35512 5010 35552
rect 5050 35512 5092 35552
rect 5132 35512 5174 35552
rect 5214 35512 5256 35552
rect 5296 35512 20048 35552
rect 20088 35512 20130 35552
rect 20170 35512 20212 35552
rect 20252 35512 20294 35552
rect 20334 35512 20376 35552
rect 20416 35512 20452 35552
rect 1152 35488 20452 35512
rect 9963 35384 10005 35393
rect 9963 35344 9964 35384
rect 10004 35344 10005 35384
rect 9963 35335 10005 35344
rect 13219 35384 13277 35385
rect 13219 35344 13228 35384
rect 13268 35344 13277 35384
rect 13219 35343 13277 35344
rect 13699 35384 13757 35385
rect 13699 35344 13708 35384
rect 13748 35344 13757 35384
rect 13699 35343 13757 35344
rect 2859 35300 2901 35309
rect 2859 35260 2860 35300
rect 2900 35260 2901 35300
rect 2859 35251 2901 35260
rect 6603 35300 6645 35309
rect 6603 35260 6604 35300
rect 6644 35260 6645 35300
rect 6603 35251 6645 35260
rect 10539 35300 10581 35309
rect 10539 35260 10540 35300
rect 10580 35260 10581 35300
rect 6883 35258 6941 35259
rect 1411 35216 1469 35217
rect 1411 35176 1420 35216
rect 1460 35176 1469 35216
rect 1411 35175 1469 35176
rect 2659 35216 2717 35217
rect 2659 35176 2668 35216
rect 2708 35176 2717 35216
rect 2659 35175 2717 35176
rect 3051 35216 3093 35225
rect 3051 35176 3052 35216
rect 3092 35176 3093 35216
rect 3051 35167 3093 35176
rect 3243 35216 3285 35225
rect 3243 35176 3244 35216
rect 3284 35176 3285 35216
rect 3243 35167 3285 35176
rect 3723 35216 3765 35225
rect 3723 35176 3724 35216
rect 3764 35176 3765 35216
rect 3723 35167 3765 35176
rect 3819 35216 3861 35225
rect 3819 35176 3820 35216
rect 3860 35176 3861 35216
rect 3819 35167 3861 35176
rect 4099 35216 4157 35217
rect 4099 35176 4108 35216
rect 4148 35176 4157 35216
rect 4099 35175 4157 35176
rect 4483 35216 4541 35217
rect 4483 35176 4492 35216
rect 4532 35176 4541 35216
rect 4483 35175 4541 35176
rect 5731 35216 5789 35217
rect 5731 35176 5740 35216
rect 5780 35176 5789 35216
rect 5731 35175 5789 35176
rect 6403 35216 6461 35217
rect 6403 35176 6412 35216
rect 6452 35176 6461 35216
rect 6403 35175 6461 35176
rect 6507 35216 6549 35225
rect 6507 35176 6508 35216
rect 6548 35176 6549 35216
rect 6507 35167 6549 35176
rect 6699 35216 6741 35225
rect 6883 35218 6892 35258
rect 6932 35218 6941 35258
rect 10539 35251 10581 35260
rect 12555 35300 12597 35309
rect 12555 35260 12556 35300
rect 12596 35260 12597 35300
rect 12555 35251 12597 35260
rect 6883 35217 6941 35218
rect 6699 35176 6700 35216
rect 6740 35176 6741 35216
rect 6699 35167 6741 35176
rect 8131 35216 8189 35217
rect 8131 35176 8140 35216
rect 8180 35176 8189 35216
rect 8131 35175 8189 35176
rect 8515 35216 8573 35217
rect 8515 35176 8524 35216
rect 8564 35176 8573 35216
rect 8515 35175 8573 35176
rect 9763 35216 9821 35217
rect 9763 35176 9772 35216
rect 9812 35176 9821 35216
rect 9763 35175 9821 35176
rect 10443 35216 10485 35225
rect 10443 35176 10444 35216
rect 10484 35176 10485 35216
rect 10443 35167 10485 35176
rect 10627 35216 10685 35217
rect 10627 35176 10636 35216
rect 10676 35176 10685 35216
rect 10627 35175 10685 35176
rect 10827 35216 10869 35225
rect 10827 35176 10828 35216
rect 10868 35176 10869 35216
rect 10827 35167 10869 35176
rect 11115 35216 11157 35225
rect 11115 35176 11116 35216
rect 11156 35176 11157 35216
rect 11115 35167 11157 35176
rect 11395 35216 11453 35217
rect 11395 35176 11404 35216
rect 11444 35176 11453 35216
rect 11395 35175 11453 35176
rect 11691 35216 11733 35225
rect 11691 35176 11692 35216
rect 11732 35176 11733 35216
rect 11691 35167 11733 35176
rect 11787 35216 11829 35225
rect 11787 35176 11788 35216
rect 11828 35176 11829 35216
rect 11787 35167 11829 35176
rect 12267 35216 12309 35225
rect 12267 35176 12268 35216
rect 12308 35176 12309 35216
rect 12267 35167 12309 35176
rect 12363 35216 12405 35225
rect 12363 35176 12364 35216
rect 12404 35176 12405 35216
rect 12363 35167 12405 35176
rect 12459 35216 12501 35225
rect 12459 35176 12460 35216
rect 12500 35176 12501 35216
rect 12459 35167 12501 35176
rect 12939 35216 12981 35225
rect 12939 35176 12940 35216
rect 12980 35176 12981 35216
rect 12939 35167 12981 35176
rect 13035 35216 13077 35225
rect 13035 35176 13036 35216
rect 13076 35176 13077 35216
rect 13035 35167 13077 35176
rect 13131 35216 13173 35225
rect 13131 35176 13132 35216
rect 13172 35176 13173 35216
rect 13131 35167 13173 35176
rect 13419 35216 13461 35225
rect 13419 35176 13420 35216
rect 13460 35176 13461 35216
rect 13419 35167 13461 35176
rect 13515 35216 13557 35225
rect 13515 35176 13516 35216
rect 13556 35176 13557 35216
rect 13515 35167 13557 35176
rect 14275 35216 14333 35217
rect 14275 35176 14284 35216
rect 14324 35176 14333 35216
rect 14275 35175 14333 35176
rect 15523 35216 15581 35217
rect 15523 35176 15532 35216
rect 15572 35176 15581 35216
rect 15523 35175 15581 35176
rect 16387 35132 16445 35133
rect 16387 35092 16396 35132
rect 16436 35092 16445 35132
rect 16387 35091 16445 35092
rect 18979 35132 19037 35133
rect 18979 35092 18988 35132
rect 19028 35092 19037 35132
rect 18979 35091 19037 35092
rect 19363 35132 19421 35133
rect 19363 35092 19372 35132
rect 19412 35092 19421 35132
rect 19363 35091 19421 35092
rect 3427 35048 3485 35049
rect 3427 35008 3436 35048
rect 3476 35008 3485 35048
rect 3427 35007 3485 35008
rect 12067 35048 12125 35049
rect 12067 35008 12076 35048
rect 12116 35008 12125 35048
rect 12067 35007 12125 35008
rect 14091 35048 14133 35057
rect 14091 35008 14092 35048
rect 14132 35008 14133 35048
rect 14091 34999 14133 35008
rect 19179 35048 19221 35057
rect 19179 35008 19180 35048
rect 19220 35008 19221 35048
rect 19179 34999 19221 35008
rect 19563 35048 19605 35057
rect 19563 35008 19564 35048
rect 19604 35008 19605 35048
rect 19563 34999 19605 35008
rect 3243 34964 3285 34973
rect 3243 34924 3244 34964
rect 3284 34924 3285 34964
rect 3243 34915 3285 34924
rect 5931 34964 5973 34973
rect 5931 34924 5932 34964
rect 5972 34924 5973 34964
rect 5931 34915 5973 34924
rect 8331 34964 8373 34973
rect 8331 34924 8332 34964
rect 8372 34924 8373 34964
rect 8331 34915 8373 34924
rect 11115 34964 11157 34973
rect 11115 34924 11116 34964
rect 11156 34924 11157 34964
rect 11115 34915 11157 34924
rect 16587 34964 16629 34973
rect 16587 34924 16588 34964
rect 16628 34924 16629 34964
rect 16587 34915 16629 34924
rect 1152 34796 20352 34820
rect 1152 34756 3688 34796
rect 3728 34756 3770 34796
rect 3810 34756 3852 34796
rect 3892 34756 3934 34796
rect 3974 34756 4016 34796
rect 4056 34756 18808 34796
rect 18848 34756 18890 34796
rect 18930 34756 18972 34796
rect 19012 34756 19054 34796
rect 19094 34756 19136 34796
rect 19176 34756 20352 34796
rect 1152 34732 20352 34756
rect 7467 34628 7509 34637
rect 7467 34588 7468 34628
rect 7508 34588 7509 34628
rect 7467 34579 7509 34588
rect 7947 34628 7989 34637
rect 7947 34588 7948 34628
rect 7988 34588 7989 34628
rect 7947 34579 7989 34588
rect 13419 34628 13461 34637
rect 13419 34588 13420 34628
rect 13460 34588 13461 34628
rect 13419 34579 13461 34588
rect 19563 34628 19605 34637
rect 19563 34588 19564 34628
rect 19604 34588 19605 34628
rect 19563 34579 19605 34588
rect 13219 34544 13277 34545
rect 13219 34504 13228 34544
rect 13268 34504 13277 34544
rect 13219 34503 13277 34504
rect 14187 34544 14229 34553
rect 14187 34504 14188 34544
rect 14228 34504 14229 34544
rect 14187 34495 14229 34504
rect 2667 34460 2709 34469
rect 2667 34420 2668 34460
rect 2708 34420 2709 34460
rect 2667 34411 2709 34420
rect 6027 34460 6069 34469
rect 6027 34420 6028 34460
rect 6068 34420 6069 34460
rect 6027 34411 6069 34420
rect 11115 34460 11157 34469
rect 11115 34420 11116 34460
rect 11156 34420 11157 34460
rect 11115 34411 11157 34420
rect 19363 34460 19421 34461
rect 19363 34420 19372 34460
rect 19412 34420 19421 34460
rect 19363 34419 19421 34420
rect 2187 34376 2229 34385
rect 2187 34336 2188 34376
rect 2228 34336 2229 34376
rect 2187 34327 2229 34336
rect 2283 34376 2325 34385
rect 2283 34336 2284 34376
rect 2324 34336 2325 34376
rect 2283 34327 2325 34336
rect 2763 34376 2805 34385
rect 3723 34381 3765 34390
rect 2763 34336 2764 34376
rect 2804 34336 2805 34376
rect 2763 34327 2805 34336
rect 3235 34376 3293 34377
rect 3235 34336 3244 34376
rect 3284 34336 3293 34376
rect 3235 34335 3293 34336
rect 3723 34341 3724 34381
rect 3764 34341 3765 34381
rect 3723 34332 3765 34341
rect 4107 34376 4149 34385
rect 4107 34336 4108 34376
rect 4148 34336 4149 34376
rect 4107 34327 4149 34336
rect 4203 34376 4245 34385
rect 4203 34336 4204 34376
rect 4244 34336 4245 34376
rect 4203 34327 4245 34336
rect 5067 34376 5109 34385
rect 5067 34336 5068 34376
rect 5108 34336 5109 34376
rect 5067 34327 5109 34336
rect 5163 34376 5205 34385
rect 5163 34336 5164 34376
rect 5204 34336 5205 34376
rect 5163 34327 5205 34336
rect 5259 34376 5301 34385
rect 5259 34336 5260 34376
rect 5300 34336 5301 34376
rect 5259 34327 5301 34336
rect 5547 34376 5589 34385
rect 5547 34336 5548 34376
rect 5588 34336 5589 34376
rect 5547 34327 5589 34336
rect 5643 34376 5685 34385
rect 5643 34336 5644 34376
rect 5684 34336 5685 34376
rect 5643 34327 5685 34336
rect 6123 34376 6165 34385
rect 7083 34381 7125 34390
rect 6123 34336 6124 34376
rect 6164 34336 6165 34376
rect 6123 34327 6165 34336
rect 6595 34376 6653 34377
rect 6595 34336 6604 34376
rect 6644 34336 6653 34376
rect 6595 34335 6653 34336
rect 7083 34341 7084 34381
rect 7124 34341 7125 34381
rect 7083 34332 7125 34341
rect 7467 34376 7509 34385
rect 7467 34336 7468 34376
rect 7508 34336 7509 34376
rect 7467 34327 7509 34336
rect 7755 34376 7797 34385
rect 7755 34336 7756 34376
rect 7796 34336 7797 34376
rect 7755 34327 7797 34336
rect 7947 34376 7989 34385
rect 7947 34336 7948 34376
rect 7988 34336 7989 34376
rect 7947 34327 7989 34336
rect 8139 34376 8181 34385
rect 8139 34336 8140 34376
rect 8180 34336 8181 34376
rect 8139 34327 8181 34336
rect 8427 34376 8469 34385
rect 8427 34336 8428 34376
rect 8468 34336 8469 34376
rect 8427 34327 8469 34336
rect 8523 34376 8565 34385
rect 8523 34336 8524 34376
rect 8564 34336 8565 34376
rect 8523 34327 8565 34336
rect 8907 34376 8949 34385
rect 8907 34336 8908 34376
rect 8948 34336 8949 34376
rect 8907 34327 8949 34336
rect 9003 34376 9045 34385
rect 9963 34381 10005 34390
rect 9003 34336 9004 34376
rect 9044 34336 9045 34376
rect 9003 34327 9045 34336
rect 9475 34376 9533 34377
rect 9475 34336 9484 34376
rect 9524 34336 9533 34376
rect 9475 34335 9533 34336
rect 9963 34341 9964 34381
rect 10004 34341 10005 34381
rect 9963 34332 10005 34341
rect 10539 34376 10581 34385
rect 10539 34336 10540 34376
rect 10580 34336 10581 34376
rect 10539 34327 10581 34336
rect 10635 34376 10677 34385
rect 10635 34336 10636 34376
rect 10676 34336 10677 34376
rect 10635 34327 10677 34336
rect 11019 34376 11061 34385
rect 12075 34381 12117 34390
rect 11019 34336 11020 34376
rect 11060 34336 11061 34376
rect 11019 34327 11061 34336
rect 11587 34376 11645 34377
rect 11587 34336 11596 34376
rect 11636 34336 11645 34376
rect 11587 34335 11645 34336
rect 12075 34341 12076 34381
rect 12116 34341 12117 34381
rect 12075 34332 12117 34341
rect 12547 34376 12605 34377
rect 12547 34336 12556 34376
rect 12596 34336 12605 34376
rect 12547 34335 12605 34336
rect 12843 34376 12885 34385
rect 12843 34336 12844 34376
rect 12884 34336 12885 34376
rect 12843 34327 12885 34336
rect 12939 34376 12981 34385
rect 12939 34336 12940 34376
rect 12980 34336 12981 34376
rect 12939 34327 12981 34336
rect 13411 34376 13469 34377
rect 13411 34336 13420 34376
rect 13460 34336 13469 34376
rect 13411 34335 13469 34336
rect 13507 34376 13565 34377
rect 13507 34336 13516 34376
rect 13556 34336 13565 34376
rect 13507 34335 13565 34336
rect 13707 34376 13749 34385
rect 13707 34336 13708 34376
rect 13748 34336 13749 34376
rect 13707 34327 13749 34336
rect 13803 34376 13845 34385
rect 13803 34336 13804 34376
rect 13844 34336 13845 34376
rect 13803 34327 13845 34336
rect 13950 34376 14008 34377
rect 13950 34336 13959 34376
rect 13999 34336 14008 34376
rect 13950 34335 14008 34336
rect 14187 34376 14229 34385
rect 14187 34336 14188 34376
rect 14228 34336 14229 34376
rect 14187 34327 14229 34336
rect 14379 34373 14421 34382
rect 14379 34333 14380 34373
rect 14420 34333 14421 34373
rect 14755 34376 14813 34377
rect 14755 34336 14764 34376
rect 14804 34336 14813 34376
rect 14755 34335 14813 34336
rect 16003 34376 16061 34377
rect 16003 34336 16012 34376
rect 16052 34336 16061 34376
rect 16003 34335 16061 34336
rect 19747 34376 19805 34377
rect 19747 34336 19756 34376
rect 19796 34336 19805 34376
rect 19747 34335 19805 34336
rect 14379 34324 14421 34333
rect 3915 34292 3957 34301
rect 3915 34252 3916 34292
rect 3956 34252 3957 34292
rect 3915 34243 3957 34252
rect 7275 34292 7317 34301
rect 7275 34252 7276 34292
rect 7316 34252 7317 34292
rect 7275 34243 7317 34252
rect 4387 34208 4445 34209
rect 4387 34168 4396 34208
rect 4436 34168 4445 34208
rect 4387 34167 4445 34168
rect 4963 34208 5021 34209
rect 4963 34168 4972 34208
rect 5012 34168 5021 34208
rect 4963 34167 5021 34168
rect 10155 34208 10197 34217
rect 10155 34168 10156 34208
rect 10196 34168 10197 34208
rect 10155 34159 10197 34168
rect 12267 34208 12309 34217
rect 12267 34168 12268 34208
rect 12308 34168 12309 34208
rect 12267 34159 12309 34168
rect 14571 34208 14613 34217
rect 14571 34168 14572 34208
rect 14612 34168 14613 34208
rect 14571 34159 14613 34168
rect 19851 34208 19893 34217
rect 19851 34168 19852 34208
rect 19892 34168 19893 34208
rect 19851 34159 19893 34168
rect 1152 34040 20452 34064
rect 1152 34000 4928 34040
rect 4968 34000 5010 34040
rect 5050 34000 5092 34040
rect 5132 34000 5174 34040
rect 5214 34000 5256 34040
rect 5296 34000 20048 34040
rect 20088 34000 20130 34040
rect 20170 34000 20212 34040
rect 20252 34000 20294 34040
rect 20334 34000 20376 34040
rect 20416 34000 20452 34040
rect 1152 33976 20452 34000
rect 3147 33872 3189 33881
rect 3147 33832 3148 33872
rect 3188 33832 3189 33872
rect 3147 33823 3189 33832
rect 6211 33872 6269 33873
rect 6211 33832 6220 33872
rect 6260 33832 6269 33872
rect 6211 33831 6269 33832
rect 7747 33872 7805 33873
rect 7747 33832 7756 33872
rect 7796 33832 7805 33872
rect 7747 33831 7805 33832
rect 9771 33872 9813 33881
rect 9771 33832 9772 33872
rect 9812 33832 9813 33872
rect 9771 33823 9813 33832
rect 11403 33872 11445 33881
rect 11403 33832 11404 33872
rect 11444 33832 11445 33872
rect 11403 33823 11445 33832
rect 11683 33872 11741 33873
rect 11683 33832 11692 33872
rect 11732 33832 11741 33872
rect 11683 33831 11741 33832
rect 12459 33872 12501 33881
rect 12459 33832 12460 33872
rect 12500 33832 12501 33872
rect 12459 33823 12501 33832
rect 12747 33872 12789 33881
rect 12747 33832 12748 33872
rect 12788 33832 12789 33872
rect 12747 33823 12789 33832
rect 14283 33872 14325 33881
rect 14283 33832 14284 33872
rect 14324 33832 14325 33872
rect 14283 33823 14325 33832
rect 14667 33872 14709 33881
rect 14667 33832 14668 33872
rect 14708 33832 14709 33872
rect 14667 33823 14709 33832
rect 5643 33788 5685 33797
rect 5643 33748 5644 33788
rect 5684 33748 5685 33788
rect 5643 33739 5685 33748
rect 6987 33788 7029 33797
rect 6987 33748 6988 33788
rect 7028 33748 7029 33788
rect 6987 33739 7029 33748
rect 1699 33704 1757 33705
rect 1699 33664 1708 33704
rect 1748 33664 1757 33704
rect 1699 33663 1757 33664
rect 2947 33704 3005 33705
rect 2947 33664 2956 33704
rect 2996 33664 3005 33704
rect 2947 33663 3005 33664
rect 3531 33704 3573 33713
rect 3531 33664 3532 33704
rect 3572 33664 3573 33704
rect 3531 33655 3573 33664
rect 3819 33704 3861 33713
rect 3819 33664 3820 33704
rect 3860 33664 3861 33704
rect 3819 33655 3861 33664
rect 4195 33704 4253 33705
rect 4195 33664 4204 33704
rect 4244 33664 4253 33704
rect 4195 33663 4253 33664
rect 5443 33704 5501 33705
rect 5443 33664 5452 33704
rect 5492 33664 5501 33704
rect 5443 33663 5501 33664
rect 6019 33704 6077 33705
rect 6019 33664 6028 33704
rect 6068 33664 6077 33704
rect 6019 33663 6077 33664
rect 6123 33704 6165 33713
rect 6123 33664 6124 33704
rect 6164 33664 6165 33704
rect 6123 33655 6165 33664
rect 6315 33704 6357 33713
rect 6315 33664 6316 33704
rect 6356 33664 6357 33704
rect 6315 33655 6357 33664
rect 6595 33704 6653 33705
rect 6595 33664 6604 33704
rect 6644 33664 6653 33704
rect 6595 33663 6653 33664
rect 6891 33704 6933 33713
rect 6891 33664 6892 33704
rect 6932 33664 6933 33704
rect 6891 33655 6933 33664
rect 7467 33704 7509 33713
rect 7467 33664 7468 33704
rect 7508 33664 7509 33704
rect 7467 33655 7509 33664
rect 7563 33704 7605 33713
rect 7563 33664 7564 33704
rect 7604 33664 7605 33704
rect 7563 33655 7605 33664
rect 8323 33704 8381 33705
rect 8323 33664 8332 33704
rect 8372 33664 8381 33704
rect 8323 33663 8381 33664
rect 9571 33704 9629 33705
rect 9571 33664 9580 33704
rect 9620 33664 9629 33704
rect 9571 33663 9629 33664
rect 9955 33704 10013 33705
rect 9955 33664 9964 33704
rect 10004 33664 10013 33704
rect 9955 33663 10013 33664
rect 11203 33704 11261 33705
rect 11203 33664 11212 33704
rect 11252 33664 11261 33704
rect 11203 33663 11261 33664
rect 11595 33704 11637 33713
rect 11595 33664 11596 33704
rect 11636 33664 11637 33704
rect 11595 33655 11637 33664
rect 11787 33704 11829 33713
rect 11787 33664 11788 33704
rect 11828 33664 11829 33704
rect 11787 33655 11829 33664
rect 11875 33704 11933 33705
rect 11875 33664 11884 33704
rect 11924 33664 11933 33704
rect 11875 33663 11933 33664
rect 12355 33704 12413 33705
rect 12355 33664 12364 33704
rect 12404 33664 12413 33704
rect 12355 33663 12413 33664
rect 12651 33704 12693 33713
rect 12651 33664 12652 33704
rect 12692 33664 12693 33704
rect 12651 33655 12693 33664
rect 12843 33704 12885 33713
rect 12843 33664 12844 33704
rect 12884 33664 12885 33704
rect 12843 33655 12885 33664
rect 12939 33704 12981 33713
rect 12939 33664 12940 33704
rect 12980 33664 12981 33704
rect 12939 33655 12981 33664
rect 13123 33704 13181 33705
rect 13123 33664 13132 33704
rect 13172 33664 13181 33704
rect 13123 33663 13181 33664
rect 13515 33704 13557 33713
rect 13515 33664 13516 33704
rect 13556 33664 13557 33704
rect 13515 33655 13557 33664
rect 13707 33704 13749 33713
rect 13707 33664 13708 33704
rect 13748 33664 13749 33704
rect 13707 33655 13749 33664
rect 13899 33704 13941 33713
rect 13899 33664 13900 33704
rect 13940 33664 13941 33704
rect 13899 33655 13941 33664
rect 13995 33704 14037 33713
rect 13995 33664 13996 33704
rect 14036 33664 14037 33704
rect 13995 33655 14037 33664
rect 14187 33704 14229 33713
rect 14187 33664 14188 33704
rect 14228 33664 14229 33704
rect 14187 33655 14229 33664
rect 14475 33704 14517 33713
rect 14475 33664 14476 33704
rect 14516 33664 14517 33704
rect 14475 33655 14517 33664
rect 14851 33704 14909 33705
rect 14851 33664 14860 33704
rect 14900 33664 14909 33704
rect 14851 33663 14909 33664
rect 16099 33704 16157 33705
rect 16099 33664 16108 33704
rect 16148 33664 16157 33704
rect 16099 33663 16157 33664
rect 13227 33620 13269 33629
rect 13227 33580 13228 33620
rect 13268 33580 13269 33620
rect 13227 33571 13269 33580
rect 13419 33620 13461 33629
rect 13419 33580 13420 33620
rect 13460 33580 13461 33620
rect 13419 33571 13461 33580
rect 13323 33536 13365 33545
rect 13323 33496 13324 33536
rect 13364 33496 13365 33536
rect 13323 33487 13365 33496
rect 13987 33536 14045 33537
rect 13987 33496 13996 33536
rect 14036 33496 14045 33536
rect 13987 33495 14045 33496
rect 3531 33452 3573 33461
rect 3531 33412 3532 33452
rect 3572 33412 3573 33452
rect 3531 33403 3573 33412
rect 7267 33452 7325 33453
rect 7267 33412 7276 33452
rect 7316 33412 7325 33452
rect 7267 33411 7325 33412
rect 1152 33284 20352 33308
rect 1152 33244 3688 33284
rect 3728 33244 3770 33284
rect 3810 33244 3852 33284
rect 3892 33244 3934 33284
rect 3974 33244 4016 33284
rect 4056 33244 18808 33284
rect 18848 33244 18890 33284
rect 18930 33244 18972 33284
rect 19012 33244 19054 33284
rect 19094 33244 19136 33284
rect 19176 33244 20352 33284
rect 1152 33220 20352 33244
rect 13707 33116 13749 33125
rect 13707 33076 13708 33116
rect 13748 33076 13749 33116
rect 13707 33067 13749 33076
rect 7939 33032 7997 33033
rect 7939 32992 7948 33032
rect 7988 32992 7997 33032
rect 7939 32991 7997 32992
rect 13411 33032 13469 33033
rect 13411 32992 13420 33032
rect 13460 32992 13469 33032
rect 13411 32991 13469 32992
rect 3147 32948 3189 32957
rect 3147 32908 3148 32948
rect 3188 32908 3189 32948
rect 3147 32899 3189 32908
rect 8427 32948 8469 32957
rect 8427 32908 8428 32948
rect 8468 32908 8469 32948
rect 8427 32899 8469 32908
rect 2763 32864 2805 32873
rect 2667 32844 2709 32853
rect 2667 32804 2668 32844
rect 2708 32804 2709 32844
rect 2763 32824 2764 32864
rect 2804 32824 2805 32864
rect 2763 32815 2805 32824
rect 3243 32864 3285 32873
rect 4203 32869 4245 32878
rect 3243 32824 3244 32864
rect 3284 32824 3285 32864
rect 3243 32815 3285 32824
rect 3715 32864 3773 32865
rect 3715 32824 3724 32864
rect 3764 32824 3773 32864
rect 3715 32823 3773 32824
rect 4203 32829 4204 32869
rect 4244 32829 4245 32869
rect 4203 32820 4245 32829
rect 6115 32864 6173 32865
rect 6115 32824 6124 32864
rect 6164 32824 6173 32864
rect 6115 32823 6173 32824
rect 7363 32864 7421 32865
rect 7363 32824 7372 32864
rect 7412 32824 7421 32864
rect 7363 32823 7421 32824
rect 7755 32864 7797 32873
rect 7755 32824 7756 32864
rect 7796 32824 7797 32864
rect 7755 32815 7797 32824
rect 7947 32860 7989 32869
rect 7947 32820 7948 32860
rect 7988 32820 7989 32860
rect 7947 32811 7989 32820
rect 8043 32864 8085 32873
rect 8043 32824 8044 32864
rect 8084 32824 8085 32864
rect 8043 32815 8085 32824
rect 8235 32857 8277 32866
rect 8235 32817 8236 32857
rect 8276 32817 8277 32857
rect 8235 32808 8277 32817
rect 8523 32864 8565 32873
rect 8523 32824 8524 32864
rect 8564 32824 8565 32864
rect 8523 32815 8565 32824
rect 12267 32864 12309 32873
rect 12267 32824 12268 32864
rect 12308 32824 12309 32864
rect 12267 32815 12309 32824
rect 12451 32864 12509 32865
rect 12451 32824 12460 32864
rect 12500 32824 12509 32864
rect 12451 32823 12509 32824
rect 13227 32864 13269 32873
rect 13227 32824 13228 32864
rect 13268 32824 13269 32864
rect 13227 32815 13269 32824
rect 13419 32864 13461 32873
rect 13419 32824 13420 32864
rect 13460 32824 13461 32864
rect 13419 32815 13461 32824
rect 13515 32864 13557 32873
rect 13515 32824 13516 32864
rect 13556 32824 13557 32864
rect 13515 32815 13557 32824
rect 13795 32864 13853 32865
rect 13795 32824 13804 32864
rect 13844 32824 13853 32864
rect 13795 32823 13853 32824
rect 13987 32864 14045 32865
rect 13987 32824 13996 32864
rect 14036 32824 14045 32864
rect 13987 32823 14045 32824
rect 15235 32864 15293 32865
rect 15235 32824 15244 32864
rect 15284 32824 15293 32864
rect 15235 32823 15293 32824
rect 16195 32864 16253 32865
rect 16195 32824 16204 32864
rect 16244 32824 16253 32864
rect 16195 32823 16253 32824
rect 17443 32864 17501 32865
rect 17443 32824 17452 32864
rect 17492 32824 17501 32864
rect 17443 32823 17501 32824
rect 2667 32795 2709 32804
rect 4395 32780 4437 32789
rect 4395 32740 4396 32780
rect 4436 32740 4437 32780
rect 4395 32731 4437 32740
rect 12363 32780 12405 32789
rect 12363 32740 12364 32780
rect 12404 32740 12405 32780
rect 12363 32731 12405 32740
rect 7563 32696 7605 32705
rect 7563 32656 7564 32696
rect 7604 32656 7605 32696
rect 7563 32647 7605 32656
rect 15435 32696 15477 32705
rect 15435 32656 15436 32696
rect 15476 32656 15477 32696
rect 15435 32647 15477 32656
rect 17643 32696 17685 32705
rect 17643 32656 17644 32696
rect 17684 32656 17685 32696
rect 17643 32647 17685 32656
rect 1152 32528 20452 32552
rect 1152 32488 4928 32528
rect 4968 32488 5010 32528
rect 5050 32488 5092 32528
rect 5132 32488 5174 32528
rect 5214 32488 5256 32528
rect 5296 32488 20048 32528
rect 20088 32488 20130 32528
rect 20170 32488 20212 32528
rect 20252 32488 20294 32528
rect 20334 32488 20376 32528
rect 20416 32488 20452 32528
rect 1152 32464 20452 32488
rect 3915 32360 3957 32369
rect 3915 32320 3916 32360
rect 3956 32320 3957 32360
rect 3915 32311 3957 32320
rect 5547 32360 5589 32369
rect 5547 32320 5548 32360
rect 5588 32320 5589 32360
rect 5547 32311 5589 32320
rect 10723 32360 10781 32361
rect 10723 32320 10732 32360
rect 10772 32320 10781 32360
rect 10723 32319 10781 32320
rect 11211 32360 11253 32369
rect 11211 32320 11212 32360
rect 11252 32320 11253 32360
rect 11211 32311 11253 32320
rect 13707 32360 13749 32369
rect 13707 32320 13708 32360
rect 13748 32320 13749 32360
rect 13707 32311 13749 32320
rect 7563 32276 7605 32285
rect 7563 32236 7564 32276
rect 7604 32236 7605 32276
rect 7563 32227 7605 32236
rect 8427 32276 8469 32285
rect 8427 32236 8428 32276
rect 8468 32236 8469 32276
rect 8427 32227 8469 32236
rect 5931 32212 5973 32221
rect 2467 32192 2525 32193
rect 2467 32152 2476 32192
rect 2516 32152 2525 32192
rect 2467 32151 2525 32152
rect 3715 32192 3773 32193
rect 3715 32152 3724 32192
rect 3764 32152 3773 32192
rect 3715 32151 3773 32152
rect 4099 32192 4157 32193
rect 4099 32152 4108 32192
rect 4148 32152 4157 32192
rect 4099 32151 4157 32152
rect 5347 32192 5405 32193
rect 5347 32152 5356 32192
rect 5396 32152 5405 32192
rect 5347 32151 5405 32152
rect 5835 32192 5877 32201
rect 5835 32152 5836 32192
rect 5876 32152 5877 32192
rect 5931 32172 5932 32212
rect 5972 32172 5973 32212
rect 5931 32163 5973 32172
rect 6883 32192 6941 32193
rect 5835 32143 5877 32152
rect 6883 32152 6892 32192
rect 6932 32152 6941 32192
rect 8035 32192 8093 32193
rect 6883 32151 6941 32152
rect 7371 32178 7413 32187
rect 7371 32138 7372 32178
rect 7412 32138 7413 32178
rect 8035 32152 8044 32192
rect 8084 32152 8093 32192
rect 8035 32151 8093 32152
rect 8331 32192 8373 32201
rect 8331 32152 8332 32192
rect 8372 32152 8373 32192
rect 8331 32143 8373 32152
rect 9283 32192 9341 32193
rect 9283 32152 9292 32192
rect 9332 32152 9341 32192
rect 9283 32151 9341 32152
rect 10531 32192 10589 32193
rect 10531 32152 10540 32192
rect 10580 32152 10589 32192
rect 10531 32151 10589 32152
rect 10923 32192 10965 32201
rect 10923 32152 10924 32192
rect 10964 32152 10965 32192
rect 10923 32143 10965 32152
rect 11019 32192 11061 32201
rect 11019 32152 11020 32192
rect 11060 32152 11061 32192
rect 11019 32143 11061 32152
rect 11395 32192 11453 32193
rect 11395 32152 11404 32192
rect 11444 32152 11453 32192
rect 11395 32151 11453 32152
rect 12643 32192 12701 32193
rect 12643 32152 12652 32192
rect 12692 32152 12701 32192
rect 12643 32151 12701 32152
rect 12835 32192 12893 32193
rect 12835 32152 12844 32192
rect 12884 32152 12893 32192
rect 12835 32151 12893 32152
rect 12939 32192 12981 32201
rect 12939 32152 12940 32192
rect 12980 32152 12981 32192
rect 12939 32143 12981 32152
rect 13123 32192 13181 32193
rect 13123 32152 13132 32192
rect 13172 32152 13181 32192
rect 13123 32151 13181 32152
rect 13795 32192 13853 32193
rect 13795 32152 13804 32192
rect 13844 32152 13853 32192
rect 13795 32151 13853 32152
rect 14371 32192 14429 32193
rect 14371 32152 14380 32192
rect 14420 32152 14429 32192
rect 14371 32151 14429 32152
rect 14475 32192 14517 32201
rect 14475 32152 14476 32192
rect 14516 32152 14517 32192
rect 14475 32143 14517 32152
rect 14667 32192 14709 32201
rect 14667 32152 14668 32192
rect 14708 32152 14709 32192
rect 14667 32143 14709 32152
rect 14859 32192 14901 32201
rect 14859 32152 14860 32192
rect 14900 32152 14901 32192
rect 14859 32143 14901 32152
rect 15147 32192 15189 32201
rect 15147 32152 15148 32192
rect 15188 32152 15189 32192
rect 15147 32143 15189 32152
rect 15331 32192 15389 32193
rect 15331 32152 15340 32192
rect 15380 32152 15389 32192
rect 15331 32151 15389 32152
rect 16579 32192 16637 32193
rect 16579 32152 16588 32192
rect 16628 32152 16637 32192
rect 16579 32151 16637 32152
rect 7371 32129 7413 32138
rect 6315 32108 6357 32117
rect 6315 32068 6316 32108
rect 6356 32068 6357 32108
rect 6315 32059 6357 32068
rect 6411 32108 6453 32117
rect 6411 32068 6412 32108
rect 6452 32068 6453 32108
rect 6411 32059 6453 32068
rect 14955 32108 14997 32117
rect 14955 32068 14956 32108
rect 14996 32068 14997 32108
rect 14955 32059 14997 32068
rect 14667 32024 14709 32033
rect 14667 31984 14668 32024
rect 14708 31984 14709 32024
rect 14667 31975 14709 31984
rect 8707 31940 8765 31941
rect 8707 31900 8716 31940
rect 8756 31900 8765 31940
rect 8707 31899 8765 31900
rect 9099 31940 9141 31949
rect 9099 31900 9100 31940
rect 9140 31900 9141 31940
rect 9099 31891 9141 31900
rect 11211 31940 11253 31949
rect 11211 31900 11212 31940
rect 11252 31900 11253 31940
rect 11211 31891 11253 31900
rect 12939 31940 12981 31949
rect 12939 31900 12940 31940
rect 12980 31900 12981 31940
rect 12939 31891 12981 31900
rect 16779 31940 16821 31949
rect 16779 31900 16780 31940
rect 16820 31900 16821 31940
rect 16779 31891 16821 31900
rect 1152 31772 20352 31796
rect 1152 31732 3688 31772
rect 3728 31732 3770 31772
rect 3810 31732 3852 31772
rect 3892 31732 3934 31772
rect 3974 31732 4016 31772
rect 4056 31732 18808 31772
rect 18848 31732 18890 31772
rect 18930 31732 18972 31772
rect 19012 31732 19054 31772
rect 19094 31732 19136 31772
rect 19176 31732 20352 31772
rect 1152 31708 20352 31732
rect 8331 31604 8373 31613
rect 8331 31564 8332 31604
rect 8372 31564 8373 31604
rect 8331 31555 8373 31564
rect 10827 31604 10869 31613
rect 10827 31564 10828 31604
rect 10868 31564 10869 31604
rect 10827 31555 10869 31564
rect 12939 31604 12981 31613
rect 12939 31564 12940 31604
rect 12980 31564 12981 31604
rect 12939 31555 12981 31564
rect 2667 31520 2709 31529
rect 2667 31480 2668 31520
rect 2708 31480 2709 31520
rect 2667 31471 2709 31480
rect 6699 31520 6741 31529
rect 6699 31480 6700 31520
rect 6740 31480 6741 31520
rect 6699 31471 6741 31480
rect 14955 31520 14997 31529
rect 14955 31480 14956 31520
rect 14996 31480 14997 31520
rect 14955 31471 14997 31480
rect 15627 31520 15669 31529
rect 15627 31480 15628 31520
rect 15668 31480 15669 31520
rect 15627 31471 15669 31480
rect 5067 31436 5109 31445
rect 5067 31396 5068 31436
rect 5108 31396 5109 31436
rect 5067 31387 5109 31396
rect 17643 31366 17685 31375
rect 3720 31362 3778 31363
rect 1219 31352 1277 31353
rect 1219 31312 1228 31352
rect 1268 31312 1277 31352
rect 1219 31311 1277 31312
rect 2467 31352 2525 31353
rect 2467 31312 2476 31352
rect 2516 31312 2525 31352
rect 2467 31311 2525 31312
rect 2851 31352 2909 31353
rect 2851 31312 2860 31352
rect 2900 31312 2909 31352
rect 2851 31311 2909 31312
rect 2947 31352 3005 31353
rect 2947 31312 2956 31352
rect 2996 31312 3005 31352
rect 2947 31311 3005 31312
rect 3147 31352 3189 31361
rect 3147 31312 3148 31352
rect 3188 31312 3189 31352
rect 3147 31303 3189 31312
rect 3243 31352 3285 31361
rect 3243 31312 3244 31352
rect 3284 31312 3285 31352
rect 3243 31303 3285 31312
rect 3336 31352 3394 31353
rect 3336 31312 3345 31352
rect 3385 31312 3394 31352
rect 3336 31311 3394 31312
rect 3627 31352 3669 31361
rect 3627 31312 3628 31352
rect 3668 31312 3669 31352
rect 3720 31322 3729 31362
rect 3769 31322 3778 31362
rect 3720 31321 3778 31322
rect 4491 31352 4533 31361
rect 3627 31303 3669 31312
rect 4491 31312 4492 31352
rect 4532 31312 4533 31352
rect 4491 31303 4533 31312
rect 4587 31352 4629 31361
rect 4587 31312 4588 31352
rect 4628 31312 4629 31352
rect 4587 31303 4629 31312
rect 4971 31352 5013 31361
rect 6027 31357 6069 31366
rect 4971 31312 4972 31352
rect 5012 31312 5013 31352
rect 4971 31303 5013 31312
rect 5539 31352 5597 31353
rect 5539 31312 5548 31352
rect 5588 31312 5597 31352
rect 5539 31311 5597 31312
rect 6027 31317 6028 31357
rect 6068 31317 6069 31357
rect 6027 31308 6069 31317
rect 6507 31352 6549 31361
rect 6507 31312 6508 31352
rect 6548 31312 6549 31352
rect 6507 31303 6549 31312
rect 6699 31352 6741 31361
rect 6699 31312 6700 31352
rect 6740 31312 6741 31352
rect 6699 31303 6741 31312
rect 6883 31352 6941 31353
rect 6883 31312 6892 31352
rect 6932 31312 6941 31352
rect 6883 31311 6941 31312
rect 8131 31352 8189 31353
rect 8131 31312 8140 31352
rect 8180 31312 8189 31352
rect 8131 31311 8189 31312
rect 9091 31352 9149 31353
rect 9091 31312 9100 31352
rect 9140 31312 9149 31352
rect 9091 31311 9149 31312
rect 9379 31352 9437 31353
rect 9379 31312 9388 31352
rect 9428 31312 9437 31352
rect 9379 31311 9437 31312
rect 10627 31352 10685 31353
rect 10627 31312 10636 31352
rect 10676 31312 10685 31352
rect 10627 31311 10685 31312
rect 11211 31352 11253 31361
rect 11211 31312 11212 31352
rect 11252 31312 11253 31352
rect 11211 31303 11253 31312
rect 11307 31352 11349 31361
rect 11307 31312 11308 31352
rect 11348 31312 11349 31352
rect 11307 31303 11349 31312
rect 11491 31352 11549 31353
rect 11491 31312 11500 31352
rect 11540 31312 11549 31352
rect 11491 31311 11549 31312
rect 12739 31352 12797 31353
rect 12739 31312 12748 31352
rect 12788 31312 12797 31352
rect 12739 31311 12797 31312
rect 13131 31352 13173 31361
rect 13131 31312 13132 31352
rect 13172 31312 13173 31352
rect 13131 31303 13173 31312
rect 13323 31352 13365 31361
rect 13323 31312 13324 31352
rect 13364 31312 13365 31352
rect 13323 31303 13365 31312
rect 13507 31352 13565 31353
rect 13507 31312 13516 31352
rect 13556 31312 13565 31352
rect 13507 31311 13565 31312
rect 14755 31352 14813 31353
rect 14755 31312 14764 31352
rect 14804 31312 14813 31352
rect 14755 31311 14813 31312
rect 15139 31352 15197 31353
rect 15139 31312 15148 31352
rect 15188 31312 15197 31352
rect 15139 31311 15197 31312
rect 15243 31352 15285 31361
rect 15243 31312 15244 31352
rect 15284 31312 15285 31352
rect 15243 31303 15285 31312
rect 15435 31352 15477 31361
rect 15435 31312 15436 31352
rect 15476 31312 15477 31352
rect 15435 31303 15477 31312
rect 15627 31352 15669 31361
rect 15627 31312 15628 31352
rect 15668 31312 15669 31352
rect 15627 31303 15669 31312
rect 15819 31352 15861 31361
rect 15819 31312 15820 31352
rect 15860 31312 15861 31352
rect 15819 31303 15861 31312
rect 16107 31352 16149 31361
rect 16107 31312 16108 31352
rect 16148 31312 16149 31352
rect 16587 31352 16629 31361
rect 16107 31303 16149 31312
rect 16203 31332 16245 31341
rect 16203 31292 16204 31332
rect 16244 31292 16245 31332
rect 16587 31312 16588 31352
rect 16628 31312 16629 31352
rect 16587 31303 16629 31312
rect 16683 31352 16725 31361
rect 16683 31312 16684 31352
rect 16724 31312 16725 31352
rect 16683 31303 16725 31312
rect 17155 31352 17213 31353
rect 17155 31312 17164 31352
rect 17204 31312 17213 31352
rect 17643 31326 17644 31366
rect 17684 31326 17685 31366
rect 17643 31317 17685 31326
rect 18211 31352 18269 31353
rect 17155 31311 17213 31312
rect 18211 31312 18220 31352
rect 18260 31312 18269 31352
rect 18211 31311 18269 31312
rect 19459 31352 19517 31353
rect 19459 31312 19468 31352
rect 19508 31312 19517 31352
rect 19459 31311 19517 31312
rect 19851 31352 19893 31361
rect 19851 31312 19852 31352
rect 19892 31312 19893 31352
rect 19851 31303 19893 31312
rect 20043 31352 20085 31361
rect 20043 31312 20044 31352
rect 20084 31312 20085 31352
rect 20043 31303 20085 31312
rect 16203 31283 16245 31292
rect 6219 31268 6261 31277
rect 6219 31228 6220 31268
rect 6260 31228 6261 31268
rect 6219 31219 6261 31228
rect 15339 31268 15381 31277
rect 15339 31228 15340 31268
rect 15380 31228 15381 31268
rect 15339 31219 15381 31228
rect 17835 31268 17877 31277
rect 17835 31228 17836 31268
rect 17876 31228 17877 31268
rect 17835 31219 17877 31228
rect 3043 31184 3101 31185
rect 3043 31144 3052 31184
rect 3092 31144 3101 31184
rect 3043 31143 3101 31144
rect 3907 31184 3965 31185
rect 3907 31144 3916 31184
rect 3956 31144 3965 31184
rect 3907 31143 3965 31144
rect 9195 31184 9237 31193
rect 9195 31144 9196 31184
rect 9236 31144 9237 31184
rect 9195 31135 9237 31144
rect 10827 31184 10869 31193
rect 10827 31144 10828 31184
rect 10868 31144 10869 31184
rect 10827 31135 10869 31144
rect 11011 31184 11069 31185
rect 11011 31144 11020 31184
rect 11060 31144 11069 31184
rect 11011 31143 11069 31144
rect 13227 31184 13269 31193
rect 13227 31144 13228 31184
rect 13268 31144 13269 31184
rect 13227 31135 13269 31144
rect 19659 31184 19701 31193
rect 19659 31144 19660 31184
rect 19700 31144 19701 31184
rect 19659 31135 19701 31144
rect 19947 31184 19989 31193
rect 19947 31144 19948 31184
rect 19988 31144 19989 31184
rect 19947 31135 19989 31144
rect 1152 31016 20452 31040
rect 1152 30976 4928 31016
rect 4968 30976 5010 31016
rect 5050 30976 5092 31016
rect 5132 30976 5174 31016
rect 5214 30976 5256 31016
rect 5296 30976 20048 31016
rect 20088 30976 20130 31016
rect 20170 30976 20212 31016
rect 20252 30976 20294 31016
rect 20334 30976 20376 31016
rect 20416 30976 20452 31016
rect 1152 30952 20452 30976
rect 1707 30848 1749 30857
rect 1707 30808 1708 30848
rect 1748 30808 1749 30848
rect 1707 30799 1749 30808
rect 1995 30848 2037 30857
rect 1995 30808 1996 30848
rect 2036 30808 2037 30848
rect 1995 30799 2037 30808
rect 3819 30848 3861 30857
rect 3819 30808 3820 30848
rect 3860 30808 3861 30848
rect 3819 30799 3861 30808
rect 13219 30848 13277 30849
rect 13219 30808 13228 30848
rect 13268 30808 13277 30848
rect 13219 30807 13277 30808
rect 15435 30848 15477 30857
rect 15435 30808 15436 30848
rect 15476 30808 15477 30848
rect 15435 30799 15477 30808
rect 15907 30848 15965 30849
rect 15907 30808 15916 30848
rect 15956 30808 15965 30848
rect 15907 30807 15965 30808
rect 19747 30848 19805 30849
rect 19747 30808 19756 30848
rect 19796 30808 19805 30848
rect 19747 30807 19805 30808
rect 5835 30764 5877 30773
rect 5835 30724 5836 30764
rect 5876 30724 5877 30764
rect 5835 30715 5877 30724
rect 8523 30764 8565 30773
rect 8523 30724 8524 30764
rect 8564 30724 8565 30764
rect 8523 30715 8565 30724
rect 10539 30764 10581 30773
rect 10539 30724 10540 30764
rect 10580 30724 10581 30764
rect 10539 30715 10581 30724
rect 11211 30764 11253 30773
rect 11211 30724 11212 30764
rect 11252 30724 11253 30764
rect 11211 30715 11253 30724
rect 12459 30764 12501 30773
rect 12459 30724 12460 30764
rect 12500 30724 12501 30764
rect 12459 30715 12501 30724
rect 18795 30764 18837 30773
rect 18795 30724 18796 30764
rect 18836 30724 18837 30764
rect 18795 30715 18837 30724
rect 1603 30680 1661 30681
rect 1603 30640 1612 30680
rect 1652 30640 1661 30680
rect 1603 30639 1661 30640
rect 1899 30680 1941 30689
rect 1899 30640 1900 30680
rect 1940 30640 1941 30680
rect 1899 30631 1941 30640
rect 2091 30680 2133 30689
rect 2091 30640 2092 30680
rect 2132 30640 2133 30680
rect 2091 30631 2133 30640
rect 2187 30680 2229 30689
rect 2187 30640 2188 30680
rect 2228 30640 2229 30680
rect 2187 30631 2229 30640
rect 2371 30680 2429 30681
rect 2371 30640 2380 30680
rect 2420 30640 2429 30680
rect 2371 30639 2429 30640
rect 3619 30680 3677 30681
rect 3619 30640 3628 30680
rect 3668 30640 3677 30680
rect 3619 30639 3677 30640
rect 4107 30680 4149 30689
rect 4107 30640 4108 30680
rect 4148 30640 4149 30680
rect 4107 30631 4149 30640
rect 4203 30680 4245 30689
rect 4203 30640 4204 30680
rect 4244 30640 4245 30680
rect 4203 30631 4245 30640
rect 4683 30680 4725 30689
rect 4683 30640 4684 30680
rect 4724 30640 4725 30680
rect 4683 30631 4725 30640
rect 5155 30680 5213 30681
rect 5155 30640 5164 30680
rect 5204 30640 5213 30680
rect 7075 30680 7133 30681
rect 5155 30639 5213 30640
rect 5643 30666 5685 30675
rect 5643 30626 5644 30666
rect 5684 30626 5685 30666
rect 7075 30640 7084 30680
rect 7124 30640 7133 30680
rect 7075 30639 7133 30640
rect 8323 30680 8381 30681
rect 8323 30640 8332 30680
rect 8372 30640 8381 30680
rect 8323 30639 8381 30640
rect 8811 30680 8853 30689
rect 8811 30640 8812 30680
rect 8852 30640 8853 30680
rect 8811 30631 8853 30640
rect 8907 30680 8949 30689
rect 8907 30640 8908 30680
rect 8948 30640 8949 30680
rect 8907 30631 8949 30640
rect 9291 30680 9333 30689
rect 9291 30640 9292 30680
rect 9332 30640 9333 30680
rect 9859 30680 9917 30681
rect 9291 30631 9333 30640
rect 9387 30638 9429 30647
rect 9859 30640 9868 30680
rect 9908 30640 9917 30680
rect 10819 30680 10877 30681
rect 9859 30639 9917 30640
rect 10347 30666 10389 30675
rect 5643 30617 5685 30626
rect 4587 30596 4629 30605
rect 4587 30556 4588 30596
rect 4628 30556 4629 30596
rect 9387 30598 9388 30638
rect 9428 30598 9429 30638
rect 10347 30626 10348 30666
rect 10388 30626 10389 30666
rect 10819 30640 10828 30680
rect 10868 30640 10877 30680
rect 10819 30639 10877 30640
rect 11115 30680 11157 30689
rect 11115 30640 11116 30680
rect 11156 30640 11157 30680
rect 11115 30631 11157 30640
rect 12067 30680 12125 30681
rect 12067 30640 12076 30680
rect 12116 30640 12125 30680
rect 12067 30639 12125 30640
rect 12363 30680 12405 30689
rect 12363 30640 12364 30680
rect 12404 30640 12405 30680
rect 12363 30631 12405 30640
rect 12939 30680 12981 30689
rect 12939 30640 12940 30680
rect 12980 30640 12981 30680
rect 12939 30631 12981 30640
rect 13035 30680 13077 30689
rect 13035 30640 13036 30680
rect 13076 30640 13077 30680
rect 13035 30631 13077 30640
rect 13707 30680 13749 30689
rect 13707 30640 13708 30680
rect 13748 30640 13749 30680
rect 13707 30631 13749 30640
rect 13803 30680 13845 30689
rect 13803 30640 13804 30680
rect 13844 30640 13845 30680
rect 13803 30631 13845 30640
rect 14187 30680 14229 30689
rect 14187 30640 14188 30680
rect 14228 30640 14229 30680
rect 14187 30631 14229 30640
rect 14755 30680 14813 30681
rect 14755 30640 14764 30680
rect 14804 30640 14813 30680
rect 14755 30639 14813 30640
rect 15243 30675 15285 30684
rect 15243 30635 15244 30675
rect 15284 30635 15285 30675
rect 15723 30680 15765 30689
rect 15243 30626 15285 30635
rect 15627 30635 15669 30644
rect 10347 30617 10389 30626
rect 9387 30589 9429 30598
rect 14283 30596 14325 30605
rect 4587 30547 4629 30556
rect 14283 30556 14284 30596
rect 14324 30556 14325 30596
rect 15627 30595 15628 30635
rect 15668 30595 15669 30635
rect 15723 30640 15724 30680
rect 15764 30640 15765 30680
rect 15723 30631 15765 30640
rect 15819 30680 15861 30689
rect 15819 30640 15820 30680
rect 15860 30640 15861 30680
rect 15819 30631 15861 30640
rect 16483 30680 16541 30681
rect 16483 30640 16492 30680
rect 16532 30640 16541 30680
rect 16483 30639 16541 30640
rect 17731 30680 17789 30681
rect 17731 30640 17740 30680
rect 17780 30640 17789 30680
rect 17731 30639 17789 30640
rect 18403 30680 18461 30681
rect 18403 30640 18412 30680
rect 18452 30640 18461 30680
rect 18403 30639 18461 30640
rect 18699 30680 18741 30689
rect 18699 30640 18700 30680
rect 18740 30640 18741 30680
rect 18699 30631 18741 30640
rect 19275 30680 19317 30689
rect 19275 30640 19276 30680
rect 19316 30640 19317 30680
rect 19275 30631 19317 30640
rect 19467 30680 19509 30689
rect 19467 30640 19468 30680
rect 19508 30640 19509 30680
rect 19467 30631 19509 30640
rect 19555 30680 19613 30681
rect 19555 30640 19564 30680
rect 19604 30640 19613 30680
rect 19555 30639 19613 30640
rect 19947 30680 19989 30689
rect 19947 30640 19948 30680
rect 19988 30640 19989 30680
rect 19947 30631 19989 30640
rect 20043 30680 20085 30689
rect 20043 30640 20044 30680
rect 20084 30640 20085 30680
rect 20043 30631 20085 30640
rect 15627 30586 15669 30595
rect 14283 30547 14325 30556
rect 11491 30512 11549 30513
rect 11491 30472 11500 30512
rect 11540 30472 11549 30512
rect 11491 30471 11549 30472
rect 12739 30512 12797 30513
rect 12739 30472 12748 30512
rect 12788 30472 12797 30512
rect 12739 30471 12797 30472
rect 19275 30512 19317 30521
rect 19275 30472 19276 30512
rect 19316 30472 19317 30512
rect 19275 30463 19317 30472
rect 17931 30428 17973 30437
rect 17931 30388 17932 30428
rect 17972 30388 17973 30428
rect 17931 30379 17973 30388
rect 19075 30428 19133 30429
rect 19075 30388 19084 30428
rect 19124 30388 19133 30428
rect 19075 30387 19133 30388
rect 1152 30260 20352 30284
rect 1152 30220 3688 30260
rect 3728 30220 3770 30260
rect 3810 30220 3852 30260
rect 3892 30220 3934 30260
rect 3974 30220 4016 30260
rect 4056 30220 18808 30260
rect 18848 30220 18890 30260
rect 18930 30220 18972 30260
rect 19012 30220 19054 30260
rect 19094 30220 19136 30260
rect 19176 30220 20352 30260
rect 1152 30196 20352 30220
rect 2667 30092 2709 30101
rect 2667 30052 2668 30092
rect 2708 30052 2709 30092
rect 2667 30043 2709 30052
rect 4395 30092 4437 30101
rect 4395 30052 4396 30092
rect 4436 30052 4437 30092
rect 4395 30043 4437 30052
rect 6027 30092 6069 30101
rect 6027 30052 6028 30092
rect 6068 30052 6069 30092
rect 6027 30043 6069 30052
rect 14667 30092 14709 30101
rect 14667 30052 14668 30092
rect 14708 30052 14709 30092
rect 14667 30043 14709 30052
rect 20227 30092 20285 30093
rect 20227 30052 20236 30092
rect 20276 30052 20285 30092
rect 20227 30051 20285 30052
rect 9195 30008 9237 30017
rect 9195 29968 9196 30008
rect 9236 29968 9237 30008
rect 9195 29959 9237 29968
rect 10147 30008 10205 30009
rect 10147 29968 10156 30008
rect 10196 29968 10205 30008
rect 10147 29967 10205 29968
rect 15619 30008 15677 30009
rect 15619 29968 15628 30008
rect 15668 29968 15677 30008
rect 15619 29967 15677 29968
rect 18123 29924 18165 29933
rect 18123 29884 18124 29924
rect 18164 29884 18165 29924
rect 18123 29875 18165 29884
rect 1219 29840 1277 29841
rect 1219 29800 1228 29840
rect 1268 29800 1277 29840
rect 1219 29799 1277 29800
rect 2467 29840 2525 29841
rect 2467 29800 2476 29840
rect 2516 29800 2525 29840
rect 2467 29799 2525 29800
rect 2947 29840 3005 29841
rect 2947 29800 2956 29840
rect 2996 29800 3005 29840
rect 2947 29799 3005 29800
rect 4195 29840 4253 29841
rect 4195 29800 4204 29840
rect 4244 29800 4253 29840
rect 4195 29799 4253 29800
rect 4579 29840 4637 29841
rect 4579 29800 4588 29840
rect 4628 29800 4637 29840
rect 4579 29799 4637 29800
rect 5827 29840 5885 29841
rect 5827 29800 5836 29840
rect 5876 29800 5885 29840
rect 5827 29799 5885 29800
rect 7075 29840 7133 29841
rect 7075 29800 7084 29840
rect 7124 29800 7133 29840
rect 7075 29799 7133 29800
rect 8323 29840 8381 29841
rect 8323 29800 8332 29840
rect 8372 29800 8381 29840
rect 8323 29799 8381 29800
rect 9003 29840 9045 29849
rect 9003 29800 9004 29840
rect 9044 29800 9045 29840
rect 9003 29791 9045 29800
rect 9195 29840 9237 29849
rect 9195 29800 9196 29840
rect 9236 29800 9237 29840
rect 9195 29791 9237 29800
rect 9475 29840 9533 29841
rect 9475 29800 9484 29840
rect 9524 29800 9533 29840
rect 9475 29799 9533 29800
rect 9771 29840 9813 29849
rect 9771 29800 9772 29840
rect 9812 29800 9813 29840
rect 9771 29791 9813 29800
rect 10443 29840 10485 29849
rect 10443 29800 10444 29840
rect 10484 29800 10485 29840
rect 10443 29791 10485 29800
rect 10635 29840 10677 29849
rect 10635 29800 10636 29840
rect 10676 29800 10677 29840
rect 10635 29791 10677 29800
rect 10723 29840 10781 29841
rect 10723 29800 10732 29840
rect 10772 29800 10781 29840
rect 10723 29799 10781 29800
rect 10915 29840 10973 29841
rect 10915 29800 10924 29840
rect 10964 29800 10973 29840
rect 10915 29799 10973 29800
rect 12163 29840 12221 29841
rect 12163 29800 12172 29840
rect 12212 29800 12221 29840
rect 12163 29799 12221 29800
rect 12651 29840 12693 29849
rect 12651 29800 12652 29840
rect 12692 29800 12693 29840
rect 12651 29791 12693 29800
rect 12939 29840 12981 29849
rect 12939 29800 12940 29840
rect 12980 29800 12981 29840
rect 12939 29791 12981 29800
rect 13219 29840 13277 29841
rect 13219 29800 13228 29840
rect 13268 29800 13277 29840
rect 13219 29799 13277 29800
rect 14467 29840 14525 29841
rect 14467 29800 14476 29840
rect 14516 29800 14525 29840
rect 14467 29799 14525 29800
rect 14947 29840 15005 29841
rect 14947 29800 14956 29840
rect 14996 29800 15005 29840
rect 14947 29799 15005 29800
rect 15243 29840 15285 29849
rect 15243 29800 15244 29840
rect 15284 29800 15285 29840
rect 15243 29791 15285 29800
rect 15819 29840 15861 29849
rect 15819 29800 15820 29840
rect 15860 29800 15861 29840
rect 15819 29791 15861 29800
rect 15915 29840 15957 29849
rect 15915 29800 15916 29840
rect 15956 29800 15957 29840
rect 15915 29791 15957 29800
rect 17547 29840 17589 29849
rect 17547 29800 17548 29840
rect 17588 29800 17589 29840
rect 17547 29791 17589 29800
rect 17643 29840 17685 29849
rect 17643 29800 17644 29840
rect 17684 29800 17685 29840
rect 17643 29791 17685 29800
rect 18027 29840 18069 29849
rect 19083 29845 19125 29854
rect 18027 29800 18028 29840
rect 18068 29800 18069 29840
rect 18027 29791 18069 29800
rect 18595 29840 18653 29841
rect 18595 29800 18604 29840
rect 18644 29800 18653 29840
rect 18595 29799 18653 29800
rect 19083 29805 19084 29845
rect 19124 29805 19125 29845
rect 19083 29796 19125 29805
rect 19555 29840 19613 29841
rect 19555 29800 19564 29840
rect 19604 29800 19613 29840
rect 19555 29799 19613 29800
rect 19851 29840 19893 29849
rect 19851 29800 19852 29840
rect 19892 29800 19893 29840
rect 19851 29791 19893 29800
rect 9867 29756 9909 29765
rect 9867 29716 9868 29756
rect 9908 29716 9909 29756
rect 9867 29707 9909 29716
rect 15339 29756 15381 29765
rect 15339 29716 15340 29756
rect 15380 29716 15381 29756
rect 15339 29707 15381 29716
rect 19275 29756 19317 29765
rect 19275 29716 19276 29756
rect 19316 29716 19317 29756
rect 19275 29707 19317 29716
rect 19947 29756 19989 29765
rect 19947 29716 19948 29756
rect 19988 29716 19989 29756
rect 19947 29707 19989 29716
rect 8523 29672 8565 29681
rect 8523 29632 8524 29672
rect 8564 29632 8565 29672
rect 8523 29623 8565 29632
rect 10531 29672 10589 29673
rect 10531 29632 10540 29672
rect 10580 29632 10589 29672
rect 10531 29631 10589 29632
rect 12363 29672 12405 29681
rect 12363 29632 12364 29672
rect 12404 29632 12405 29672
rect 12363 29623 12405 29632
rect 12747 29672 12789 29681
rect 12747 29632 12748 29672
rect 12788 29632 12789 29672
rect 12747 29623 12789 29632
rect 16099 29672 16157 29673
rect 16099 29632 16108 29672
rect 16148 29632 16157 29672
rect 16099 29631 16157 29632
rect 1152 29504 20452 29528
rect 1152 29464 4928 29504
rect 4968 29464 5010 29504
rect 5050 29464 5092 29504
rect 5132 29464 5174 29504
rect 5214 29464 5256 29504
rect 5296 29464 20048 29504
rect 20088 29464 20130 29504
rect 20170 29464 20212 29504
rect 20252 29464 20294 29504
rect 20334 29464 20376 29504
rect 20416 29464 20452 29504
rect 1152 29440 20452 29464
rect 1899 29336 1941 29345
rect 1899 29296 1900 29336
rect 1940 29296 1941 29336
rect 1899 29287 1941 29296
rect 3819 29336 3861 29345
rect 3819 29296 3820 29336
rect 3860 29296 3861 29336
rect 3819 29287 3861 29296
rect 10723 29336 10781 29337
rect 10723 29296 10732 29336
rect 10772 29296 10781 29336
rect 10723 29295 10781 29296
rect 11395 29336 11453 29337
rect 11395 29296 11404 29336
rect 11444 29296 11453 29336
rect 11395 29295 11453 29296
rect 13611 29336 13653 29345
rect 13611 29296 13612 29336
rect 13652 29296 13653 29336
rect 13611 29287 13653 29296
rect 16299 29336 16341 29345
rect 16299 29296 16300 29336
rect 16340 29296 16341 29336
rect 16299 29287 16341 29296
rect 17731 29336 17789 29337
rect 17731 29296 17740 29336
rect 17780 29296 17789 29336
rect 17731 29295 17789 29296
rect 20035 29336 20093 29337
rect 20035 29296 20044 29336
rect 20084 29296 20093 29336
rect 20035 29295 20093 29296
rect 6603 29252 6645 29261
rect 6603 29212 6604 29252
rect 6644 29212 6645 29252
rect 6603 29203 6645 29212
rect 8619 29252 8661 29261
rect 8619 29212 8620 29252
rect 8660 29212 8661 29252
rect 8619 29203 8661 29212
rect 11883 29188 11925 29197
rect 2371 29168 2429 29169
rect 2371 29128 2380 29168
rect 2420 29128 2429 29168
rect 2371 29127 2429 29128
rect 3619 29168 3677 29169
rect 3619 29128 3628 29168
rect 3668 29128 3677 29168
rect 3619 29127 3677 29128
rect 4003 29168 4061 29169
rect 4003 29128 4012 29168
rect 4052 29128 4061 29168
rect 4003 29127 4061 29128
rect 4203 29168 4245 29177
rect 4203 29128 4204 29168
rect 4244 29128 4245 29168
rect 4203 29119 4245 29128
rect 5155 29168 5213 29169
rect 5155 29128 5164 29168
rect 5204 29128 5213 29168
rect 5155 29127 5213 29128
rect 6403 29168 6461 29169
rect 6403 29128 6412 29168
rect 6452 29128 6461 29168
rect 6403 29127 6461 29128
rect 6891 29168 6933 29177
rect 6891 29128 6892 29168
rect 6932 29128 6933 29168
rect 6891 29119 6933 29128
rect 6987 29168 7029 29177
rect 6987 29128 6988 29168
rect 7028 29128 7029 29168
rect 6987 29119 7029 29128
rect 7371 29168 7413 29177
rect 7371 29128 7372 29168
rect 7412 29128 7413 29168
rect 7371 29119 7413 29128
rect 7939 29168 7997 29169
rect 7939 29128 7948 29168
rect 7988 29128 7997 29168
rect 8995 29168 9053 29169
rect 7939 29127 7997 29128
rect 8475 29158 8517 29167
rect 8475 29118 8476 29158
rect 8516 29118 8517 29158
rect 8995 29128 9004 29168
rect 9044 29128 9053 29168
rect 8995 29127 9053 29128
rect 10243 29168 10301 29169
rect 10243 29128 10252 29168
rect 10292 29128 10301 29168
rect 10243 29127 10301 29128
rect 10635 29168 10677 29177
rect 10635 29128 10636 29168
rect 10676 29128 10677 29168
rect 10635 29119 10677 29128
rect 10827 29168 10869 29177
rect 10827 29128 10828 29168
rect 10868 29128 10869 29168
rect 10827 29119 10869 29128
rect 10915 29168 10973 29169
rect 10915 29128 10924 29168
rect 10964 29128 10973 29168
rect 10915 29127 10973 29128
rect 11115 29168 11157 29177
rect 11115 29128 11116 29168
rect 11156 29128 11157 29168
rect 11115 29119 11157 29128
rect 11211 29168 11253 29177
rect 11211 29128 11212 29168
rect 11252 29128 11253 29168
rect 11883 29148 11884 29188
rect 11924 29148 11925 29188
rect 11883 29139 11925 29148
rect 11979 29168 12021 29177
rect 11211 29119 11253 29128
rect 11979 29128 11980 29168
rect 12020 29128 12021 29168
rect 11979 29119 12021 29128
rect 12363 29168 12405 29177
rect 12363 29128 12364 29168
rect 12404 29128 12405 29168
rect 12363 29119 12405 29128
rect 12459 29168 12501 29177
rect 12459 29128 12460 29168
rect 12500 29128 12501 29168
rect 12459 29119 12501 29128
rect 12931 29168 12989 29169
rect 12931 29128 12940 29168
rect 12980 29128 12989 29168
rect 14467 29168 14525 29169
rect 12931 29127 12989 29128
rect 13467 29126 13509 29135
rect 14467 29128 14476 29168
rect 14516 29128 14525 29168
rect 14467 29127 14525 29128
rect 15715 29168 15773 29169
rect 15715 29128 15724 29168
rect 15764 29128 15773 29168
rect 15715 29127 15773 29128
rect 16203 29168 16245 29177
rect 16203 29128 16204 29168
rect 16244 29128 16245 29168
rect 8475 29109 8517 29118
rect 2083 29084 2141 29085
rect 2083 29044 2092 29084
rect 2132 29044 2141 29084
rect 2083 29043 2141 29044
rect 7467 29084 7509 29093
rect 7467 29044 7468 29084
rect 7508 29044 7509 29084
rect 13467 29086 13468 29126
rect 13508 29086 13509 29126
rect 16203 29119 16245 29128
rect 16395 29168 16437 29177
rect 16395 29128 16396 29168
rect 16436 29128 16437 29168
rect 16395 29119 16437 29128
rect 16491 29168 16533 29177
rect 16491 29128 16492 29168
rect 16532 29128 16533 29168
rect 16491 29119 16533 29128
rect 16675 29168 16733 29169
rect 16675 29128 16684 29168
rect 16724 29128 16733 29168
rect 16675 29127 16733 29128
rect 16771 29168 16829 29169
rect 16771 29128 16780 29168
rect 16820 29128 16829 29168
rect 16771 29127 16829 29128
rect 16971 29168 17013 29177
rect 16971 29128 16972 29168
rect 17012 29128 17013 29168
rect 16971 29119 17013 29128
rect 17067 29168 17109 29177
rect 17067 29128 17068 29168
rect 17108 29128 17109 29168
rect 17067 29119 17109 29128
rect 17211 29168 17269 29169
rect 17211 29128 17220 29168
rect 17260 29128 17269 29168
rect 17211 29127 17269 29128
rect 17451 29168 17493 29177
rect 17451 29128 17452 29168
rect 17492 29128 17493 29168
rect 17451 29119 17493 29128
rect 17547 29168 17589 29177
rect 17547 29128 17548 29168
rect 17588 29128 17589 29168
rect 17547 29119 17589 29128
rect 18027 29168 18069 29177
rect 18027 29128 18028 29168
rect 18068 29128 18069 29168
rect 18027 29119 18069 29128
rect 18115 29168 18173 29169
rect 18115 29128 18124 29168
rect 18164 29128 18173 29168
rect 18115 29127 18173 29128
rect 18307 29168 18365 29169
rect 18307 29128 18316 29168
rect 18356 29128 18365 29168
rect 18307 29127 18365 29128
rect 19555 29168 19613 29169
rect 19555 29128 19564 29168
rect 19604 29128 19613 29168
rect 19555 29127 19613 29128
rect 19947 29168 19989 29177
rect 19947 29128 19948 29168
rect 19988 29128 19989 29168
rect 19947 29119 19989 29128
rect 20139 29168 20181 29177
rect 20139 29128 20140 29168
rect 20180 29128 20181 29168
rect 20139 29119 20181 29128
rect 20227 29168 20285 29169
rect 20227 29128 20236 29168
rect 20276 29128 20285 29168
rect 20227 29127 20285 29128
rect 13467 29077 13509 29086
rect 7467 29035 7509 29044
rect 19755 29000 19797 29009
rect 19755 28960 19756 29000
rect 19796 28960 19797 29000
rect 19755 28951 19797 28960
rect 4107 28916 4149 28925
rect 4107 28876 4108 28916
rect 4148 28876 4149 28916
rect 4107 28867 4149 28876
rect 10443 28916 10485 28925
rect 10443 28876 10444 28916
rect 10484 28876 10485 28916
rect 10443 28867 10485 28876
rect 15915 28916 15957 28925
rect 15915 28876 15916 28916
rect 15956 28876 15957 28916
rect 15915 28867 15957 28876
rect 16683 28916 16725 28925
rect 16683 28876 16684 28916
rect 16724 28876 16725 28916
rect 16683 28867 16725 28876
rect 1152 28748 20352 28772
rect 1152 28708 3688 28748
rect 3728 28708 3770 28748
rect 3810 28708 3852 28748
rect 3892 28708 3934 28748
rect 3974 28708 4016 28748
rect 4056 28708 18808 28748
rect 18848 28708 18890 28748
rect 18930 28708 18972 28748
rect 19012 28708 19054 28748
rect 19094 28708 19136 28748
rect 19176 28708 20352 28748
rect 1152 28684 20352 28708
rect 2667 28580 2709 28589
rect 2667 28540 2668 28580
rect 2708 28540 2709 28580
rect 2667 28531 2709 28540
rect 13515 28580 13557 28589
rect 13515 28540 13516 28580
rect 13556 28540 13557 28580
rect 13515 28531 13557 28540
rect 16395 28580 16437 28589
rect 16395 28540 16396 28580
rect 16436 28540 16437 28580
rect 16395 28531 16437 28540
rect 5547 28496 5589 28505
rect 5547 28456 5548 28496
rect 5588 28456 5589 28496
rect 5547 28447 5589 28456
rect 6411 28412 6453 28421
rect 6411 28372 6412 28412
rect 6452 28372 6453 28412
rect 6411 28363 6453 28372
rect 15051 28412 15093 28421
rect 15051 28372 15052 28412
rect 15092 28372 15093 28412
rect 15051 28363 15093 28372
rect 16011 28342 16053 28351
rect 1219 28328 1277 28329
rect 1219 28288 1228 28328
rect 1268 28288 1277 28328
rect 1219 28287 1277 28288
rect 2467 28328 2525 28329
rect 2467 28288 2476 28328
rect 2516 28288 2525 28328
rect 2467 28287 2525 28288
rect 3147 28328 3189 28337
rect 3147 28288 3148 28328
rect 3188 28288 3189 28328
rect 3147 28279 3189 28288
rect 3243 28328 3285 28337
rect 3243 28288 3244 28328
rect 3284 28288 3285 28328
rect 3243 28279 3285 28288
rect 3619 28328 3677 28329
rect 3619 28288 3628 28328
rect 3668 28288 3677 28328
rect 3619 28287 3677 28288
rect 3723 28328 3765 28337
rect 3723 28288 3724 28328
rect 3764 28288 3765 28328
rect 3723 28279 3765 28288
rect 3907 28328 3965 28329
rect 3907 28288 3916 28328
rect 3956 28288 3965 28328
rect 3907 28287 3965 28288
rect 4099 28328 4157 28329
rect 4099 28288 4108 28328
rect 4148 28288 4157 28328
rect 4099 28287 4157 28288
rect 5347 28328 5405 28329
rect 5347 28288 5356 28328
rect 5396 28288 5405 28328
rect 5347 28287 5405 28288
rect 5835 28328 5877 28337
rect 5835 28288 5836 28328
rect 5876 28288 5877 28328
rect 5835 28279 5877 28288
rect 5931 28328 5973 28337
rect 5931 28288 5932 28328
rect 5972 28288 5973 28328
rect 5931 28279 5973 28288
rect 6315 28328 6357 28337
rect 7371 28333 7413 28342
rect 6315 28288 6316 28328
rect 6356 28288 6357 28328
rect 6315 28279 6357 28288
rect 6883 28328 6941 28329
rect 6883 28288 6892 28328
rect 6932 28288 6941 28328
rect 6883 28287 6941 28288
rect 7371 28293 7372 28333
rect 7412 28293 7413 28333
rect 7371 28284 7413 28293
rect 8035 28328 8093 28329
rect 8035 28288 8044 28328
rect 8084 28288 8093 28328
rect 8035 28287 8093 28288
rect 9283 28328 9341 28329
rect 9283 28288 9292 28328
rect 9332 28288 9341 28328
rect 9283 28287 9341 28288
rect 9859 28328 9917 28329
rect 9859 28288 9868 28328
rect 9908 28288 9917 28328
rect 9859 28287 9917 28288
rect 11107 28328 11165 28329
rect 11107 28288 11116 28328
rect 11156 28288 11165 28328
rect 11107 28287 11165 28288
rect 11499 28328 11541 28337
rect 11499 28288 11500 28328
rect 11540 28288 11541 28328
rect 11499 28279 11541 28288
rect 11595 28328 11637 28337
rect 11595 28288 11596 28328
rect 11636 28288 11637 28328
rect 11595 28279 11637 28288
rect 11691 28328 11733 28337
rect 11691 28288 11692 28328
rect 11732 28288 11733 28328
rect 11691 28279 11733 28288
rect 12067 28328 12125 28329
rect 12067 28288 12076 28328
rect 12116 28288 12125 28328
rect 12067 28287 12125 28288
rect 13315 28328 13373 28329
rect 13315 28288 13324 28328
rect 13364 28288 13373 28328
rect 13315 28287 13373 28288
rect 14475 28328 14517 28337
rect 14475 28288 14476 28328
rect 14516 28288 14517 28328
rect 14475 28279 14517 28288
rect 14571 28328 14613 28337
rect 14571 28288 14572 28328
rect 14612 28288 14613 28328
rect 14571 28279 14613 28288
rect 14955 28328 14997 28337
rect 14955 28288 14956 28328
rect 14996 28288 14997 28328
rect 14955 28279 14997 28288
rect 15523 28328 15581 28329
rect 15523 28288 15532 28328
rect 15572 28288 15581 28328
rect 16011 28302 16012 28342
rect 16052 28302 16053 28342
rect 16011 28293 16053 28302
rect 16579 28328 16637 28329
rect 15523 28287 15581 28288
rect 16579 28288 16588 28328
rect 16628 28288 16637 28328
rect 16579 28287 16637 28288
rect 17827 28328 17885 28329
rect 17827 28288 17836 28328
rect 17876 28288 17885 28328
rect 17827 28287 17885 28288
rect 18211 28328 18269 28329
rect 18211 28288 18220 28328
rect 18260 28288 18269 28328
rect 18211 28287 18269 28288
rect 19459 28328 19517 28329
rect 19459 28288 19468 28328
rect 19508 28288 19517 28328
rect 19459 28287 19517 28288
rect 19851 28328 19893 28337
rect 19851 28288 19852 28328
rect 19892 28288 19893 28328
rect 19851 28279 19893 28288
rect 19947 28328 19989 28337
rect 19947 28288 19948 28328
rect 19988 28288 19989 28328
rect 19947 28279 19989 28288
rect 20043 28328 20085 28337
rect 20043 28288 20044 28328
rect 20084 28288 20085 28328
rect 20043 28279 20085 28288
rect 3427 28160 3485 28161
rect 3427 28120 3436 28160
rect 3476 28120 3485 28160
rect 3427 28119 3485 28120
rect 3915 28160 3957 28169
rect 3915 28120 3916 28160
rect 3956 28120 3957 28160
rect 3915 28111 3957 28120
rect 7563 28160 7605 28169
rect 7563 28120 7564 28160
rect 7604 28120 7605 28160
rect 7563 28111 7605 28120
rect 9483 28160 9525 28169
rect 9483 28120 9484 28160
rect 9524 28120 9525 28160
rect 9483 28111 9525 28120
rect 11307 28160 11349 28169
rect 11307 28120 11308 28160
rect 11348 28120 11349 28160
rect 11307 28111 11349 28120
rect 11779 28160 11837 28161
rect 11779 28120 11788 28160
rect 11828 28120 11837 28160
rect 11779 28119 11837 28120
rect 16203 28160 16245 28169
rect 16203 28120 16204 28160
rect 16244 28120 16245 28160
rect 16203 28111 16245 28120
rect 19659 28160 19701 28169
rect 19659 28120 19660 28160
rect 19700 28120 19701 28160
rect 19659 28111 19701 28120
rect 20131 28160 20189 28161
rect 20131 28120 20140 28160
rect 20180 28120 20189 28160
rect 20131 28119 20189 28120
rect 1152 27992 20452 28016
rect 1152 27952 4928 27992
rect 4968 27952 5010 27992
rect 5050 27952 5092 27992
rect 5132 27952 5174 27992
rect 5214 27952 5256 27992
rect 5296 27952 20048 27992
rect 20088 27952 20130 27992
rect 20170 27952 20212 27992
rect 20252 27952 20294 27992
rect 20334 27952 20376 27992
rect 20416 27952 20452 27992
rect 1152 27928 20452 27952
rect 4483 27824 4541 27825
rect 4483 27784 4492 27824
rect 4532 27784 4541 27824
rect 4483 27783 4541 27784
rect 7371 27824 7413 27833
rect 7371 27784 7372 27824
rect 7412 27784 7413 27824
rect 7371 27775 7413 27784
rect 14475 27824 14517 27833
rect 14475 27784 14476 27824
rect 14516 27784 14517 27824
rect 14475 27775 14517 27784
rect 17355 27824 17397 27833
rect 17355 27784 17356 27824
rect 17396 27784 17397 27824
rect 17355 27775 17397 27784
rect 20035 27824 20093 27825
rect 20035 27784 20044 27824
rect 20084 27784 20093 27824
rect 20035 27783 20093 27784
rect 2667 27740 2709 27749
rect 2667 27700 2668 27740
rect 2708 27700 2709 27740
rect 2667 27691 2709 27700
rect 4299 27740 4341 27749
rect 4299 27700 4300 27740
rect 4340 27700 4341 27740
rect 4299 27691 4341 27700
rect 10347 27740 10389 27749
rect 10347 27700 10348 27740
rect 10388 27700 10389 27740
rect 10347 27691 10389 27700
rect 1219 27656 1277 27657
rect 1219 27616 1228 27656
rect 1268 27616 1277 27656
rect 1219 27615 1277 27616
rect 2467 27656 2525 27657
rect 2467 27616 2476 27656
rect 2516 27616 2525 27656
rect 2467 27615 2525 27616
rect 2851 27656 2909 27657
rect 2851 27616 2860 27656
rect 2900 27616 2909 27656
rect 2851 27615 2909 27616
rect 4099 27656 4157 27657
rect 4099 27616 4108 27656
rect 4148 27616 4157 27656
rect 4099 27615 4157 27616
rect 4683 27656 4725 27665
rect 4683 27616 4684 27656
rect 4724 27616 4725 27656
rect 4683 27607 4725 27616
rect 4779 27656 4821 27665
rect 4779 27616 4780 27656
rect 4820 27616 4821 27656
rect 4779 27607 4821 27616
rect 4971 27656 5013 27665
rect 4971 27616 4972 27656
rect 5012 27616 5013 27656
rect 4971 27607 5013 27616
rect 5259 27656 5301 27665
rect 5259 27616 5260 27656
rect 5300 27616 5301 27656
rect 5259 27607 5301 27616
rect 5451 27656 5493 27665
rect 5451 27616 5452 27656
rect 5492 27616 5493 27656
rect 5451 27607 5493 27616
rect 5643 27656 5685 27665
rect 5643 27616 5644 27656
rect 5684 27616 5685 27656
rect 5643 27607 5685 27616
rect 5923 27656 5981 27657
rect 5923 27616 5932 27656
rect 5972 27616 5981 27656
rect 5923 27615 5981 27616
rect 7171 27656 7229 27657
rect 7171 27616 7180 27656
rect 7220 27616 7229 27656
rect 7171 27615 7229 27616
rect 8619 27656 8661 27665
rect 8619 27616 8620 27656
rect 8660 27616 8661 27656
rect 8619 27607 8661 27616
rect 8715 27656 8757 27665
rect 8715 27616 8716 27656
rect 8756 27616 8757 27656
rect 8715 27607 8757 27616
rect 9099 27656 9141 27665
rect 9099 27616 9100 27656
rect 9140 27616 9141 27656
rect 9099 27607 9141 27616
rect 9667 27656 9725 27657
rect 9667 27616 9676 27656
rect 9716 27616 9725 27656
rect 10915 27656 10973 27657
rect 9667 27615 9725 27616
rect 10203 27646 10245 27655
rect 10203 27606 10204 27646
rect 10244 27606 10245 27646
rect 10915 27616 10924 27656
rect 10964 27616 10973 27656
rect 10915 27615 10973 27616
rect 12163 27656 12221 27657
rect 12163 27616 12172 27656
rect 12212 27616 12221 27656
rect 12163 27615 12221 27616
rect 13027 27656 13085 27657
rect 13027 27616 13036 27656
rect 13076 27616 13085 27656
rect 13027 27615 13085 27616
rect 14275 27656 14333 27657
rect 14275 27616 14284 27656
rect 14324 27616 14333 27656
rect 14275 27615 14333 27616
rect 15619 27656 15677 27657
rect 15619 27616 15628 27656
rect 15668 27616 15677 27656
rect 15619 27615 15677 27616
rect 15723 27656 15765 27665
rect 19755 27657 19797 27666
rect 15723 27616 15724 27656
rect 15764 27616 15765 27656
rect 15723 27607 15765 27616
rect 15907 27656 15965 27657
rect 15907 27616 15916 27656
rect 15956 27616 15965 27656
rect 15907 27615 15965 27616
rect 17155 27656 17213 27657
rect 17155 27616 17164 27656
rect 17204 27616 17213 27656
rect 17155 27615 17213 27616
rect 18115 27656 18173 27657
rect 18115 27616 18124 27656
rect 18164 27616 18173 27656
rect 18115 27615 18173 27616
rect 19363 27635 19421 27636
rect 10203 27597 10245 27606
rect 19363 27595 19372 27635
rect 19412 27595 19421 27635
rect 19755 27617 19756 27657
rect 19796 27617 19797 27657
rect 19755 27608 19797 27617
rect 19851 27656 19893 27665
rect 19851 27616 19852 27656
rect 19892 27616 19893 27656
rect 19851 27607 19893 27616
rect 19363 27594 19421 27595
rect 9195 27572 9237 27581
rect 9195 27532 9196 27572
rect 9236 27532 9237 27572
rect 9195 27523 9237 27532
rect 5451 27488 5493 27497
rect 5451 27448 5452 27488
rect 5492 27448 5493 27488
rect 5451 27439 5493 27448
rect 5259 27404 5301 27413
rect 5259 27364 5260 27404
rect 5300 27364 5301 27404
rect 5259 27355 5301 27364
rect 12363 27404 12405 27413
rect 12363 27364 12364 27404
rect 12404 27364 12405 27404
rect 12363 27355 12405 27364
rect 19563 27404 19605 27413
rect 19563 27364 19564 27404
rect 19604 27364 19605 27404
rect 19563 27355 19605 27364
rect 1152 27236 20352 27260
rect 1152 27196 3688 27236
rect 3728 27196 3770 27236
rect 3810 27196 3852 27236
rect 3892 27196 3934 27236
rect 3974 27196 4016 27236
rect 4056 27196 18808 27236
rect 18848 27196 18890 27236
rect 18930 27196 18972 27236
rect 19012 27196 19054 27236
rect 19094 27196 19136 27236
rect 19176 27196 20352 27236
rect 1152 27172 20352 27196
rect 4099 27068 4157 27069
rect 4099 27028 4108 27068
rect 4148 27028 4157 27068
rect 4099 27027 4157 27028
rect 1995 26900 2037 26909
rect 1995 26860 1996 26900
rect 2036 26860 2037 26900
rect 1995 26851 2037 26860
rect 6795 26900 6837 26909
rect 6795 26860 6796 26900
rect 6836 26860 6837 26900
rect 6795 26851 6837 26860
rect 17835 26900 17877 26909
rect 17835 26860 17836 26900
rect 17876 26860 17877 26900
rect 17835 26851 17877 26860
rect 3003 26825 3045 26834
rect 1419 26816 1461 26825
rect 1419 26776 1420 26816
rect 1460 26776 1461 26816
rect 1419 26767 1461 26776
rect 1515 26816 1557 26825
rect 1515 26776 1516 26816
rect 1556 26776 1557 26816
rect 1515 26767 1557 26776
rect 1899 26816 1941 26825
rect 1899 26776 1900 26816
rect 1940 26776 1941 26816
rect 1899 26767 1941 26776
rect 2467 26816 2525 26817
rect 2467 26776 2476 26816
rect 2516 26776 2525 26816
rect 3003 26785 3004 26825
rect 3044 26785 3045 26825
rect 3003 26776 3045 26785
rect 3427 26816 3485 26817
rect 3427 26776 3436 26816
rect 3476 26776 3485 26816
rect 2467 26775 2525 26776
rect 3427 26775 3485 26776
rect 3723 26816 3765 26825
rect 3723 26776 3724 26816
rect 3764 26776 3765 26816
rect 3723 26767 3765 26776
rect 4483 26816 4541 26817
rect 4483 26776 4492 26816
rect 4532 26776 4541 26816
rect 4483 26775 4541 26776
rect 5731 26816 5789 26817
rect 5731 26776 5740 26816
rect 5780 26776 5789 26816
rect 5731 26775 5789 26776
rect 6219 26816 6261 26825
rect 6219 26776 6220 26816
rect 6260 26776 6261 26816
rect 6219 26767 6261 26776
rect 6315 26816 6357 26825
rect 6315 26776 6316 26816
rect 6356 26776 6357 26816
rect 6315 26767 6357 26776
rect 6699 26816 6741 26825
rect 7755 26821 7797 26830
rect 13371 26825 13413 26834
rect 18939 26825 18981 26834
rect 6699 26776 6700 26816
rect 6740 26776 6741 26816
rect 6699 26767 6741 26776
rect 7267 26816 7325 26817
rect 7267 26776 7276 26816
rect 7316 26776 7325 26816
rect 7267 26775 7325 26776
rect 7755 26781 7756 26821
rect 7796 26781 7797 26821
rect 7755 26772 7797 26781
rect 8323 26816 8381 26817
rect 8323 26776 8332 26816
rect 8372 26776 8381 26816
rect 8323 26775 8381 26776
rect 9571 26816 9629 26817
rect 9571 26776 9580 26816
rect 9620 26776 9629 26816
rect 9571 26775 9629 26776
rect 10059 26816 10101 26825
rect 10059 26776 10060 26816
rect 10100 26776 10101 26816
rect 10059 26767 10101 26776
rect 10155 26816 10197 26825
rect 10155 26776 10156 26816
rect 10196 26776 10197 26816
rect 10155 26767 10197 26776
rect 10251 26816 10293 26825
rect 10251 26776 10252 26816
rect 10292 26776 10293 26816
rect 10251 26767 10293 26776
rect 10539 26816 10581 26825
rect 10539 26776 10540 26816
rect 10580 26776 10581 26816
rect 10539 26767 10581 26776
rect 10635 26816 10677 26825
rect 10635 26776 10636 26816
rect 10676 26776 10677 26816
rect 10635 26767 10677 26776
rect 11019 26816 11061 26825
rect 11019 26776 11020 26816
rect 11060 26776 11061 26816
rect 11019 26767 11061 26776
rect 11115 26816 11157 26825
rect 11115 26776 11116 26816
rect 11156 26776 11157 26816
rect 11115 26767 11157 26776
rect 11787 26816 11829 26825
rect 11787 26776 11788 26816
rect 11828 26776 11829 26816
rect 11787 26767 11829 26776
rect 11883 26816 11925 26825
rect 11883 26776 11884 26816
rect 11924 26776 11925 26816
rect 11883 26767 11925 26776
rect 12267 26816 12309 26825
rect 12267 26776 12268 26816
rect 12308 26776 12309 26816
rect 12267 26767 12309 26776
rect 12363 26816 12405 26825
rect 12363 26776 12364 26816
rect 12404 26776 12405 26816
rect 12363 26767 12405 26776
rect 12835 26816 12893 26817
rect 12835 26776 12844 26816
rect 12884 26776 12893 26816
rect 13371 26785 13372 26825
rect 13412 26785 13413 26825
rect 13371 26776 13413 26785
rect 14179 26816 14237 26817
rect 14179 26776 14188 26816
rect 14228 26776 14237 26816
rect 12835 26775 12893 26776
rect 14179 26775 14237 26776
rect 15427 26816 15485 26817
rect 15427 26776 15436 26816
rect 15476 26776 15485 26816
rect 15427 26775 15485 26776
rect 15819 26816 15861 26825
rect 15819 26776 15820 26816
rect 15860 26776 15861 26816
rect 15819 26767 15861 26776
rect 16011 26816 16053 26825
rect 16011 26776 16012 26816
rect 16052 26776 16053 26816
rect 16011 26767 16053 26776
rect 16107 26816 16149 26825
rect 16107 26776 16108 26816
rect 16148 26776 16149 26816
rect 16107 26767 16149 26776
rect 17355 26816 17397 26825
rect 17355 26776 17356 26816
rect 17396 26776 17397 26816
rect 17355 26767 17397 26776
rect 17451 26816 17493 26825
rect 17451 26776 17452 26816
rect 17492 26776 17493 26816
rect 17451 26767 17493 26776
rect 17931 26816 17973 26825
rect 17931 26776 17932 26816
rect 17972 26776 17973 26816
rect 17931 26767 17973 26776
rect 18403 26816 18461 26817
rect 18403 26776 18412 26816
rect 18452 26776 18461 26816
rect 18939 26785 18940 26825
rect 18980 26785 18981 26825
rect 18939 26776 18981 26785
rect 19275 26816 19317 26825
rect 19275 26776 19276 26816
rect 19316 26776 19317 26816
rect 18403 26775 18461 26776
rect 19275 26767 19317 26776
rect 19371 26816 19413 26825
rect 19371 26776 19372 26816
rect 19412 26776 19413 26816
rect 19371 26767 19413 26776
rect 19467 26816 19509 26825
rect 19467 26776 19468 26816
rect 19508 26776 19509 26816
rect 19467 26767 19509 26776
rect 19755 26816 19797 26825
rect 19755 26776 19756 26816
rect 19796 26776 19797 26816
rect 19755 26767 19797 26776
rect 19851 26816 19893 26825
rect 19851 26776 19852 26816
rect 19892 26776 19893 26816
rect 19851 26767 19893 26776
rect 3147 26732 3189 26741
rect 3147 26692 3148 26732
rect 3188 26692 3189 26732
rect 3147 26683 3189 26692
rect 3819 26732 3861 26741
rect 3819 26692 3820 26732
rect 3860 26692 3861 26732
rect 3819 26683 3861 26692
rect 5931 26732 5973 26741
rect 5931 26692 5932 26732
rect 5972 26692 5973 26732
rect 5931 26683 5973 26692
rect 7947 26732 7989 26741
rect 7947 26692 7948 26732
rect 7988 26692 7989 26732
rect 7947 26683 7989 26692
rect 8139 26732 8181 26741
rect 8139 26692 8140 26732
rect 8180 26692 8181 26732
rect 8139 26683 8181 26692
rect 10347 26732 10389 26741
rect 10347 26692 10348 26732
rect 10388 26692 10389 26732
rect 10347 26683 10389 26692
rect 15627 26732 15669 26741
rect 15627 26692 15628 26732
rect 15668 26692 15669 26732
rect 15627 26683 15669 26692
rect 10819 26648 10877 26649
rect 10819 26608 10828 26648
rect 10868 26608 10877 26648
rect 10819 26607 10877 26608
rect 11299 26648 11357 26649
rect 11299 26608 11308 26648
rect 11348 26608 11357 26648
rect 11299 26607 11357 26608
rect 13515 26648 13557 26657
rect 13515 26608 13516 26648
rect 13556 26608 13557 26648
rect 13515 26599 13557 26608
rect 15915 26648 15957 26657
rect 15915 26608 15916 26648
rect 15956 26608 15957 26648
rect 15915 26599 15957 26608
rect 19083 26648 19125 26657
rect 19083 26608 19084 26648
rect 19124 26608 19125 26648
rect 19083 26599 19125 26608
rect 19555 26648 19613 26649
rect 19555 26608 19564 26648
rect 19604 26608 19613 26648
rect 19555 26607 19613 26608
rect 20035 26648 20093 26649
rect 20035 26608 20044 26648
rect 20084 26608 20093 26648
rect 20035 26607 20093 26608
rect 1152 26480 20452 26504
rect 1152 26440 4928 26480
rect 4968 26440 5010 26480
rect 5050 26440 5092 26480
rect 5132 26440 5174 26480
rect 5214 26440 5256 26480
rect 5296 26440 20048 26480
rect 20088 26440 20130 26480
rect 20170 26440 20212 26480
rect 20252 26440 20294 26480
rect 20334 26440 20376 26480
rect 20416 26440 20452 26480
rect 1152 26416 20452 26440
rect 2955 26312 2997 26321
rect 2955 26272 2956 26312
rect 2996 26272 2997 26312
rect 2955 26263 2997 26272
rect 5443 26312 5501 26313
rect 5443 26272 5452 26312
rect 5492 26272 5501 26312
rect 5443 26271 5501 26272
rect 11211 26312 11253 26321
rect 11211 26272 11212 26312
rect 11252 26272 11253 26312
rect 11211 26263 11253 26272
rect 13419 26312 13461 26321
rect 13419 26272 13420 26312
rect 13460 26272 13461 26312
rect 13419 26263 13461 26272
rect 17643 26312 17685 26321
rect 17643 26272 17644 26312
rect 17684 26272 17685 26312
rect 17643 26263 17685 26272
rect 19267 26312 19325 26313
rect 19267 26272 19276 26312
rect 19316 26272 19325 26312
rect 19267 26271 19325 26272
rect 15819 26228 15861 26237
rect 15819 26188 15820 26228
rect 15860 26188 15861 26228
rect 15819 26179 15861 26188
rect 1507 26144 1565 26145
rect 1507 26104 1516 26144
rect 1556 26104 1565 26144
rect 1507 26103 1565 26104
rect 2755 26144 2813 26145
rect 2755 26104 2764 26144
rect 2804 26104 2813 26144
rect 2755 26103 2813 26104
rect 3523 26144 3581 26145
rect 3523 26104 3532 26144
rect 3572 26104 3581 26144
rect 3523 26103 3581 26104
rect 4771 26144 4829 26145
rect 4771 26104 4780 26144
rect 4820 26104 4829 26144
rect 4771 26103 4829 26104
rect 5163 26144 5205 26153
rect 5163 26104 5164 26144
rect 5204 26104 5205 26144
rect 5163 26095 5205 26104
rect 5259 26144 5301 26153
rect 5259 26104 5260 26144
rect 5300 26104 5301 26144
rect 5259 26095 5301 26104
rect 6115 26144 6173 26145
rect 6115 26104 6124 26144
rect 6164 26104 6173 26144
rect 6115 26103 6173 26104
rect 7363 26144 7421 26145
rect 7363 26104 7372 26144
rect 7412 26104 7421 26144
rect 7363 26103 7421 26104
rect 7747 26144 7805 26145
rect 7747 26104 7756 26144
rect 7796 26104 7805 26144
rect 7747 26103 7805 26104
rect 8995 26144 9053 26145
rect 8995 26104 9004 26144
rect 9044 26104 9053 26144
rect 8995 26103 9053 26104
rect 9483 26144 9525 26153
rect 9483 26104 9484 26144
rect 9524 26104 9525 26144
rect 9483 26095 9525 26104
rect 9579 26144 9621 26153
rect 9579 26104 9580 26144
rect 9620 26104 9621 26144
rect 9579 26095 9621 26104
rect 10531 26144 10589 26145
rect 10531 26104 10540 26144
rect 10580 26104 10589 26144
rect 11971 26144 12029 26145
rect 10531 26103 10589 26104
rect 11067 26134 11109 26143
rect 11067 26094 11068 26134
rect 11108 26094 11109 26134
rect 11971 26104 11980 26144
rect 12020 26104 12029 26144
rect 11971 26103 12029 26104
rect 13219 26144 13277 26145
rect 13219 26104 13228 26144
rect 13268 26104 13277 26144
rect 13219 26103 13277 26104
rect 14091 26144 14133 26153
rect 14091 26104 14092 26144
rect 14132 26104 14133 26144
rect 14091 26095 14133 26104
rect 14187 26144 14229 26153
rect 14187 26104 14188 26144
rect 14228 26104 14229 26144
rect 14187 26095 14229 26104
rect 14667 26144 14709 26153
rect 14667 26104 14668 26144
rect 14708 26104 14709 26144
rect 14667 26095 14709 26104
rect 15139 26144 15197 26145
rect 15139 26104 15148 26144
rect 15188 26104 15197 26144
rect 15139 26103 15197 26104
rect 15627 26139 15669 26148
rect 15627 26099 15628 26139
rect 15668 26099 15669 26139
rect 16195 26144 16253 26145
rect 16195 26104 16204 26144
rect 16244 26104 16253 26144
rect 16195 26103 16253 26104
rect 17443 26144 17501 26145
rect 17443 26104 17452 26144
rect 17492 26104 17501 26144
rect 17443 26103 17501 26104
rect 17827 26144 17885 26145
rect 17827 26104 17836 26144
rect 17876 26104 17885 26144
rect 17827 26103 17885 26104
rect 19075 26144 19133 26145
rect 19075 26104 19084 26144
rect 19124 26104 19133 26144
rect 19075 26103 19133 26104
rect 19467 26144 19509 26153
rect 19467 26104 19468 26144
rect 19508 26104 19509 26144
rect 11067 26085 11109 26094
rect 15627 26090 15669 26099
rect 19467 26095 19509 26104
rect 19563 26144 19605 26153
rect 19563 26104 19564 26144
rect 19604 26104 19605 26144
rect 19563 26095 19605 26104
rect 9963 26060 10005 26069
rect 9963 26020 9964 26060
rect 10004 26020 10005 26060
rect 9963 26011 10005 26020
rect 10059 26060 10101 26069
rect 10059 26020 10060 26060
rect 10100 26020 10101 26060
rect 10059 26011 10101 26020
rect 14571 26060 14613 26069
rect 14571 26020 14572 26060
rect 14612 26020 14613 26060
rect 14571 26011 14613 26020
rect 4971 25892 5013 25901
rect 4971 25852 4972 25892
rect 5012 25852 5013 25892
rect 4971 25843 5013 25852
rect 7563 25892 7605 25901
rect 7563 25852 7564 25892
rect 7604 25852 7605 25892
rect 7563 25843 7605 25852
rect 9195 25892 9237 25901
rect 9195 25852 9196 25892
rect 9236 25852 9237 25892
rect 9195 25843 9237 25852
rect 16011 25892 16053 25901
rect 16011 25852 16012 25892
rect 16052 25852 16053 25892
rect 16011 25843 16053 25852
rect 1152 25724 20352 25748
rect 1152 25684 3688 25724
rect 3728 25684 3770 25724
rect 3810 25684 3852 25724
rect 3892 25684 3934 25724
rect 3974 25684 4016 25724
rect 4056 25684 18808 25724
rect 18848 25684 18890 25724
rect 18930 25684 18972 25724
rect 19012 25684 19054 25724
rect 19094 25684 19136 25724
rect 19176 25684 20352 25724
rect 1152 25660 20352 25684
rect 11211 25556 11253 25565
rect 11211 25516 11212 25556
rect 11252 25516 11253 25556
rect 11211 25507 11253 25516
rect 14571 25556 14613 25565
rect 14571 25516 14572 25556
rect 14612 25516 14613 25556
rect 14571 25507 14613 25516
rect 15147 25556 15189 25565
rect 15147 25516 15148 25556
rect 15188 25516 15189 25556
rect 15147 25507 15189 25516
rect 15627 25556 15669 25565
rect 15627 25516 15628 25556
rect 15668 25516 15669 25556
rect 15627 25507 15669 25516
rect 16291 25472 16349 25473
rect 16291 25432 16300 25472
rect 16340 25432 16349 25472
rect 16291 25431 16349 25432
rect 17347 25472 17405 25473
rect 17347 25432 17356 25472
rect 17396 25432 17405 25472
rect 17347 25431 17405 25432
rect 7755 25318 7797 25327
rect 2379 25304 2421 25313
rect 2379 25264 2380 25304
rect 2420 25264 2421 25304
rect 2379 25255 2421 25264
rect 2475 25304 2517 25313
rect 2475 25264 2476 25304
rect 2516 25264 2517 25304
rect 2475 25255 2517 25264
rect 2763 25304 2805 25313
rect 2763 25264 2764 25304
rect 2804 25264 2805 25304
rect 2763 25255 2805 25264
rect 2859 25304 2901 25313
rect 2859 25264 2860 25304
rect 2900 25264 2901 25304
rect 2859 25255 2901 25264
rect 3243 25304 3285 25313
rect 3243 25264 3244 25304
rect 3284 25264 3285 25304
rect 3243 25255 3285 25264
rect 3339 25304 3381 25313
rect 4299 25309 4341 25318
rect 3339 25264 3340 25304
rect 3380 25264 3381 25304
rect 3339 25255 3381 25264
rect 3811 25304 3869 25305
rect 3811 25264 3820 25304
rect 3860 25264 3869 25304
rect 3811 25263 3869 25264
rect 4299 25269 4300 25309
rect 4340 25269 4341 25309
rect 4299 25260 4341 25269
rect 4683 25304 4725 25313
rect 4683 25264 4684 25304
rect 4724 25264 4725 25304
rect 4683 25255 4725 25264
rect 4779 25304 4821 25313
rect 4779 25264 4780 25304
rect 4820 25264 4821 25304
rect 4779 25255 4821 25264
rect 4875 25304 4917 25313
rect 4875 25264 4876 25304
rect 4916 25264 4917 25304
rect 4875 25255 4917 25264
rect 5163 25304 5205 25313
rect 5163 25264 5164 25304
rect 5204 25264 5205 25304
rect 5163 25255 5205 25264
rect 5259 25304 5301 25313
rect 5259 25264 5260 25304
rect 5300 25264 5301 25304
rect 5259 25255 5301 25264
rect 5355 25304 5397 25313
rect 5355 25264 5356 25304
rect 5396 25264 5397 25304
rect 5835 25304 5877 25313
rect 5355 25255 5397 25264
rect 5451 25283 5493 25292
rect 5451 25243 5452 25283
rect 5492 25243 5493 25283
rect 5835 25264 5836 25304
rect 5876 25264 5877 25304
rect 5835 25255 5877 25264
rect 5931 25304 5973 25313
rect 5931 25264 5932 25304
rect 5972 25264 5973 25304
rect 5931 25255 5973 25264
rect 6219 25304 6261 25313
rect 6219 25264 6220 25304
rect 6260 25264 6261 25304
rect 6219 25255 6261 25264
rect 6315 25304 6357 25313
rect 6315 25264 6316 25304
rect 6356 25264 6357 25304
rect 6315 25255 6357 25264
rect 6699 25304 6741 25313
rect 6699 25264 6700 25304
rect 6740 25264 6741 25304
rect 6699 25255 6741 25264
rect 6795 25304 6837 25313
rect 6795 25264 6796 25304
rect 6836 25264 6837 25304
rect 6795 25255 6837 25264
rect 7267 25304 7325 25305
rect 7267 25264 7276 25304
rect 7316 25264 7325 25304
rect 7755 25278 7756 25318
rect 7796 25278 7797 25318
rect 7755 25269 7797 25278
rect 8139 25304 8181 25313
rect 7267 25263 7325 25264
rect 8139 25264 8140 25304
rect 8180 25264 8181 25304
rect 8139 25255 8181 25264
rect 8235 25304 8277 25313
rect 8235 25264 8236 25304
rect 8276 25264 8277 25304
rect 8235 25255 8277 25264
rect 9763 25304 9821 25305
rect 9763 25264 9772 25304
rect 9812 25264 9821 25304
rect 9763 25263 9821 25264
rect 11011 25304 11069 25305
rect 11011 25264 11020 25304
rect 11060 25264 11069 25304
rect 11011 25263 11069 25264
rect 13123 25304 13181 25305
rect 13123 25264 13132 25304
rect 13172 25264 13181 25304
rect 13123 25263 13181 25264
rect 14371 25304 14429 25305
rect 14371 25264 14380 25304
rect 14420 25264 14429 25304
rect 14371 25263 14429 25264
rect 14955 25304 14997 25313
rect 14955 25264 14956 25304
rect 14996 25264 14997 25304
rect 14955 25255 14997 25264
rect 15147 25304 15189 25313
rect 15147 25264 15148 25304
rect 15188 25264 15189 25304
rect 15147 25255 15189 25264
rect 15339 25304 15381 25313
rect 15339 25264 15340 25304
rect 15380 25264 15381 25304
rect 15339 25255 15381 25264
rect 15627 25304 15669 25313
rect 15627 25264 15628 25304
rect 15668 25264 15669 25304
rect 15627 25255 15669 25264
rect 15915 25304 15957 25313
rect 15915 25264 15916 25304
rect 15956 25264 15957 25304
rect 15915 25255 15957 25264
rect 16011 25304 16053 25313
rect 16011 25264 16012 25304
rect 16052 25264 16053 25304
rect 16011 25255 16053 25264
rect 16107 25304 16149 25313
rect 16107 25264 16108 25304
rect 16148 25264 16149 25304
rect 16107 25255 16149 25264
rect 16675 25304 16733 25305
rect 16675 25264 16684 25304
rect 16724 25264 16733 25304
rect 16675 25263 16733 25264
rect 16971 25304 17013 25313
rect 16971 25264 16972 25304
rect 17012 25264 17013 25304
rect 16971 25255 17013 25264
rect 17067 25304 17109 25313
rect 17067 25264 17068 25304
rect 17108 25264 17109 25304
rect 17067 25255 17109 25264
rect 5451 25234 5493 25243
rect 4491 25220 4533 25229
rect 4491 25180 4492 25220
rect 4532 25180 4533 25220
rect 4491 25171 4533 25180
rect 7947 25220 7989 25229
rect 7947 25180 7948 25220
rect 7988 25180 7989 25220
rect 7947 25171 7989 25180
rect 2179 25136 2237 25137
rect 2179 25096 2188 25136
rect 2228 25096 2237 25136
rect 2179 25095 2237 25096
rect 4963 25136 5021 25137
rect 4963 25096 4972 25136
rect 5012 25096 5021 25136
rect 4963 25095 5021 25096
rect 5635 25136 5693 25137
rect 5635 25096 5644 25136
rect 5684 25096 5693 25136
rect 5635 25095 5693 25096
rect 8419 25136 8477 25137
rect 8419 25096 8428 25136
rect 8468 25096 8477 25136
rect 8419 25095 8477 25096
rect 1152 24968 20452 24992
rect 1152 24928 4928 24968
rect 4968 24928 5010 24968
rect 5050 24928 5092 24968
rect 5132 24928 5174 24968
rect 5214 24928 5256 24968
rect 5296 24928 20048 24968
rect 20088 24928 20130 24968
rect 20170 24928 20212 24968
rect 20252 24928 20294 24968
rect 20334 24928 20376 24968
rect 20416 24928 20452 24968
rect 1152 24904 20452 24928
rect 11019 24842 11061 24851
rect 2763 24800 2805 24809
rect 2763 24760 2764 24800
rect 2804 24760 2805 24800
rect 2763 24751 2805 24760
rect 2955 24800 2997 24809
rect 2955 24760 2956 24800
rect 2996 24760 2997 24800
rect 2955 24751 2997 24760
rect 6315 24800 6357 24809
rect 6315 24760 6316 24800
rect 6356 24760 6357 24800
rect 11019 24802 11020 24842
rect 11060 24802 11061 24842
rect 11019 24793 11061 24802
rect 16779 24800 16821 24809
rect 6315 24751 6357 24760
rect 16779 24760 16780 24800
rect 16820 24760 16821 24800
rect 16779 24751 16821 24760
rect 9003 24716 9045 24725
rect 9003 24676 9004 24716
rect 9044 24676 9045 24716
rect 9003 24667 9045 24676
rect 1315 24632 1373 24633
rect 1315 24592 1324 24632
rect 1364 24592 1373 24632
rect 1315 24591 1373 24592
rect 2563 24632 2621 24633
rect 2563 24592 2572 24632
rect 2612 24592 2621 24632
rect 2563 24591 2621 24592
rect 3139 24632 3197 24633
rect 3139 24592 3148 24632
rect 3188 24592 3197 24632
rect 3139 24591 3197 24592
rect 4387 24632 4445 24633
rect 4387 24592 4396 24632
rect 4436 24592 4445 24632
rect 4387 24591 4445 24592
rect 4867 24632 4925 24633
rect 4867 24592 4876 24632
rect 4916 24592 4925 24632
rect 4867 24591 4925 24592
rect 6115 24632 6173 24633
rect 6115 24592 6124 24632
rect 6164 24592 6173 24632
rect 6115 24591 6173 24592
rect 6691 24632 6749 24633
rect 6691 24592 6700 24632
rect 6740 24592 6749 24632
rect 6691 24591 6749 24592
rect 6987 24632 7029 24641
rect 6987 24592 6988 24632
rect 7028 24592 7029 24632
rect 6987 24583 7029 24592
rect 7083 24632 7125 24641
rect 7083 24592 7084 24632
rect 7124 24592 7125 24632
rect 7083 24583 7125 24592
rect 7555 24632 7613 24633
rect 7555 24592 7564 24632
rect 7604 24592 7613 24632
rect 7555 24591 7613 24592
rect 8803 24632 8861 24633
rect 8803 24592 8812 24632
rect 8852 24592 8861 24632
rect 9867 24632 9909 24641
rect 8803 24591 8861 24592
rect 9291 24613 9333 24622
rect 9291 24573 9292 24613
rect 9332 24573 9333 24613
rect 9291 24564 9333 24573
rect 9387 24613 9429 24622
rect 9387 24573 9388 24613
rect 9428 24573 9429 24613
rect 9867 24592 9868 24632
rect 9908 24592 9909 24632
rect 9867 24583 9909 24592
rect 10339 24632 10397 24633
rect 10339 24592 10348 24632
rect 10388 24592 10397 24632
rect 11395 24632 11453 24633
rect 10339 24591 10397 24592
rect 10827 24618 10869 24627
rect 9387 24564 9429 24573
rect 10827 24578 10828 24618
rect 10868 24578 10869 24618
rect 11395 24592 11404 24632
rect 11444 24592 11453 24632
rect 11395 24591 11453 24592
rect 12643 24632 12701 24633
rect 12643 24592 12652 24632
rect 12692 24592 12701 24632
rect 12643 24591 12701 24592
rect 13123 24632 13181 24633
rect 13123 24592 13132 24632
rect 13172 24592 13181 24632
rect 13123 24591 13181 24592
rect 14371 24632 14429 24633
rect 14371 24592 14380 24632
rect 14420 24592 14429 24632
rect 14371 24591 14429 24592
rect 15331 24632 15389 24633
rect 15331 24592 15340 24632
rect 15380 24592 15389 24632
rect 15331 24591 15389 24592
rect 16579 24632 16637 24633
rect 16579 24592 16588 24632
rect 16628 24592 16637 24632
rect 16579 24591 16637 24592
rect 16971 24632 17013 24641
rect 16971 24592 16972 24632
rect 17012 24592 17013 24632
rect 16971 24583 17013 24592
rect 17067 24632 17109 24641
rect 17067 24592 17068 24632
rect 17108 24592 17109 24632
rect 17067 24583 17109 24592
rect 17163 24632 17205 24641
rect 17163 24592 17164 24632
rect 17204 24592 17205 24632
rect 17163 24583 17205 24592
rect 17259 24632 17301 24641
rect 17259 24592 17260 24632
rect 17300 24592 17301 24632
rect 17259 24583 17301 24592
rect 18211 24632 18269 24633
rect 18211 24592 18220 24632
rect 18260 24592 18269 24632
rect 18211 24591 18269 24592
rect 19459 24632 19517 24633
rect 19459 24592 19468 24632
rect 19508 24592 19517 24632
rect 19459 24591 19517 24592
rect 10827 24569 10869 24578
rect 9771 24548 9813 24557
rect 9771 24508 9772 24548
rect 9812 24508 9813 24548
rect 9771 24499 9813 24508
rect 7363 24464 7421 24465
rect 7363 24424 7372 24464
rect 7412 24424 7421 24464
rect 7363 24423 7421 24424
rect 11211 24380 11253 24389
rect 11211 24340 11212 24380
rect 11252 24340 11253 24380
rect 11211 24331 11253 24340
rect 14571 24380 14613 24389
rect 14571 24340 14572 24380
rect 14612 24340 14613 24380
rect 14571 24331 14613 24340
rect 18027 24380 18069 24389
rect 18027 24340 18028 24380
rect 18068 24340 18069 24380
rect 18027 24331 18069 24340
rect 1152 24212 20352 24236
rect 1152 24172 3688 24212
rect 3728 24172 3770 24212
rect 3810 24172 3852 24212
rect 3892 24172 3934 24212
rect 3974 24172 4016 24212
rect 4056 24172 18808 24212
rect 18848 24172 18890 24212
rect 18930 24172 18972 24212
rect 19012 24172 19054 24212
rect 19094 24172 19136 24212
rect 19176 24172 20352 24212
rect 1152 24148 20352 24172
rect 1227 24044 1269 24053
rect 1227 24004 1228 24044
rect 1268 24004 1269 24044
rect 1227 23995 1269 24004
rect 3811 24044 3869 24045
rect 3811 24004 3820 24044
rect 3860 24004 3869 24044
rect 3811 24003 3869 24004
rect 10923 24044 10965 24053
rect 10923 24004 10924 24044
rect 10964 24004 10965 24044
rect 10923 23995 10965 24004
rect 12363 24044 12405 24053
rect 12363 24004 12364 24044
rect 12404 24004 12405 24044
rect 12363 23995 12405 24004
rect 15627 24044 15669 24053
rect 15627 24004 15628 24044
rect 15668 24004 15669 24044
rect 15627 23995 15669 24004
rect 8419 23960 8477 23961
rect 8419 23920 8428 23960
rect 8468 23920 8477 23960
rect 8419 23919 8477 23920
rect 9099 23960 9141 23969
rect 9099 23920 9100 23960
rect 9140 23920 9141 23960
rect 9099 23911 9141 23920
rect 11691 23960 11733 23969
rect 11691 23920 11692 23960
rect 11732 23920 11733 23960
rect 11691 23911 11733 23920
rect 6219 23876 6261 23885
rect 6219 23836 6220 23876
rect 6260 23836 6261 23876
rect 6219 23827 6261 23836
rect 6315 23876 6357 23885
rect 6315 23836 6316 23876
rect 6356 23836 6357 23876
rect 6315 23827 6357 23836
rect 16491 23876 16533 23885
rect 16491 23836 16492 23876
rect 16532 23836 16533 23876
rect 16491 23827 16533 23836
rect 7275 23806 7317 23815
rect 1411 23792 1469 23793
rect 1411 23752 1420 23792
rect 1460 23752 1469 23792
rect 1411 23751 1469 23752
rect 2659 23792 2717 23793
rect 2659 23752 2668 23792
rect 2708 23752 2717 23792
rect 2659 23751 2717 23752
rect 3139 23792 3197 23793
rect 3139 23752 3148 23792
rect 3188 23752 3197 23792
rect 3139 23751 3197 23752
rect 3435 23792 3477 23801
rect 3435 23752 3436 23792
rect 3476 23752 3477 23792
rect 3435 23743 3477 23752
rect 4003 23792 4061 23793
rect 4003 23752 4012 23792
rect 4052 23752 4061 23792
rect 4003 23751 4061 23752
rect 5251 23792 5309 23793
rect 5251 23752 5260 23792
rect 5300 23752 5309 23792
rect 5251 23751 5309 23752
rect 5739 23792 5781 23801
rect 5739 23752 5740 23792
rect 5780 23752 5781 23792
rect 5739 23743 5781 23752
rect 5835 23792 5877 23801
rect 5835 23752 5836 23792
rect 5876 23752 5877 23792
rect 5835 23743 5877 23752
rect 6787 23792 6845 23793
rect 6787 23752 6796 23792
rect 6836 23752 6845 23792
rect 7275 23766 7276 23806
rect 7316 23766 7317 23806
rect 7275 23757 7317 23766
rect 7747 23792 7805 23793
rect 6787 23751 6845 23752
rect 7747 23752 7756 23792
rect 7796 23752 7805 23792
rect 7747 23751 7805 23752
rect 8043 23792 8085 23801
rect 8043 23752 8044 23792
rect 8084 23752 8085 23792
rect 8043 23743 8085 23752
rect 8611 23792 8669 23793
rect 8611 23752 8620 23792
rect 8660 23752 8669 23792
rect 8611 23751 8669 23752
rect 8715 23792 8757 23801
rect 8715 23752 8716 23792
rect 8756 23752 8757 23792
rect 8715 23743 8757 23752
rect 8907 23792 8949 23801
rect 8907 23752 8908 23792
rect 8948 23752 8949 23792
rect 8907 23743 8949 23752
rect 9099 23792 9141 23801
rect 9099 23752 9100 23792
rect 9140 23752 9141 23792
rect 9099 23743 9141 23752
rect 9291 23792 9333 23801
rect 9291 23752 9292 23792
rect 9332 23752 9333 23792
rect 9291 23743 9333 23752
rect 9475 23792 9533 23793
rect 9475 23752 9484 23792
rect 9524 23752 9533 23792
rect 9475 23751 9533 23752
rect 10723 23792 10781 23793
rect 10723 23752 10732 23792
rect 10772 23752 10781 23792
rect 10723 23751 10781 23752
rect 11499 23792 11541 23801
rect 11499 23752 11500 23792
rect 11540 23752 11541 23792
rect 11499 23743 11541 23752
rect 11691 23792 11733 23801
rect 11691 23752 11692 23792
rect 11732 23752 11733 23792
rect 11691 23743 11733 23752
rect 11883 23792 11925 23801
rect 11883 23752 11884 23792
rect 11924 23752 11925 23792
rect 11883 23743 11925 23752
rect 12075 23792 12117 23801
rect 12075 23752 12076 23792
rect 12116 23752 12117 23792
rect 12075 23743 12117 23752
rect 12171 23792 12213 23801
rect 12171 23752 12172 23792
rect 12212 23752 12213 23792
rect 12171 23743 12213 23752
rect 12363 23792 12405 23801
rect 12363 23752 12364 23792
rect 12404 23752 12405 23792
rect 12363 23743 12405 23752
rect 12555 23792 12597 23801
rect 12555 23752 12556 23792
rect 12596 23752 12597 23792
rect 12555 23743 12597 23752
rect 12643 23792 12701 23793
rect 12643 23752 12652 23792
rect 12692 23752 12701 23792
rect 12643 23751 12701 23752
rect 13035 23792 13077 23801
rect 13035 23752 13036 23792
rect 13076 23752 13077 23792
rect 13035 23743 13077 23752
rect 13131 23792 13173 23801
rect 13131 23752 13132 23792
rect 13172 23752 13173 23792
rect 13131 23743 13173 23752
rect 13515 23792 13557 23801
rect 13515 23752 13516 23792
rect 13556 23752 13557 23792
rect 13515 23743 13557 23752
rect 13611 23792 13653 23801
rect 13611 23752 13612 23792
rect 13652 23752 13653 23792
rect 13611 23743 13653 23752
rect 13995 23792 14037 23801
rect 13995 23752 13996 23792
rect 14036 23752 14037 23792
rect 13995 23743 14037 23752
rect 14091 23792 14133 23801
rect 15051 23797 15093 23806
rect 14091 23752 14092 23792
rect 14132 23752 14133 23792
rect 14091 23743 14133 23752
rect 14563 23792 14621 23793
rect 14563 23752 14572 23792
rect 14612 23752 14621 23792
rect 14563 23751 14621 23752
rect 15051 23757 15052 23797
rect 15092 23757 15093 23797
rect 15915 23792 15957 23801
rect 15051 23748 15093 23757
rect 15523 23781 15581 23782
rect 15523 23741 15532 23781
rect 15572 23741 15581 23781
rect 15915 23752 15916 23792
rect 15956 23752 15957 23792
rect 15915 23743 15957 23752
rect 16011 23792 16053 23801
rect 16011 23752 16012 23792
rect 16052 23752 16053 23792
rect 16011 23743 16053 23752
rect 16395 23792 16437 23801
rect 17451 23797 17493 23806
rect 16395 23752 16396 23792
rect 16436 23752 16437 23792
rect 16395 23743 16437 23752
rect 16963 23792 17021 23793
rect 16963 23752 16972 23792
rect 17012 23752 17021 23792
rect 16963 23751 17021 23752
rect 17451 23757 17452 23797
rect 17492 23757 17493 23797
rect 17451 23748 17493 23757
rect 18115 23792 18173 23793
rect 18115 23752 18124 23792
rect 18164 23752 18173 23792
rect 18115 23751 18173 23752
rect 19363 23792 19421 23793
rect 19363 23752 19372 23792
rect 19412 23752 19421 23792
rect 19363 23751 19421 23752
rect 19755 23792 19797 23801
rect 19755 23752 19756 23792
rect 19796 23752 19797 23792
rect 19755 23743 19797 23752
rect 19851 23792 19893 23801
rect 19851 23752 19852 23792
rect 19892 23752 19893 23792
rect 19851 23743 19893 23752
rect 15523 23740 15581 23741
rect 3531 23708 3573 23717
rect 3531 23668 3532 23708
rect 3572 23668 3573 23708
rect 3531 23659 3573 23668
rect 5451 23708 5493 23717
rect 5451 23668 5452 23708
rect 5492 23668 5493 23708
rect 5451 23659 5493 23668
rect 7467 23708 7509 23717
rect 7467 23668 7468 23708
rect 7508 23668 7509 23708
rect 7467 23659 7509 23668
rect 8139 23708 8181 23717
rect 8139 23668 8140 23708
rect 8180 23668 8181 23708
rect 8139 23659 8181 23668
rect 15243 23708 15285 23717
rect 15243 23668 15244 23708
rect 15284 23668 15285 23708
rect 15243 23659 15285 23668
rect 17643 23708 17685 23717
rect 17643 23668 17644 23708
rect 17684 23668 17685 23708
rect 17643 23659 17685 23668
rect 8803 23624 8861 23625
rect 8803 23584 8812 23624
rect 8852 23584 8861 23624
rect 8803 23583 8861 23584
rect 12835 23624 12893 23625
rect 12835 23584 12844 23624
rect 12884 23584 12893 23624
rect 12835 23583 12893 23584
rect 19563 23624 19605 23633
rect 19563 23584 19564 23624
rect 19604 23584 19605 23624
rect 19563 23575 19605 23584
rect 20035 23624 20093 23625
rect 20035 23584 20044 23624
rect 20084 23584 20093 23624
rect 20035 23583 20093 23584
rect 1152 23456 20452 23480
rect 1152 23416 4928 23456
rect 4968 23416 5010 23456
rect 5050 23416 5092 23456
rect 5132 23416 5174 23456
rect 5214 23416 5256 23456
rect 5296 23416 20048 23456
rect 20088 23416 20130 23456
rect 20170 23416 20212 23456
rect 20252 23416 20294 23456
rect 20334 23416 20376 23456
rect 20416 23416 20452 23456
rect 1152 23392 20452 23416
rect 3723 23288 3765 23297
rect 3723 23248 3724 23288
rect 3764 23248 3765 23288
rect 3723 23239 3765 23248
rect 7083 23288 7125 23297
rect 7083 23248 7084 23288
rect 7124 23248 7125 23288
rect 7083 23239 7125 23248
rect 11691 23288 11733 23297
rect 11691 23248 11692 23288
rect 11732 23248 11733 23288
rect 11691 23239 11733 23248
rect 15435 23288 15477 23297
rect 15435 23248 15436 23288
rect 15476 23248 15477 23288
rect 15435 23239 15477 23248
rect 18219 23288 18261 23297
rect 18219 23248 18220 23288
rect 18260 23248 18261 23288
rect 18219 23239 18261 23248
rect 19459 23288 19517 23289
rect 19459 23248 19468 23288
rect 19508 23248 19517 23288
rect 19459 23247 19517 23248
rect 19939 23288 19997 23289
rect 19939 23248 19948 23288
rect 19988 23248 19997 23288
rect 19939 23247 19997 23248
rect 8715 23204 8757 23213
rect 8715 23164 8716 23204
rect 8756 23164 8757 23204
rect 8715 23155 8757 23164
rect 11499 23204 11541 23213
rect 11499 23164 11500 23204
rect 11540 23164 11541 23204
rect 11499 23155 11541 23164
rect 16011 23147 16053 23156
rect 1419 23120 1461 23129
rect 1419 23080 1420 23120
rect 1460 23080 1461 23120
rect 1419 23071 1461 23080
rect 1707 23120 1749 23129
rect 1707 23080 1708 23120
rect 1748 23080 1749 23120
rect 1707 23071 1749 23080
rect 1995 23120 2037 23129
rect 1995 23080 1996 23120
rect 2036 23080 2037 23120
rect 1995 23071 2037 23080
rect 2091 23120 2133 23129
rect 2091 23080 2092 23120
rect 2132 23080 2133 23120
rect 2091 23071 2133 23080
rect 2475 23120 2517 23129
rect 2475 23080 2476 23120
rect 2516 23080 2517 23120
rect 2475 23071 2517 23080
rect 2571 23120 2613 23129
rect 2571 23080 2572 23120
rect 2612 23080 2613 23120
rect 2571 23071 2613 23080
rect 3043 23120 3101 23121
rect 3043 23080 3052 23120
rect 3092 23080 3101 23120
rect 3907 23120 3965 23121
rect 3043 23079 3101 23080
rect 3531 23106 3573 23115
rect 3531 23066 3532 23106
rect 3572 23066 3573 23106
rect 3907 23080 3916 23120
rect 3956 23080 3965 23120
rect 3907 23079 3965 23080
rect 5155 23120 5213 23121
rect 5155 23080 5164 23120
rect 5204 23080 5213 23120
rect 5155 23079 5213 23080
rect 5635 23120 5693 23121
rect 5635 23080 5644 23120
rect 5684 23080 5693 23120
rect 5635 23079 5693 23080
rect 6883 23120 6941 23121
rect 6883 23080 6892 23120
rect 6932 23080 6941 23120
rect 6883 23079 6941 23080
rect 7267 23120 7325 23121
rect 7267 23080 7276 23120
rect 7316 23080 7325 23120
rect 7267 23079 7325 23080
rect 8515 23120 8573 23121
rect 8515 23080 8524 23120
rect 8564 23080 8573 23120
rect 8515 23079 8573 23080
rect 8995 23120 9053 23121
rect 8995 23080 9004 23120
rect 9044 23080 9053 23120
rect 8995 23079 9053 23080
rect 10051 23120 10109 23121
rect 10051 23080 10060 23120
rect 10100 23080 10109 23120
rect 10051 23079 10109 23080
rect 11299 23120 11357 23121
rect 11299 23080 11308 23120
rect 11348 23080 11357 23120
rect 12355 23120 12413 23121
rect 11299 23079 11357 23080
rect 11883 23106 11925 23115
rect 3531 23057 3573 23066
rect 11883 23066 11884 23106
rect 11924 23066 11925 23106
rect 12355 23080 12364 23120
rect 12404 23080 12413 23120
rect 12355 23079 12413 23080
rect 12843 23120 12885 23129
rect 12843 23080 12844 23120
rect 12884 23080 12885 23120
rect 12843 23071 12885 23080
rect 13323 23120 13365 23129
rect 13323 23080 13324 23120
rect 13364 23080 13365 23120
rect 13323 23071 13365 23080
rect 13419 23120 13461 23129
rect 13419 23080 13420 23120
rect 13460 23080 13461 23120
rect 13419 23071 13461 23080
rect 13987 23120 14045 23121
rect 13987 23080 13996 23120
rect 14036 23080 14045 23120
rect 13987 23079 14045 23080
rect 15235 23120 15293 23121
rect 15235 23080 15244 23120
rect 15284 23080 15293 23120
rect 15235 23079 15293 23080
rect 15715 23120 15773 23121
rect 15715 23080 15724 23120
rect 15764 23080 15773 23120
rect 16011 23107 16012 23147
rect 16052 23107 16053 23147
rect 16011 23098 16053 23107
rect 16771 23120 16829 23121
rect 15715 23079 15773 23080
rect 16771 23080 16780 23120
rect 16820 23080 16829 23120
rect 16771 23079 16829 23080
rect 18019 23120 18077 23121
rect 18019 23080 18028 23120
rect 18068 23080 18077 23120
rect 18019 23079 18077 23080
rect 18411 23120 18453 23129
rect 18411 23080 18412 23120
rect 18452 23080 18453 23120
rect 16099 23078 16157 23079
rect 11883 23057 11925 23066
rect 12939 23036 12981 23045
rect 16099 23038 16108 23078
rect 16148 23038 16157 23078
rect 18411 23071 18453 23080
rect 18507 23120 18549 23129
rect 18507 23080 18508 23120
rect 18548 23080 18549 23120
rect 18507 23071 18549 23080
rect 18603 23120 18645 23129
rect 18603 23080 18604 23120
rect 18644 23080 18645 23120
rect 18603 23071 18645 23080
rect 18699 23120 18741 23129
rect 18699 23080 18700 23120
rect 18740 23080 18741 23120
rect 18699 23071 18741 23080
rect 19179 23120 19221 23129
rect 19179 23080 19180 23120
rect 19220 23080 19221 23120
rect 19179 23071 19221 23080
rect 19275 23120 19317 23129
rect 19275 23080 19276 23120
rect 19316 23080 19317 23120
rect 19275 23071 19317 23080
rect 19659 23120 19701 23129
rect 19659 23080 19660 23120
rect 19700 23080 19701 23120
rect 19659 23071 19701 23080
rect 19755 23120 19797 23129
rect 19755 23080 19756 23120
rect 19796 23080 19797 23120
rect 19755 23071 19797 23080
rect 19851 23120 19893 23129
rect 19851 23080 19852 23120
rect 19892 23080 19893 23120
rect 19851 23071 19893 23080
rect 16099 23037 16157 23038
rect 12939 22996 12940 23036
rect 12980 22996 12981 23036
rect 12939 22987 12981 22996
rect 16387 22952 16445 22953
rect 16387 22912 16396 22952
rect 16436 22912 16445 22952
rect 16387 22911 16445 22912
rect 1707 22868 1749 22877
rect 1707 22828 1708 22868
rect 1748 22828 1749 22868
rect 1707 22819 1749 22828
rect 5355 22868 5397 22877
rect 5355 22828 5356 22868
rect 5396 22828 5397 22868
rect 5355 22819 5397 22828
rect 7083 22868 7125 22877
rect 7083 22828 7084 22868
rect 7124 22828 7125 22868
rect 7083 22819 7125 22828
rect 8907 22868 8949 22877
rect 8907 22828 8908 22868
rect 8948 22828 8949 22868
rect 8907 22819 8949 22828
rect 1152 22700 20352 22724
rect 1152 22660 3688 22700
rect 3728 22660 3770 22700
rect 3810 22660 3852 22700
rect 3892 22660 3934 22700
rect 3974 22660 4016 22700
rect 4056 22660 18808 22700
rect 18848 22660 18890 22700
rect 18930 22660 18972 22700
rect 19012 22660 19054 22700
rect 19094 22660 19136 22700
rect 19176 22660 20352 22700
rect 1152 22636 20352 22660
rect 2667 22532 2709 22541
rect 2667 22492 2668 22532
rect 2708 22492 2709 22532
rect 2667 22483 2709 22492
rect 2859 22532 2901 22541
rect 2859 22492 2860 22532
rect 2900 22492 2901 22532
rect 2859 22483 2901 22492
rect 8331 22532 8373 22541
rect 8331 22492 8332 22532
rect 8372 22492 8373 22532
rect 8331 22483 8373 22492
rect 12835 22532 12893 22533
rect 12835 22492 12844 22532
rect 12884 22492 12893 22532
rect 12835 22491 12893 22492
rect 6115 22448 6173 22449
rect 6115 22408 6124 22448
rect 6164 22408 6173 22448
rect 6115 22407 6173 22408
rect 1219 22280 1277 22281
rect 1219 22240 1228 22280
rect 1268 22240 1277 22280
rect 1219 22239 1277 22240
rect 2467 22280 2525 22281
rect 2467 22240 2476 22280
rect 2516 22240 2525 22280
rect 2467 22239 2525 22240
rect 3043 22280 3101 22281
rect 3043 22240 3052 22280
rect 3092 22240 3101 22280
rect 3043 22239 3101 22240
rect 4291 22280 4349 22281
rect 4291 22240 4300 22280
rect 4340 22240 4349 22280
rect 4291 22239 4349 22240
rect 4483 22280 4541 22281
rect 4483 22240 4492 22280
rect 4532 22240 4541 22280
rect 4483 22239 4541 22240
rect 5731 22280 5789 22281
rect 5731 22240 5740 22280
rect 5780 22240 5789 22280
rect 5731 22239 5789 22240
rect 6123 22280 6165 22289
rect 6123 22240 6124 22280
rect 6164 22240 6165 22280
rect 6123 22231 6165 22240
rect 6219 22280 6261 22289
rect 6219 22240 6220 22280
rect 6260 22240 6261 22280
rect 6219 22231 6261 22240
rect 6411 22280 6453 22289
rect 6411 22240 6412 22280
rect 6452 22240 6453 22280
rect 6411 22231 6453 22240
rect 6603 22280 6645 22289
rect 6603 22240 6604 22280
rect 6644 22240 6645 22280
rect 6603 22231 6645 22240
rect 6795 22280 6837 22289
rect 6795 22240 6796 22280
rect 6836 22240 6837 22280
rect 6795 22231 6837 22240
rect 8035 22280 8093 22281
rect 8035 22240 8044 22280
rect 8084 22240 8093 22280
rect 8035 22239 8093 22240
rect 8139 22280 8181 22289
rect 8139 22240 8140 22280
rect 8180 22240 8181 22280
rect 8139 22231 8181 22240
rect 8331 22280 8373 22289
rect 8331 22240 8332 22280
rect 8372 22240 8373 22280
rect 8331 22231 8373 22240
rect 11595 22280 11637 22289
rect 11595 22240 11596 22280
rect 11636 22240 11637 22280
rect 11595 22231 11637 22240
rect 11691 22280 11733 22289
rect 11691 22240 11692 22280
rect 11732 22240 11733 22280
rect 11691 22231 11733 22240
rect 11787 22280 11829 22289
rect 11787 22240 11788 22280
rect 11828 22240 11829 22280
rect 11787 22231 11829 22240
rect 11883 22280 11925 22289
rect 11883 22240 11884 22280
rect 11924 22240 11925 22280
rect 11883 22231 11925 22240
rect 12163 22280 12221 22281
rect 12163 22240 12172 22280
rect 12212 22240 12221 22280
rect 12163 22239 12221 22240
rect 12459 22280 12501 22289
rect 12459 22240 12460 22280
rect 12500 22240 12501 22280
rect 12459 22231 12501 22240
rect 13035 22280 13077 22289
rect 13035 22240 13036 22280
rect 13076 22240 13077 22280
rect 13035 22231 13077 22240
rect 13227 22280 13269 22289
rect 13227 22240 13228 22280
rect 13268 22240 13269 22280
rect 13227 22231 13269 22240
rect 13315 22280 13373 22281
rect 13315 22240 13324 22280
rect 13364 22240 13373 22280
rect 13315 22239 13373 22240
rect 13699 22280 13757 22281
rect 13699 22240 13708 22280
rect 13748 22240 13757 22280
rect 13699 22239 13757 22240
rect 14947 22280 15005 22281
rect 14947 22240 14956 22280
rect 14996 22240 15005 22280
rect 14947 22239 15005 22240
rect 16963 22280 17021 22281
rect 16963 22240 16972 22280
rect 17012 22240 17021 22280
rect 16963 22239 17021 22240
rect 17451 22280 17493 22289
rect 17451 22240 17452 22280
rect 17492 22240 17493 22280
rect 17451 22231 17493 22240
rect 17547 22280 17589 22289
rect 17547 22240 17548 22280
rect 17588 22240 17589 22280
rect 17547 22231 17589 22240
rect 6699 22196 6741 22205
rect 6699 22156 6700 22196
rect 6740 22156 6741 22196
rect 6699 22147 6741 22156
rect 12555 22196 12597 22205
rect 12555 22156 12556 22196
rect 12596 22156 12597 22196
rect 12555 22147 12597 22156
rect 13131 22196 13173 22205
rect 13131 22156 13132 22196
rect 13172 22156 13173 22196
rect 13131 22147 13173 22156
rect 5931 22112 5973 22121
rect 5931 22072 5932 22112
rect 5972 22072 5973 22112
rect 5931 22063 5973 22072
rect 15147 22112 15189 22121
rect 15147 22072 15148 22112
rect 15188 22072 15189 22112
rect 15147 22063 15189 22072
rect 17067 22112 17109 22121
rect 17067 22072 17068 22112
rect 17108 22072 17109 22112
rect 17067 22063 17109 22072
rect 17731 22112 17789 22113
rect 17731 22072 17740 22112
rect 17780 22072 17789 22112
rect 17731 22071 17789 22072
rect 1152 21944 20452 21968
rect 1152 21904 4928 21944
rect 4968 21904 5010 21944
rect 5050 21904 5092 21944
rect 5132 21904 5174 21944
rect 5214 21904 5256 21944
rect 5296 21904 20048 21944
rect 20088 21904 20130 21944
rect 20170 21904 20212 21944
rect 20252 21904 20294 21944
rect 20334 21904 20376 21944
rect 20416 21904 20452 21944
rect 1152 21880 20452 21904
rect 3147 21776 3189 21785
rect 3147 21736 3148 21776
rect 3188 21736 3189 21776
rect 3147 21727 3189 21736
rect 6979 21776 7037 21777
rect 6979 21736 6988 21776
rect 7028 21736 7037 21776
rect 6979 21735 7037 21736
rect 12843 21776 12885 21785
rect 12843 21736 12844 21776
rect 12884 21736 12885 21776
rect 12843 21727 12885 21736
rect 15243 21776 15285 21785
rect 15243 21736 15244 21776
rect 15284 21736 15285 21776
rect 15243 21727 15285 21736
rect 5355 21692 5397 21701
rect 5355 21652 5356 21692
rect 5396 21652 5397 21692
rect 5355 21643 5397 21652
rect 5931 21692 5973 21701
rect 5931 21652 5932 21692
rect 5972 21652 5973 21692
rect 5931 21643 5973 21652
rect 9003 21692 9045 21701
rect 9003 21652 9004 21692
rect 9044 21652 9045 21692
rect 9003 21643 9045 21652
rect 11019 21692 11061 21701
rect 11019 21652 11020 21692
rect 11060 21652 11061 21692
rect 11019 21643 11061 21652
rect 17355 21692 17397 21701
rect 17355 21652 17356 21692
rect 17396 21652 17397 21692
rect 17355 21643 17397 21652
rect 1699 21608 1757 21609
rect 1699 21568 1708 21608
rect 1748 21568 1757 21608
rect 1699 21567 1757 21568
rect 2947 21608 3005 21609
rect 2947 21568 2956 21608
rect 2996 21568 3005 21608
rect 2947 21567 3005 21568
rect 3627 21608 3669 21617
rect 3627 21568 3628 21608
rect 3668 21568 3669 21608
rect 3627 21559 3669 21568
rect 3723 21608 3765 21617
rect 3723 21568 3724 21608
rect 3764 21568 3765 21608
rect 3723 21559 3765 21568
rect 4107 21608 4149 21617
rect 4107 21568 4108 21608
rect 4148 21568 4149 21608
rect 4107 21559 4149 21568
rect 4203 21608 4245 21617
rect 4203 21568 4204 21608
rect 4244 21568 4245 21608
rect 4203 21559 4245 21568
rect 4675 21608 4733 21609
rect 4675 21568 4684 21608
rect 4724 21568 4733 21608
rect 4675 21567 4733 21568
rect 5163 21603 5205 21612
rect 5163 21563 5164 21603
rect 5204 21563 5205 21603
rect 5731 21608 5789 21609
rect 5731 21568 5740 21608
rect 5780 21568 5789 21608
rect 5731 21567 5789 21568
rect 5835 21608 5877 21617
rect 5835 21568 5836 21608
rect 5876 21568 5877 21608
rect 5163 21554 5205 21563
rect 5835 21559 5877 21568
rect 6027 21608 6069 21617
rect 6027 21568 6028 21608
rect 6068 21568 6069 21608
rect 6027 21559 6069 21568
rect 6219 21608 6261 21617
rect 6219 21568 6220 21608
rect 6260 21568 6261 21608
rect 6219 21559 6261 21568
rect 6315 21608 6357 21617
rect 6315 21568 6316 21608
rect 6356 21568 6357 21608
rect 6315 21559 6357 21568
rect 6507 21608 6549 21617
rect 6507 21568 6508 21608
rect 6548 21568 6549 21608
rect 6507 21559 6549 21568
rect 6699 21608 6741 21617
rect 6699 21568 6700 21608
rect 6740 21568 6741 21608
rect 6699 21559 6741 21568
rect 6795 21608 6837 21617
rect 6795 21568 6796 21608
rect 6836 21568 6837 21608
rect 6795 21559 6837 21568
rect 6891 21608 6933 21617
rect 6891 21568 6892 21608
rect 6932 21568 6933 21608
rect 6891 21559 6933 21568
rect 7179 21608 7221 21617
rect 7179 21568 7180 21608
rect 7220 21568 7221 21608
rect 7179 21559 7221 21568
rect 7371 21608 7413 21617
rect 7371 21568 7372 21608
rect 7412 21568 7413 21608
rect 7371 21559 7413 21568
rect 7555 21608 7613 21609
rect 7555 21568 7564 21608
rect 7604 21568 7613 21608
rect 7555 21567 7613 21568
rect 8803 21608 8861 21609
rect 8803 21568 8812 21608
rect 8852 21568 8861 21608
rect 8803 21567 8861 21568
rect 9291 21608 9333 21617
rect 9291 21568 9292 21608
rect 9332 21568 9333 21608
rect 9291 21559 9333 21568
rect 9387 21608 9429 21617
rect 9387 21568 9388 21608
rect 9428 21568 9429 21608
rect 9387 21559 9429 21568
rect 9771 21608 9813 21617
rect 9771 21568 9772 21608
rect 9812 21568 9813 21608
rect 9771 21559 9813 21568
rect 9867 21608 9909 21617
rect 9867 21568 9868 21608
rect 9908 21568 9909 21608
rect 9867 21559 9909 21568
rect 10339 21608 10397 21609
rect 10339 21568 10348 21608
rect 10388 21568 10397 21608
rect 11395 21608 11453 21609
rect 10339 21567 10397 21568
rect 10875 21598 10917 21607
rect 10875 21558 10876 21598
rect 10916 21558 10917 21598
rect 11395 21568 11404 21608
rect 11444 21568 11453 21608
rect 11395 21567 11453 21568
rect 12643 21608 12701 21609
rect 12643 21568 12652 21608
rect 12692 21568 12701 21608
rect 12643 21567 12701 21568
rect 13515 21608 13557 21617
rect 13515 21568 13516 21608
rect 13556 21568 13557 21608
rect 13515 21559 13557 21568
rect 13611 21608 13653 21617
rect 13611 21568 13612 21608
rect 13652 21568 13653 21608
rect 13611 21559 13653 21568
rect 13995 21608 14037 21617
rect 13995 21568 13996 21608
rect 14036 21568 14037 21608
rect 13995 21559 14037 21568
rect 14091 21608 14133 21617
rect 14091 21568 14092 21608
rect 14132 21568 14133 21608
rect 14091 21559 14133 21568
rect 14563 21608 14621 21609
rect 14563 21568 14572 21608
rect 14612 21568 14621 21608
rect 15627 21608 15669 21617
rect 14563 21567 14621 21568
rect 15099 21598 15141 21607
rect 10875 21549 10917 21558
rect 15099 21558 15100 21598
rect 15140 21558 15141 21598
rect 15627 21568 15628 21608
rect 15668 21568 15669 21608
rect 15627 21559 15669 21568
rect 15723 21608 15765 21617
rect 15723 21568 15724 21608
rect 15764 21568 15765 21608
rect 15723 21559 15765 21568
rect 16107 21608 16149 21617
rect 16107 21568 16108 21608
rect 16148 21568 16149 21608
rect 16107 21559 16149 21568
rect 16203 21608 16245 21617
rect 16203 21568 16204 21608
rect 16244 21568 16245 21608
rect 16203 21559 16245 21568
rect 16675 21608 16733 21609
rect 16675 21568 16684 21608
rect 16724 21568 16733 21608
rect 17731 21608 17789 21609
rect 16675 21567 16733 21568
rect 17163 21594 17205 21603
rect 15099 21549 15141 21558
rect 17163 21554 17164 21594
rect 17204 21554 17205 21594
rect 17731 21568 17740 21608
rect 17780 21568 17789 21608
rect 17731 21567 17789 21568
rect 18979 21608 19037 21609
rect 18979 21568 18988 21608
rect 19028 21568 19037 21608
rect 18979 21567 19037 21568
rect 17163 21545 17205 21554
rect 7179 21440 7221 21449
rect 7179 21400 7180 21440
rect 7220 21400 7221 21440
rect 7179 21391 7221 21400
rect 17547 21440 17589 21449
rect 17547 21400 17548 21440
rect 17588 21400 17589 21440
rect 17547 21391 17589 21400
rect 1152 21188 20352 21212
rect 1152 21148 3688 21188
rect 3728 21148 3770 21188
rect 3810 21148 3852 21188
rect 3892 21148 3934 21188
rect 3974 21148 4016 21188
rect 4056 21148 18808 21188
rect 18848 21148 18890 21188
rect 18930 21148 18972 21188
rect 19012 21148 19054 21188
rect 19094 21148 19136 21188
rect 19176 21148 20352 21188
rect 1152 21124 20352 21148
rect 4875 21020 4917 21029
rect 4875 20980 4876 21020
rect 4916 20980 4917 21020
rect 4875 20971 4917 20980
rect 11019 21020 11061 21029
rect 11019 20980 11020 21020
rect 11060 20980 11061 21020
rect 11019 20971 11061 20980
rect 13707 21020 13749 21029
rect 13707 20980 13708 21020
rect 13748 20980 13749 21020
rect 13707 20971 13749 20980
rect 15819 21020 15861 21029
rect 15819 20980 15820 21020
rect 15860 20980 15861 21020
rect 15819 20971 15861 20980
rect 16867 20936 16925 20937
rect 16867 20896 16876 20936
rect 16916 20896 16925 20936
rect 16867 20895 16925 20896
rect 17827 20936 17885 20937
rect 17827 20896 17836 20936
rect 17876 20896 17885 20936
rect 17827 20895 17885 20896
rect 1995 20852 2037 20861
rect 1995 20812 1996 20852
rect 2036 20812 2037 20852
rect 1995 20803 2037 20812
rect 2091 20852 2133 20861
rect 2091 20812 2092 20852
rect 2132 20812 2133 20852
rect 2091 20803 2133 20812
rect 7755 20852 7797 20861
rect 7755 20812 7756 20852
rect 7796 20812 7797 20852
rect 7755 20803 7797 20812
rect 7851 20852 7893 20861
rect 7851 20812 7852 20852
rect 7892 20812 7893 20852
rect 7851 20803 7893 20812
rect 1515 20768 1557 20777
rect 1515 20728 1516 20768
rect 1556 20728 1557 20768
rect 1515 20719 1557 20728
rect 1611 20768 1653 20777
rect 3051 20773 3093 20782
rect 8859 20777 8901 20786
rect 1611 20728 1612 20768
rect 1652 20728 1653 20768
rect 1611 20719 1653 20728
rect 2563 20768 2621 20769
rect 2563 20728 2572 20768
rect 2612 20728 2621 20768
rect 2563 20727 2621 20728
rect 3051 20733 3052 20773
rect 3092 20733 3093 20773
rect 3051 20724 3093 20733
rect 3427 20768 3485 20769
rect 3427 20728 3436 20768
rect 3476 20728 3485 20768
rect 3427 20727 3485 20728
rect 4675 20768 4733 20769
rect 4675 20728 4684 20768
rect 4724 20728 4733 20768
rect 4675 20727 4733 20728
rect 5067 20768 5109 20777
rect 5067 20728 5068 20768
rect 5108 20728 5109 20768
rect 5067 20719 5109 20728
rect 5163 20768 5205 20777
rect 5163 20728 5164 20768
rect 5204 20728 5205 20768
rect 5163 20719 5205 20728
rect 5539 20768 5597 20769
rect 5539 20728 5548 20768
rect 5588 20728 5597 20768
rect 5539 20727 5597 20728
rect 6787 20768 6845 20769
rect 6787 20728 6796 20768
rect 6836 20728 6845 20768
rect 6787 20727 6845 20728
rect 7275 20768 7317 20777
rect 7275 20728 7276 20768
rect 7316 20728 7317 20768
rect 7275 20719 7317 20728
rect 7371 20768 7413 20777
rect 7371 20728 7372 20768
rect 7412 20728 7413 20768
rect 7371 20719 7413 20728
rect 8323 20768 8381 20769
rect 8323 20728 8332 20768
rect 8372 20728 8381 20768
rect 8859 20737 8860 20777
rect 8900 20737 8901 20777
rect 8859 20728 8901 20737
rect 9571 20768 9629 20769
rect 9571 20728 9580 20768
rect 9620 20728 9629 20768
rect 8323 20727 8381 20728
rect 9571 20727 9629 20728
rect 10819 20768 10877 20769
rect 10819 20728 10828 20768
rect 10868 20728 10877 20768
rect 10819 20727 10877 20728
rect 12259 20768 12317 20769
rect 12259 20728 12268 20768
rect 12308 20728 12317 20768
rect 12259 20727 12317 20728
rect 13507 20768 13565 20769
rect 13507 20728 13516 20768
rect 13556 20728 13565 20768
rect 13507 20727 13565 20728
rect 14371 20768 14429 20769
rect 14371 20728 14380 20768
rect 14420 20728 14429 20768
rect 14371 20727 14429 20728
rect 15619 20768 15677 20769
rect 15619 20728 15628 20768
rect 15668 20728 15677 20768
rect 15619 20727 15677 20728
rect 16195 20768 16253 20769
rect 16195 20728 16204 20768
rect 16244 20728 16253 20768
rect 16195 20727 16253 20728
rect 16491 20768 16533 20777
rect 16491 20728 16492 20768
rect 16532 20728 16533 20768
rect 16491 20719 16533 20728
rect 16587 20768 16629 20777
rect 16587 20728 16588 20768
rect 16628 20728 16629 20768
rect 16587 20719 16629 20728
rect 17155 20768 17213 20769
rect 17155 20728 17164 20768
rect 17204 20728 17213 20768
rect 17155 20727 17213 20728
rect 17451 20768 17493 20777
rect 17451 20728 17452 20768
rect 17492 20728 17493 20768
rect 17451 20719 17493 20728
rect 18027 20768 18069 20777
rect 18027 20728 18028 20768
rect 18068 20728 18069 20768
rect 18027 20719 18069 20728
rect 18123 20768 18165 20777
rect 18123 20728 18124 20768
rect 18164 20728 18165 20768
rect 18123 20719 18165 20728
rect 18507 20768 18549 20777
rect 18507 20728 18508 20768
rect 18548 20728 18549 20768
rect 18507 20719 18549 20728
rect 18699 20768 18741 20777
rect 18699 20728 18700 20768
rect 18740 20728 18741 20768
rect 18699 20719 18741 20728
rect 17547 20684 17589 20693
rect 17547 20644 17548 20684
rect 17588 20644 17589 20684
rect 5347 20642 5405 20643
rect 3243 20600 3285 20609
rect 5347 20602 5356 20642
rect 5396 20602 5405 20642
rect 17547 20635 17589 20644
rect 5347 20601 5405 20602
rect 3243 20560 3244 20600
rect 3284 20560 3285 20600
rect 3243 20551 3285 20560
rect 6987 20600 7029 20609
rect 6987 20560 6988 20600
rect 7028 20560 7029 20600
rect 6987 20551 7029 20560
rect 9003 20600 9045 20609
rect 9003 20560 9004 20600
rect 9044 20560 9045 20600
rect 9003 20551 9045 20560
rect 18307 20600 18365 20601
rect 18307 20560 18316 20600
rect 18356 20560 18365 20600
rect 18307 20559 18365 20560
rect 18603 20600 18645 20609
rect 18603 20560 18604 20600
rect 18644 20560 18645 20600
rect 18603 20551 18645 20560
rect 1152 20432 20452 20456
rect 1152 20392 4928 20432
rect 4968 20392 5010 20432
rect 5050 20392 5092 20432
rect 5132 20392 5174 20432
rect 5214 20392 5256 20432
rect 5296 20392 20048 20432
rect 20088 20392 20130 20432
rect 20170 20392 20212 20432
rect 20252 20392 20294 20432
rect 20334 20392 20376 20432
rect 20416 20392 20452 20432
rect 1152 20368 20452 20392
rect 8907 20264 8949 20273
rect 8907 20224 8908 20264
rect 8948 20224 8949 20264
rect 8907 20215 8949 20224
rect 3915 20180 3957 20189
rect 3915 20140 3916 20180
rect 3956 20140 3957 20180
rect 3915 20131 3957 20140
rect 5163 20180 5205 20189
rect 5163 20140 5164 20180
rect 5204 20140 5205 20180
rect 5163 20131 5205 20140
rect 10539 20180 10581 20189
rect 10539 20140 10540 20180
rect 10580 20140 10581 20180
rect 10539 20131 10581 20140
rect 12555 20180 12597 20189
rect 12555 20140 12556 20180
rect 12596 20140 12597 20180
rect 12555 20131 12597 20140
rect 2467 20096 2525 20097
rect 2467 20056 2476 20096
rect 2516 20056 2525 20096
rect 2467 20055 2525 20056
rect 3715 20096 3773 20097
rect 3715 20056 3724 20096
rect 3764 20056 3773 20096
rect 3715 20055 3773 20056
rect 4387 20096 4445 20097
rect 4387 20056 4396 20096
rect 4436 20056 4445 20096
rect 4387 20055 4445 20056
rect 4491 20096 4533 20105
rect 4491 20056 4492 20096
rect 4532 20056 4533 20096
rect 4491 20047 4533 20056
rect 4683 20096 4725 20105
rect 4683 20056 4684 20096
rect 4724 20056 4725 20096
rect 4683 20047 4725 20056
rect 5259 20096 5301 20105
rect 5259 20056 5260 20096
rect 5300 20056 5301 20096
rect 5259 20047 5301 20056
rect 5539 20096 5597 20097
rect 5539 20056 5548 20096
rect 5588 20056 5597 20096
rect 5539 20055 5597 20056
rect 5827 20096 5885 20097
rect 5827 20056 5836 20096
rect 5876 20056 5885 20096
rect 5827 20055 5885 20056
rect 7075 20096 7133 20097
rect 7075 20056 7084 20096
rect 7124 20056 7133 20096
rect 7075 20055 7133 20056
rect 7459 20096 7517 20097
rect 7459 20056 7468 20096
rect 7508 20056 7517 20096
rect 7459 20055 7517 20056
rect 8707 20096 8765 20097
rect 8707 20056 8716 20096
rect 8756 20056 8765 20096
rect 8707 20055 8765 20056
rect 9091 20096 9149 20097
rect 9091 20056 9100 20096
rect 9140 20056 9149 20096
rect 9091 20055 9149 20056
rect 10339 20096 10397 20097
rect 10339 20056 10348 20096
rect 10388 20056 10397 20096
rect 10339 20055 10397 20056
rect 10827 20096 10869 20105
rect 10827 20056 10828 20096
rect 10868 20056 10869 20096
rect 10827 20047 10869 20056
rect 10923 20096 10965 20105
rect 10923 20056 10924 20096
rect 10964 20056 10965 20096
rect 10923 20047 10965 20056
rect 11403 20096 11445 20105
rect 11403 20056 11404 20096
rect 11444 20056 11445 20096
rect 12739 20096 12797 20097
rect 11403 20047 11445 20056
rect 12363 20086 12405 20095
rect 11875 20054 11933 20055
rect 11307 20012 11349 20021
rect 11875 20014 11884 20054
rect 11924 20014 11933 20054
rect 12363 20046 12364 20086
rect 12404 20046 12405 20086
rect 12739 20056 12748 20096
rect 12788 20056 12797 20096
rect 12739 20055 12797 20056
rect 13987 20096 14045 20097
rect 13987 20056 13996 20096
rect 14036 20056 14045 20096
rect 13987 20055 14045 20056
rect 14371 20096 14429 20097
rect 14371 20056 14380 20096
rect 14420 20056 14429 20096
rect 14371 20055 14429 20056
rect 15619 20096 15677 20097
rect 15619 20056 15628 20096
rect 15668 20056 15677 20096
rect 15619 20055 15677 20056
rect 16867 20096 16925 20097
rect 16867 20056 16876 20096
rect 16916 20056 16925 20096
rect 16867 20055 16925 20056
rect 17259 20096 17301 20105
rect 17259 20056 17260 20096
rect 17300 20056 17301 20096
rect 17739 20096 17781 20105
rect 17259 20047 17301 20056
rect 17443 20082 17501 20083
rect 12363 20037 12405 20046
rect 17443 20042 17452 20082
rect 17492 20042 17501 20082
rect 17443 20041 17501 20042
rect 17543 20077 17601 20078
rect 17543 20037 17552 20077
rect 17592 20037 17601 20077
rect 17739 20056 17740 20096
rect 17780 20056 17781 20096
rect 17739 20047 17781 20056
rect 17931 20096 17973 20105
rect 17931 20056 17932 20096
rect 17972 20056 17973 20096
rect 17931 20047 17973 20056
rect 18019 20096 18077 20097
rect 18019 20056 18028 20096
rect 18068 20056 18077 20096
rect 18019 20055 18077 20056
rect 17543 20036 17601 20037
rect 11875 20013 11933 20014
rect 11307 19972 11308 20012
rect 11348 19972 11349 20012
rect 11307 19963 11349 19972
rect 4683 19928 4725 19937
rect 4683 19888 4684 19928
rect 4724 19888 4725 19928
rect 4683 19879 4725 19888
rect 4867 19928 4925 19929
rect 4867 19888 4876 19928
rect 4916 19888 4925 19928
rect 4867 19887 4925 19888
rect 17067 19928 17109 19937
rect 17067 19888 17068 19928
rect 17108 19888 17109 19928
rect 17067 19879 17109 19888
rect 7275 19844 7317 19853
rect 7275 19804 7276 19844
rect 7316 19804 7317 19844
rect 7275 19795 7317 19804
rect 14187 19844 14229 19853
rect 14187 19804 14188 19844
rect 14228 19804 14229 19844
rect 14187 19795 14229 19804
rect 14475 19844 14517 19853
rect 14475 19804 14476 19844
rect 14516 19804 14517 19844
rect 14475 19795 14517 19804
rect 17259 19844 17301 19853
rect 17259 19804 17260 19844
rect 17300 19804 17301 19844
rect 17259 19795 17301 19804
rect 17739 19844 17781 19853
rect 17739 19804 17740 19844
rect 17780 19804 17781 19844
rect 17739 19795 17781 19804
rect 1152 19676 20352 19700
rect 1152 19636 3688 19676
rect 3728 19636 3770 19676
rect 3810 19636 3852 19676
rect 3892 19636 3934 19676
rect 3974 19636 4016 19676
rect 4056 19636 18808 19676
rect 18848 19636 18890 19676
rect 18930 19636 18972 19676
rect 19012 19636 19054 19676
rect 19094 19636 19136 19676
rect 19176 19636 20352 19676
rect 1152 19612 20352 19636
rect 2763 19508 2805 19517
rect 2763 19468 2764 19508
rect 2804 19468 2805 19508
rect 2763 19459 2805 19468
rect 12651 19508 12693 19517
rect 12651 19468 12652 19508
rect 12692 19468 12693 19508
rect 12651 19459 12693 19468
rect 6507 19340 6549 19349
rect 6507 19300 6508 19340
rect 6548 19300 6549 19340
rect 6507 19291 6549 19300
rect 9099 19340 9141 19349
rect 9099 19300 9100 19340
rect 9140 19300 9141 19340
rect 9099 19291 9141 19300
rect 13995 19340 14037 19349
rect 13995 19300 13996 19340
rect 14036 19300 14037 19340
rect 13995 19291 14037 19300
rect 7467 19270 7509 19279
rect 1315 19256 1373 19257
rect 1315 19216 1324 19256
rect 1364 19216 1373 19256
rect 1315 19215 1373 19216
rect 2563 19256 2621 19257
rect 2563 19216 2572 19256
rect 2612 19216 2621 19256
rect 2563 19215 2621 19216
rect 4195 19256 4253 19257
rect 4195 19216 4204 19256
rect 4244 19216 4253 19256
rect 4195 19215 4253 19216
rect 5443 19256 5501 19257
rect 5443 19216 5452 19256
rect 5492 19216 5501 19256
rect 5443 19215 5501 19216
rect 5931 19256 5973 19265
rect 5931 19216 5932 19256
rect 5972 19216 5973 19256
rect 5931 19207 5973 19216
rect 6027 19256 6069 19265
rect 6027 19216 6028 19256
rect 6068 19216 6069 19256
rect 6027 19207 6069 19216
rect 6411 19256 6453 19265
rect 6411 19216 6412 19256
rect 6452 19216 6453 19256
rect 6411 19207 6453 19216
rect 6979 19256 7037 19257
rect 6979 19216 6988 19256
rect 7028 19216 7037 19256
rect 7467 19230 7468 19270
rect 7508 19230 7509 19270
rect 10203 19265 10245 19274
rect 15099 19265 15141 19274
rect 7467 19221 7509 19230
rect 8619 19256 8661 19265
rect 6979 19215 7037 19216
rect 8619 19216 8620 19256
rect 8660 19216 8661 19256
rect 8619 19207 8661 19216
rect 8715 19256 8757 19265
rect 8715 19216 8716 19256
rect 8756 19216 8757 19256
rect 8715 19207 8757 19216
rect 9195 19256 9237 19265
rect 9195 19216 9196 19256
rect 9236 19216 9237 19256
rect 9195 19207 9237 19216
rect 9667 19256 9725 19257
rect 9667 19216 9676 19256
rect 9716 19216 9725 19256
rect 10203 19225 10204 19265
rect 10244 19225 10245 19265
rect 10203 19216 10245 19225
rect 11203 19256 11261 19257
rect 11203 19216 11212 19256
rect 11252 19216 11261 19256
rect 9667 19215 9725 19216
rect 11203 19215 11261 19216
rect 12451 19256 12509 19257
rect 12451 19216 12460 19256
rect 12500 19216 12509 19256
rect 12451 19215 12509 19216
rect 13515 19256 13557 19265
rect 13515 19216 13516 19256
rect 13556 19216 13557 19256
rect 13515 19207 13557 19216
rect 13611 19256 13653 19265
rect 13611 19216 13612 19256
rect 13652 19216 13653 19256
rect 13611 19207 13653 19216
rect 14091 19256 14133 19265
rect 14091 19216 14092 19256
rect 14132 19216 14133 19256
rect 14091 19207 14133 19216
rect 14563 19256 14621 19257
rect 14563 19216 14572 19256
rect 14612 19216 14621 19256
rect 15099 19225 15100 19265
rect 15140 19225 15141 19265
rect 15099 19216 15141 19225
rect 17443 19256 17501 19257
rect 17443 19216 17452 19256
rect 17492 19216 17501 19256
rect 14563 19215 14621 19216
rect 17443 19215 17501 19216
rect 18691 19256 18749 19257
rect 18691 19216 18700 19256
rect 18740 19216 18749 19256
rect 18691 19215 18749 19216
rect 5643 19088 5685 19097
rect 5643 19048 5644 19088
rect 5684 19048 5685 19088
rect 5643 19039 5685 19048
rect 7659 19088 7701 19097
rect 7659 19048 7660 19088
rect 7700 19048 7701 19088
rect 7659 19039 7701 19048
rect 10347 19088 10389 19097
rect 10347 19048 10348 19088
rect 10388 19048 10389 19088
rect 10347 19039 10389 19048
rect 15243 19088 15285 19097
rect 15243 19048 15244 19088
rect 15284 19048 15285 19088
rect 15243 19039 15285 19048
rect 18891 19088 18933 19097
rect 18891 19048 18892 19088
rect 18932 19048 18933 19088
rect 18891 19039 18933 19048
rect 1152 18920 20452 18944
rect 1152 18880 4928 18920
rect 4968 18880 5010 18920
rect 5050 18880 5092 18920
rect 5132 18880 5174 18920
rect 5214 18880 5256 18920
rect 5296 18880 20048 18920
rect 20088 18880 20130 18920
rect 20170 18880 20212 18920
rect 20252 18880 20294 18920
rect 20334 18880 20376 18920
rect 20416 18880 20452 18920
rect 1152 18856 20452 18880
rect 2667 18752 2709 18761
rect 2667 18712 2668 18752
rect 2708 18712 2709 18752
rect 2667 18703 2709 18712
rect 3139 18752 3197 18753
rect 3139 18712 3148 18752
rect 3188 18712 3197 18752
rect 3139 18711 3197 18712
rect 15243 18752 15285 18761
rect 15243 18712 15244 18752
rect 15284 18712 15285 18752
rect 15243 18703 15285 18712
rect 15715 18752 15773 18753
rect 15715 18712 15724 18752
rect 15764 18712 15773 18752
rect 15715 18711 15773 18712
rect 7755 18668 7797 18677
rect 7755 18628 7756 18668
rect 7796 18628 7797 18668
rect 7755 18619 7797 18628
rect 10731 18668 10773 18677
rect 10731 18628 10732 18668
rect 10772 18628 10773 18668
rect 10731 18619 10773 18628
rect 12747 18668 12789 18677
rect 12747 18628 12748 18668
rect 12788 18628 12789 18668
rect 12747 18619 12789 18628
rect 18699 18668 18741 18677
rect 18699 18628 18700 18668
rect 18740 18628 18741 18668
rect 18699 18619 18741 18628
rect 1219 18584 1277 18585
rect 1219 18544 1228 18584
rect 1268 18544 1277 18584
rect 1219 18543 1277 18544
rect 2467 18584 2525 18585
rect 2467 18544 2476 18584
rect 2516 18544 2525 18584
rect 2467 18543 2525 18544
rect 2859 18584 2901 18593
rect 2859 18544 2860 18584
rect 2900 18544 2901 18584
rect 2859 18535 2901 18544
rect 2955 18584 2997 18593
rect 2955 18544 2956 18584
rect 2996 18544 2997 18584
rect 2955 18535 2997 18544
rect 4291 18584 4349 18585
rect 4291 18544 4300 18584
rect 4340 18544 4349 18584
rect 4291 18543 4349 18544
rect 5539 18584 5597 18585
rect 5539 18544 5548 18584
rect 5588 18544 5597 18584
rect 5539 18543 5597 18544
rect 6027 18584 6069 18593
rect 6027 18544 6028 18584
rect 6068 18544 6069 18584
rect 6027 18535 6069 18544
rect 6123 18584 6165 18593
rect 6123 18544 6124 18584
rect 6164 18544 6165 18584
rect 6123 18535 6165 18544
rect 6507 18584 6549 18593
rect 6507 18544 6508 18584
rect 6548 18544 6549 18584
rect 6507 18535 6549 18544
rect 6603 18584 6645 18593
rect 6603 18544 6604 18584
rect 6644 18544 6645 18584
rect 6603 18535 6645 18544
rect 7075 18584 7133 18585
rect 7075 18544 7084 18584
rect 7124 18544 7133 18584
rect 9283 18584 9341 18585
rect 7075 18543 7133 18544
rect 7563 18570 7605 18579
rect 7563 18530 7564 18570
rect 7604 18530 7605 18570
rect 9283 18544 9292 18584
rect 9332 18544 9341 18584
rect 9283 18543 9341 18544
rect 10531 18584 10589 18585
rect 10531 18544 10540 18584
rect 10580 18544 10589 18584
rect 10531 18543 10589 18544
rect 11019 18584 11061 18593
rect 11019 18544 11020 18584
rect 11060 18544 11061 18584
rect 11019 18535 11061 18544
rect 11115 18584 11157 18593
rect 11115 18544 11116 18584
rect 11156 18544 11157 18584
rect 11115 18535 11157 18544
rect 11499 18584 11541 18593
rect 11499 18544 11500 18584
rect 11540 18544 11541 18584
rect 11499 18535 11541 18544
rect 12067 18584 12125 18585
rect 12067 18544 12076 18584
rect 12116 18544 12125 18584
rect 13795 18584 13853 18585
rect 12067 18543 12125 18544
rect 12555 18570 12597 18579
rect 7563 18521 7605 18530
rect 12555 18530 12556 18570
rect 12596 18530 12597 18570
rect 13795 18544 13804 18584
rect 13844 18544 13853 18584
rect 13795 18543 13853 18544
rect 15043 18584 15101 18585
rect 15043 18544 15052 18584
rect 15092 18544 15101 18584
rect 15043 18543 15101 18544
rect 15427 18584 15485 18585
rect 15427 18544 15436 18584
rect 15476 18544 15485 18584
rect 15723 18584 15765 18593
rect 15427 18543 15485 18544
rect 15531 18569 15573 18578
rect 12555 18521 12597 18530
rect 15531 18529 15532 18569
rect 15572 18529 15573 18569
rect 15723 18544 15724 18584
rect 15764 18544 15765 18584
rect 15723 18535 15765 18544
rect 15819 18584 15861 18593
rect 15819 18544 15820 18584
rect 15860 18544 15861 18584
rect 15819 18535 15861 18544
rect 15912 18584 15970 18585
rect 15912 18544 15921 18584
rect 15961 18544 15970 18584
rect 15912 18543 15970 18544
rect 16971 18584 17013 18593
rect 16971 18544 16972 18584
rect 17012 18544 17013 18584
rect 16971 18535 17013 18544
rect 17067 18584 17109 18593
rect 17067 18544 17068 18584
rect 17108 18544 17109 18584
rect 17067 18535 17109 18544
rect 17547 18584 17589 18593
rect 17547 18544 17548 18584
rect 17588 18544 17589 18584
rect 17547 18535 17589 18544
rect 18019 18584 18077 18585
rect 18019 18544 18028 18584
rect 18068 18544 18077 18584
rect 18019 18543 18077 18544
rect 18555 18574 18597 18583
rect 15531 18520 15573 18529
rect 18555 18534 18556 18574
rect 18596 18534 18597 18574
rect 18555 18525 18597 18534
rect 11595 18500 11637 18509
rect 11595 18460 11596 18500
rect 11636 18460 11637 18500
rect 11595 18451 11637 18460
rect 17451 18500 17493 18509
rect 17451 18460 17452 18500
rect 17492 18460 17493 18500
rect 17451 18451 17493 18460
rect 5739 18416 5781 18425
rect 5739 18376 5740 18416
rect 5780 18376 5781 18416
rect 5739 18367 5781 18376
rect 1152 18164 20352 18188
rect 1152 18124 3688 18164
rect 3728 18124 3770 18164
rect 3810 18124 3852 18164
rect 3892 18124 3934 18164
rect 3974 18124 4016 18164
rect 4056 18124 18808 18164
rect 18848 18124 18890 18164
rect 18930 18124 18972 18164
rect 19012 18124 19054 18164
rect 19094 18124 19136 18164
rect 19176 18124 20352 18164
rect 1152 18100 20352 18124
rect 7083 17996 7125 18005
rect 7083 17956 7084 17996
rect 7124 17956 7125 17996
rect 7083 17947 7125 17956
rect 8715 17996 8757 18005
rect 8715 17956 8716 17996
rect 8756 17956 8757 17996
rect 8715 17947 8757 17956
rect 10347 17996 10389 18005
rect 10347 17956 10348 17996
rect 10388 17956 10389 17996
rect 10347 17947 10389 17956
rect 12939 17996 12981 18005
rect 12939 17956 12940 17996
rect 12980 17956 12981 17996
rect 12939 17947 12981 17956
rect 14955 17996 14997 18005
rect 14955 17956 14956 17996
rect 14996 17956 14997 17996
rect 14955 17947 14997 17956
rect 17067 17996 17109 18005
rect 17067 17956 17068 17996
rect 17108 17956 17109 17996
rect 17067 17947 17109 17956
rect 4107 17828 4149 17837
rect 4107 17788 4108 17828
rect 4148 17788 4149 17828
rect 4107 17779 4149 17788
rect 4579 17786 4637 17787
rect 1323 17744 1365 17753
rect 1323 17704 1324 17744
rect 1364 17704 1365 17744
rect 1323 17695 1365 17704
rect 1515 17744 1557 17753
rect 1515 17704 1516 17744
rect 1556 17704 1557 17744
rect 1515 17695 1557 17704
rect 1611 17744 1653 17753
rect 1611 17704 1612 17744
rect 1652 17704 1653 17744
rect 1611 17695 1653 17704
rect 1795 17744 1853 17745
rect 1795 17704 1804 17744
rect 1844 17704 1853 17744
rect 1795 17703 1853 17704
rect 3043 17744 3101 17745
rect 3043 17704 3052 17744
rect 3092 17704 3101 17744
rect 3043 17703 3101 17704
rect 3531 17744 3573 17753
rect 3531 17704 3532 17744
rect 3572 17704 3573 17744
rect 3531 17695 3573 17704
rect 3627 17744 3669 17753
rect 3627 17704 3628 17744
rect 3668 17704 3669 17744
rect 3627 17695 3669 17704
rect 4011 17744 4053 17753
rect 4579 17746 4588 17786
rect 4628 17746 4637 17786
rect 4579 17745 4637 17746
rect 5067 17749 5109 17758
rect 4011 17704 4012 17744
rect 4052 17704 4053 17744
rect 4011 17695 4053 17704
rect 5067 17709 5068 17749
rect 5108 17709 5109 17749
rect 5067 17700 5109 17709
rect 5635 17744 5693 17745
rect 5635 17704 5644 17744
rect 5684 17704 5693 17744
rect 5635 17703 5693 17704
rect 6883 17744 6941 17745
rect 6883 17704 6892 17744
rect 6932 17704 6941 17744
rect 6883 17703 6941 17704
rect 7267 17744 7325 17745
rect 7267 17704 7276 17744
rect 7316 17704 7325 17744
rect 7267 17703 7325 17704
rect 8515 17744 8573 17745
rect 8515 17704 8524 17744
rect 8564 17704 8573 17744
rect 8515 17703 8573 17704
rect 8899 17744 8957 17745
rect 8899 17704 8908 17744
rect 8948 17704 8957 17744
rect 8899 17703 8957 17704
rect 10147 17744 10205 17745
rect 10147 17704 10156 17744
rect 10196 17704 10205 17744
rect 10147 17703 10205 17704
rect 11491 17744 11549 17745
rect 11491 17704 11500 17744
rect 11540 17704 11549 17744
rect 11491 17703 11549 17704
rect 12739 17744 12797 17745
rect 12739 17704 12748 17744
rect 12788 17704 12797 17744
rect 12739 17703 12797 17704
rect 13507 17744 13565 17745
rect 13507 17704 13516 17744
rect 13556 17704 13565 17744
rect 13507 17703 13565 17704
rect 14755 17744 14813 17745
rect 14755 17704 14764 17744
rect 14804 17704 14813 17744
rect 14755 17703 14813 17704
rect 15147 17744 15189 17753
rect 15147 17704 15148 17744
rect 15188 17704 15189 17744
rect 15147 17695 15189 17704
rect 15243 17744 15285 17753
rect 15243 17704 15244 17744
rect 15284 17704 15285 17744
rect 15243 17695 15285 17704
rect 15619 17744 15677 17745
rect 15619 17704 15628 17744
rect 15668 17704 15677 17744
rect 15619 17703 15677 17704
rect 16867 17744 16925 17745
rect 16867 17704 16876 17744
rect 16916 17704 16925 17744
rect 16867 17703 16925 17704
rect 17635 17744 17693 17745
rect 17635 17704 17644 17744
rect 17684 17704 17693 17744
rect 17635 17703 17693 17704
rect 18883 17744 18941 17745
rect 18883 17704 18892 17744
rect 18932 17704 18941 17744
rect 18883 17703 18941 17704
rect 3243 17660 3285 17669
rect 3243 17620 3244 17660
rect 3284 17620 3285 17660
rect 3243 17611 3285 17620
rect 19083 17660 19125 17669
rect 19083 17620 19084 17660
rect 19124 17620 19125 17660
rect 19083 17611 19125 17620
rect 1419 17576 1461 17585
rect 1419 17536 1420 17576
rect 1460 17536 1461 17576
rect 1419 17527 1461 17536
rect 5259 17576 5301 17585
rect 5259 17536 5260 17576
rect 5300 17536 5301 17576
rect 5259 17527 5301 17536
rect 14955 17576 14997 17585
rect 14955 17536 14956 17576
rect 14996 17536 14997 17576
rect 14955 17527 14997 17536
rect 15427 17576 15485 17577
rect 15427 17536 15436 17576
rect 15476 17536 15485 17576
rect 15427 17535 15485 17536
rect 1152 17408 20452 17432
rect 1152 17368 4928 17408
rect 4968 17368 5010 17408
rect 5050 17368 5092 17408
rect 5132 17368 5174 17408
rect 5214 17368 5256 17408
rect 5296 17368 20048 17408
rect 20088 17368 20130 17408
rect 20170 17368 20212 17408
rect 20252 17368 20294 17408
rect 20334 17368 20376 17408
rect 20416 17368 20452 17408
rect 1152 17344 20452 17368
rect 2667 17240 2709 17249
rect 2667 17200 2668 17240
rect 2708 17200 2709 17240
rect 2667 17191 2709 17200
rect 15051 17240 15093 17249
rect 15051 17200 15052 17240
rect 15092 17200 15093 17240
rect 15051 17191 15093 17200
rect 5163 17156 5205 17165
rect 5163 17116 5164 17156
rect 5204 17116 5205 17156
rect 5163 17107 5205 17116
rect 9099 17156 9141 17165
rect 9099 17116 9100 17156
rect 9140 17116 9141 17156
rect 9099 17107 9141 17116
rect 11115 17156 11157 17165
rect 11115 17116 11116 17156
rect 11156 17116 11157 17156
rect 11115 17107 11157 17116
rect 11307 17156 11349 17165
rect 11307 17116 11308 17156
rect 11348 17116 11349 17156
rect 11307 17107 11349 17116
rect 18699 17156 18741 17165
rect 18699 17116 18700 17156
rect 18740 17116 18741 17156
rect 18699 17107 18741 17116
rect 1219 17072 1277 17073
rect 1219 17032 1228 17072
rect 1268 17032 1277 17072
rect 1219 17031 1277 17032
rect 2467 17072 2525 17073
rect 2467 17032 2476 17072
rect 2516 17032 2525 17072
rect 2467 17031 2525 17032
rect 2851 17072 2909 17073
rect 2851 17032 2860 17072
rect 2900 17032 2909 17072
rect 2851 17031 2909 17032
rect 2947 17072 3005 17073
rect 2947 17032 2956 17072
rect 2996 17032 3005 17072
rect 2947 17031 3005 17032
rect 3147 17072 3189 17081
rect 3147 17032 3148 17072
rect 3188 17032 3189 17072
rect 3147 17023 3189 17032
rect 3243 17072 3285 17081
rect 3243 17032 3244 17072
rect 3284 17032 3285 17072
rect 3243 17023 3285 17032
rect 3336 17072 3394 17073
rect 3336 17032 3345 17072
rect 3385 17032 3394 17072
rect 3336 17031 3394 17032
rect 3715 17072 3773 17073
rect 3715 17032 3724 17072
rect 3764 17032 3773 17072
rect 3715 17031 3773 17032
rect 4963 17072 5021 17073
rect 4963 17032 4972 17072
rect 5012 17032 5021 17072
rect 4963 17031 5021 17032
rect 6019 17072 6077 17073
rect 6019 17032 6028 17072
rect 6068 17032 6077 17072
rect 6019 17031 6077 17032
rect 7267 17072 7325 17073
rect 7267 17032 7276 17072
rect 7316 17032 7325 17072
rect 7267 17031 7325 17032
rect 7651 17072 7709 17073
rect 7651 17032 7660 17072
rect 7700 17032 7709 17072
rect 7651 17031 7709 17032
rect 8899 17072 8957 17073
rect 8899 17032 8908 17072
rect 8948 17032 8957 17072
rect 8899 17031 8957 17032
rect 9387 17072 9429 17081
rect 9387 17032 9388 17072
rect 9428 17032 9429 17072
rect 9387 17023 9429 17032
rect 9483 17072 9525 17081
rect 9483 17032 9484 17072
rect 9524 17032 9525 17072
rect 9483 17023 9525 17032
rect 9867 17072 9909 17081
rect 9867 17032 9868 17072
rect 9908 17032 9909 17072
rect 9867 17023 9909 17032
rect 9963 17072 10005 17081
rect 9963 17032 9964 17072
rect 10004 17032 10005 17072
rect 9963 17023 10005 17032
rect 10435 17072 10493 17073
rect 10435 17032 10444 17072
rect 10484 17032 10493 17072
rect 10435 17031 10493 17032
rect 10923 17067 10965 17076
rect 10923 17027 10924 17067
rect 10964 17027 10965 17067
rect 11491 17072 11549 17073
rect 11491 17032 11500 17072
rect 11540 17032 11549 17072
rect 11491 17031 11549 17032
rect 12739 17072 12797 17073
rect 12739 17032 12748 17072
rect 12788 17032 12797 17072
rect 12739 17031 12797 17032
rect 13603 17072 13661 17073
rect 13603 17032 13612 17072
rect 13652 17032 13661 17072
rect 13603 17031 13661 17032
rect 14851 17072 14909 17073
rect 14851 17032 14860 17072
rect 14900 17032 14909 17072
rect 14851 17031 14909 17032
rect 15235 17072 15293 17073
rect 15235 17032 15244 17072
rect 15284 17032 15293 17072
rect 15235 17031 15293 17032
rect 16483 17072 16541 17073
rect 16483 17032 16492 17072
rect 16532 17032 16541 17072
rect 16483 17031 16541 17032
rect 16971 17072 17013 17081
rect 16971 17032 16972 17072
rect 17012 17032 17013 17072
rect 10923 17018 10965 17027
rect 16971 17023 17013 17032
rect 17067 17072 17109 17081
rect 17067 17032 17068 17072
rect 17108 17032 17109 17072
rect 17067 17023 17109 17032
rect 18019 17072 18077 17073
rect 18019 17032 18028 17072
rect 18068 17032 18077 17072
rect 18019 17031 18077 17032
rect 18507 17067 18549 17076
rect 18507 17027 18508 17067
rect 18548 17027 18549 17067
rect 18507 17018 18549 17027
rect 17451 16988 17493 16997
rect 17451 16948 17452 16988
rect 17492 16948 17493 16988
rect 17451 16939 17493 16948
rect 17547 16988 17589 16997
rect 17547 16948 17548 16988
rect 17588 16948 17589 16988
rect 17547 16939 17589 16948
rect 16683 16904 16725 16913
rect 16683 16864 16684 16904
rect 16724 16864 16725 16904
rect 16683 16855 16725 16864
rect 2859 16820 2901 16829
rect 2859 16780 2860 16820
rect 2900 16780 2901 16820
rect 2859 16771 2901 16780
rect 7467 16820 7509 16829
rect 7467 16780 7468 16820
rect 7508 16780 7509 16820
rect 7467 16771 7509 16780
rect 15051 16820 15093 16829
rect 15051 16780 15052 16820
rect 15092 16780 15093 16820
rect 15051 16771 15093 16780
rect 1152 16652 20352 16676
rect 1152 16612 3688 16652
rect 3728 16612 3770 16652
rect 3810 16612 3852 16652
rect 3892 16612 3934 16652
rect 3974 16612 4016 16652
rect 4056 16612 18808 16652
rect 18848 16612 18890 16652
rect 18930 16612 18972 16652
rect 19012 16612 19054 16652
rect 19094 16612 19136 16652
rect 19176 16612 20352 16652
rect 1152 16588 20352 16612
rect 2667 16484 2709 16493
rect 2667 16444 2668 16484
rect 2708 16444 2709 16484
rect 2667 16435 2709 16444
rect 5547 16400 5589 16409
rect 5547 16360 5548 16400
rect 5588 16360 5589 16400
rect 5547 16351 5589 16360
rect 14659 16400 14717 16401
rect 14659 16360 14668 16400
rect 14708 16360 14717 16400
rect 14659 16359 14717 16360
rect 6411 16316 6453 16325
rect 3043 16303 3101 16304
rect 3043 16263 3052 16303
rect 3092 16263 3101 16303
rect 6411 16276 6412 16316
rect 6452 16276 6453 16316
rect 9867 16316 9909 16325
rect 6411 16267 6453 16276
rect 7419 16274 7461 16283
rect 3043 16262 3101 16263
rect 5835 16251 5877 16260
rect 1219 16232 1277 16233
rect 1219 16192 1228 16232
rect 1268 16192 1277 16232
rect 1219 16191 1277 16192
rect 2467 16232 2525 16233
rect 2467 16192 2476 16232
rect 2516 16192 2525 16232
rect 2467 16191 2525 16192
rect 3243 16232 3285 16241
rect 3243 16192 3244 16232
rect 3284 16192 3285 16232
rect 3243 16183 3285 16192
rect 3339 16232 3381 16241
rect 3339 16192 3340 16232
rect 3380 16192 3381 16232
rect 3339 16183 3381 16192
rect 3531 16232 3573 16241
rect 3531 16192 3532 16232
rect 3572 16192 3573 16232
rect 3531 16183 3573 16192
rect 4099 16232 4157 16233
rect 4099 16192 4108 16232
rect 4148 16192 4157 16232
rect 4099 16191 4157 16192
rect 5347 16232 5405 16233
rect 5347 16192 5356 16232
rect 5396 16192 5405 16232
rect 5835 16211 5836 16251
rect 5876 16211 5877 16251
rect 5835 16202 5877 16211
rect 5931 16232 5973 16241
rect 5347 16191 5405 16192
rect 5931 16192 5932 16232
rect 5972 16192 5973 16232
rect 5931 16183 5973 16192
rect 6315 16232 6357 16241
rect 7419 16234 7420 16274
rect 7460 16234 7461 16274
rect 9867 16276 9868 16316
rect 9908 16276 9909 16316
rect 9867 16267 9909 16276
rect 10875 16241 10917 16250
rect 6315 16192 6316 16232
rect 6356 16192 6357 16232
rect 6315 16183 6357 16192
rect 6883 16232 6941 16233
rect 6883 16192 6892 16232
rect 6932 16192 6941 16232
rect 7419 16225 7461 16234
rect 9291 16232 9333 16241
rect 6883 16191 6941 16192
rect 9291 16192 9292 16232
rect 9332 16192 9333 16232
rect 9291 16183 9333 16192
rect 9387 16232 9429 16241
rect 9387 16192 9388 16232
rect 9428 16192 9429 16232
rect 9387 16183 9429 16192
rect 9771 16232 9813 16241
rect 9771 16192 9772 16232
rect 9812 16192 9813 16232
rect 9771 16183 9813 16192
rect 10339 16232 10397 16233
rect 10339 16192 10348 16232
rect 10388 16192 10397 16232
rect 10875 16201 10876 16241
rect 10916 16201 10917 16241
rect 10875 16192 10917 16201
rect 12451 16232 12509 16233
rect 12451 16192 12460 16232
rect 12500 16192 12509 16232
rect 10339 16191 10397 16192
rect 12451 16191 12509 16192
rect 13699 16232 13757 16233
rect 13699 16192 13708 16232
rect 13748 16192 13757 16232
rect 13699 16191 13757 16192
rect 14475 16232 14517 16241
rect 14475 16192 14476 16232
rect 14516 16192 14517 16232
rect 14475 16183 14517 16192
rect 14667 16232 14709 16241
rect 14667 16192 14668 16232
rect 14708 16192 14709 16232
rect 14667 16183 14709 16192
rect 14763 16232 14805 16241
rect 14763 16192 14764 16232
rect 14804 16192 14805 16232
rect 14763 16183 14805 16192
rect 14947 16232 15005 16233
rect 14947 16192 14956 16232
rect 14996 16192 15005 16232
rect 14947 16191 15005 16192
rect 16195 16232 16253 16233
rect 16195 16192 16204 16232
rect 16244 16192 16253 16232
rect 16195 16191 16253 16192
rect 16683 16232 16725 16241
rect 16683 16192 16684 16232
rect 16724 16192 16725 16232
rect 16683 16183 16725 16192
rect 16779 16232 16821 16241
rect 16779 16192 16780 16232
rect 16820 16192 16821 16232
rect 16779 16183 16821 16192
rect 17163 16232 17205 16241
rect 17163 16192 17164 16232
rect 17204 16192 17205 16232
rect 17163 16183 17205 16192
rect 17259 16232 17301 16241
rect 18219 16237 18261 16246
rect 17259 16192 17260 16232
rect 17300 16192 17301 16232
rect 17259 16183 17301 16192
rect 17731 16232 17789 16233
rect 17731 16192 17740 16232
rect 17780 16192 17789 16232
rect 17731 16191 17789 16192
rect 18219 16197 18220 16237
rect 18260 16197 18261 16237
rect 18219 16188 18261 16197
rect 16395 16148 16437 16157
rect 16395 16108 16396 16148
rect 16436 16108 16437 16148
rect 16395 16099 16437 16108
rect 18411 16148 18453 16157
rect 18411 16108 18412 16148
rect 18452 16108 18453 16148
rect 18411 16099 18453 16108
rect 2859 16064 2901 16073
rect 2859 16024 2860 16064
rect 2900 16024 2901 16064
rect 2859 16015 2901 16024
rect 3435 16064 3477 16073
rect 3435 16024 3436 16064
rect 3476 16024 3477 16064
rect 3435 16015 3477 16024
rect 7563 16064 7605 16073
rect 7563 16024 7564 16064
rect 7604 16024 7605 16064
rect 7563 16015 7605 16024
rect 11019 16064 11061 16073
rect 11019 16024 11020 16064
rect 11060 16024 11061 16064
rect 11019 16015 11061 16024
rect 13899 16064 13941 16073
rect 13899 16024 13900 16064
rect 13940 16024 13941 16064
rect 13899 16015 13941 16024
rect 1152 15896 20452 15920
rect 1152 15856 4928 15896
rect 4968 15856 5010 15896
rect 5050 15856 5092 15896
rect 5132 15856 5174 15896
rect 5214 15856 5256 15896
rect 5296 15856 20048 15896
rect 20088 15856 20130 15896
rect 20170 15856 20212 15896
rect 20252 15856 20294 15896
rect 20334 15856 20376 15896
rect 20416 15856 20452 15896
rect 1152 15832 20452 15856
rect 14091 15728 14133 15737
rect 14091 15688 14092 15728
rect 14132 15688 14133 15728
rect 14091 15679 14133 15688
rect 18027 15728 18069 15737
rect 18027 15688 18028 15728
rect 18068 15688 18069 15728
rect 18027 15679 18069 15688
rect 8715 15644 8757 15653
rect 8715 15604 8716 15644
rect 8756 15604 8757 15644
rect 1795 15602 1853 15603
rect 1795 15562 1804 15602
rect 1844 15562 1853 15602
rect 8715 15595 8757 15604
rect 12075 15644 12117 15653
rect 12075 15604 12076 15644
rect 12116 15604 12117 15644
rect 12075 15595 12117 15604
rect 1795 15561 1853 15562
rect 3043 15560 3101 15561
rect 3043 15520 3052 15560
rect 3092 15520 3101 15560
rect 3043 15519 3101 15520
rect 3435 15556 3477 15565
rect 3435 15516 3436 15556
rect 3476 15516 3477 15556
rect 3523 15560 3581 15561
rect 3523 15520 3532 15560
rect 3572 15520 3581 15560
rect 3523 15519 3581 15520
rect 3723 15560 3765 15569
rect 3723 15520 3724 15560
rect 3764 15520 3765 15560
rect 3435 15507 3477 15516
rect 3723 15511 3765 15520
rect 3819 15560 3861 15569
rect 3819 15520 3820 15560
rect 3860 15520 3861 15560
rect 3819 15511 3861 15520
rect 3966 15560 4024 15561
rect 3966 15520 3975 15560
rect 4015 15520 4024 15560
rect 3966 15519 4024 15520
rect 5251 15560 5309 15561
rect 5251 15520 5260 15560
rect 5300 15520 5309 15560
rect 5251 15519 5309 15520
rect 6499 15560 6557 15561
rect 6499 15520 6508 15560
rect 6548 15520 6557 15560
rect 6499 15519 6557 15520
rect 6987 15560 7029 15569
rect 6987 15520 6988 15560
rect 7028 15520 7029 15560
rect 6987 15511 7029 15520
rect 7083 15560 7125 15569
rect 7083 15520 7084 15560
rect 7124 15520 7125 15560
rect 7083 15511 7125 15520
rect 7467 15560 7509 15569
rect 7467 15520 7468 15560
rect 7508 15520 7509 15560
rect 7467 15511 7509 15520
rect 8035 15560 8093 15561
rect 8035 15520 8044 15560
rect 8084 15520 8093 15560
rect 10627 15560 10685 15561
rect 8035 15519 8093 15520
rect 8571 15518 8613 15527
rect 10627 15520 10636 15560
rect 10676 15520 10685 15560
rect 10627 15519 10685 15520
rect 11875 15560 11933 15561
rect 11875 15520 11884 15560
rect 11924 15520 11933 15560
rect 11875 15519 11933 15520
rect 12363 15560 12405 15569
rect 12363 15520 12364 15560
rect 12404 15520 12405 15560
rect 1603 15476 1661 15477
rect 1603 15436 1612 15476
rect 1652 15436 1661 15476
rect 1603 15435 1661 15436
rect 4387 15476 4445 15477
rect 4387 15436 4396 15476
rect 4436 15436 4445 15476
rect 4387 15435 4445 15436
rect 7563 15476 7605 15485
rect 7563 15436 7564 15476
rect 7604 15436 7605 15476
rect 8571 15478 8572 15518
rect 8612 15478 8613 15518
rect 12363 15511 12405 15520
rect 12459 15560 12501 15569
rect 12459 15520 12460 15560
rect 12500 15520 12501 15560
rect 12459 15511 12501 15520
rect 13411 15560 13469 15561
rect 13411 15520 13420 15560
rect 13460 15520 13469 15560
rect 13411 15519 13469 15520
rect 13899 15555 13941 15564
rect 13899 15515 13900 15555
rect 13940 15515 13941 15555
rect 14275 15560 14333 15561
rect 14275 15520 14284 15560
rect 14324 15520 14333 15560
rect 14275 15519 14333 15520
rect 15523 15560 15581 15561
rect 15523 15520 15532 15560
rect 15572 15520 15581 15560
rect 15523 15519 15581 15520
rect 16579 15560 16637 15561
rect 16579 15520 16588 15560
rect 16628 15520 16637 15560
rect 16579 15519 16637 15520
rect 17827 15560 17885 15561
rect 17827 15520 17836 15560
rect 17876 15520 17885 15560
rect 17827 15519 17885 15520
rect 13899 15506 13941 15515
rect 8571 15469 8613 15478
rect 12843 15476 12885 15485
rect 7563 15427 7605 15436
rect 12843 15436 12844 15476
rect 12884 15436 12885 15476
rect 12843 15427 12885 15436
rect 12939 15476 12981 15485
rect 12939 15436 12940 15476
rect 12980 15436 12981 15476
rect 12939 15427 12981 15436
rect 1419 15392 1461 15401
rect 1419 15352 1420 15392
rect 1460 15352 1461 15392
rect 1419 15343 1461 15352
rect 6699 15392 6741 15401
rect 6699 15352 6700 15392
rect 6740 15352 6741 15392
rect 6699 15343 6741 15352
rect 3243 15308 3285 15317
rect 3243 15268 3244 15308
rect 3284 15268 3285 15308
rect 3243 15259 3285 15268
rect 3435 15308 3477 15317
rect 3435 15268 3436 15308
rect 3476 15268 3477 15308
rect 3435 15259 3477 15268
rect 4203 15308 4245 15317
rect 4203 15268 4204 15308
rect 4244 15268 4245 15308
rect 4203 15259 4245 15268
rect 15723 15308 15765 15317
rect 15723 15268 15724 15308
rect 15764 15268 15765 15308
rect 15723 15259 15765 15268
rect 1152 15140 20352 15164
rect 1152 15100 3688 15140
rect 3728 15100 3770 15140
rect 3810 15100 3852 15140
rect 3892 15100 3934 15140
rect 3974 15100 4016 15140
rect 4056 15100 18808 15140
rect 18848 15100 18890 15140
rect 18930 15100 18972 15140
rect 19012 15100 19054 15140
rect 19094 15100 19136 15140
rect 19176 15100 20352 15140
rect 1152 15076 20352 15100
rect 1419 14972 1461 14981
rect 1419 14932 1420 14972
rect 1460 14932 1461 14972
rect 1419 14923 1461 14932
rect 3243 14972 3285 14981
rect 3243 14932 3244 14972
rect 3284 14932 3285 14972
rect 3243 14923 3285 14932
rect 9483 14972 9525 14981
rect 9483 14932 9484 14972
rect 9524 14932 9525 14972
rect 9483 14923 9525 14932
rect 11211 14972 11253 14981
rect 11211 14932 11212 14972
rect 11252 14932 11253 14972
rect 11211 14923 11253 14932
rect 7659 14888 7701 14897
rect 7659 14848 7660 14888
rect 7700 14848 7701 14888
rect 7659 14839 7701 14848
rect 1603 14804 1661 14805
rect 1603 14764 1612 14804
rect 1652 14764 1661 14804
rect 1603 14763 1661 14764
rect 4587 14804 4629 14813
rect 4587 14764 4588 14804
rect 4628 14764 4629 14804
rect 4587 14755 4629 14764
rect 4683 14804 4725 14813
rect 4683 14764 4684 14804
rect 4724 14764 4725 14804
rect 4683 14755 4725 14764
rect 7843 14804 7901 14805
rect 7843 14764 7852 14804
rect 7892 14764 7901 14804
rect 7843 14763 7901 14764
rect 13995 14804 14037 14813
rect 13995 14764 13996 14804
rect 14036 14764 14037 14804
rect 13995 14755 14037 14764
rect 17547 14804 17589 14813
rect 17547 14764 17548 14804
rect 17588 14764 17589 14804
rect 17547 14755 17589 14764
rect 15051 14734 15093 14743
rect 1795 14720 1853 14721
rect 1795 14680 1804 14720
rect 1844 14680 1853 14720
rect 1795 14679 1853 14680
rect 3043 14720 3101 14721
rect 3043 14680 3052 14720
rect 3092 14680 3101 14720
rect 3043 14679 3101 14680
rect 3435 14720 3477 14729
rect 3435 14680 3436 14720
rect 3476 14680 3477 14720
rect 3435 14671 3477 14680
rect 3531 14720 3573 14729
rect 3531 14680 3532 14720
rect 3572 14680 3573 14720
rect 3531 14671 3573 14680
rect 4107 14720 4149 14729
rect 4107 14680 4108 14720
rect 4148 14680 4149 14720
rect 4107 14671 4149 14680
rect 4203 14720 4245 14729
rect 5643 14725 5685 14734
rect 4203 14680 4204 14720
rect 4244 14680 4245 14720
rect 4203 14671 4245 14680
rect 5155 14720 5213 14721
rect 5155 14680 5164 14720
rect 5204 14680 5213 14720
rect 5155 14679 5213 14680
rect 5643 14685 5644 14725
rect 5684 14685 5685 14725
rect 5643 14676 5685 14685
rect 8035 14720 8093 14721
rect 8035 14680 8044 14720
rect 8084 14680 8093 14720
rect 8035 14679 8093 14680
rect 9283 14720 9341 14721
rect 9283 14680 9292 14720
rect 9332 14680 9341 14720
rect 9283 14679 9341 14680
rect 9763 14720 9821 14721
rect 9763 14680 9772 14720
rect 9812 14680 9821 14720
rect 9763 14679 9821 14680
rect 11011 14720 11069 14721
rect 11011 14680 11020 14720
rect 11060 14680 11069 14720
rect 11011 14679 11069 14680
rect 11779 14720 11837 14721
rect 11779 14680 11788 14720
rect 11828 14680 11837 14720
rect 11779 14679 11837 14680
rect 13027 14720 13085 14721
rect 13027 14680 13036 14720
rect 13076 14680 13085 14720
rect 13027 14679 13085 14680
rect 13515 14720 13557 14729
rect 13515 14680 13516 14720
rect 13556 14680 13557 14720
rect 13515 14671 13557 14680
rect 13611 14720 13653 14729
rect 13611 14680 13612 14720
rect 13652 14680 13653 14720
rect 13611 14671 13653 14680
rect 14091 14720 14133 14729
rect 14091 14680 14092 14720
rect 14132 14680 14133 14720
rect 14091 14671 14133 14680
rect 14563 14720 14621 14721
rect 14563 14680 14572 14720
rect 14612 14680 14621 14720
rect 15051 14694 15052 14734
rect 15092 14694 15093 14734
rect 15051 14685 15093 14694
rect 17067 14720 17109 14729
rect 14563 14679 14621 14680
rect 17067 14680 17068 14720
rect 17108 14680 17109 14720
rect 17067 14671 17109 14680
rect 17163 14720 17205 14729
rect 17163 14680 17164 14720
rect 17204 14680 17205 14720
rect 17163 14671 17205 14680
rect 17643 14720 17685 14729
rect 18603 14725 18645 14734
rect 17643 14680 17644 14720
rect 17684 14680 17685 14720
rect 17643 14671 17685 14680
rect 18115 14720 18173 14721
rect 18115 14680 18124 14720
rect 18164 14680 18173 14720
rect 18115 14679 18173 14680
rect 18603 14685 18604 14725
rect 18644 14685 18645 14725
rect 18603 14676 18645 14685
rect 5835 14636 5877 14645
rect 5835 14596 5836 14636
rect 5876 14596 5877 14636
rect 5835 14587 5877 14596
rect 13227 14636 13269 14645
rect 13227 14596 13228 14636
rect 13268 14596 13269 14636
rect 13227 14587 13269 14596
rect 15243 14636 15285 14645
rect 15243 14596 15244 14636
rect 15284 14596 15285 14636
rect 15243 14587 15285 14596
rect 3715 14552 3773 14553
rect 3715 14512 3724 14552
rect 3764 14512 3773 14552
rect 3715 14511 3773 14512
rect 18795 14552 18837 14561
rect 18795 14512 18796 14552
rect 18836 14512 18837 14552
rect 18795 14503 18837 14512
rect 1152 14384 20452 14408
rect 1152 14344 4928 14384
rect 4968 14344 5010 14384
rect 5050 14344 5092 14384
rect 5132 14344 5174 14384
rect 5214 14344 5256 14384
rect 5296 14344 20048 14384
rect 20088 14344 20130 14384
rect 20170 14344 20212 14384
rect 20252 14344 20294 14384
rect 20334 14344 20376 14384
rect 20416 14344 20452 14384
rect 1152 14320 20452 14344
rect 1323 14216 1365 14225
rect 1323 14176 1324 14216
rect 1364 14176 1365 14216
rect 1323 14167 1365 14176
rect 4011 14216 4053 14225
rect 4011 14176 4012 14216
rect 4052 14176 4053 14216
rect 4011 14167 4053 14176
rect 5643 14216 5685 14225
rect 5643 14176 5644 14216
rect 5684 14176 5685 14216
rect 5643 14167 5685 14176
rect 8811 14216 8853 14225
rect 8811 14176 8812 14216
rect 8852 14176 8853 14216
rect 8811 14167 8853 14176
rect 17355 14216 17397 14225
rect 17355 14176 17356 14216
rect 17396 14176 17397 14216
rect 17355 14167 17397 14176
rect 19179 14216 19221 14225
rect 19179 14176 19180 14216
rect 19220 14176 19221 14216
rect 19179 14167 19221 14176
rect 11115 14132 11157 14141
rect 11115 14092 11116 14132
rect 11156 14092 11157 14132
rect 11115 14083 11157 14092
rect 15339 14132 15381 14141
rect 15339 14092 15340 14132
rect 15380 14092 15381 14132
rect 15339 14083 15381 14092
rect 2091 14048 2133 14057
rect 2091 14008 2092 14048
rect 2132 14008 2133 14048
rect 2091 13999 2133 14008
rect 2283 14048 2325 14057
rect 2283 14008 2284 14048
rect 2324 14008 2325 14048
rect 2283 13999 2325 14008
rect 2379 14048 2421 14057
rect 2379 14008 2380 14048
rect 2420 14008 2421 14048
rect 2379 13999 2421 14008
rect 2563 14048 2621 14049
rect 2563 14008 2572 14048
rect 2612 14008 2621 14048
rect 2563 14007 2621 14008
rect 3811 14048 3869 14049
rect 3811 14008 3820 14048
rect 3860 14008 3869 14048
rect 3811 14007 3869 14008
rect 5443 14048 5501 14049
rect 5443 14008 5452 14048
rect 5492 14008 5501 14048
rect 5443 14007 5501 14008
rect 7363 14048 7421 14049
rect 7363 14008 7372 14048
rect 7412 14008 7421 14048
rect 7363 14007 7421 14008
rect 8611 14048 8669 14049
rect 8611 14008 8620 14048
rect 8660 14008 8669 14048
rect 8611 14007 8669 14008
rect 9387 14048 9429 14057
rect 9387 14008 9388 14048
rect 9428 14008 9429 14048
rect 4195 14006 4253 14007
rect 4195 13966 4204 14006
rect 4244 13966 4253 14006
rect 9387 13999 9429 14008
rect 9483 14048 9525 14057
rect 9483 14008 9484 14048
rect 9524 14008 9525 14048
rect 9483 13999 9525 14008
rect 9867 14048 9909 14057
rect 9867 14008 9868 14048
rect 9908 14008 9909 14048
rect 9867 13999 9909 14008
rect 9963 14048 10005 14057
rect 9963 14008 9964 14048
rect 10004 14008 10005 14048
rect 9963 13999 10005 14008
rect 10435 14048 10493 14049
rect 10435 14008 10444 14048
rect 10484 14008 10493 14048
rect 11875 14048 11933 14049
rect 10435 14007 10493 14008
rect 10971 14006 11013 14015
rect 11875 14008 11884 14048
rect 11924 14008 11933 14048
rect 11875 14007 11933 14008
rect 13123 14048 13181 14049
rect 13123 14008 13132 14048
rect 13172 14008 13181 14048
rect 13123 14007 13181 14008
rect 13891 14048 13949 14049
rect 13891 14008 13900 14048
rect 13940 14008 13949 14048
rect 13891 14007 13949 14008
rect 15139 14048 15197 14049
rect 15139 14008 15148 14048
rect 15188 14008 15197 14048
rect 15139 14007 15197 14008
rect 15627 14048 15669 14057
rect 15627 14008 15628 14048
rect 15668 14008 15669 14048
rect 4195 13965 4253 13966
rect 10971 13966 10972 14006
rect 11012 13966 11013 14006
rect 15627 13999 15669 14008
rect 15723 14048 15765 14057
rect 15723 14008 15724 14048
rect 15764 14008 15765 14048
rect 15723 13999 15765 14008
rect 16107 14048 16149 14057
rect 16107 14008 16108 14048
rect 16148 14008 16149 14048
rect 16107 13999 16149 14008
rect 16675 14048 16733 14049
rect 16675 14008 16684 14048
rect 16724 14008 16733 14048
rect 17731 14048 17789 14049
rect 16675 14007 16733 14008
rect 17211 14038 17253 14047
rect 17211 13998 17212 14038
rect 17252 13998 17253 14038
rect 17731 14008 17740 14048
rect 17780 14008 17789 14048
rect 17731 14007 17789 14008
rect 18979 14048 19037 14049
rect 18979 14008 18988 14048
rect 19028 14008 19037 14048
rect 18979 14007 19037 14008
rect 17211 13989 17253 13998
rect 1507 13964 1565 13965
rect 1507 13924 1516 13964
rect 1556 13924 1565 13964
rect 1507 13923 1565 13924
rect 1891 13964 1949 13965
rect 1891 13924 1900 13964
rect 1940 13924 1949 13964
rect 10971 13957 11013 13966
rect 16203 13964 16245 13973
rect 1891 13923 1949 13924
rect 16203 13924 16204 13964
rect 16244 13924 16245 13964
rect 16203 13915 16245 13924
rect 2187 13880 2229 13889
rect 2187 13840 2188 13880
rect 2228 13840 2229 13880
rect 2187 13831 2229 13840
rect 1707 13796 1749 13805
rect 1707 13756 1708 13796
rect 1748 13756 1749 13796
rect 1707 13747 1749 13756
rect 13323 13796 13365 13805
rect 13323 13756 13324 13796
rect 13364 13756 13365 13796
rect 13323 13747 13365 13756
rect 1152 13628 20352 13652
rect 1152 13588 3688 13628
rect 3728 13588 3770 13628
rect 3810 13588 3852 13628
rect 3892 13588 3934 13628
rect 3974 13588 4016 13628
rect 4056 13588 18808 13628
rect 18848 13588 18890 13628
rect 18930 13588 18972 13628
rect 19012 13588 19054 13628
rect 19094 13588 19136 13628
rect 19176 13588 20352 13628
rect 1152 13564 20352 13588
rect 2667 13460 2709 13469
rect 2667 13420 2668 13460
rect 2708 13420 2709 13460
rect 2667 13411 2709 13420
rect 11211 13460 11253 13469
rect 11211 13420 11212 13460
rect 11252 13420 11253 13460
rect 11211 13411 11253 13420
rect 17355 13460 17397 13469
rect 17355 13420 17356 13460
rect 17396 13420 17397 13460
rect 17355 13411 17397 13420
rect 5067 13292 5109 13301
rect 5067 13252 5068 13292
rect 5108 13252 5109 13292
rect 5067 13243 5109 13252
rect 8043 13292 8085 13301
rect 8043 13252 8044 13292
rect 8084 13252 8085 13292
rect 8043 13243 8085 13252
rect 13803 13292 13845 13301
rect 13803 13252 13804 13292
rect 13844 13252 13845 13292
rect 13803 13243 13845 13252
rect 13899 13292 13941 13301
rect 13899 13252 13900 13292
rect 13940 13252 13941 13292
rect 13899 13243 13941 13252
rect 11011 13229 11069 13230
rect 1219 13208 1277 13209
rect 1219 13168 1228 13208
rect 1268 13168 1277 13208
rect 1219 13167 1277 13168
rect 2467 13208 2525 13209
rect 2467 13168 2476 13208
rect 2516 13168 2525 13208
rect 2467 13167 2525 13168
rect 2851 13208 2909 13209
rect 2851 13168 2860 13208
rect 2900 13168 2909 13208
rect 2851 13167 2909 13168
rect 4099 13208 4157 13209
rect 4099 13168 4108 13208
rect 4148 13168 4157 13208
rect 4099 13167 4157 13168
rect 4587 13208 4629 13217
rect 4587 13168 4588 13208
rect 4628 13168 4629 13208
rect 4587 13159 4629 13168
rect 4683 13208 4725 13217
rect 4683 13168 4684 13208
rect 4724 13168 4725 13208
rect 4683 13159 4725 13168
rect 5163 13208 5205 13217
rect 6123 13213 6165 13222
rect 5163 13168 5164 13208
rect 5204 13168 5205 13208
rect 5163 13159 5205 13168
rect 5635 13208 5693 13209
rect 5635 13168 5644 13208
rect 5684 13168 5693 13208
rect 5635 13167 5693 13168
rect 6123 13173 6124 13213
rect 6164 13173 6165 13213
rect 6123 13164 6165 13173
rect 6987 13213 7029 13222
rect 6987 13173 6988 13213
rect 7028 13173 7029 13213
rect 6987 13164 7029 13173
rect 7459 13208 7517 13209
rect 7459 13168 7468 13208
rect 7508 13168 7517 13208
rect 7459 13167 7517 13168
rect 7947 13208 7989 13217
rect 7947 13168 7948 13208
rect 7988 13168 7989 13208
rect 7947 13159 7989 13168
rect 8427 13208 8469 13217
rect 8427 13168 8428 13208
rect 8468 13168 8469 13208
rect 8427 13159 8469 13168
rect 8523 13208 8565 13217
rect 8523 13168 8524 13208
rect 8564 13168 8565 13208
rect 8523 13159 8565 13168
rect 9763 13208 9821 13209
rect 9763 13168 9772 13208
rect 9812 13168 9821 13208
rect 11011 13189 11020 13229
rect 11060 13189 11069 13229
rect 14907 13217 14949 13226
rect 11011 13188 11069 13189
rect 13323 13208 13365 13217
rect 9763 13167 9821 13168
rect 13323 13168 13324 13208
rect 13364 13168 13365 13208
rect 13323 13159 13365 13168
rect 13419 13208 13461 13217
rect 13419 13168 13420 13208
rect 13460 13168 13461 13208
rect 13419 13159 13461 13168
rect 14371 13208 14429 13209
rect 14371 13168 14380 13208
rect 14420 13168 14429 13208
rect 14907 13177 14908 13217
rect 14948 13177 14949 13217
rect 14907 13168 14949 13177
rect 15907 13208 15965 13209
rect 15907 13168 15916 13208
rect 15956 13168 15965 13208
rect 14371 13167 14429 13168
rect 15907 13167 15965 13168
rect 17155 13208 17213 13209
rect 17155 13168 17164 13208
rect 17204 13168 17213 13208
rect 17155 13167 17213 13168
rect 4299 13124 4341 13133
rect 4299 13084 4300 13124
rect 4340 13084 4341 13124
rect 4299 13075 4341 13084
rect 6795 13124 6837 13133
rect 6795 13084 6796 13124
rect 6836 13084 6837 13124
rect 6795 13075 6837 13084
rect 6315 13040 6357 13049
rect 6315 13000 6316 13040
rect 6356 13000 6357 13040
rect 6315 12991 6357 13000
rect 15051 13040 15093 13049
rect 15051 13000 15052 13040
rect 15092 13000 15093 13040
rect 15051 12991 15093 13000
rect 1152 12872 20452 12896
rect 1152 12832 4928 12872
rect 4968 12832 5010 12872
rect 5050 12832 5092 12872
rect 5132 12832 5174 12872
rect 5214 12832 5256 12872
rect 5296 12832 20048 12872
rect 20088 12832 20130 12872
rect 20170 12832 20212 12872
rect 20252 12832 20294 12872
rect 20334 12832 20376 12872
rect 20416 12832 20452 12872
rect 1152 12808 20452 12832
rect 2667 12704 2709 12713
rect 2667 12664 2668 12704
rect 2708 12664 2709 12704
rect 2667 12655 2709 12664
rect 3907 12704 3965 12705
rect 3907 12664 3916 12704
rect 3956 12664 3965 12704
rect 3907 12663 3965 12664
rect 6027 12704 6069 12713
rect 6027 12664 6028 12704
rect 6068 12664 6069 12704
rect 6027 12655 6069 12664
rect 7659 12620 7701 12629
rect 7659 12580 7660 12620
rect 7700 12580 7701 12620
rect 7659 12571 7701 12580
rect 9291 12620 9333 12629
rect 9291 12580 9292 12620
rect 9332 12580 9333 12620
rect 9291 12571 9333 12580
rect 12939 12620 12981 12629
rect 12939 12580 12940 12620
rect 12980 12580 12981 12620
rect 12939 12571 12981 12580
rect 15147 12620 15189 12629
rect 15147 12580 15148 12620
rect 15188 12580 15189 12620
rect 15147 12571 15189 12580
rect 17451 12620 17493 12629
rect 17451 12580 17452 12620
rect 17492 12580 17493 12620
rect 17451 12571 17493 12580
rect 1219 12536 1277 12537
rect 1219 12496 1228 12536
rect 1268 12496 1277 12536
rect 1219 12495 1277 12496
rect 2467 12536 2525 12537
rect 2467 12496 2476 12536
rect 2516 12496 2525 12536
rect 2467 12495 2525 12496
rect 2851 12536 2909 12537
rect 2851 12496 2860 12536
rect 2900 12496 2909 12536
rect 2851 12495 2909 12496
rect 2947 12536 3005 12537
rect 2947 12496 2956 12536
rect 2996 12496 3005 12536
rect 2947 12495 3005 12496
rect 3147 12536 3189 12545
rect 3147 12496 3148 12536
rect 3188 12496 3189 12536
rect 3147 12487 3189 12496
rect 3243 12536 3285 12545
rect 3243 12496 3244 12536
rect 3284 12496 3285 12536
rect 3243 12487 3285 12496
rect 3336 12536 3394 12537
rect 3336 12496 3345 12536
rect 3385 12496 3394 12536
rect 3336 12495 3394 12496
rect 3627 12536 3669 12545
rect 3627 12496 3628 12536
rect 3668 12496 3669 12536
rect 3627 12487 3669 12496
rect 3723 12536 3765 12545
rect 3723 12496 3724 12536
rect 3764 12496 3765 12536
rect 3723 12487 3765 12496
rect 4579 12536 4637 12537
rect 4579 12496 4588 12536
rect 4628 12496 4637 12536
rect 4579 12495 4637 12496
rect 5827 12536 5885 12537
rect 5827 12496 5836 12536
rect 5876 12496 5885 12536
rect 5827 12495 5885 12496
rect 6211 12536 6269 12537
rect 6211 12496 6220 12536
rect 6260 12496 6269 12536
rect 6211 12495 6269 12496
rect 7459 12536 7517 12537
rect 7459 12496 7468 12536
rect 7508 12496 7517 12536
rect 7459 12495 7517 12496
rect 7843 12536 7901 12537
rect 7843 12496 7852 12536
rect 7892 12496 7901 12536
rect 7843 12495 7901 12496
rect 9091 12536 9149 12537
rect 9091 12496 9100 12536
rect 9140 12496 9149 12536
rect 9091 12495 9149 12496
rect 9475 12536 9533 12537
rect 9475 12496 9484 12536
rect 9524 12496 9533 12536
rect 9475 12495 9533 12496
rect 10723 12536 10781 12537
rect 10723 12496 10732 12536
rect 10772 12496 10781 12536
rect 10723 12495 10781 12496
rect 11211 12536 11253 12545
rect 11211 12496 11212 12536
rect 11252 12496 11253 12536
rect 11211 12487 11253 12496
rect 11307 12536 11349 12545
rect 11307 12496 11308 12536
rect 11348 12496 11349 12536
rect 11307 12487 11349 12496
rect 12259 12536 12317 12537
rect 12259 12496 12268 12536
rect 12308 12496 12317 12536
rect 13699 12536 13757 12537
rect 12259 12495 12317 12496
rect 12747 12522 12789 12531
rect 12747 12482 12748 12522
rect 12788 12482 12789 12522
rect 13699 12496 13708 12536
rect 13748 12496 13757 12536
rect 13699 12495 13757 12496
rect 14947 12536 15005 12537
rect 14947 12496 14956 12536
rect 14996 12496 15005 12536
rect 14947 12495 15005 12496
rect 16003 12536 16061 12537
rect 16003 12496 16012 12536
rect 16052 12496 16061 12536
rect 16003 12495 16061 12496
rect 17251 12536 17309 12537
rect 17251 12496 17260 12536
rect 17300 12496 17309 12536
rect 17251 12495 17309 12496
rect 18307 12536 18365 12537
rect 18307 12496 18316 12536
rect 18356 12496 18365 12536
rect 18307 12495 18365 12496
rect 19555 12536 19613 12537
rect 19555 12496 19564 12536
rect 19604 12496 19613 12536
rect 19555 12495 19613 12496
rect 12747 12473 12789 12482
rect 11691 12452 11733 12461
rect 11691 12412 11692 12452
rect 11732 12412 11733 12452
rect 11691 12403 11733 12412
rect 11787 12452 11829 12461
rect 11787 12412 11788 12452
rect 11828 12412 11829 12452
rect 11787 12403 11829 12412
rect 17827 12452 17885 12453
rect 17827 12412 17836 12452
rect 17876 12412 17885 12452
rect 17827 12411 17885 12412
rect 17643 12368 17685 12377
rect 17643 12328 17644 12368
rect 17684 12328 17685 12368
rect 17643 12319 17685 12328
rect 2859 12284 2901 12293
rect 2859 12244 2860 12284
rect 2900 12244 2901 12284
rect 2859 12235 2901 12244
rect 10923 12284 10965 12293
rect 10923 12244 10924 12284
rect 10964 12244 10965 12284
rect 10923 12235 10965 12244
rect 18123 12284 18165 12293
rect 18123 12244 18124 12284
rect 18164 12244 18165 12284
rect 18123 12235 18165 12244
rect 1152 12116 20352 12140
rect 1152 12076 3688 12116
rect 3728 12076 3770 12116
rect 3810 12076 3852 12116
rect 3892 12076 3934 12116
rect 3974 12076 4016 12116
rect 4056 12076 18808 12116
rect 18848 12076 18890 12116
rect 18930 12076 18972 12116
rect 19012 12076 19054 12116
rect 19094 12076 19136 12116
rect 19176 12076 20352 12116
rect 1152 12052 20352 12076
rect 1803 11948 1845 11957
rect 1803 11908 1804 11948
rect 1844 11908 1845 11948
rect 1803 11899 1845 11908
rect 7275 11948 7317 11957
rect 7275 11908 7276 11948
rect 7316 11908 7317 11948
rect 7275 11899 7317 11908
rect 7467 11948 7509 11957
rect 7467 11908 7468 11948
rect 7508 11908 7509 11948
rect 7467 11899 7509 11908
rect 12651 11948 12693 11957
rect 12651 11908 12652 11948
rect 12692 11908 12693 11948
rect 12651 11899 12693 11908
rect 1603 11780 1661 11781
rect 1603 11740 1612 11780
rect 1652 11740 1661 11780
rect 1603 11739 1661 11740
rect 1987 11780 2045 11781
rect 1987 11740 1996 11780
rect 2036 11740 2045 11780
rect 1987 11739 2045 11740
rect 4395 11780 4437 11789
rect 4395 11740 4396 11780
rect 4436 11740 4437 11780
rect 4395 11731 4437 11740
rect 4491 11780 4533 11789
rect 4491 11740 4492 11780
rect 4532 11740 4533 11780
rect 4491 11731 4533 11740
rect 7651 11780 7709 11781
rect 7651 11740 7660 11780
rect 7700 11740 7709 11780
rect 7651 11739 7709 11740
rect 8811 11780 8853 11789
rect 8811 11740 8812 11780
rect 8852 11740 8853 11780
rect 5827 11738 5885 11739
rect 5499 11705 5541 11714
rect 2179 11696 2237 11697
rect 2179 11656 2188 11696
rect 2228 11656 2237 11696
rect 2179 11655 2237 11656
rect 3427 11696 3485 11697
rect 3427 11656 3436 11696
rect 3476 11656 3485 11696
rect 3427 11655 3485 11656
rect 3915 11696 3957 11705
rect 3915 11656 3916 11696
rect 3956 11656 3957 11696
rect 3915 11647 3957 11656
rect 4011 11696 4053 11705
rect 4011 11656 4012 11696
rect 4052 11656 4053 11696
rect 4011 11647 4053 11656
rect 4963 11696 5021 11697
rect 4963 11656 4972 11696
rect 5012 11656 5021 11696
rect 5499 11665 5500 11705
rect 5540 11665 5541 11705
rect 5827 11698 5836 11738
rect 5876 11698 5885 11738
rect 8811 11731 8853 11740
rect 8907 11780 8949 11789
rect 8907 11740 8908 11780
rect 8948 11740 8949 11780
rect 8907 11731 8949 11740
rect 10723 11780 10781 11781
rect 10723 11740 10732 11780
rect 10772 11740 10781 11780
rect 10723 11739 10781 11740
rect 13611 11780 13653 11789
rect 13611 11740 13612 11780
rect 13652 11740 13653 11780
rect 13611 11731 13653 11740
rect 13707 11780 13749 11789
rect 13707 11740 13708 11780
rect 13748 11740 13749 11780
rect 13707 11731 13749 11740
rect 16395 11780 16437 11789
rect 16395 11740 16396 11780
rect 16436 11740 16437 11780
rect 16395 11731 16437 11740
rect 16491 11780 16533 11789
rect 16491 11740 16492 11780
rect 16532 11740 16533 11780
rect 16491 11731 16533 11740
rect 5827 11697 5885 11698
rect 5499 11656 5541 11665
rect 7075 11696 7133 11697
rect 7075 11656 7084 11696
rect 7124 11656 7133 11696
rect 4963 11655 5021 11656
rect 7075 11655 7133 11656
rect 8331 11696 8373 11705
rect 8331 11656 8332 11696
rect 8372 11656 8373 11696
rect 8331 11647 8373 11656
rect 8427 11696 8469 11705
rect 9867 11701 9909 11710
rect 14715 11705 14757 11714
rect 8427 11656 8428 11696
rect 8468 11656 8469 11696
rect 8427 11647 8469 11656
rect 9379 11696 9437 11697
rect 9379 11656 9388 11696
rect 9428 11656 9437 11696
rect 9379 11655 9437 11656
rect 9867 11661 9868 11701
rect 9908 11661 9909 11701
rect 9867 11652 9909 11661
rect 11203 11696 11261 11697
rect 11203 11656 11212 11696
rect 11252 11656 11261 11696
rect 11203 11655 11261 11656
rect 12451 11696 12509 11697
rect 12451 11656 12460 11696
rect 12500 11656 12509 11696
rect 12451 11655 12509 11656
rect 13131 11696 13173 11705
rect 13131 11656 13132 11696
rect 13172 11656 13173 11696
rect 13131 11647 13173 11656
rect 13227 11696 13269 11705
rect 13227 11656 13228 11696
rect 13268 11656 13269 11696
rect 13227 11647 13269 11656
rect 14179 11696 14237 11697
rect 14179 11656 14188 11696
rect 14228 11656 14237 11696
rect 14715 11665 14716 11705
rect 14756 11665 14757 11705
rect 14715 11656 14757 11665
rect 15915 11696 15957 11705
rect 15915 11656 15916 11696
rect 15956 11656 15957 11696
rect 14179 11655 14237 11656
rect 15915 11647 15957 11656
rect 16011 11696 16053 11705
rect 17451 11701 17493 11710
rect 16011 11656 16012 11696
rect 16052 11656 16053 11696
rect 16011 11647 16053 11656
rect 16963 11696 17021 11697
rect 16963 11656 16972 11696
rect 17012 11656 17021 11696
rect 16963 11655 17021 11656
rect 17451 11661 17452 11701
rect 17492 11661 17493 11701
rect 17451 11652 17493 11661
rect 18019 11696 18077 11697
rect 18019 11656 18028 11696
rect 18068 11656 18077 11696
rect 18019 11655 18077 11656
rect 19267 11696 19325 11697
rect 19267 11656 19276 11696
rect 19316 11656 19325 11696
rect 19267 11655 19325 11656
rect 3627 11612 3669 11621
rect 3627 11572 3628 11612
rect 3668 11572 3669 11612
rect 17835 11612 17877 11621
rect 3627 11563 3669 11572
rect 5643 11570 5685 11579
rect 1419 11528 1461 11537
rect 1419 11488 1420 11528
rect 1460 11488 1461 11528
rect 5643 11530 5644 11570
rect 5684 11530 5685 11570
rect 17835 11572 17836 11612
rect 17876 11572 17877 11612
rect 17835 11563 17877 11572
rect 5643 11521 5685 11530
rect 10059 11528 10101 11537
rect 1419 11479 1461 11488
rect 10059 11488 10060 11528
rect 10100 11488 10101 11528
rect 10059 11479 10101 11488
rect 10539 11528 10581 11537
rect 10539 11488 10540 11528
rect 10580 11488 10581 11528
rect 10539 11479 10581 11488
rect 14859 11528 14901 11537
rect 14859 11488 14860 11528
rect 14900 11488 14901 11528
rect 14859 11479 14901 11488
rect 17643 11528 17685 11537
rect 17643 11488 17644 11528
rect 17684 11488 17685 11528
rect 17643 11479 17685 11488
rect 1152 11360 20452 11384
rect 1152 11320 4928 11360
rect 4968 11320 5010 11360
rect 5050 11320 5092 11360
rect 5132 11320 5174 11360
rect 5214 11320 5256 11360
rect 5296 11320 20048 11360
rect 20088 11320 20130 11360
rect 20170 11320 20212 11360
rect 20252 11320 20294 11360
rect 20334 11320 20376 11360
rect 20416 11320 20452 11360
rect 1152 11296 20452 11320
rect 1707 11192 1749 11201
rect 1707 11152 1708 11192
rect 1748 11152 1749 11192
rect 1707 11143 1749 11152
rect 5739 11192 5781 11201
rect 5739 11152 5740 11192
rect 5780 11152 5781 11192
rect 5739 11143 5781 11152
rect 10155 11192 10197 11201
rect 10155 11152 10156 11192
rect 10196 11152 10197 11192
rect 10155 11143 10197 11152
rect 10627 11192 10685 11193
rect 10627 11152 10636 11192
rect 10676 11152 10685 11192
rect 10627 11151 10685 11152
rect 13131 11192 13173 11201
rect 13131 11152 13132 11192
rect 13172 11152 13173 11192
rect 13131 11143 13173 11152
rect 14859 11192 14901 11201
rect 14859 11152 14860 11192
rect 14900 11152 14901 11192
rect 14859 11143 14901 11152
rect 16491 11192 16533 11201
rect 16491 11152 16492 11192
rect 16532 11152 16533 11192
rect 16491 11143 16533 11152
rect 7755 11108 7797 11117
rect 7755 11068 7756 11108
rect 7796 11068 7797 11108
rect 7755 11059 7797 11068
rect 17739 11108 17781 11117
rect 17739 11068 17740 11108
rect 17780 11068 17781 11108
rect 17739 11059 17781 11068
rect 2083 11024 2141 11025
rect 2083 10984 2092 11024
rect 2132 10984 2141 11024
rect 2083 10983 2141 10984
rect 3331 11024 3389 11025
rect 3331 10984 3340 11024
rect 3380 10984 3389 11024
rect 3331 10983 3389 10984
rect 4291 11024 4349 11025
rect 4291 10984 4300 11024
rect 4340 10984 4349 11024
rect 4291 10983 4349 10984
rect 5539 11024 5597 11025
rect 5539 10984 5548 11024
rect 5588 10984 5597 11024
rect 5539 10983 5597 10984
rect 6027 11024 6069 11033
rect 6027 10984 6028 11024
rect 6068 10984 6069 11024
rect 6027 10975 6069 10984
rect 6123 11024 6165 11033
rect 6123 10984 6124 11024
rect 6164 10984 6165 11024
rect 6123 10975 6165 10984
rect 6507 11024 6549 11033
rect 6507 10984 6508 11024
rect 6548 10984 6549 11024
rect 6507 10975 6549 10984
rect 7075 11024 7133 11025
rect 7075 10984 7084 11024
rect 7124 10984 7133 11024
rect 8707 11024 8765 11025
rect 7075 10983 7133 10984
rect 7611 10982 7653 10991
rect 8707 10984 8716 11024
rect 8756 10984 8765 11024
rect 8707 10983 8765 10984
rect 9955 11024 10013 11025
rect 9955 10984 9964 11024
rect 10004 10984 10013 11024
rect 9955 10983 10013 10984
rect 10347 11024 10389 11033
rect 10347 10984 10348 11024
rect 10388 10984 10389 11024
rect 1891 10940 1949 10941
rect 1517 10929 1575 10930
rect 1517 10889 1526 10929
rect 1566 10889 1575 10929
rect 1891 10900 1900 10940
rect 1940 10900 1949 10940
rect 1891 10899 1949 10900
rect 6603 10940 6645 10949
rect 6603 10900 6604 10940
rect 6644 10900 6645 10940
rect 7611 10942 7612 10982
rect 7652 10942 7653 10982
rect 10347 10975 10389 10984
rect 10443 11024 10485 11033
rect 10443 10984 10444 11024
rect 10484 10984 10485 11024
rect 10443 10975 10485 10984
rect 11683 11024 11741 11025
rect 11683 10984 11692 11024
rect 11732 10984 11741 11024
rect 11683 10983 11741 10984
rect 12931 11024 12989 11025
rect 12931 10984 12940 11024
rect 12980 10984 12989 11024
rect 12931 10983 12989 10984
rect 13411 11024 13469 11025
rect 13411 10984 13420 11024
rect 13460 10984 13469 11024
rect 13411 10983 13469 10984
rect 14659 11024 14717 11025
rect 14659 10984 14668 11024
rect 14708 10984 14717 11024
rect 14659 10983 14717 10984
rect 15043 11024 15101 11025
rect 15043 10984 15052 11024
rect 15092 10984 15101 11024
rect 15043 10983 15101 10984
rect 16291 11024 16349 11025
rect 16291 10984 16300 11024
rect 16340 10984 16349 11024
rect 16291 10983 16349 10984
rect 17931 11019 17973 11028
rect 17931 10979 17932 11019
rect 17972 10979 17973 11019
rect 18403 11024 18461 11025
rect 18403 10984 18412 11024
rect 18452 10984 18461 11024
rect 18403 10983 18461 10984
rect 18987 11024 19029 11033
rect 18987 10984 18988 11024
rect 19028 10984 19029 11024
rect 17931 10970 17973 10979
rect 18987 10975 19029 10984
rect 19371 11024 19413 11033
rect 19371 10984 19372 11024
rect 19412 10984 19413 11024
rect 19371 10975 19413 10984
rect 19467 11024 19509 11033
rect 19467 10984 19468 11024
rect 19508 10984 19509 11024
rect 19467 10975 19509 10984
rect 7611 10933 7653 10942
rect 8131 10940 8189 10941
rect 6603 10891 6645 10900
rect 8131 10900 8140 10940
rect 8180 10900 8189 10940
rect 8131 10899 8189 10900
rect 18891 10940 18933 10949
rect 18891 10900 18892 10940
rect 18932 10900 18933 10940
rect 18891 10891 18933 10900
rect 1517 10888 1575 10889
rect 1323 10772 1365 10781
rect 1323 10732 1324 10772
rect 1364 10732 1365 10772
rect 1323 10723 1365 10732
rect 3531 10772 3573 10781
rect 3531 10732 3532 10772
rect 3572 10732 3573 10772
rect 3531 10723 3573 10732
rect 7947 10772 7989 10781
rect 7947 10732 7948 10772
rect 7988 10732 7989 10772
rect 7947 10723 7989 10732
rect 1152 10604 20352 10628
rect 1152 10564 3688 10604
rect 3728 10564 3770 10604
rect 3810 10564 3852 10604
rect 3892 10564 3934 10604
rect 3974 10564 4016 10604
rect 4056 10564 18808 10604
rect 18848 10564 18890 10604
rect 18930 10564 18972 10604
rect 19012 10564 19054 10604
rect 19094 10564 19136 10604
rect 19176 10564 20352 10604
rect 1152 10540 20352 10564
rect 1419 10436 1461 10445
rect 1419 10396 1420 10436
rect 1460 10396 1461 10436
rect 1419 10387 1461 10396
rect 6123 10436 6165 10445
rect 6123 10396 6124 10436
rect 6164 10396 6165 10436
rect 6123 10387 6165 10396
rect 8523 10436 8565 10445
rect 8523 10396 8524 10436
rect 8564 10396 8565 10436
rect 8523 10387 8565 10396
rect 18699 10436 18741 10445
rect 18699 10396 18700 10436
rect 18740 10396 18741 10436
rect 18699 10387 18741 10396
rect 3243 10352 3285 10361
rect 3243 10312 3244 10352
rect 3284 10312 3285 10352
rect 3243 10303 3285 10312
rect 10539 10352 10581 10361
rect 10539 10312 10540 10352
rect 10580 10312 10581 10352
rect 10539 10303 10581 10312
rect 1603 10268 1661 10269
rect 1603 10228 1612 10268
rect 1652 10228 1661 10268
rect 1603 10227 1661 10228
rect 11883 10268 11925 10277
rect 11883 10228 11884 10268
rect 11924 10228 11925 10268
rect 11883 10219 11925 10228
rect 13707 10268 13749 10277
rect 13707 10228 13708 10268
rect 13748 10228 13749 10268
rect 13707 10219 13749 10228
rect 15819 10268 15861 10277
rect 15819 10228 15820 10268
rect 15860 10228 15861 10268
rect 15819 10219 15861 10228
rect 3976 10199 4018 10208
rect 1795 10184 1853 10185
rect 1795 10144 1804 10184
rect 1844 10144 1853 10184
rect 1795 10143 1853 10144
rect 3043 10184 3101 10185
rect 3043 10144 3052 10184
rect 3092 10144 3101 10184
rect 3043 10143 3101 10144
rect 3427 10184 3485 10185
rect 3427 10144 3436 10184
rect 3476 10144 3485 10184
rect 3427 10143 3485 10144
rect 3523 10184 3581 10185
rect 3523 10144 3532 10184
rect 3572 10144 3581 10184
rect 3523 10143 3581 10144
rect 3723 10184 3765 10193
rect 3723 10144 3724 10184
rect 3764 10144 3765 10184
rect 3723 10135 3765 10144
rect 3819 10184 3861 10193
rect 3819 10144 3820 10184
rect 3860 10144 3861 10184
rect 3976 10159 3977 10199
rect 4017 10159 4018 10199
rect 10875 10193 10917 10202
rect 14811 10193 14853 10202
rect 16923 10193 16965 10202
rect 3976 10150 4018 10159
rect 4203 10184 4245 10193
rect 3819 10135 3861 10144
rect 4203 10144 4204 10184
rect 4244 10144 4245 10184
rect 4203 10135 4245 10144
rect 4299 10184 4341 10193
rect 4299 10144 4300 10184
rect 4340 10144 4341 10184
rect 4299 10135 4341 10144
rect 4675 10184 4733 10185
rect 4675 10144 4684 10184
rect 4724 10144 4733 10184
rect 4675 10143 4733 10144
rect 5923 10184 5981 10185
rect 5923 10144 5932 10184
rect 5972 10144 5981 10184
rect 5923 10143 5981 10144
rect 7075 10184 7133 10185
rect 7075 10144 7084 10184
rect 7124 10144 7133 10184
rect 7075 10143 7133 10144
rect 8323 10184 8381 10185
rect 8323 10144 8332 10184
rect 8372 10144 8381 10184
rect 8323 10143 8381 10144
rect 9091 10184 9149 10185
rect 9091 10144 9100 10184
rect 9140 10144 9149 10184
rect 9091 10143 9149 10144
rect 10339 10184 10397 10185
rect 10339 10144 10348 10184
rect 10388 10144 10397 10184
rect 10875 10153 10876 10193
rect 10916 10153 10917 10193
rect 10875 10144 10917 10153
rect 11395 10184 11453 10185
rect 11395 10144 11404 10184
rect 11444 10144 11453 10184
rect 10339 10143 10397 10144
rect 11395 10143 11453 10144
rect 11979 10184 12021 10193
rect 11979 10144 11980 10184
rect 12020 10144 12021 10184
rect 11979 10135 12021 10144
rect 12363 10184 12405 10193
rect 12363 10144 12364 10184
rect 12404 10144 12405 10184
rect 12363 10135 12405 10144
rect 12459 10184 12501 10193
rect 12459 10144 12460 10184
rect 12500 10144 12501 10184
rect 12459 10135 12501 10144
rect 13227 10184 13269 10193
rect 13227 10144 13228 10184
rect 13268 10144 13269 10184
rect 13227 10135 13269 10144
rect 13323 10184 13365 10193
rect 13323 10144 13324 10184
rect 13364 10144 13365 10184
rect 13323 10135 13365 10144
rect 13803 10184 13845 10193
rect 13803 10144 13804 10184
rect 13844 10144 13845 10184
rect 13803 10135 13845 10144
rect 14275 10184 14333 10185
rect 14275 10144 14284 10184
rect 14324 10144 14333 10184
rect 14811 10153 14812 10193
rect 14852 10153 14853 10193
rect 14811 10144 14853 10153
rect 15339 10184 15381 10193
rect 15339 10144 15340 10184
rect 15380 10144 15381 10184
rect 14275 10143 14333 10144
rect 15339 10135 15381 10144
rect 15435 10184 15477 10193
rect 15435 10144 15436 10184
rect 15476 10144 15477 10184
rect 15435 10135 15477 10144
rect 15915 10184 15957 10193
rect 15915 10144 15916 10184
rect 15956 10144 15957 10184
rect 15915 10135 15957 10144
rect 16387 10184 16445 10185
rect 16387 10144 16396 10184
rect 16436 10144 16445 10184
rect 16923 10153 16924 10193
rect 16964 10153 16965 10193
rect 16923 10144 16965 10153
rect 17251 10184 17309 10185
rect 17251 10144 17260 10184
rect 17300 10144 17309 10184
rect 16387 10143 16445 10144
rect 17251 10143 17309 10144
rect 18499 10184 18557 10185
rect 18499 10144 18508 10184
rect 18548 10144 18557 10184
rect 18499 10143 18557 10144
rect 17067 10058 17109 10067
rect 3619 10016 3677 10017
rect 3619 9976 3628 10016
rect 3668 9976 3677 10016
rect 3619 9975 3677 9976
rect 4483 10016 4541 10017
rect 4483 9976 4492 10016
rect 4532 9976 4541 10016
rect 4483 9975 4541 9976
rect 10731 10016 10773 10025
rect 10731 9976 10732 10016
rect 10772 9976 10773 10016
rect 10731 9967 10773 9976
rect 14955 10016 14997 10025
rect 14955 9976 14956 10016
rect 14996 9976 14997 10016
rect 17067 10018 17068 10058
rect 17108 10018 17109 10058
rect 17067 10009 17109 10018
rect 14955 9967 14997 9976
rect 1152 9848 20452 9872
rect 1152 9808 4928 9848
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 5296 9808 20048 9848
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20416 9808 20452 9848
rect 1152 9784 20452 9808
rect 1899 9680 1941 9689
rect 1899 9640 1900 9680
rect 1940 9640 1941 9680
rect 1899 9631 1941 9640
rect 2283 9680 2325 9689
rect 2283 9640 2284 9680
rect 2324 9640 2325 9680
rect 2283 9631 2325 9640
rect 3339 9680 3381 9689
rect 3339 9640 3340 9680
rect 3380 9640 3381 9680
rect 3339 9631 3381 9640
rect 7755 9680 7797 9689
rect 7755 9640 7756 9680
rect 7796 9640 7797 9680
rect 7755 9631 7797 9640
rect 10347 9680 10389 9689
rect 10347 9640 10348 9680
rect 10388 9640 10389 9680
rect 10347 9631 10389 9640
rect 13419 9680 13461 9689
rect 13419 9640 13420 9680
rect 13460 9640 13461 9680
rect 13419 9631 13461 9640
rect 15051 9680 15093 9689
rect 15051 9640 15052 9680
rect 15092 9640 15093 9680
rect 15051 9631 15093 9640
rect 17259 9680 17301 9689
rect 17259 9640 17260 9680
rect 17300 9640 17301 9680
rect 17259 9631 17301 9640
rect 2763 9512 2805 9521
rect 2763 9472 2764 9512
rect 2804 9472 2805 9512
rect 2763 9463 2805 9472
rect 2859 9512 2901 9521
rect 2859 9472 2860 9512
rect 2900 9472 2901 9512
rect 2859 9463 2901 9472
rect 3051 9512 3093 9521
rect 3051 9472 3052 9512
rect 3092 9472 3093 9512
rect 3051 9463 3093 9472
rect 3243 9512 3285 9521
rect 3243 9472 3244 9512
rect 3284 9472 3285 9512
rect 3243 9463 3285 9472
rect 3435 9512 3477 9521
rect 3435 9472 3436 9512
rect 3476 9472 3477 9512
rect 3435 9463 3477 9472
rect 3531 9512 3573 9521
rect 3531 9472 3532 9512
rect 3572 9472 3573 9512
rect 3531 9463 3573 9472
rect 4107 9512 4149 9521
rect 4107 9472 4108 9512
rect 4148 9472 4149 9512
rect 4107 9463 4149 9472
rect 4299 9512 4341 9521
rect 4299 9472 4300 9512
rect 4340 9472 4341 9512
rect 4299 9463 4341 9472
rect 4395 9512 4437 9521
rect 4395 9472 4396 9512
rect 4436 9472 4437 9512
rect 4395 9463 4437 9472
rect 4579 9512 4637 9513
rect 4579 9472 4588 9512
rect 4628 9472 4637 9512
rect 4579 9471 4637 9472
rect 4675 9512 4733 9513
rect 4675 9472 4684 9512
rect 4724 9472 4733 9512
rect 4675 9471 4733 9472
rect 4875 9512 4917 9521
rect 4875 9472 4876 9512
rect 4916 9472 4917 9512
rect 4875 9463 4917 9472
rect 4971 9512 5013 9521
rect 4971 9472 4972 9512
rect 5012 9472 5013 9512
rect 4971 9463 5013 9472
rect 5064 9512 5122 9513
rect 5064 9472 5073 9512
rect 5113 9472 5122 9512
rect 5064 9471 5122 9472
rect 6307 9512 6365 9513
rect 6307 9472 6316 9512
rect 6356 9472 6365 9512
rect 6307 9471 6365 9472
rect 7555 9512 7613 9513
rect 7555 9472 7564 9512
rect 7604 9472 7613 9512
rect 7555 9471 7613 9472
rect 7947 9512 7989 9521
rect 7947 9472 7948 9512
rect 7988 9472 7989 9512
rect 7947 9463 7989 9472
rect 8139 9512 8181 9521
rect 8139 9472 8140 9512
rect 8180 9472 8181 9512
rect 8139 9463 8181 9472
rect 8235 9512 8277 9521
rect 8235 9472 8236 9512
rect 8276 9472 8277 9512
rect 8235 9463 8277 9472
rect 8611 9512 8669 9513
rect 8611 9472 8620 9512
rect 8660 9472 8669 9512
rect 8611 9471 8669 9472
rect 9859 9512 9917 9513
rect 9859 9472 9868 9512
rect 9908 9472 9917 9512
rect 9859 9471 9917 9472
rect 10531 9512 10589 9513
rect 10531 9472 10540 9512
rect 10580 9472 10589 9512
rect 10531 9471 10589 9472
rect 11779 9512 11837 9513
rect 11779 9472 11788 9512
rect 11828 9472 11837 9512
rect 11779 9471 11837 9472
rect 13219 9512 13277 9513
rect 13219 9472 13228 9512
rect 13268 9472 13277 9512
rect 13219 9471 13277 9472
rect 13603 9512 13661 9513
rect 13603 9472 13612 9512
rect 13652 9472 13661 9512
rect 13603 9471 13661 9472
rect 14851 9512 14909 9513
rect 14851 9472 14860 9512
rect 14900 9472 14909 9512
rect 14851 9471 14909 9472
rect 15811 9512 15869 9513
rect 15811 9472 15820 9512
rect 15860 9472 15869 9512
rect 15811 9471 15869 9472
rect 17059 9512 17117 9513
rect 17059 9472 17068 9512
rect 17108 9472 17117 9512
rect 17059 9471 17117 9472
rect 17731 9512 17789 9513
rect 17731 9472 17740 9512
rect 17780 9472 17789 9512
rect 17731 9471 17789 9472
rect 18979 9512 19037 9513
rect 18979 9472 18988 9512
rect 19028 9472 19037 9512
rect 18979 9471 19037 9472
rect 11971 9470 12029 9471
rect 11971 9430 11980 9470
rect 12020 9430 12029 9470
rect 11971 9429 12029 9430
rect 1699 9428 1757 9429
rect 1699 9388 1708 9428
rect 1748 9388 1757 9428
rect 1699 9387 1757 9388
rect 2083 9428 2141 9429
rect 2083 9388 2092 9428
rect 2132 9388 2141 9428
rect 2083 9387 2141 9388
rect 2467 9428 2525 9429
rect 2467 9388 2476 9428
rect 2516 9388 2525 9428
rect 2467 9387 2525 9388
rect 2955 9344 2997 9353
rect 2955 9304 2956 9344
rect 2996 9304 2997 9344
rect 2955 9295 2997 9304
rect 4387 9344 4445 9345
rect 4387 9304 4396 9344
rect 4436 9304 4445 9344
rect 4387 9303 4445 9304
rect 8227 9344 8285 9345
rect 8227 9304 8236 9344
rect 8276 9304 8285 9344
rect 8227 9303 8285 9304
rect 1515 9260 1557 9269
rect 1515 9220 1516 9260
rect 1556 9220 1557 9260
rect 1515 9211 1557 9220
rect 4587 9260 4629 9269
rect 4587 9220 4588 9260
rect 4628 9220 4629 9260
rect 4587 9211 4629 9220
rect 8427 9260 8469 9269
rect 8427 9220 8428 9260
rect 8468 9220 8469 9260
rect 8427 9211 8469 9220
rect 19179 9260 19221 9269
rect 19179 9220 19180 9260
rect 19220 9220 19221 9260
rect 19179 9211 19221 9220
rect 1152 9092 20352 9116
rect 1152 9052 3688 9092
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 4056 9052 18808 9092
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 19176 9052 20352 9092
rect 1152 9028 20352 9052
rect 3723 8840 3765 8849
rect 3723 8800 3724 8840
rect 3764 8800 3765 8840
rect 3723 8791 3765 8800
rect 8331 8840 8373 8849
rect 8331 8800 8332 8840
rect 8372 8800 8373 8840
rect 8331 8791 8373 8800
rect 15627 8840 15669 8849
rect 15627 8800 15628 8840
rect 15668 8800 15669 8840
rect 15627 8791 15669 8800
rect 1699 8756 1757 8757
rect 1699 8716 1708 8756
rect 1748 8716 1757 8756
rect 1699 8715 1757 8716
rect 2083 8756 2141 8757
rect 2083 8716 2092 8756
rect 2132 8716 2141 8756
rect 2083 8715 2141 8716
rect 3907 8756 3965 8757
rect 3907 8716 3916 8756
rect 3956 8716 3965 8756
rect 3907 8715 3965 8716
rect 6987 8756 7029 8765
rect 6987 8716 6988 8756
rect 7028 8716 7029 8756
rect 6987 8707 7029 8716
rect 17931 8756 17973 8765
rect 17931 8716 17932 8756
rect 17972 8716 17973 8756
rect 17931 8707 17973 8716
rect 18027 8756 18069 8765
rect 18027 8716 18028 8756
rect 18068 8716 18069 8756
rect 18027 8707 18069 8716
rect 10504 8687 10546 8696
rect 2667 8672 2709 8681
rect 2667 8632 2668 8672
rect 2708 8632 2709 8672
rect 2667 8623 2709 8632
rect 2763 8672 2805 8681
rect 2763 8632 2764 8672
rect 2804 8632 2805 8672
rect 2763 8623 2805 8632
rect 2947 8672 3005 8673
rect 2947 8632 2956 8672
rect 2996 8632 3005 8672
rect 2947 8631 3005 8632
rect 3043 8672 3101 8673
rect 3043 8632 3052 8672
rect 3092 8632 3101 8672
rect 3043 8631 3101 8632
rect 3243 8672 3285 8681
rect 3243 8632 3244 8672
rect 3284 8632 3285 8672
rect 3243 8623 3285 8632
rect 3339 8672 3381 8681
rect 5931 8677 5973 8686
rect 3339 8632 3340 8672
rect 3380 8632 3381 8672
rect 3339 8623 3381 8632
rect 3459 8672 3517 8673
rect 3459 8632 3468 8672
rect 3508 8632 3517 8672
rect 3459 8631 3517 8632
rect 4099 8672 4157 8673
rect 4099 8632 4108 8672
rect 4148 8632 4157 8672
rect 4099 8631 4157 8632
rect 5347 8672 5405 8673
rect 5347 8632 5356 8672
rect 5396 8632 5405 8672
rect 5347 8631 5405 8632
rect 5931 8637 5932 8677
rect 5972 8637 5973 8677
rect 5931 8628 5973 8637
rect 6403 8672 6461 8673
rect 6403 8632 6412 8672
rect 6452 8632 6461 8672
rect 6403 8631 6461 8632
rect 6891 8672 6933 8681
rect 6891 8632 6892 8672
rect 6932 8632 6933 8672
rect 6891 8623 6933 8632
rect 7371 8672 7413 8681
rect 7371 8632 7372 8672
rect 7412 8632 7413 8672
rect 7371 8623 7413 8632
rect 7467 8672 7509 8681
rect 7467 8632 7468 8672
rect 7508 8632 7509 8672
rect 7467 8623 7509 8632
rect 8515 8672 8573 8673
rect 8515 8632 8524 8672
rect 8564 8632 8573 8672
rect 8515 8631 8573 8632
rect 9763 8672 9821 8673
rect 9763 8632 9772 8672
rect 9812 8632 9821 8672
rect 9763 8631 9821 8632
rect 9955 8672 10013 8673
rect 9955 8632 9964 8672
rect 10004 8632 10013 8672
rect 9955 8631 10013 8632
rect 10051 8672 10109 8673
rect 10051 8632 10060 8672
rect 10100 8632 10109 8672
rect 10051 8631 10109 8632
rect 10251 8672 10293 8681
rect 10251 8632 10252 8672
rect 10292 8632 10293 8672
rect 10251 8623 10293 8632
rect 10347 8672 10389 8681
rect 10347 8632 10348 8672
rect 10388 8632 10389 8672
rect 10504 8647 10505 8687
rect 10545 8647 10546 8687
rect 12411 8681 12453 8690
rect 19035 8681 19077 8690
rect 10504 8638 10546 8647
rect 10827 8672 10869 8681
rect 10347 8623 10389 8632
rect 10827 8632 10828 8672
rect 10868 8632 10869 8672
rect 10827 8623 10869 8632
rect 10923 8672 10965 8681
rect 10923 8632 10924 8672
rect 10964 8632 10965 8672
rect 10923 8623 10965 8632
rect 11307 8672 11349 8681
rect 11307 8632 11308 8672
rect 11348 8632 11349 8672
rect 11307 8623 11349 8632
rect 11403 8672 11445 8681
rect 11403 8632 11404 8672
rect 11444 8632 11445 8672
rect 11403 8623 11445 8632
rect 11875 8672 11933 8673
rect 11875 8632 11884 8672
rect 11924 8632 11933 8672
rect 12411 8641 12412 8681
rect 12452 8641 12453 8681
rect 12411 8632 12453 8641
rect 14179 8672 14237 8673
rect 14179 8632 14188 8672
rect 14228 8632 14237 8672
rect 11875 8631 11933 8632
rect 14179 8631 14237 8632
rect 15427 8672 15485 8673
rect 15427 8632 15436 8672
rect 15476 8632 15485 8672
rect 15427 8631 15485 8632
rect 17451 8672 17493 8681
rect 17451 8632 17452 8672
rect 17492 8632 17493 8672
rect 17451 8623 17493 8632
rect 17547 8672 17589 8681
rect 17547 8632 17548 8672
rect 17588 8632 17589 8672
rect 17547 8623 17589 8632
rect 18499 8672 18557 8673
rect 18499 8632 18508 8672
rect 18548 8632 18557 8672
rect 19035 8641 19036 8681
rect 19076 8641 19077 8681
rect 19035 8632 19077 8641
rect 18499 8631 18557 8632
rect 5547 8588 5589 8597
rect 5547 8548 5548 8588
rect 5588 8548 5589 8588
rect 5547 8539 5589 8548
rect 12555 8588 12597 8597
rect 12555 8548 12556 8588
rect 12596 8548 12597 8588
rect 12555 8539 12597 8548
rect 1515 8504 1557 8513
rect 1515 8464 1516 8504
rect 1556 8464 1557 8504
rect 1515 8455 1557 8464
rect 1899 8504 1941 8513
rect 1899 8464 1900 8504
rect 1940 8464 1941 8504
rect 1899 8455 1941 8464
rect 2467 8504 2525 8505
rect 2467 8464 2476 8504
rect 2516 8464 2525 8504
rect 2467 8463 2525 8464
rect 3427 8504 3485 8505
rect 3427 8464 3436 8504
rect 3476 8464 3485 8504
rect 3427 8463 3485 8464
rect 5739 8504 5781 8513
rect 5739 8464 5740 8504
rect 5780 8464 5781 8504
rect 5739 8455 5781 8464
rect 10147 8504 10205 8505
rect 10147 8464 10156 8504
rect 10196 8464 10205 8504
rect 10147 8463 10205 8464
rect 19179 8504 19221 8513
rect 19179 8464 19180 8504
rect 19220 8464 19221 8504
rect 19179 8455 19221 8464
rect 1152 8336 20452 8360
rect 1152 8296 4928 8336
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 5296 8296 20048 8336
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20416 8296 20452 8336
rect 1152 8272 20452 8296
rect 1227 8168 1269 8177
rect 1227 8128 1228 8168
rect 1268 8128 1269 8168
rect 1227 8119 1269 8128
rect 3051 8168 3093 8177
rect 3051 8128 3052 8168
rect 3092 8128 3093 8168
rect 3051 8119 3093 8128
rect 5067 8168 5109 8177
rect 5067 8128 5068 8168
rect 5108 8128 5109 8168
rect 5067 8119 5109 8128
rect 6699 8168 6741 8177
rect 6699 8128 6700 8168
rect 6740 8128 6741 8168
rect 6699 8119 6741 8128
rect 10635 8168 10677 8177
rect 10635 8128 10636 8168
rect 10676 8128 10677 8168
rect 10635 8119 10677 8128
rect 12459 8168 12501 8177
rect 12459 8128 12460 8168
rect 12500 8128 12501 8168
rect 12459 8119 12501 8128
rect 14571 8168 14613 8177
rect 14571 8128 14572 8168
rect 14612 8128 14613 8168
rect 14571 8119 14613 8128
rect 16779 8168 16821 8177
rect 16779 8128 16780 8168
rect 16820 8128 16821 8168
rect 16779 8119 16821 8128
rect 16971 8168 17013 8177
rect 16971 8128 16972 8168
rect 17012 8128 17013 8168
rect 16971 8119 17013 8128
rect 8715 8084 8757 8093
rect 8715 8044 8716 8084
rect 8756 8044 8757 8084
rect 8715 8035 8757 8044
rect 1603 8000 1661 8001
rect 1603 7960 1612 8000
rect 1652 7960 1661 8000
rect 1603 7959 1661 7960
rect 2851 8000 2909 8001
rect 2851 7960 2860 8000
rect 2900 7960 2909 8000
rect 2851 7959 2909 7960
rect 3619 8000 3677 8001
rect 3619 7960 3628 8000
rect 3668 7960 3677 8000
rect 3619 7959 3677 7960
rect 4867 8000 4925 8001
rect 4867 7960 4876 8000
rect 4916 7960 4925 8000
rect 4867 7959 4925 7960
rect 5251 8000 5309 8001
rect 5251 7960 5260 8000
rect 5300 7960 5309 8000
rect 5251 7959 5309 7960
rect 6499 8000 6557 8001
rect 6499 7960 6508 8000
rect 6548 7960 6557 8000
rect 6499 7959 6557 7960
rect 6987 8000 7029 8009
rect 6987 7960 6988 8000
rect 7028 7960 7029 8000
rect 6987 7951 7029 7960
rect 7083 8000 7125 8009
rect 7083 7960 7084 8000
rect 7124 7960 7125 8000
rect 7083 7951 7125 7960
rect 7467 8000 7509 8009
rect 7467 7960 7468 8000
rect 7508 7960 7509 8000
rect 7467 7951 7509 7960
rect 7563 8000 7605 8009
rect 7563 7960 7564 8000
rect 7604 7960 7605 8000
rect 7563 7951 7605 7960
rect 8035 8000 8093 8001
rect 8035 7960 8044 8000
rect 8084 7960 8093 8000
rect 9187 8000 9245 8001
rect 8035 7959 8093 7960
rect 8571 7958 8613 7967
rect 9187 7960 9196 8000
rect 9236 7960 9245 8000
rect 9187 7959 9245 7960
rect 10435 8000 10493 8001
rect 10435 7960 10444 8000
rect 10484 7960 10493 8000
rect 10435 7959 10493 7960
rect 11011 8000 11069 8001
rect 11011 7960 11020 8000
rect 11060 7960 11069 8000
rect 11011 7959 11069 7960
rect 12259 8000 12317 8001
rect 12259 7960 12268 8000
rect 12308 7960 12317 8000
rect 12259 7959 12317 7960
rect 12843 8000 12885 8009
rect 12843 7960 12844 8000
rect 12884 7960 12885 8000
rect 8571 7918 8572 7958
rect 8612 7918 8613 7958
rect 12843 7951 12885 7960
rect 12939 8000 12981 8009
rect 12939 7960 12940 8000
rect 12980 7960 12981 8000
rect 12939 7951 12981 7960
rect 13891 8000 13949 8001
rect 13891 7960 13900 8000
rect 13940 7960 13949 8000
rect 15051 8000 15093 8009
rect 13891 7959 13949 7960
rect 14427 7958 14469 7967
rect 1411 7916 1469 7917
rect 1411 7876 1420 7916
rect 1460 7876 1469 7916
rect 1411 7875 1469 7876
rect 3427 7916 3485 7917
rect 3427 7876 3436 7916
rect 3476 7876 3485 7916
rect 8571 7909 8613 7918
rect 13323 7916 13365 7925
rect 3427 7875 3485 7876
rect 13323 7876 13324 7916
rect 13364 7876 13365 7916
rect 13323 7867 13365 7876
rect 13419 7916 13461 7925
rect 13419 7876 13420 7916
rect 13460 7876 13461 7916
rect 14427 7918 14428 7958
rect 14468 7918 14469 7958
rect 15051 7960 15052 8000
rect 15092 7960 15093 8000
rect 15051 7951 15093 7960
rect 15147 8000 15189 8009
rect 15147 7960 15148 8000
rect 15188 7960 15189 8000
rect 15147 7951 15189 7960
rect 16099 8000 16157 8001
rect 16099 7960 16108 8000
rect 16148 7960 16157 8000
rect 17155 8000 17213 8001
rect 16099 7959 16157 7960
rect 16635 7958 16677 7967
rect 17155 7960 17164 8000
rect 17204 7960 17213 8000
rect 17155 7959 17213 7960
rect 18403 8000 18461 8001
rect 18403 7960 18412 8000
rect 18452 7960 18461 8000
rect 18403 7959 18461 7960
rect 14427 7909 14469 7918
rect 15531 7916 15573 7925
rect 13419 7867 13461 7876
rect 15531 7876 15532 7916
rect 15572 7876 15573 7916
rect 15531 7867 15573 7876
rect 15627 7916 15669 7925
rect 15627 7876 15628 7916
rect 15668 7876 15669 7916
rect 16635 7918 16636 7958
rect 16676 7918 16677 7958
rect 16635 7909 16677 7918
rect 18787 7916 18845 7917
rect 15627 7867 15669 7876
rect 18787 7876 18796 7916
rect 18836 7876 18845 7916
rect 18787 7875 18845 7876
rect 3243 7832 3285 7841
rect 3243 7792 3244 7832
rect 3284 7792 3285 7832
rect 3243 7783 3285 7792
rect 18603 7748 18645 7757
rect 18603 7708 18604 7748
rect 18644 7708 18645 7748
rect 18603 7699 18645 7708
rect 1152 7580 20352 7604
rect 1152 7540 3688 7580
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 4056 7540 18808 7580
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 19176 7540 20352 7580
rect 1152 7516 20352 7540
rect 2955 7412 2997 7421
rect 2955 7372 2956 7412
rect 2996 7372 2997 7412
rect 2955 7363 2997 7372
rect 7179 7412 7221 7421
rect 7179 7372 7180 7412
rect 7220 7372 7221 7412
rect 7179 7363 7221 7372
rect 8811 7412 8853 7421
rect 8811 7372 8812 7412
rect 8852 7372 8853 7412
rect 8811 7363 8853 7372
rect 12939 7412 12981 7421
rect 12939 7372 12940 7412
rect 12980 7372 12981 7412
rect 12939 7363 12981 7372
rect 14571 7412 14613 7421
rect 14571 7372 14572 7412
rect 14612 7372 14613 7412
rect 14571 7363 14613 7372
rect 14763 7412 14805 7421
rect 14763 7372 14764 7412
rect 14804 7372 14805 7412
rect 14763 7363 14805 7372
rect 10635 7328 10677 7337
rect 10635 7288 10636 7328
rect 10676 7288 10677 7328
rect 10635 7279 10677 7288
rect 3331 7244 3389 7245
rect 3331 7204 3340 7244
rect 3380 7204 3389 7244
rect 3331 7203 3389 7204
rect 1507 7160 1565 7161
rect 1507 7120 1516 7160
rect 1556 7120 1565 7160
rect 1507 7119 1565 7120
rect 2755 7160 2813 7161
rect 2755 7120 2764 7160
rect 2804 7120 2813 7160
rect 2755 7119 2813 7120
rect 3523 7160 3581 7161
rect 3523 7120 3532 7160
rect 3572 7120 3581 7160
rect 3523 7119 3581 7120
rect 4771 7160 4829 7161
rect 4771 7120 4780 7160
rect 4820 7120 4829 7160
rect 4771 7119 4829 7120
rect 5163 7160 5205 7169
rect 5163 7120 5164 7160
rect 5204 7120 5205 7160
rect 5163 7111 5205 7120
rect 5259 7160 5301 7169
rect 10834 7165 10876 7174
rect 11122 7165 11164 7174
rect 5259 7120 5260 7160
rect 5300 7120 5301 7160
rect 5259 7111 5301 7120
rect 5731 7160 5789 7161
rect 5731 7120 5740 7160
rect 5780 7120 5789 7160
rect 5731 7119 5789 7120
rect 6979 7160 7037 7161
rect 6979 7120 6988 7160
rect 7028 7120 7037 7160
rect 6979 7119 7037 7120
rect 7363 7160 7421 7161
rect 7363 7120 7372 7160
rect 7412 7120 7421 7160
rect 7363 7119 7421 7120
rect 8611 7160 8669 7161
rect 8611 7120 8620 7160
rect 8660 7120 8669 7160
rect 8611 7119 8669 7120
rect 9187 7160 9245 7161
rect 9187 7120 9196 7160
rect 9236 7120 9245 7160
rect 9187 7119 9245 7120
rect 10435 7160 10493 7161
rect 10435 7120 10444 7160
rect 10484 7120 10493 7160
rect 10435 7119 10493 7120
rect 10834 7125 10835 7165
rect 10875 7125 10876 7165
rect 10834 7116 10876 7125
rect 10930 7156 10972 7165
rect 10930 7116 10931 7156
rect 10971 7116 10972 7156
rect 11122 7125 11123 7165
rect 11163 7125 11164 7165
rect 11122 7116 11164 7125
rect 11491 7160 11549 7161
rect 11491 7120 11500 7160
rect 11540 7120 11549 7160
rect 11491 7119 11549 7120
rect 12739 7160 12797 7161
rect 12739 7120 12748 7160
rect 12788 7120 12797 7160
rect 12739 7119 12797 7120
rect 13123 7160 13181 7161
rect 13123 7120 13132 7160
rect 13172 7120 13181 7160
rect 13123 7119 13181 7120
rect 14371 7160 14429 7161
rect 14371 7120 14380 7160
rect 14420 7120 14429 7160
rect 14371 7119 14429 7120
rect 14947 7160 15005 7161
rect 14947 7120 14956 7160
rect 14996 7120 15005 7160
rect 14947 7119 15005 7120
rect 16195 7160 16253 7161
rect 16195 7120 16204 7160
rect 16244 7120 16253 7160
rect 16195 7119 16253 7120
rect 10930 7107 10972 7116
rect 3147 6992 3189 7001
rect 3147 6952 3148 6992
rect 3188 6952 3189 6992
rect 3147 6943 3189 6952
rect 4971 6992 5013 7001
rect 4971 6952 4972 6992
rect 5012 6952 5013 6992
rect 4971 6943 5013 6952
rect 5443 6992 5501 6993
rect 5443 6952 5452 6992
rect 5492 6952 5501 6992
rect 5443 6951 5501 6952
rect 11019 6992 11061 7001
rect 11019 6952 11020 6992
rect 11060 6952 11061 6992
rect 11019 6943 11061 6952
rect 1152 6824 20452 6848
rect 1152 6784 4928 6824
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 5296 6784 20048 6824
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20416 6784 20452 6824
rect 1152 6760 20452 6784
rect 1323 6656 1365 6665
rect 1323 6616 1324 6656
rect 1364 6616 1365 6656
rect 1323 6607 1365 6616
rect 1707 6656 1749 6665
rect 1707 6616 1708 6656
rect 1748 6616 1749 6656
rect 1707 6607 1749 6616
rect 4291 6656 4349 6657
rect 4291 6616 4300 6656
rect 4340 6616 4349 6656
rect 4291 6615 4349 6616
rect 6787 6656 6845 6657
rect 6787 6616 6796 6656
rect 6836 6616 6845 6656
rect 6787 6615 6845 6616
rect 8707 6656 8765 6657
rect 8707 6616 8716 6656
rect 8756 6616 8765 6656
rect 8707 6615 8765 6616
rect 11683 6656 11741 6657
rect 11683 6616 11692 6656
rect 11732 6616 11741 6656
rect 11683 6615 11741 6616
rect 14283 6656 14325 6665
rect 14283 6616 14284 6656
rect 14324 6616 14325 6656
rect 14283 6607 14325 6616
rect 16875 6656 16917 6665
rect 16875 6616 16876 6656
rect 16916 6616 16917 6656
rect 16875 6607 16917 6616
rect 2187 6572 2229 6581
rect 2187 6532 2188 6572
rect 2228 6532 2229 6572
rect 2187 6523 2229 6532
rect 9195 6572 9237 6581
rect 9195 6532 9196 6572
rect 9236 6532 9237 6572
rect 9195 6523 9237 6532
rect 2091 6488 2133 6497
rect 2091 6448 2092 6488
rect 2132 6448 2133 6488
rect 2091 6439 2133 6448
rect 2283 6488 2325 6497
rect 2283 6448 2284 6488
rect 2324 6448 2325 6488
rect 2283 6439 2325 6448
rect 2379 6488 2421 6497
rect 2379 6448 2380 6488
rect 2420 6448 2421 6488
rect 2379 6439 2421 6448
rect 2563 6488 2621 6489
rect 2563 6448 2572 6488
rect 2612 6448 2621 6488
rect 2563 6447 2621 6448
rect 2659 6488 2717 6489
rect 2659 6448 2668 6488
rect 2708 6448 2717 6488
rect 2659 6447 2717 6448
rect 2859 6488 2901 6497
rect 2859 6448 2860 6488
rect 2900 6448 2901 6488
rect 2859 6439 2901 6448
rect 2955 6488 2997 6497
rect 2955 6448 2956 6488
rect 2996 6448 2997 6488
rect 2955 6439 2997 6448
rect 3048 6488 3106 6489
rect 3048 6448 3057 6488
rect 3097 6448 3106 6488
rect 3048 6447 3106 6448
rect 3627 6488 3669 6497
rect 3627 6448 3628 6488
rect 3668 6448 3669 6488
rect 3627 6439 3669 6448
rect 3819 6488 3861 6497
rect 3819 6448 3820 6488
rect 3860 6448 3861 6488
rect 3819 6439 3861 6448
rect 3915 6488 3957 6497
rect 3915 6448 3916 6488
rect 3956 6448 3957 6488
rect 3915 6439 3957 6448
rect 4099 6488 4157 6489
rect 4099 6448 4108 6488
rect 4148 6448 4157 6488
rect 4099 6447 4157 6448
rect 4195 6488 4253 6489
rect 4195 6448 4204 6488
rect 4244 6448 4253 6488
rect 4195 6447 4253 6448
rect 4395 6488 4437 6497
rect 4395 6448 4396 6488
rect 4436 6448 4437 6488
rect 4395 6439 4437 6448
rect 4491 6488 4533 6497
rect 4491 6448 4492 6488
rect 4532 6448 4533 6488
rect 4491 6439 4533 6448
rect 4584 6488 4642 6489
rect 4584 6448 4593 6488
rect 4633 6448 4642 6488
rect 4584 6447 4642 6448
rect 4867 6488 4925 6489
rect 4867 6448 4876 6488
rect 4916 6448 4925 6488
rect 4867 6447 4925 6448
rect 6115 6488 6173 6489
rect 6115 6448 6124 6488
rect 6164 6448 6173 6488
rect 6115 6447 6173 6448
rect 6507 6488 6549 6497
rect 6507 6448 6508 6488
rect 6548 6448 6549 6488
rect 6507 6439 6549 6448
rect 6603 6488 6645 6497
rect 6603 6448 6604 6488
rect 6644 6448 6645 6488
rect 6603 6439 6645 6448
rect 6979 6488 7037 6489
rect 6979 6448 6988 6488
rect 7028 6448 7037 6488
rect 6979 6447 7037 6448
rect 8227 6488 8285 6489
rect 8227 6448 8236 6488
rect 8276 6448 8285 6488
rect 8227 6447 8285 6448
rect 8907 6488 8949 6497
rect 8907 6448 8908 6488
rect 8948 6448 8949 6488
rect 8907 6439 8949 6448
rect 9003 6488 9045 6497
rect 9003 6448 9004 6488
rect 9044 6448 9045 6488
rect 9003 6439 9045 6448
rect 9379 6488 9437 6489
rect 9379 6448 9388 6488
rect 9428 6448 9437 6488
rect 9379 6447 9437 6448
rect 10627 6488 10685 6489
rect 10627 6448 10636 6488
rect 10676 6448 10685 6488
rect 10627 6447 10685 6448
rect 10819 6488 10877 6489
rect 10819 6448 10828 6488
rect 10868 6448 10877 6488
rect 10819 6447 10877 6448
rect 10915 6488 10973 6489
rect 10915 6448 10924 6488
rect 10964 6448 10973 6488
rect 10915 6447 10973 6448
rect 11115 6488 11157 6497
rect 11115 6448 11116 6488
rect 11156 6448 11157 6488
rect 11115 6439 11157 6448
rect 11211 6488 11253 6497
rect 11211 6448 11212 6488
rect 11252 6448 11253 6488
rect 11211 6439 11253 6448
rect 11368 6481 11410 6490
rect 11787 6488 11829 6497
rect 11368 6441 11369 6481
rect 11409 6441 11410 6481
rect 11368 6432 11410 6441
rect 11629 6473 11671 6482
rect 11629 6433 11630 6473
rect 11670 6433 11671 6473
rect 11787 6448 11788 6488
rect 11828 6448 11829 6488
rect 11787 6439 11829 6448
rect 11883 6488 11925 6497
rect 11883 6448 11884 6488
rect 11924 6448 11925 6488
rect 11883 6439 11925 6448
rect 12067 6488 12125 6489
rect 12067 6448 12076 6488
rect 12116 6448 12125 6488
rect 12067 6447 12125 6448
rect 12163 6488 12221 6489
rect 12163 6448 12172 6488
rect 12212 6448 12221 6488
rect 12163 6447 12221 6448
rect 12555 6488 12597 6497
rect 12555 6448 12556 6488
rect 12596 6448 12597 6488
rect 12555 6439 12597 6448
rect 12651 6488 12693 6497
rect 12651 6448 12652 6488
rect 12692 6448 12693 6488
rect 12651 6439 12693 6448
rect 13131 6488 13173 6497
rect 13131 6448 13132 6488
rect 13172 6448 13173 6488
rect 13131 6439 13173 6448
rect 13603 6488 13661 6489
rect 13603 6448 13612 6488
rect 13652 6448 13661 6488
rect 15427 6488 15485 6489
rect 13603 6447 13661 6448
rect 14139 6478 14181 6487
rect 11629 6424 11671 6433
rect 14139 6438 14140 6478
rect 14180 6438 14181 6478
rect 15427 6448 15436 6488
rect 15476 6448 15485 6488
rect 15427 6447 15485 6448
rect 16675 6488 16733 6489
rect 16675 6448 16684 6488
rect 16724 6448 16733 6488
rect 16675 6447 16733 6448
rect 17155 6488 17213 6489
rect 17155 6448 17164 6488
rect 17204 6448 17213 6488
rect 17155 6447 17213 6448
rect 18403 6488 18461 6489
rect 18403 6448 18412 6488
rect 18452 6448 18461 6488
rect 18403 6447 18461 6448
rect 14139 6429 14181 6438
rect 1507 6404 1565 6405
rect 1507 6364 1516 6404
rect 1556 6364 1565 6404
rect 1507 6363 1565 6364
rect 1891 6404 1949 6405
rect 1891 6364 1900 6404
rect 1940 6364 1949 6404
rect 1891 6363 1949 6364
rect 13035 6404 13077 6413
rect 13035 6364 13036 6404
rect 13076 6364 13077 6404
rect 13035 6355 13077 6364
rect 3907 6320 3965 6321
rect 3907 6280 3916 6320
rect 3956 6280 3965 6320
rect 3907 6279 3965 6280
rect 2571 6236 2613 6245
rect 2571 6196 2572 6236
rect 2612 6196 2613 6236
rect 2571 6187 2613 6196
rect 6315 6236 6357 6245
rect 6315 6196 6316 6236
rect 6356 6196 6357 6236
rect 6315 6187 6357 6196
rect 8427 6236 8469 6245
rect 8427 6196 8428 6236
rect 8468 6196 8469 6236
rect 8427 6187 8469 6196
rect 10827 6236 10869 6245
rect 10827 6196 10828 6236
rect 10868 6196 10869 6236
rect 10827 6187 10869 6196
rect 18603 6236 18645 6245
rect 18603 6196 18604 6236
rect 18644 6196 18645 6236
rect 18603 6187 18645 6196
rect 1152 6068 20352 6092
rect 1152 6028 3688 6068
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 4056 6028 18808 6068
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 19176 6028 20352 6068
rect 1152 6004 20352 6028
rect 4587 5900 4629 5909
rect 4587 5860 4588 5900
rect 4628 5860 4629 5900
rect 4587 5851 4629 5860
rect 6219 5900 6261 5909
rect 6219 5860 6220 5900
rect 6260 5860 6261 5900
rect 6219 5851 6261 5860
rect 12747 5900 12789 5909
rect 12747 5860 12748 5900
rect 12788 5860 12789 5900
rect 12747 5851 12789 5860
rect 14379 5900 14421 5909
rect 14379 5860 14380 5900
rect 14420 5860 14421 5900
rect 14379 5851 14421 5860
rect 2859 5816 2901 5825
rect 2859 5776 2860 5816
rect 2900 5776 2901 5816
rect 2859 5767 2901 5776
rect 6987 5732 7029 5741
rect 6987 5692 6988 5732
rect 7028 5692 7029 5732
rect 6987 5683 7029 5692
rect 7083 5732 7125 5741
rect 7083 5692 7084 5732
rect 7124 5692 7125 5732
rect 7083 5683 7125 5692
rect 17643 5732 17685 5741
rect 17643 5692 17644 5732
rect 17684 5692 17685 5732
rect 17643 5683 17685 5692
rect 17739 5732 17781 5741
rect 17739 5692 17740 5732
rect 17780 5692 17781 5732
rect 17739 5683 17781 5692
rect 8043 5662 8085 5671
rect 1411 5648 1469 5649
rect 1411 5608 1420 5648
rect 1460 5608 1469 5648
rect 1411 5607 1469 5608
rect 2659 5648 2717 5649
rect 2659 5608 2668 5648
rect 2708 5608 2717 5648
rect 2659 5607 2717 5608
rect 3139 5648 3197 5649
rect 3139 5608 3148 5648
rect 3188 5608 3197 5648
rect 3139 5607 3197 5608
rect 4387 5648 4445 5649
rect 4387 5608 4396 5648
rect 4436 5608 4445 5648
rect 4387 5607 4445 5608
rect 4771 5648 4829 5649
rect 4771 5608 4780 5648
rect 4820 5608 4829 5648
rect 4771 5607 4829 5608
rect 6019 5648 6077 5649
rect 6019 5608 6028 5648
rect 6068 5608 6077 5648
rect 6019 5607 6077 5608
rect 6507 5648 6549 5657
rect 6507 5608 6508 5648
rect 6548 5608 6549 5648
rect 6507 5599 6549 5608
rect 6603 5648 6645 5657
rect 6603 5608 6604 5648
rect 6644 5608 6645 5648
rect 6603 5599 6645 5608
rect 7555 5648 7613 5649
rect 7555 5608 7564 5648
rect 7604 5608 7613 5648
rect 8043 5622 8044 5662
rect 8084 5622 8085 5662
rect 10696 5663 10738 5672
rect 8043 5613 8085 5622
rect 8515 5648 8573 5649
rect 7555 5607 7613 5608
rect 8515 5608 8524 5648
rect 8564 5608 8573 5648
rect 8515 5607 8573 5608
rect 9763 5648 9821 5649
rect 9763 5608 9772 5648
rect 9812 5608 9821 5648
rect 9763 5607 9821 5608
rect 10147 5648 10205 5649
rect 10147 5608 10156 5648
rect 10196 5608 10205 5648
rect 10147 5607 10205 5608
rect 10243 5648 10301 5649
rect 10243 5608 10252 5648
rect 10292 5608 10301 5648
rect 10243 5607 10301 5608
rect 10443 5648 10485 5657
rect 10443 5608 10444 5648
rect 10484 5608 10485 5648
rect 10443 5599 10485 5608
rect 10539 5648 10581 5657
rect 10539 5608 10540 5648
rect 10580 5608 10581 5648
rect 10696 5623 10697 5663
rect 10737 5623 10738 5663
rect 16731 5657 16773 5666
rect 18699 5662 18741 5671
rect 10696 5614 10738 5623
rect 11299 5648 11357 5649
rect 10539 5599 10581 5608
rect 11299 5608 11308 5648
rect 11348 5608 11357 5648
rect 11299 5607 11357 5608
rect 12547 5648 12605 5649
rect 12547 5608 12556 5648
rect 12596 5608 12605 5648
rect 12547 5607 12605 5608
rect 12931 5648 12989 5649
rect 12931 5608 12940 5648
rect 12980 5608 12989 5648
rect 12931 5607 12989 5608
rect 14179 5648 14237 5649
rect 14179 5608 14188 5648
rect 14228 5608 14237 5648
rect 14179 5607 14237 5608
rect 15147 5648 15189 5657
rect 15147 5608 15148 5648
rect 15188 5608 15189 5648
rect 15147 5599 15189 5608
rect 15243 5648 15285 5657
rect 15243 5608 15244 5648
rect 15284 5608 15285 5648
rect 15243 5599 15285 5608
rect 15627 5648 15669 5657
rect 15627 5608 15628 5648
rect 15668 5608 15669 5648
rect 15627 5599 15669 5608
rect 15723 5648 15765 5657
rect 15723 5608 15724 5648
rect 15764 5608 15765 5648
rect 15723 5599 15765 5608
rect 16195 5648 16253 5649
rect 16195 5608 16204 5648
rect 16244 5608 16253 5648
rect 16731 5617 16732 5657
rect 16772 5617 16773 5657
rect 16731 5608 16773 5617
rect 17163 5648 17205 5657
rect 17163 5608 17164 5648
rect 17204 5608 17205 5648
rect 16195 5607 16253 5608
rect 17163 5599 17205 5608
rect 17259 5648 17301 5657
rect 17259 5608 17260 5648
rect 17300 5608 17301 5648
rect 17259 5599 17301 5608
rect 18211 5648 18269 5649
rect 18211 5608 18220 5648
rect 18260 5608 18269 5648
rect 18699 5622 18700 5662
rect 18740 5622 18741 5662
rect 18699 5613 18741 5622
rect 18211 5607 18269 5608
rect 16875 5564 16917 5573
rect 16875 5524 16876 5564
rect 16916 5524 16917 5564
rect 16875 5515 16917 5524
rect 6219 5480 6261 5489
rect 6219 5440 6220 5480
rect 6260 5440 6261 5480
rect 6219 5431 6261 5440
rect 8235 5480 8277 5489
rect 8235 5440 8236 5480
rect 8276 5440 8277 5480
rect 8235 5431 8277 5440
rect 9963 5480 10005 5489
rect 9963 5440 9964 5480
rect 10004 5440 10005 5480
rect 9963 5431 10005 5440
rect 10627 5480 10685 5481
rect 10627 5440 10636 5480
rect 10676 5440 10685 5480
rect 10627 5439 10685 5440
rect 18891 5480 18933 5489
rect 18891 5440 18892 5480
rect 18932 5440 18933 5480
rect 18891 5431 18933 5440
rect 1152 5312 20452 5336
rect 1152 5272 4928 5312
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 5296 5272 20048 5312
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20416 5272 20452 5312
rect 1152 5248 20452 5272
rect 2859 5144 2901 5153
rect 2859 5104 2860 5144
rect 2900 5104 2901 5144
rect 2859 5095 2901 5104
rect 5347 5144 5405 5145
rect 5347 5104 5356 5144
rect 5396 5104 5405 5144
rect 5347 5103 5405 5104
rect 10339 5144 10397 5145
rect 10339 5104 10348 5144
rect 10388 5104 10397 5144
rect 10339 5103 10397 5104
rect 12259 5144 12317 5145
rect 12259 5104 12268 5144
rect 12308 5104 12317 5144
rect 12259 5103 12317 5104
rect 15243 5144 15285 5153
rect 15243 5104 15244 5144
rect 15284 5104 15285 5144
rect 15243 5095 15285 5104
rect 16971 5144 17013 5153
rect 16971 5104 16972 5144
rect 17012 5104 17013 5144
rect 16971 5095 17013 5104
rect 4875 5060 4917 5069
rect 4875 5020 4876 5060
rect 4916 5020 4917 5060
rect 4875 5011 4917 5020
rect 7179 5060 7221 5069
rect 7179 5020 7180 5060
rect 7220 5020 7221 5060
rect 7179 5011 7221 5020
rect 9867 5060 9909 5069
rect 9867 5020 9868 5060
rect 9908 5020 9909 5060
rect 9867 5011 9909 5020
rect 12939 5060 12981 5069
rect 12939 5020 12940 5060
rect 12980 5020 12981 5060
rect 12939 5011 12981 5020
rect 1411 4976 1469 4977
rect 1411 4936 1420 4976
rect 1460 4936 1469 4976
rect 1411 4935 1469 4936
rect 2659 4976 2717 4977
rect 2659 4936 2668 4976
rect 2708 4936 2717 4976
rect 2659 4935 2717 4936
rect 3427 4976 3485 4977
rect 3427 4936 3436 4976
rect 3476 4936 3485 4976
rect 3427 4935 3485 4936
rect 5067 4976 5109 4985
rect 5067 4936 5068 4976
rect 5108 4936 5109 4976
rect 4675 4934 4733 4935
rect 4675 4894 4684 4934
rect 4724 4894 4733 4934
rect 5067 4927 5109 4936
rect 5163 4976 5205 4985
rect 5163 4936 5164 4976
rect 5204 4936 5205 4976
rect 5163 4927 5205 4936
rect 5731 4976 5789 4977
rect 5731 4936 5740 4976
rect 5780 4936 5789 4976
rect 5731 4935 5789 4936
rect 6979 4976 7037 4977
rect 6979 4936 6988 4976
rect 7028 4936 7037 4976
rect 6979 4935 7037 4936
rect 7363 4976 7421 4977
rect 7363 4936 7372 4976
rect 7412 4936 7421 4976
rect 7363 4935 7421 4936
rect 7459 4976 7517 4977
rect 7459 4936 7468 4976
rect 7508 4936 7517 4976
rect 7459 4935 7517 4936
rect 7659 4976 7701 4985
rect 7659 4936 7660 4976
rect 7700 4936 7701 4976
rect 7659 4927 7701 4936
rect 7755 4976 7797 4985
rect 7755 4936 7756 4976
rect 7796 4936 7797 4976
rect 7755 4927 7797 4936
rect 7848 4976 7906 4977
rect 7848 4936 7857 4976
rect 7897 4936 7906 4976
rect 7848 4935 7906 4936
rect 8419 4976 8477 4977
rect 8419 4936 8428 4976
rect 8468 4936 8477 4976
rect 8419 4935 8477 4936
rect 9667 4976 9725 4977
rect 9667 4936 9676 4976
rect 9716 4936 9725 4976
rect 9667 4935 9725 4936
rect 10059 4976 10101 4985
rect 10059 4936 10060 4976
rect 10100 4936 10101 4976
rect 10059 4927 10101 4936
rect 10155 4976 10197 4985
rect 10155 4936 10156 4976
rect 10196 4936 10197 4976
rect 10155 4927 10197 4936
rect 10627 4976 10685 4977
rect 10627 4936 10636 4976
rect 10676 4936 10685 4976
rect 10627 4935 10685 4936
rect 11875 4976 11933 4977
rect 11875 4936 11884 4976
rect 11924 4936 11933 4976
rect 11875 4935 11933 4936
rect 12459 4976 12501 4985
rect 12459 4936 12460 4976
rect 12500 4936 12501 4976
rect 12459 4927 12501 4936
rect 12555 4976 12597 4985
rect 12555 4936 12556 4976
rect 12596 4936 12597 4976
rect 12555 4927 12597 4936
rect 12747 4976 12789 4985
rect 12747 4936 12748 4976
rect 12788 4936 12789 4976
rect 12747 4927 12789 4936
rect 12843 4976 12885 4985
rect 12843 4936 12844 4976
rect 12884 4936 12885 4976
rect 12843 4927 12885 4936
rect 13035 4976 13077 4985
rect 13035 4936 13036 4976
rect 13076 4936 13077 4976
rect 13035 4927 13077 4936
rect 13795 4976 13853 4977
rect 13795 4936 13804 4976
rect 13844 4936 13853 4976
rect 13795 4935 13853 4936
rect 15043 4976 15101 4977
rect 15043 4936 15052 4976
rect 15092 4936 15101 4976
rect 15043 4935 15101 4936
rect 15523 4976 15581 4977
rect 15523 4936 15532 4976
rect 15572 4936 15581 4976
rect 15523 4935 15581 4936
rect 16771 4976 16829 4977
rect 16771 4936 16780 4976
rect 16820 4936 16829 4976
rect 16771 4935 16829 4936
rect 4675 4893 4733 4894
rect 3235 4892 3293 4893
rect 3235 4852 3244 4892
rect 3284 4852 3293 4892
rect 3235 4851 3293 4852
rect 3051 4808 3093 4817
rect 3051 4768 3052 4808
rect 3092 4768 3093 4808
rect 3051 4759 3093 4768
rect 12075 4808 12117 4817
rect 12075 4768 12076 4808
rect 12116 4768 12117 4808
rect 12075 4759 12117 4768
rect 7371 4724 7413 4733
rect 7371 4684 7372 4724
rect 7412 4684 7413 4724
rect 7371 4675 7413 4684
rect 1152 4556 20352 4580
rect 1152 4516 3688 4556
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 4056 4516 18808 4556
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 19176 4516 20352 4556
rect 1152 4492 20352 4516
rect 1515 4388 1557 4397
rect 1515 4348 1516 4388
rect 1556 4348 1557 4388
rect 1515 4339 1557 4348
rect 1899 4388 1941 4397
rect 1899 4348 1900 4388
rect 1940 4348 1941 4388
rect 1899 4339 1941 4348
rect 2283 4388 2325 4397
rect 2283 4348 2284 4388
rect 2324 4348 2325 4388
rect 2283 4339 2325 4348
rect 12171 4388 12213 4397
rect 12171 4348 12172 4388
rect 12212 4348 12213 4388
rect 12171 4339 12213 4348
rect 9763 4304 9821 4305
rect 9763 4264 9772 4304
rect 9812 4264 9821 4304
rect 9763 4263 9821 4264
rect 1699 4220 1757 4221
rect 1699 4180 1708 4220
rect 1748 4180 1757 4220
rect 1699 4179 1757 4180
rect 2083 4220 2141 4221
rect 2083 4180 2092 4220
rect 2132 4180 2141 4220
rect 2083 4179 2141 4180
rect 2467 4220 2525 4221
rect 2467 4180 2476 4220
rect 2516 4180 2525 4220
rect 2467 4179 2525 4180
rect 16251 4145 16293 4154
rect 3051 4136 3093 4145
rect 3051 4096 3052 4136
rect 3092 4096 3093 4136
rect 3051 4087 3093 4096
rect 3147 4136 3189 4145
rect 3147 4096 3148 4136
rect 3188 4096 3189 4136
rect 3147 4087 3189 4096
rect 3619 4136 3677 4137
rect 3619 4096 3628 4136
rect 3668 4096 3677 4136
rect 3619 4095 3677 4096
rect 4867 4136 4925 4137
rect 4867 4096 4876 4136
rect 4916 4096 4925 4136
rect 4867 4095 4925 4096
rect 5739 4136 5781 4145
rect 5739 4096 5740 4136
rect 5780 4096 5781 4136
rect 5739 4087 5781 4096
rect 5835 4136 5877 4145
rect 5835 4096 5836 4136
rect 5876 4096 5877 4136
rect 5835 4087 5877 4096
rect 6891 4136 6933 4145
rect 6891 4096 6892 4136
rect 6932 4096 6933 4136
rect 6891 4087 6933 4096
rect 7083 4136 7125 4145
rect 7083 4096 7084 4136
rect 7124 4096 7125 4136
rect 7083 4087 7125 4096
rect 7179 4136 7221 4145
rect 7179 4096 7180 4136
rect 7220 4096 7221 4136
rect 7179 4087 7221 4096
rect 7363 4136 7421 4137
rect 7363 4096 7372 4136
rect 7412 4096 7421 4136
rect 7363 4095 7421 4096
rect 7459 4136 7517 4137
rect 7459 4096 7468 4136
rect 7508 4096 7517 4136
rect 7459 4095 7517 4096
rect 7659 4136 7701 4145
rect 7659 4096 7660 4136
rect 7700 4096 7701 4136
rect 7659 4087 7701 4096
rect 7755 4136 7797 4145
rect 7755 4096 7756 4136
rect 7796 4096 7797 4136
rect 7755 4087 7797 4096
rect 7875 4136 7933 4137
rect 7875 4096 7884 4136
rect 7924 4096 7933 4136
rect 7875 4095 7933 4096
rect 9579 4136 9621 4145
rect 9579 4096 9580 4136
rect 9620 4096 9621 4136
rect 9579 4087 9621 4096
rect 9771 4136 9813 4145
rect 9771 4096 9772 4136
rect 9812 4096 9813 4136
rect 9771 4087 9813 4096
rect 9867 4136 9909 4145
rect 9867 4096 9868 4136
rect 9908 4096 9909 4136
rect 9867 4087 9909 4096
rect 10347 4136 10389 4145
rect 10347 4096 10348 4136
rect 10388 4096 10389 4136
rect 10347 4087 10389 4096
rect 10443 4136 10485 4145
rect 10443 4096 10444 4136
rect 10484 4096 10485 4136
rect 10443 4087 10485 4096
rect 10723 4136 10781 4137
rect 10723 4096 10732 4136
rect 10772 4096 10781 4136
rect 10723 4095 10781 4096
rect 11971 4136 12029 4137
rect 11971 4096 11980 4136
rect 12020 4096 12029 4136
rect 11971 4095 12029 4096
rect 12931 4136 12989 4137
rect 12931 4096 12940 4136
rect 12980 4096 12989 4136
rect 12931 4095 12989 4096
rect 14179 4136 14237 4137
rect 14179 4096 14188 4136
rect 14228 4096 14237 4136
rect 14179 4095 14237 4096
rect 14667 4136 14709 4145
rect 14667 4096 14668 4136
rect 14708 4096 14709 4136
rect 14667 4087 14709 4096
rect 14763 4136 14805 4145
rect 14763 4096 14764 4136
rect 14804 4096 14805 4136
rect 14763 4087 14805 4096
rect 15147 4136 15189 4145
rect 15147 4096 15148 4136
rect 15188 4096 15189 4136
rect 15147 4087 15189 4096
rect 15243 4136 15285 4145
rect 15243 4096 15244 4136
rect 15284 4096 15285 4136
rect 15243 4087 15285 4096
rect 15715 4136 15773 4137
rect 15715 4096 15724 4136
rect 15764 4096 15773 4136
rect 16251 4105 16252 4145
rect 16292 4105 16293 4145
rect 16251 4096 16293 4105
rect 15715 4095 15773 4096
rect 14379 4052 14421 4061
rect 14379 4012 14380 4052
rect 14420 4012 14421 4052
rect 14379 4003 14421 4012
rect 16395 4052 16437 4061
rect 16395 4012 16396 4052
rect 16436 4012 16437 4052
rect 16395 4003 16437 4012
rect 2851 3968 2909 3969
rect 2851 3928 2860 3968
rect 2900 3928 2909 3968
rect 2851 3927 2909 3928
rect 5067 3968 5109 3977
rect 5067 3928 5068 3968
rect 5108 3928 5109 3968
rect 5067 3919 5109 3928
rect 5539 3968 5597 3969
rect 5539 3928 5548 3968
rect 5588 3928 5597 3968
rect 5539 3927 5597 3928
rect 6987 3968 7029 3977
rect 6987 3928 6988 3968
rect 7028 3928 7029 3968
rect 6987 3919 7029 3928
rect 7555 3968 7613 3969
rect 7555 3928 7564 3968
rect 7604 3928 7613 3968
rect 7555 3927 7613 3928
rect 10147 3968 10205 3969
rect 10147 3928 10156 3968
rect 10196 3928 10205 3968
rect 10147 3927 10205 3928
rect 1152 3800 20452 3824
rect 1152 3760 4928 3800
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 5296 3760 20048 3800
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20416 3760 20452 3800
rect 1152 3736 20452 3760
rect 1515 3632 1557 3641
rect 1515 3592 1516 3632
rect 1556 3592 1557 3632
rect 1515 3583 1557 3592
rect 1899 3632 1941 3641
rect 1899 3592 1900 3632
rect 1940 3592 1941 3632
rect 1899 3583 1941 3592
rect 2283 3632 2325 3641
rect 2283 3592 2284 3632
rect 2324 3592 2325 3632
rect 2283 3583 2325 3592
rect 2667 3632 2709 3641
rect 2667 3592 2668 3632
rect 2708 3592 2709 3632
rect 2667 3583 2709 3592
rect 7851 3632 7893 3641
rect 7851 3592 7852 3632
rect 7892 3592 7893 3632
rect 7851 3583 7893 3592
rect 8323 3632 8381 3633
rect 8323 3592 8332 3632
rect 8372 3592 8381 3632
rect 8323 3591 8381 3592
rect 16875 3632 16917 3641
rect 16875 3592 16876 3632
rect 16916 3592 16917 3632
rect 16875 3583 16917 3592
rect 5251 3548 5309 3549
rect 5251 3508 5260 3548
rect 5300 3508 5309 3548
rect 5251 3507 5309 3508
rect 12555 3548 12597 3557
rect 12555 3508 12556 3548
rect 12596 3508 12597 3548
rect 12555 3499 12597 3508
rect 14571 3548 14613 3557
rect 14571 3508 14572 3548
rect 14612 3508 14613 3548
rect 14571 3499 14613 3508
rect 3619 3464 3677 3465
rect 3619 3424 3628 3464
rect 3668 3424 3677 3464
rect 3619 3423 3677 3424
rect 4867 3464 4925 3465
rect 4867 3424 4876 3464
rect 4916 3424 4925 3464
rect 5347 3464 5405 3465
rect 4867 3423 4925 3424
rect 5259 3441 5301 3450
rect 5259 3401 5260 3441
rect 5300 3401 5301 3441
rect 5347 3424 5356 3464
rect 5396 3424 5405 3464
rect 5347 3423 5405 3424
rect 5547 3464 5589 3473
rect 5547 3424 5548 3464
rect 5588 3424 5589 3464
rect 5547 3415 5589 3424
rect 5643 3464 5685 3473
rect 5643 3424 5644 3464
rect 5684 3424 5685 3464
rect 6403 3464 6461 3465
rect 5643 3415 5685 3424
rect 5763 3461 5821 3462
rect 5763 3421 5772 3461
rect 5812 3421 5821 3461
rect 6403 3424 6412 3464
rect 6452 3424 6461 3464
rect 6403 3423 6461 3424
rect 7651 3464 7709 3465
rect 7651 3424 7660 3464
rect 7700 3424 7709 3464
rect 7651 3423 7709 3424
rect 8043 3464 8085 3473
rect 8043 3424 8044 3464
rect 8084 3424 8085 3464
rect 5763 3420 5821 3421
rect 8043 3415 8085 3424
rect 8139 3464 8181 3473
rect 8139 3424 8140 3464
rect 8180 3424 8181 3464
rect 8139 3415 8181 3424
rect 8611 3464 8669 3465
rect 8611 3424 8620 3464
rect 8660 3424 8669 3464
rect 8611 3423 8669 3424
rect 9859 3464 9917 3465
rect 9859 3424 9868 3464
rect 9908 3424 9917 3464
rect 9859 3423 9917 3424
rect 10251 3464 10293 3473
rect 10251 3424 10252 3464
rect 10292 3424 10293 3464
rect 10251 3415 10293 3424
rect 10539 3464 10581 3473
rect 10539 3424 10540 3464
rect 10580 3424 10581 3464
rect 10539 3415 10581 3424
rect 10723 3464 10781 3465
rect 10723 3424 10732 3464
rect 10772 3424 10781 3464
rect 10723 3423 10781 3424
rect 10923 3464 10965 3473
rect 10923 3424 10924 3464
rect 10964 3424 10965 3464
rect 10923 3415 10965 3424
rect 11107 3464 11165 3465
rect 11107 3424 11116 3464
rect 11156 3424 11165 3464
rect 11107 3423 11165 3424
rect 12355 3464 12413 3465
rect 12355 3424 12364 3464
rect 12404 3424 12413 3464
rect 12355 3423 12413 3424
rect 12843 3464 12885 3473
rect 12843 3424 12844 3464
rect 12884 3424 12885 3464
rect 12843 3415 12885 3424
rect 12939 3464 12981 3473
rect 12939 3424 12940 3464
rect 12980 3424 12981 3464
rect 12939 3415 12981 3424
rect 13323 3464 13365 3473
rect 13323 3424 13324 3464
rect 13364 3424 13365 3464
rect 13323 3415 13365 3424
rect 13419 3464 13461 3473
rect 13419 3424 13420 3464
rect 13460 3424 13461 3464
rect 13419 3415 13461 3424
rect 13891 3464 13949 3465
rect 13891 3424 13900 3464
rect 13940 3424 13949 3464
rect 15427 3464 15485 3465
rect 13891 3423 13949 3424
rect 14379 3450 14421 3459
rect 14379 3410 14380 3450
rect 14420 3410 14421 3450
rect 15427 3424 15436 3464
rect 15476 3424 15485 3464
rect 15427 3423 15485 3424
rect 16675 3464 16733 3465
rect 16675 3424 16684 3464
rect 16724 3424 16733 3464
rect 16675 3423 16733 3424
rect 14379 3401 14421 3410
rect 5259 3392 5301 3401
rect 1699 3380 1757 3381
rect 1699 3340 1708 3380
rect 1748 3340 1757 3380
rect 1699 3339 1757 3340
rect 2083 3380 2141 3381
rect 2083 3340 2092 3380
rect 2132 3340 2141 3380
rect 2083 3339 2141 3340
rect 2467 3380 2525 3381
rect 2467 3340 2476 3380
rect 2516 3340 2525 3380
rect 2467 3339 2525 3340
rect 2851 3380 2909 3381
rect 2851 3340 2860 3380
rect 2900 3340 2909 3380
rect 2851 3339 2909 3340
rect 3235 3380 3293 3381
rect 3235 3340 3244 3380
rect 3284 3340 3293 3380
rect 3235 3339 3293 3340
rect 10539 3296 10581 3305
rect 10539 3256 10540 3296
rect 10580 3256 10581 3296
rect 10539 3247 10581 3256
rect 10827 3296 10869 3305
rect 10827 3256 10828 3296
rect 10868 3256 10869 3296
rect 10827 3247 10869 3256
rect 3051 3212 3093 3221
rect 3051 3172 3052 3212
rect 3092 3172 3093 3212
rect 3051 3163 3093 3172
rect 5067 3212 5109 3221
rect 5067 3172 5068 3212
rect 5108 3172 5109 3212
rect 5067 3163 5109 3172
rect 7851 3212 7893 3221
rect 7851 3172 7852 3212
rect 7892 3172 7893 3212
rect 7851 3163 7893 3172
rect 10059 3212 10101 3221
rect 10059 3172 10060 3212
rect 10100 3172 10101 3212
rect 10059 3163 10101 3172
rect 1152 3044 20352 3068
rect 1152 3004 3688 3044
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 4056 3004 18808 3044
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 19176 3004 20352 3044
rect 1152 2980 20352 3004
rect 1515 2876 1557 2885
rect 1515 2836 1516 2876
rect 1556 2836 1557 2876
rect 1515 2827 1557 2836
rect 1899 2876 1941 2885
rect 1899 2836 1900 2876
rect 1940 2836 1941 2876
rect 1899 2827 1941 2836
rect 4971 2876 5013 2885
rect 4971 2836 4972 2876
rect 5012 2836 5013 2876
rect 4971 2827 5013 2836
rect 5163 2876 5205 2885
rect 5163 2836 5164 2876
rect 5204 2836 5205 2876
rect 5163 2827 5205 2836
rect 7755 2876 7797 2885
rect 7755 2836 7756 2876
rect 7796 2836 7797 2876
rect 7755 2827 7797 2836
rect 14379 2876 14421 2885
rect 14379 2836 14380 2876
rect 14420 2836 14421 2876
rect 14379 2827 14421 2836
rect 16299 2876 16341 2885
rect 16299 2836 16300 2876
rect 16340 2836 16341 2876
rect 16299 2827 16341 2836
rect 9579 2792 9621 2801
rect 9579 2752 9580 2792
rect 9620 2752 9621 2792
rect 9579 2743 9621 2752
rect 10531 2792 10589 2793
rect 10531 2752 10540 2792
rect 10580 2752 10589 2792
rect 10531 2751 10589 2752
rect 1699 2708 1757 2709
rect 1699 2668 1708 2708
rect 1748 2668 1757 2708
rect 1699 2667 1757 2668
rect 2083 2708 2141 2709
rect 2083 2668 2092 2708
rect 2132 2668 2141 2708
rect 2083 2667 2141 2668
rect 2563 2708 2621 2709
rect 2563 2668 2572 2708
rect 2612 2668 2621 2708
rect 2563 2667 2621 2668
rect 10827 2708 10869 2717
rect 10827 2668 10828 2708
rect 10868 2668 10869 2708
rect 10827 2659 10869 2668
rect 11299 2708 11357 2709
rect 11299 2668 11308 2708
rect 11348 2668 11357 2708
rect 11299 2667 11357 2668
rect 5163 2647 5205 2656
rect 3523 2624 3581 2625
rect 3523 2584 3532 2624
rect 3572 2584 3581 2624
rect 3523 2583 3581 2584
rect 4771 2624 4829 2625
rect 4771 2584 4780 2624
rect 4820 2584 4829 2624
rect 5163 2607 5164 2647
rect 5204 2607 5205 2647
rect 5704 2639 5746 2648
rect 5163 2598 5205 2607
rect 5251 2624 5309 2625
rect 4771 2583 4829 2584
rect 5251 2584 5260 2624
rect 5300 2584 5309 2624
rect 5251 2583 5309 2584
rect 5451 2624 5493 2633
rect 5451 2584 5452 2624
rect 5492 2584 5493 2624
rect 5451 2575 5493 2584
rect 5547 2624 5589 2633
rect 5547 2584 5548 2624
rect 5588 2584 5589 2624
rect 5704 2599 5705 2639
rect 5745 2599 5746 2639
rect 10923 2637 10965 2646
rect 5704 2590 5746 2599
rect 6307 2624 6365 2625
rect 5547 2575 5589 2584
rect 6307 2584 6316 2624
rect 6356 2584 6365 2624
rect 6307 2583 6365 2584
rect 7555 2624 7613 2625
rect 7555 2584 7564 2624
rect 7604 2584 7613 2624
rect 7555 2583 7613 2584
rect 8131 2624 8189 2625
rect 8131 2584 8140 2624
rect 8180 2584 8189 2624
rect 8131 2583 8189 2584
rect 9379 2624 9437 2625
rect 9379 2584 9388 2624
rect 9428 2584 9437 2624
rect 9379 2583 9437 2584
rect 9859 2624 9917 2625
rect 9859 2584 9868 2624
rect 9908 2584 9917 2624
rect 9859 2583 9917 2584
rect 10155 2624 10197 2633
rect 10155 2584 10156 2624
rect 10196 2584 10197 2624
rect 10155 2575 10197 2584
rect 10731 2624 10773 2633
rect 10731 2584 10732 2624
rect 10772 2584 10773 2624
rect 10923 2597 10924 2637
rect 10964 2597 10965 2637
rect 10923 2588 10965 2597
rect 12931 2624 12989 2625
rect 10731 2575 10773 2584
rect 12931 2584 12940 2624
rect 12980 2584 12989 2624
rect 12931 2583 12989 2584
rect 14179 2624 14237 2625
rect 14179 2584 14188 2624
rect 14228 2584 14237 2624
rect 14179 2583 14237 2584
rect 14851 2624 14909 2625
rect 14851 2584 14860 2624
rect 14900 2584 14909 2624
rect 14851 2583 14909 2584
rect 16099 2624 16157 2625
rect 16099 2584 16108 2624
rect 16148 2584 16157 2624
rect 16099 2583 16157 2584
rect 10251 2540 10293 2549
rect 10251 2500 10252 2540
rect 10292 2500 10293 2540
rect 10251 2491 10293 2500
rect 2379 2456 2421 2465
rect 2379 2416 2380 2456
rect 2420 2416 2421 2456
rect 2379 2407 2421 2416
rect 11115 2456 11157 2465
rect 11115 2416 11116 2456
rect 11156 2416 11157 2456
rect 11115 2407 11157 2416
rect 1152 2288 20452 2312
rect 1152 2248 4928 2288
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 5296 2248 20048 2288
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20416 2248 20452 2288
rect 1152 2224 20452 2248
rect 1899 2120 1941 2129
rect 1899 2080 1900 2120
rect 1940 2080 1941 2120
rect 1899 2071 1941 2080
rect 5355 2120 5397 2129
rect 5355 2080 5356 2120
rect 5396 2080 5397 2120
rect 5355 2071 5397 2080
rect 5923 2120 5981 2121
rect 5923 2080 5932 2120
rect 5972 2080 5981 2120
rect 5923 2079 5981 2080
rect 6603 2120 6645 2129
rect 6603 2080 6604 2120
rect 6644 2080 6645 2120
rect 6603 2071 6645 2080
rect 6987 2120 7029 2129
rect 6987 2080 6988 2120
rect 7028 2080 7029 2120
rect 6987 2071 7029 2080
rect 7467 2120 7509 2129
rect 7467 2080 7468 2120
rect 7508 2080 7509 2120
rect 7467 2071 7509 2080
rect 9667 2120 9725 2121
rect 9667 2080 9676 2120
rect 9716 2080 9725 2120
rect 9667 2079 9725 2080
rect 10155 2120 10197 2129
rect 10155 2080 10156 2120
rect 10196 2080 10197 2120
rect 10155 2071 10197 2080
rect 3523 1952 3581 1953
rect 3523 1912 3532 1952
rect 3572 1912 3581 1952
rect 3523 1911 3581 1912
rect 4771 1952 4829 1953
rect 4771 1912 4780 1952
rect 4820 1912 4829 1952
rect 4771 1911 4829 1912
rect 5163 1952 5205 1961
rect 5163 1912 5164 1952
rect 5204 1912 5205 1952
rect 5163 1903 5205 1912
rect 5259 1952 5301 1961
rect 5259 1912 5260 1952
rect 5300 1912 5301 1952
rect 5259 1903 5301 1912
rect 5451 1952 5493 1961
rect 5451 1912 5452 1952
rect 5492 1912 5493 1952
rect 5451 1903 5493 1912
rect 5643 1952 5685 1961
rect 5643 1912 5644 1952
rect 5684 1912 5685 1952
rect 5643 1903 5685 1912
rect 5739 1952 5781 1961
rect 5739 1912 5740 1952
rect 5780 1912 5781 1952
rect 5739 1903 5781 1912
rect 7371 1952 7413 1961
rect 7371 1912 7372 1952
rect 7412 1912 7413 1952
rect 7371 1903 7413 1912
rect 7563 1952 7605 1961
rect 7563 1912 7564 1952
rect 7604 1912 7605 1952
rect 7563 1903 7605 1912
rect 7659 1952 7701 1961
rect 7659 1912 7660 1952
rect 7700 1912 7701 1952
rect 7659 1903 7701 1912
rect 9387 1952 9429 1961
rect 9387 1912 9388 1952
rect 9428 1912 9429 1952
rect 9387 1903 9429 1912
rect 9483 1952 9525 1961
rect 9483 1912 9484 1952
rect 9524 1912 9525 1952
rect 9483 1903 9525 1912
rect 9859 1952 9917 1953
rect 9859 1912 9868 1952
rect 9908 1912 9917 1952
rect 9859 1911 9917 1912
rect 9963 1952 10005 1961
rect 9963 1912 9964 1952
rect 10004 1912 10005 1952
rect 9963 1903 10005 1912
rect 10147 1952 10205 1953
rect 10147 1912 10156 1952
rect 10196 1912 10205 1952
rect 10147 1911 10205 1912
rect 1699 1868 1757 1869
rect 1699 1828 1708 1868
rect 1748 1828 1757 1868
rect 1699 1827 1757 1828
rect 2083 1868 2141 1869
rect 2083 1828 2092 1868
rect 2132 1828 2141 1868
rect 2083 1827 2141 1828
rect 2467 1868 2525 1869
rect 2467 1828 2476 1868
rect 2516 1828 2525 1868
rect 2467 1827 2525 1828
rect 2851 1868 2909 1869
rect 2851 1828 2860 1868
rect 2900 1828 2909 1868
rect 2851 1827 2909 1828
rect 3139 1868 3197 1869
rect 3139 1828 3148 1868
rect 3188 1828 3197 1868
rect 3139 1827 3197 1828
rect 6403 1868 6461 1869
rect 6403 1828 6412 1868
rect 6452 1828 6461 1868
rect 7171 1868 7229 1869
rect 6403 1827 6461 1828
rect 6787 1857 6845 1858
rect 6787 1817 6796 1857
rect 6836 1817 6845 1857
rect 7171 1828 7180 1868
rect 7220 1828 7229 1868
rect 7171 1827 7229 1828
rect 7843 1868 7901 1869
rect 7843 1828 7852 1868
rect 7892 1828 7901 1868
rect 7843 1827 7901 1828
rect 8227 1868 8285 1869
rect 8227 1828 8236 1868
rect 8276 1828 8285 1868
rect 8227 1827 8285 1828
rect 8611 1868 8669 1869
rect 8611 1828 8620 1868
rect 8660 1828 8669 1868
rect 8611 1827 8669 1828
rect 8995 1868 9053 1869
rect 8995 1828 9004 1868
rect 9044 1828 9053 1868
rect 8995 1827 9053 1828
rect 10531 1868 10589 1869
rect 10531 1828 10540 1868
rect 10580 1828 10589 1868
rect 10531 1827 10589 1828
rect 10915 1868 10973 1869
rect 10915 1828 10924 1868
rect 10964 1828 10973 1868
rect 10915 1827 10973 1828
rect 11299 1868 11357 1869
rect 11299 1828 11308 1868
rect 11348 1828 11357 1868
rect 11299 1827 11357 1828
rect 11875 1868 11933 1869
rect 11875 1828 11884 1868
rect 11924 1828 11933 1868
rect 11875 1827 11933 1828
rect 12259 1868 12317 1869
rect 12259 1828 12268 1868
rect 12308 1828 12317 1868
rect 12259 1827 12317 1828
rect 12931 1868 12989 1869
rect 12931 1828 12940 1868
rect 12980 1828 12989 1868
rect 12931 1827 12989 1828
rect 13219 1868 13277 1869
rect 13219 1828 13228 1868
rect 13268 1828 13277 1868
rect 13219 1827 13277 1828
rect 13891 1868 13949 1869
rect 13891 1828 13900 1868
rect 13940 1828 13949 1868
rect 13891 1827 13949 1828
rect 14275 1868 14333 1869
rect 14275 1828 14284 1868
rect 14324 1828 14333 1868
rect 14275 1827 14333 1828
rect 14659 1868 14717 1869
rect 14659 1828 14668 1868
rect 14708 1828 14717 1868
rect 14659 1827 14717 1828
rect 15235 1868 15293 1869
rect 15235 1828 15244 1868
rect 15284 1828 15293 1868
rect 15235 1827 15293 1828
rect 15619 1868 15677 1869
rect 15619 1828 15628 1868
rect 15668 1828 15677 1868
rect 15619 1827 15677 1828
rect 16003 1868 16061 1869
rect 16003 1828 16012 1868
rect 16052 1828 16061 1868
rect 16003 1827 16061 1828
rect 16387 1868 16445 1869
rect 16387 1828 16396 1868
rect 16436 1828 16445 1868
rect 16387 1827 16445 1828
rect 6787 1816 6845 1817
rect 1515 1784 1557 1793
rect 1515 1744 1516 1784
rect 1556 1744 1557 1784
rect 1515 1735 1557 1744
rect 4971 1784 5013 1793
rect 4971 1744 4972 1784
rect 5012 1744 5013 1784
rect 4971 1735 5013 1744
rect 2283 1700 2325 1709
rect 2283 1660 2284 1700
rect 2324 1660 2325 1700
rect 2283 1651 2325 1660
rect 2667 1700 2709 1709
rect 2667 1660 2668 1700
rect 2708 1660 2709 1700
rect 2667 1651 2709 1660
rect 3339 1700 3381 1709
rect 3339 1660 3340 1700
rect 3380 1660 3381 1700
rect 3339 1651 3381 1660
rect 6219 1700 6261 1709
rect 6219 1660 6220 1700
rect 6260 1660 6261 1700
rect 6219 1651 6261 1660
rect 8043 1700 8085 1709
rect 8043 1660 8044 1700
rect 8084 1660 8085 1700
rect 8043 1651 8085 1660
rect 8427 1700 8469 1709
rect 8427 1660 8428 1700
rect 8468 1660 8469 1700
rect 8427 1651 8469 1660
rect 8811 1700 8853 1709
rect 8811 1660 8812 1700
rect 8852 1660 8853 1700
rect 8811 1651 8853 1660
rect 9195 1700 9237 1709
rect 9195 1660 9196 1700
rect 9236 1660 9237 1700
rect 9195 1651 9237 1660
rect 10731 1700 10773 1709
rect 10731 1660 10732 1700
rect 10772 1660 10773 1700
rect 10731 1651 10773 1660
rect 11115 1700 11157 1709
rect 11115 1660 11116 1700
rect 11156 1660 11157 1700
rect 11115 1651 11157 1660
rect 11499 1700 11541 1709
rect 11499 1660 11500 1700
rect 11540 1660 11541 1700
rect 11499 1651 11541 1660
rect 11691 1700 11733 1709
rect 11691 1660 11692 1700
rect 11732 1660 11733 1700
rect 11691 1651 11733 1660
rect 12075 1700 12117 1709
rect 12075 1660 12076 1700
rect 12116 1660 12117 1700
rect 12075 1651 12117 1660
rect 12747 1700 12789 1709
rect 12747 1660 12748 1700
rect 12788 1660 12789 1700
rect 12747 1651 12789 1660
rect 13419 1700 13461 1709
rect 13419 1660 13420 1700
rect 13460 1660 13461 1700
rect 13419 1651 13461 1660
rect 14091 1700 14133 1709
rect 14091 1660 14092 1700
rect 14132 1660 14133 1700
rect 14091 1651 14133 1660
rect 14475 1700 14517 1709
rect 14475 1660 14476 1700
rect 14516 1660 14517 1700
rect 14475 1651 14517 1660
rect 14859 1700 14901 1709
rect 14859 1660 14860 1700
rect 14900 1660 14901 1700
rect 14859 1651 14901 1660
rect 15051 1700 15093 1709
rect 15051 1660 15052 1700
rect 15092 1660 15093 1700
rect 15051 1651 15093 1660
rect 15435 1700 15477 1709
rect 15435 1660 15436 1700
rect 15476 1660 15477 1700
rect 15435 1651 15477 1660
rect 15819 1700 15861 1709
rect 15819 1660 15820 1700
rect 15860 1660 15861 1700
rect 15819 1651 15861 1660
rect 16203 1700 16245 1709
rect 16203 1660 16204 1700
rect 16244 1660 16245 1700
rect 16203 1651 16245 1660
rect 1152 1532 20352 1556
rect 1152 1492 3688 1532
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 4056 1492 18808 1532
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 19176 1492 20352 1532
rect 1152 1468 20352 1492
rect 5355 1280 5397 1289
rect 5355 1240 5356 1280
rect 5396 1240 5397 1280
rect 5355 1231 5397 1240
rect 6699 1280 6741 1289
rect 6699 1240 6700 1280
rect 6740 1240 6741 1280
rect 6699 1231 6741 1240
rect 7371 1280 7413 1289
rect 7371 1240 7372 1280
rect 7412 1240 7413 1280
rect 7371 1231 7413 1240
rect 7755 1280 7797 1289
rect 7755 1240 7756 1280
rect 7796 1240 7797 1280
rect 7755 1231 7797 1240
rect 1699 1196 1757 1197
rect 1699 1156 1708 1196
rect 1748 1156 1757 1196
rect 1699 1155 1757 1156
rect 2083 1196 2141 1197
rect 2083 1156 2092 1196
rect 2132 1156 2141 1196
rect 2083 1155 2141 1156
rect 2467 1196 2525 1197
rect 2467 1156 2476 1196
rect 2516 1156 2525 1196
rect 2467 1155 2525 1156
rect 6115 1196 6173 1197
rect 6115 1156 6124 1196
rect 6164 1156 6173 1196
rect 6115 1155 6173 1156
rect 6499 1196 6557 1197
rect 6499 1156 6508 1196
rect 6548 1156 6557 1196
rect 6499 1155 6557 1156
rect 6883 1196 6941 1197
rect 6883 1156 6892 1196
rect 6932 1156 6941 1196
rect 6883 1155 6941 1156
rect 7555 1196 7613 1197
rect 7555 1156 7564 1196
rect 7604 1156 7613 1196
rect 7555 1155 7613 1156
rect 7939 1196 7997 1197
rect 7939 1156 7948 1196
rect 7988 1156 7997 1196
rect 7939 1155 7997 1156
rect 8995 1196 9053 1197
rect 8995 1156 9004 1196
rect 9044 1156 9053 1196
rect 8995 1155 9053 1156
rect 9379 1196 9437 1197
rect 9379 1156 9388 1196
rect 9428 1156 9437 1196
rect 9379 1155 9437 1156
rect 9763 1196 9821 1197
rect 9763 1156 9772 1196
rect 9812 1156 9821 1196
rect 9763 1155 9821 1156
rect 10147 1196 10205 1197
rect 10147 1156 10156 1196
rect 10196 1156 10205 1196
rect 10147 1155 10205 1156
rect 10531 1196 10589 1197
rect 10531 1156 10540 1196
rect 10580 1156 10589 1196
rect 10531 1155 10589 1156
rect 10915 1196 10973 1197
rect 10915 1156 10924 1196
rect 10964 1156 10973 1196
rect 10915 1155 10973 1156
rect 15139 1196 15197 1197
rect 15139 1156 15148 1196
rect 15188 1156 15197 1196
rect 15139 1155 15197 1156
rect 16003 1196 16061 1197
rect 16003 1156 16012 1196
rect 16052 1156 16061 1196
rect 16003 1155 16061 1156
rect 5163 1112 5205 1121
rect 5163 1072 5164 1112
rect 5204 1072 5205 1112
rect 5163 1063 5205 1072
rect 5259 1112 5301 1121
rect 5259 1072 5260 1112
rect 5300 1072 5301 1112
rect 5259 1063 5301 1072
rect 5451 1112 5493 1121
rect 5451 1072 5452 1112
rect 5492 1072 5493 1112
rect 5451 1063 5493 1072
rect 1515 944 1557 953
rect 1515 904 1516 944
rect 1556 904 1557 944
rect 1515 895 1557 904
rect 1899 944 1941 953
rect 1899 904 1900 944
rect 1940 904 1941 944
rect 1899 895 1941 904
rect 2283 944 2325 953
rect 2283 904 2284 944
rect 2324 904 2325 944
rect 2283 895 2325 904
rect 5931 944 5973 953
rect 5931 904 5932 944
rect 5972 904 5973 944
rect 5931 895 5973 904
rect 6315 944 6357 953
rect 6315 904 6316 944
rect 6356 904 6357 944
rect 6315 895 6357 904
rect 9195 944 9237 953
rect 9195 904 9196 944
rect 9236 904 9237 944
rect 9195 895 9237 904
rect 9579 944 9621 953
rect 9579 904 9580 944
rect 9620 904 9621 944
rect 9579 895 9621 904
rect 9963 944 10005 953
rect 9963 904 9964 944
rect 10004 904 10005 944
rect 9963 895 10005 904
rect 10347 944 10389 953
rect 10347 904 10348 944
rect 10388 904 10389 944
rect 10347 895 10389 904
rect 10731 944 10773 953
rect 10731 904 10732 944
rect 10772 904 10773 944
rect 10731 895 10773 904
rect 11115 944 11157 953
rect 11115 904 11116 944
rect 11156 904 11157 944
rect 11115 895 11157 904
rect 14955 944 14997 953
rect 14955 904 14956 944
rect 14996 904 14997 944
rect 14955 895 14997 904
rect 15819 944 15861 953
rect 15819 904 15820 944
rect 15860 904 15861 944
rect 15819 895 15861 904
rect 1152 776 20452 800
rect 1152 736 4928 776
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 5296 736 20048 776
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20416 736 20452 776
rect 1152 712 20452 736
<< via1 >>
rect 3688 84652 3728 84692
rect 3770 84652 3810 84692
rect 3852 84652 3892 84692
rect 3934 84652 3974 84692
rect 4016 84652 4056 84692
rect 18808 84652 18848 84692
rect 18890 84652 18930 84692
rect 18972 84652 19012 84692
rect 19054 84652 19094 84692
rect 19136 84652 19176 84692
rect 3052 84400 3092 84440
rect 3436 84400 3476 84440
rect 3244 84316 3284 84356
rect 3628 84316 3668 84356
rect 18124 84064 18164 84104
rect 18508 84064 18548 84104
rect 18988 84064 19028 84104
rect 19276 84064 19316 84104
rect 4928 83896 4968 83936
rect 5010 83896 5050 83936
rect 5092 83896 5132 83936
rect 5174 83896 5214 83936
rect 5256 83896 5296 83936
rect 20048 83896 20088 83936
rect 20130 83896 20170 83936
rect 20212 83896 20252 83936
rect 20294 83896 20334 83936
rect 20376 83896 20416 83936
rect 1900 83728 1940 83768
rect 2284 83728 2324 83768
rect 2668 83728 2708 83768
rect 3052 83728 3092 83768
rect 3436 83728 3476 83768
rect 3820 83728 3860 83768
rect 4204 83728 4244 83768
rect 5356 83728 5396 83768
rect 5548 83728 5588 83768
rect 6220 83728 6260 83768
rect 6412 83728 6452 83768
rect 6988 83728 7028 83768
rect 7564 83728 7604 83768
rect 8428 83728 8468 83768
rect 8812 83728 8852 83768
rect 9580 83728 9620 83768
rect 10060 83728 10100 83768
rect 10444 83728 10484 83768
rect 11308 83728 11348 83768
rect 15724 83728 15764 83768
rect 16780 83728 16820 83768
rect 17356 83728 17396 83768
rect 17740 83728 17780 83768
rect 18892 83728 18932 83768
rect 19660 83728 19700 83768
rect 20044 83728 20084 83768
rect 1708 83476 1748 83516
rect 2092 83476 2132 83516
rect 2476 83476 2516 83516
rect 2860 83476 2900 83516
rect 3244 83476 3284 83516
rect 3628 83476 3668 83516
rect 4012 83476 4052 83516
rect 4396 83476 4436 83516
rect 4972 83476 5012 83516
rect 5164 83476 5204 83516
rect 5740 83476 5780 83516
rect 6028 83476 6068 83516
rect 6604 83476 6644 83516
rect 6796 83476 6836 83516
rect 7180 83476 7220 83516
rect 7756 83476 7796 83516
rect 8140 83476 8180 83516
rect 8620 83476 8660 83516
rect 9004 83476 9044 83516
rect 9772 83476 9812 83516
rect 10252 83476 10292 83516
rect 10636 83476 10676 83516
rect 11500 83476 11540 83516
rect 13324 83476 13364 83516
rect 13708 83476 13748 83516
rect 14092 83476 14132 83516
rect 14476 83476 14516 83516
rect 14860 83476 14900 83516
rect 15244 83476 15284 83516
rect 15916 83476 15956 83516
rect 16588 83476 16628 83516
rect 17164 83476 17204 83516
rect 17548 83476 17588 83516
rect 17932 83476 17972 83516
rect 18316 83476 18356 83516
rect 18700 83476 18740 83516
rect 19084 83476 19124 83516
rect 19468 83476 19508 83516
rect 19852 83476 19892 83516
rect 20236 83476 20276 83516
rect 4588 83392 4628 83432
rect 7372 83392 7412 83432
rect 4780 83308 4820 83348
rect 7948 83308 7988 83348
rect 13132 83308 13172 83348
rect 13516 83308 13556 83348
rect 13900 83308 13940 83348
rect 14284 83308 14324 83348
rect 14668 83308 14708 83348
rect 15052 83308 15092 83348
rect 16972 83308 17012 83348
rect 18124 83308 18164 83348
rect 18508 83308 18548 83348
rect 19276 83308 19316 83348
rect 3688 83140 3728 83180
rect 3770 83140 3810 83180
rect 3852 83140 3892 83180
rect 3934 83140 3974 83180
rect 4016 83140 4056 83180
rect 18808 83140 18848 83180
rect 18890 83140 18930 83180
rect 18972 83140 19012 83180
rect 19054 83140 19094 83180
rect 19136 83140 19176 83180
rect 3628 82972 3668 83012
rect 7468 82972 7508 83012
rect 18220 82972 18260 83012
rect 18604 82972 18644 83012
rect 18988 82972 19028 83012
rect 17452 82888 17492 82928
rect 17836 82888 17876 82928
rect 19372 82888 19412 82928
rect 19756 82888 19796 82928
rect 20140 82888 20180 82928
rect 3820 82804 3860 82844
rect 7276 82804 7316 82844
rect 14380 82804 14420 82844
rect 14764 82804 14804 82844
rect 18028 82804 18068 82844
rect 18412 82804 18452 82844
rect 18796 82804 18836 82844
rect 19180 82804 19220 82844
rect 1900 82720 1940 82760
rect 3148 82720 3188 82760
rect 4108 82720 4148 82760
rect 5356 82720 5396 82760
rect 3340 82552 3380 82592
rect 5548 82552 5588 82592
rect 14188 82552 14228 82592
rect 14572 82552 14612 82592
rect 17356 82552 17396 82592
rect 17740 82552 17780 82592
rect 19660 82552 19700 82592
rect 20044 82552 20084 82592
rect 4928 82384 4968 82424
rect 5010 82384 5050 82424
rect 5092 82384 5132 82424
rect 5174 82384 5214 82424
rect 5256 82384 5296 82424
rect 20048 82384 20088 82424
rect 20130 82384 20170 82424
rect 20212 82384 20252 82424
rect 20294 82384 20334 82424
rect 20376 82384 20416 82424
rect 18028 82216 18068 82256
rect 18412 82216 18452 82256
rect 19180 82216 19220 82256
rect 1228 82048 1268 82088
rect 2476 82048 2516 82088
rect 3724 82048 3764 82088
rect 4972 82048 5012 82088
rect 18796 81964 18836 82004
rect 18124 81880 18164 81920
rect 18508 81880 18548 81920
rect 19276 81880 19316 81920
rect 2668 81796 2708 81836
rect 5164 81796 5204 81836
rect 3688 81628 3728 81668
rect 3770 81628 3810 81668
rect 3852 81628 3892 81668
rect 3934 81628 3974 81668
rect 4016 81628 4056 81668
rect 18808 81628 18848 81668
rect 18890 81628 18930 81668
rect 18972 81628 19012 81668
rect 19054 81628 19094 81668
rect 19136 81628 19176 81668
rect 15820 81460 15860 81500
rect 15628 81292 15668 81332
rect 1420 81208 1460 81248
rect 2668 81208 2708 81248
rect 2860 81208 2900 81248
rect 4108 81208 4148 81248
rect 4492 81208 4532 81248
rect 5740 81208 5780 81248
rect 6124 81208 6164 81248
rect 7372 81208 7412 81248
rect 1228 81124 1268 81164
rect 4300 81040 4340 81080
rect 5932 81040 5972 81080
rect 7564 81040 7604 81080
rect 4928 80872 4968 80912
rect 5010 80872 5050 80912
rect 5092 80872 5132 80912
rect 5174 80872 5214 80912
rect 5256 80872 5296 80912
rect 20048 80872 20088 80912
rect 20130 80872 20170 80912
rect 20212 80872 20252 80912
rect 20294 80872 20334 80912
rect 20376 80872 20416 80912
rect 7180 80620 7220 80660
rect 1612 80536 1652 80576
rect 2860 80536 2900 80576
rect 3724 80536 3764 80576
rect 4972 80536 5012 80576
rect 5452 80536 5492 80576
rect 5548 80536 5588 80576
rect 6508 80536 6548 80576
rect 6988 80531 7028 80571
rect 5932 80452 5972 80492
rect 6028 80452 6068 80492
rect 3052 80284 3092 80324
rect 5164 80284 5204 80324
rect 3688 80116 3728 80156
rect 3770 80116 3810 80156
rect 3852 80116 3892 80156
rect 3934 80116 3974 80156
rect 4016 80116 4056 80156
rect 18808 80116 18848 80156
rect 18890 80116 18930 80156
rect 18972 80116 19012 80156
rect 19054 80116 19094 80156
rect 19136 80116 19176 80156
rect 16012 79948 16052 79988
rect 4108 79780 4148 79820
rect 7276 79780 7316 79820
rect 15820 79780 15860 79820
rect 1420 79696 1460 79736
rect 2668 79696 2708 79736
rect 3628 79696 3668 79736
rect 3724 79696 3764 79736
rect 4204 79696 4244 79736
rect 4684 79696 4724 79736
rect 5212 79705 5252 79745
rect 5548 79696 5588 79736
rect 6796 79696 6836 79736
rect 7180 79696 7220 79736
rect 7372 79696 7412 79736
rect 7948 79696 7988 79736
rect 9196 79696 9236 79736
rect 1228 79528 1268 79568
rect 5356 79528 5396 79568
rect 6988 79528 7028 79568
rect 9388 79528 9428 79568
rect 4928 79360 4968 79400
rect 5010 79360 5050 79400
rect 5092 79360 5132 79400
rect 5174 79360 5214 79400
rect 5256 79360 5296 79400
rect 20048 79360 20088 79400
rect 20130 79360 20170 79400
rect 20212 79360 20252 79400
rect 20294 79360 20334 79400
rect 20376 79360 20416 79400
rect 5932 79192 5972 79232
rect 7948 79192 7988 79232
rect 16972 79192 17012 79232
rect 1900 79024 1940 79064
rect 3148 79024 3188 79064
rect 4204 79024 4244 79064
rect 5452 79024 5492 79064
rect 5836 79024 5876 79064
rect 6028 79024 6068 79064
rect 6220 79024 6260 79064
rect 7468 79024 7508 79064
rect 7852 79024 7892 79064
rect 8044 79024 8084 79064
rect 8140 79024 8180 79064
rect 8908 79024 8948 79064
rect 10156 79024 10196 79064
rect 16780 78940 16820 78980
rect 3340 78772 3380 78812
rect 5644 78772 5684 78812
rect 7660 78772 7700 78812
rect 10348 78772 10388 78812
rect 3688 78604 3728 78644
rect 3770 78604 3810 78644
rect 3852 78604 3892 78644
rect 3934 78604 3974 78644
rect 4016 78604 4056 78644
rect 18808 78604 18848 78644
rect 18890 78604 18930 78644
rect 18972 78604 19012 78644
rect 19054 78604 19094 78644
rect 19136 78604 19176 78644
rect 9004 78268 9044 78308
rect 1228 78184 1268 78224
rect 2476 78184 2516 78224
rect 3340 78184 3380 78224
rect 4588 78184 4628 78224
rect 5164 78184 5204 78224
rect 6412 78184 6452 78224
rect 6700 78184 6740 78224
rect 7948 78184 7988 78224
rect 8428 78184 8468 78224
rect 8524 78184 8564 78224
rect 8908 78184 8948 78224
rect 9484 78184 9524 78224
rect 9964 78198 10004 78238
rect 2668 78100 2708 78140
rect 8140 78100 8180 78140
rect 10156 78100 10196 78140
rect 4780 78016 4820 78056
rect 4972 78016 5012 78056
rect 4928 77848 4968 77888
rect 5010 77848 5050 77888
rect 5092 77848 5132 77888
rect 5174 77848 5214 77888
rect 5256 77848 5296 77888
rect 20048 77848 20088 77888
rect 20130 77848 20170 77888
rect 20212 77848 20252 77888
rect 20294 77848 20334 77888
rect 20376 77848 20416 77888
rect 4588 77596 4628 77636
rect 9484 77596 9524 77636
rect 2860 77512 2900 77552
rect 2956 77512 2996 77552
rect 3340 77512 3380 77552
rect 3916 77512 3956 77552
rect 4396 77507 4436 77547
rect 5164 77512 5204 77552
rect 5452 77512 5492 77552
rect 5548 77512 5588 77552
rect 6028 77512 6068 77552
rect 7276 77512 7316 77552
rect 7756 77512 7796 77552
rect 7852 77512 7892 77552
rect 8812 77512 8852 77552
rect 9340 77502 9380 77542
rect 3436 77428 3476 77468
rect 8236 77428 8276 77468
rect 8332 77428 8372 77468
rect 5836 77344 5876 77384
rect 7468 77260 7508 77300
rect 3688 77092 3728 77132
rect 3770 77092 3810 77132
rect 3852 77092 3892 77132
rect 3934 77092 3974 77132
rect 4016 77092 4056 77132
rect 18808 77092 18848 77132
rect 18890 77092 18930 77132
rect 18972 77092 19012 77132
rect 19054 77092 19094 77132
rect 19136 77092 19176 77132
rect 17164 76840 17204 76880
rect 9004 76756 9044 76796
rect 16972 76756 17012 76796
rect 2092 76672 2132 76712
rect 3340 76672 3380 76712
rect 4396 76672 4436 76712
rect 5644 76672 5684 76712
rect 6028 76672 6068 76712
rect 6124 76672 6164 76712
rect 6700 76672 6740 76712
rect 7948 76672 7988 76712
rect 8428 76672 8468 76712
rect 8524 76672 8564 76712
rect 8908 76672 8948 76712
rect 9484 76672 9524 76712
rect 10012 76681 10052 76721
rect 10540 76672 10580 76712
rect 11788 76672 11828 76712
rect 10348 76588 10388 76628
rect 3532 76504 3572 76544
rect 5836 76504 5876 76544
rect 6316 76504 6356 76544
rect 8140 76504 8180 76544
rect 10156 76504 10196 76544
rect 4928 76336 4968 76376
rect 5010 76336 5050 76376
rect 5092 76336 5132 76376
rect 5174 76336 5214 76376
rect 5256 76336 5296 76376
rect 20048 76336 20088 76376
rect 20130 76336 20170 76376
rect 20212 76336 20252 76376
rect 20294 76336 20334 76376
rect 20376 76336 20416 76376
rect 3244 76168 3284 76208
rect 6700 76168 6740 76208
rect 7660 76168 7700 76208
rect 9868 76168 9908 76208
rect 10444 76168 10484 76208
rect 11020 76084 11060 76124
rect 1516 76000 1556 76040
rect 1612 76000 1652 76040
rect 2572 76000 2612 76040
rect 3052 75995 3092 76035
rect 4972 76000 5012 76040
rect 5068 76000 5108 76040
rect 6028 76000 6068 76040
rect 6508 75995 6548 76035
rect 6892 76000 6932 76040
rect 6988 76000 7028 76040
rect 7084 76000 7124 76040
rect 7180 76000 7220 76040
rect 7372 76000 7412 76040
rect 7468 76000 7508 76040
rect 7564 76000 7604 76040
rect 8140 76000 8180 76040
rect 8236 76000 8276 76040
rect 8716 76000 8756 76040
rect 9196 76000 9236 76040
rect 9676 75995 9716 76035
rect 10348 76000 10388 76040
rect 10540 76000 10580 76040
rect 11212 76000 11252 76040
rect 12460 76000 12500 76040
rect 1996 75916 2036 75956
rect 2092 75916 2132 75956
rect 5452 75916 5492 75956
rect 5548 75916 5588 75956
rect 8620 75916 8660 75956
rect 10828 75832 10868 75872
rect 3688 75580 3728 75620
rect 3770 75580 3810 75620
rect 3852 75580 3892 75620
rect 3934 75580 3974 75620
rect 4016 75580 4056 75620
rect 18808 75580 18848 75620
rect 18890 75580 18930 75620
rect 18972 75580 19012 75620
rect 19054 75580 19094 75620
rect 19136 75580 19176 75620
rect 4780 75244 4820 75284
rect 11308 75244 11348 75284
rect 11404 75244 11444 75284
rect 1228 75160 1268 75200
rect 2476 75160 2516 75200
rect 4300 75160 4340 75200
rect 4396 75160 4436 75200
rect 4876 75160 4916 75200
rect 5356 75160 5396 75200
rect 5836 75174 5876 75214
rect 6220 75160 6260 75200
rect 7468 75160 7508 75200
rect 9100 75160 9140 75200
rect 10348 75160 10388 75200
rect 10828 75160 10868 75200
rect 10924 75160 10964 75200
rect 11884 75160 11924 75200
rect 12412 75169 12452 75209
rect 6028 75076 6068 75116
rect 10540 75076 10580 75116
rect 2668 74992 2708 75032
rect 7660 74992 7700 75032
rect 12556 74992 12596 75032
rect 4928 74824 4968 74864
rect 5010 74824 5050 74864
rect 5092 74824 5132 74864
rect 5174 74824 5214 74864
rect 5256 74824 5296 74864
rect 20048 74824 20088 74864
rect 20130 74824 20170 74864
rect 20212 74824 20252 74864
rect 20294 74824 20334 74864
rect 20376 74824 20416 74864
rect 8908 74698 8948 74738
rect 7372 74656 7412 74696
rect 9580 74656 9620 74696
rect 12748 74656 12788 74696
rect 9868 74572 9908 74612
rect 1420 74488 1460 74528
rect 2668 74488 2708 74528
rect 2860 74488 2900 74528
rect 4108 74488 4148 74528
rect 5452 74488 5492 74528
rect 5740 74488 5780 74528
rect 6988 74488 7028 74528
rect 7564 74488 7604 74528
rect 7660 74488 7700 74528
rect 8620 74488 8660 74528
rect 8716 74488 8756 74528
rect 9100 74488 9140 74528
rect 9196 74488 9236 74528
rect 9292 74488 9332 74528
rect 9388 74488 9428 74528
rect 9676 74488 9716 74528
rect 10060 74488 10100 74528
rect 10156 74488 10196 74528
rect 10252 74488 10292 74528
rect 10348 74488 10388 74528
rect 11308 74488 11348 74528
rect 12556 74488 12596 74528
rect 5548 74320 5588 74360
rect 10732 74320 10772 74360
rect 1228 74236 1268 74276
rect 4300 74236 4340 74276
rect 7180 74236 7220 74276
rect 3688 74068 3728 74108
rect 3770 74068 3810 74108
rect 3852 74068 3892 74108
rect 3934 74068 3974 74108
rect 4016 74068 4056 74108
rect 18808 74068 18848 74108
rect 18890 74068 18930 74108
rect 18972 74068 19012 74108
rect 19054 74068 19094 74108
rect 19136 74068 19176 74108
rect 6796 73900 6836 73940
rect 10828 73900 10868 73940
rect 5260 73732 5300 73772
rect 5356 73732 5396 73772
rect 1804 73648 1844 73688
rect 1900 73648 1940 73688
rect 2284 73648 2324 73688
rect 2380 73648 2420 73688
rect 2860 73648 2900 73688
rect 3340 73662 3380 73702
rect 4780 73648 4820 73688
rect 4876 73648 4916 73688
rect 5836 73648 5876 73688
rect 6316 73662 6356 73702
rect 6796 73648 6836 73688
rect 6892 73648 6932 73688
rect 7084 73648 7124 73688
rect 7180 73648 7220 73688
rect 7281 73648 7321 73688
rect 7756 73648 7796 73688
rect 7852 73648 7892 73688
rect 8236 73648 8276 73688
rect 9484 73648 9524 73688
rect 10060 73648 10100 73688
rect 10156 73648 10196 73688
rect 10252 73648 10292 73688
rect 10348 73648 10388 73688
rect 10540 73648 10580 73688
rect 11020 73648 11060 73688
rect 12268 73648 12308 73688
rect 3532 73564 3572 73604
rect 6508 73480 6548 73520
rect 8044 73480 8084 73520
rect 9676 73480 9716 73520
rect 10636 73480 10676 73520
rect 4928 73312 4968 73352
rect 5010 73312 5050 73352
rect 5092 73312 5132 73352
rect 5174 73312 5214 73352
rect 5256 73312 5296 73352
rect 20048 73312 20088 73352
rect 20130 73312 20170 73352
rect 20212 73312 20252 73352
rect 20294 73312 20334 73352
rect 20376 73312 20416 73352
rect 8236 73060 8276 73100
rect 10252 73060 10292 73100
rect 1228 72976 1268 73016
rect 2476 72976 2516 73016
rect 3052 72976 3092 73016
rect 4300 72976 4340 73016
rect 4492 72976 4532 73016
rect 5740 72976 5780 73016
rect 6316 72976 6356 73016
rect 6508 72976 6548 73016
rect 6604 72980 6644 73020
rect 6796 72976 6836 73016
rect 8044 72976 8084 73016
rect 8524 72976 8564 73016
rect 8620 72976 8660 73016
rect 9580 72976 9620 73016
rect 10060 72971 10100 73011
rect 10444 72976 10484 73016
rect 10540 72976 10580 73016
rect 10924 73018 10964 73058
rect 10732 72976 10772 73016
rect 12172 72976 12212 73016
rect 9004 72892 9044 72932
rect 9100 72892 9140 72932
rect 16012 72892 16052 72932
rect 6508 72808 6548 72848
rect 16204 72808 16244 72848
rect 2668 72724 2708 72764
rect 2860 72724 2900 72764
rect 5932 72724 5972 72764
rect 10732 72724 10772 72764
rect 12364 72724 12404 72764
rect 3688 72556 3728 72596
rect 3770 72556 3810 72596
rect 3852 72556 3892 72596
rect 3934 72556 3974 72596
rect 4016 72556 4056 72596
rect 18808 72556 18848 72596
rect 18890 72556 18930 72596
rect 18972 72556 19012 72596
rect 19054 72556 19094 72596
rect 19136 72556 19176 72596
rect 2572 72220 2612 72260
rect 1996 72136 2036 72176
rect 2092 72136 2132 72176
rect 2476 72136 2516 72176
rect 3052 72136 3092 72176
rect 3532 72150 3572 72190
rect 4588 72136 4628 72176
rect 5836 72136 5876 72176
rect 6220 72136 6260 72176
rect 6316 72136 6356 72176
rect 6412 72136 6452 72176
rect 6796 72136 6836 72176
rect 6988 72136 7028 72176
rect 8236 72136 8276 72176
rect 8620 72136 8660 72176
rect 8812 72136 8852 72176
rect 8908 72136 8948 72176
rect 9100 72136 9140 72176
rect 9196 72136 9236 72176
rect 9292 72136 9332 72176
rect 9388 72136 9428 72176
rect 9580 72136 9620 72176
rect 9772 72136 9812 72176
rect 9868 72136 9908 72176
rect 10060 72136 10100 72176
rect 10348 72136 10388 72176
rect 11884 72136 11924 72176
rect 11980 72136 12020 72176
rect 12364 72136 12404 72176
rect 12460 72136 12500 72176
rect 12940 72136 12980 72176
rect 13468 72145 13508 72185
rect 13996 72136 14036 72176
rect 15244 72136 15284 72176
rect 15724 72136 15764 72176
rect 15820 72136 15860 72176
rect 16204 72136 16244 72176
rect 16300 72136 16340 72176
rect 16780 72136 16820 72176
rect 17308 72145 17348 72185
rect 15436 72052 15476 72092
rect 17452 72052 17492 72092
rect 3724 71968 3764 72008
rect 6028 71968 6068 72008
rect 6508 71968 6548 72008
rect 6700 71968 6740 72008
rect 8428 71968 8468 72008
rect 9676 71968 9716 72008
rect 10252 71968 10292 72008
rect 13612 71968 13652 72008
rect 4928 71800 4968 71840
rect 5010 71800 5050 71840
rect 5092 71800 5132 71840
rect 5174 71800 5214 71840
rect 5256 71800 5296 71840
rect 20048 71800 20088 71840
rect 20130 71800 20170 71840
rect 20212 71800 20252 71840
rect 20294 71800 20334 71840
rect 20376 71800 20416 71840
rect 5644 71632 5684 71672
rect 9196 71632 9236 71672
rect 13612 71632 13652 71672
rect 17356 71632 17396 71672
rect 15244 71548 15284 71588
rect 1228 71464 1268 71504
rect 2476 71464 2516 71504
rect 2860 71464 2900 71504
rect 4108 71464 4148 71504
rect 5452 71464 5492 71504
rect 5548 71464 5588 71504
rect 5740 71464 5780 71504
rect 5932 71464 5972 71504
rect 7180 71464 7220 71504
rect 7756 71464 7796 71504
rect 9004 71464 9044 71504
rect 9580 71464 9620 71504
rect 10828 71464 10868 71504
rect 12172 71464 12212 71504
rect 13420 71464 13460 71504
rect 13804 71464 13844 71504
rect 15052 71464 15092 71504
rect 15532 71464 15572 71504
rect 15724 71464 15764 71504
rect 15916 71464 15956 71504
rect 17164 71464 17204 71504
rect 17548 71464 17588 71504
rect 18796 71464 18836 71504
rect 19372 71464 19412 71504
rect 7372 71296 7412 71336
rect 9388 71296 9428 71336
rect 2668 71212 2708 71252
rect 4300 71212 4340 71252
rect 15724 71212 15764 71252
rect 18988 71212 19028 71252
rect 19468 71212 19508 71252
rect 3688 71044 3728 71084
rect 3770 71044 3810 71084
rect 3852 71044 3892 71084
rect 3934 71044 3974 71084
rect 4016 71044 4056 71084
rect 18808 71044 18848 71084
rect 18890 71044 18930 71084
rect 18972 71044 19012 71084
rect 19054 71044 19094 71084
rect 19136 71044 19176 71084
rect 16396 70876 16436 70916
rect 7468 70792 7508 70832
rect 10348 70792 10388 70832
rect 10540 70792 10580 70832
rect 15052 70792 15092 70832
rect 2956 70708 2996 70748
rect 3052 70708 3092 70748
rect 5644 70708 5684 70748
rect 2476 70624 2516 70664
rect 2572 70624 2612 70664
rect 3532 70624 3572 70664
rect 4012 70638 4052 70678
rect 5068 70624 5108 70664
rect 5164 70624 5204 70664
rect 5548 70624 5588 70664
rect 6124 70615 6164 70655
rect 6604 70638 6644 70678
rect 6988 70624 7028 70664
rect 7084 70624 7124 70664
rect 7276 70624 7316 70664
rect 7468 70624 7508 70664
rect 7660 70624 7700 70664
rect 8044 70624 8084 70664
rect 8140 70624 8180 70664
rect 8524 70624 8564 70664
rect 8620 70624 8660 70664
rect 9087 70637 9127 70677
rect 9628 70666 9668 70706
rect 10348 70624 10388 70664
rect 10732 70624 10772 70664
rect 11980 70624 12020 70664
rect 13036 70624 13076 70664
rect 14284 70624 14324 70664
rect 14764 70624 14804 70664
rect 14860 70624 14900 70664
rect 15052 70624 15092 70664
rect 15244 70624 15284 70664
rect 15340 70624 15380 70664
rect 15436 70624 15476 70664
rect 15532 70624 15572 70664
rect 15724 70624 15764 70664
rect 15916 70624 15956 70664
rect 16972 70624 17012 70664
rect 17644 70624 17684 70664
rect 18892 70624 18932 70664
rect 19276 70624 19316 70664
rect 19372 70624 19412 70664
rect 19468 70624 19508 70664
rect 19852 70624 19892 70664
rect 4204 70540 4244 70580
rect 6796 70540 6836 70580
rect 7180 70540 7220 70580
rect 9772 70540 9812 70580
rect 15820 70540 15860 70580
rect 20044 70540 20084 70580
rect 12172 70456 12212 70496
rect 14476 70456 14516 70496
rect 19084 70456 19124 70496
rect 19564 70456 19604 70496
rect 19756 70456 19796 70496
rect 4928 70288 4968 70328
rect 5010 70288 5050 70328
rect 5092 70288 5132 70328
rect 5174 70288 5214 70328
rect 5256 70288 5296 70328
rect 20048 70288 20088 70328
rect 20130 70288 20170 70328
rect 20212 70288 20252 70328
rect 20294 70288 20334 70328
rect 20376 70288 20416 70328
rect 16204 70120 16244 70160
rect 16396 70120 16436 70160
rect 16876 70120 16916 70160
rect 13324 70036 13364 70076
rect 19372 70036 19412 70076
rect 1228 69952 1268 69992
rect 2476 69952 2516 69992
rect 3052 69952 3092 69992
rect 4300 69952 4340 69992
rect 4684 69952 4724 69992
rect 5932 69952 5972 69992
rect 6124 69952 6164 69992
rect 6220 69952 6260 69992
rect 6316 69952 6356 69992
rect 6412 69952 6452 69992
rect 6796 69952 6836 69992
rect 6988 69952 7028 69992
rect 8236 69952 8276 69992
rect 9484 69952 9524 69992
rect 9868 69952 9908 69992
rect 11116 69952 11156 69992
rect 11596 69952 11636 69992
rect 11692 69952 11732 69992
rect 12652 69952 12692 69992
rect 13180 69942 13220 69982
rect 14476 69952 14516 69992
rect 14572 69952 14612 69992
rect 15532 69952 15572 69992
rect 16012 69938 16052 69978
rect 16492 69952 16532 69992
rect 16588 69952 16628 69992
rect 16684 69952 16724 69992
rect 17068 69952 17108 69992
rect 17164 69952 17204 69992
rect 17644 69952 17684 69992
rect 17740 69952 17780 69992
rect 18124 69952 18164 69992
rect 18700 69952 18740 69992
rect 19180 69947 19220 69987
rect 19564 69952 19604 69992
rect 19660 69952 19700 69992
rect 19852 69952 19892 69992
rect 20044 69952 20084 69992
rect 20236 69952 20276 69992
rect 6892 69868 6932 69908
rect 12076 69868 12116 69908
rect 12172 69868 12212 69908
rect 14956 69868 14996 69908
rect 15052 69868 15092 69908
rect 18220 69868 18260 69908
rect 20044 69784 20084 69824
rect 2668 69700 2708 69740
rect 2860 69700 2900 69740
rect 4492 69700 4532 69740
rect 9676 69700 9716 69740
rect 11308 69700 11348 69740
rect 19852 69700 19892 69740
rect 3688 69532 3728 69572
rect 3770 69532 3810 69572
rect 3852 69532 3892 69572
rect 3934 69532 3974 69572
rect 4016 69532 4056 69572
rect 18808 69532 18848 69572
rect 18890 69532 18930 69572
rect 18972 69532 19012 69572
rect 19054 69532 19094 69572
rect 19136 69532 19176 69572
rect 13420 69364 13460 69404
rect 15148 69364 15188 69404
rect 17836 69364 17876 69404
rect 5452 69280 5492 69320
rect 15340 69280 15380 69320
rect 2476 69196 2516 69236
rect 10444 69196 10484 69236
rect 1900 69112 1940 69152
rect 1996 69112 2036 69152
rect 2380 69112 2420 69152
rect 2956 69112 2996 69152
rect 3436 69126 3476 69166
rect 4012 69112 4052 69152
rect 5260 69112 5300 69152
rect 5644 69112 5684 69152
rect 6892 69112 6932 69152
rect 7084 69112 7124 69152
rect 7180 69112 7220 69152
rect 7372 69112 7412 69152
rect 8236 69112 8276 69152
rect 9484 69112 9524 69152
rect 9964 69112 10004 69152
rect 10060 69112 10100 69152
rect 10540 69112 10580 69152
rect 11020 69112 11060 69152
rect 11500 69117 11540 69157
rect 11980 69112 12020 69152
rect 13228 69112 13268 69152
rect 13708 69112 13748 69152
rect 14956 69112 14996 69152
rect 15724 69112 15764 69152
rect 16012 69112 16052 69152
rect 16396 69112 16436 69152
rect 17644 69112 17684 69152
rect 18220 69112 18260 69152
rect 18316 69091 18356 69131
rect 18412 69112 18452 69152
rect 18700 69112 18740 69152
rect 18796 69112 18836 69152
rect 18892 69112 18932 69152
rect 18988 69112 19028 69152
rect 19180 69112 19220 69152
rect 19276 69112 19316 69152
rect 19660 69112 19700 69152
rect 19756 69112 19796 69152
rect 3628 69028 3668 69068
rect 15628 69028 15668 69068
rect 3820 68944 3860 68984
rect 7276 68944 7316 68984
rect 9676 68944 9716 68984
rect 11692 68944 11732 68984
rect 18508 68944 18548 68984
rect 19468 68944 19508 68984
rect 19948 68944 19988 68984
rect 4928 68776 4968 68816
rect 5010 68776 5050 68816
rect 5092 68776 5132 68816
rect 5174 68776 5214 68816
rect 5256 68776 5296 68816
rect 20048 68776 20088 68816
rect 20130 68776 20170 68816
rect 20212 68776 20252 68816
rect 20294 68776 20334 68816
rect 20376 68776 20416 68816
rect 6412 68608 6452 68648
rect 10348 68608 10388 68648
rect 8332 68524 8372 68564
rect 2380 68440 2420 68480
rect 3628 68440 3668 68480
rect 4108 68440 4148 68480
rect 4204 68440 4244 68480
rect 4396 68440 4436 68480
rect 4684 68440 4724 68480
rect 4780 68440 4820 68480
rect 5164 68440 5204 68480
rect 5740 68440 5780 68480
rect 6220 68435 6260 68475
rect 6591 68451 6631 68491
rect 6892 68440 6932 68480
rect 8140 68440 8180 68480
rect 8620 68440 8660 68480
rect 8716 68440 8756 68480
rect 9196 68440 9236 68480
rect 9676 68440 9716 68480
rect 10156 68435 10196 68475
rect 11500 68440 11540 68480
rect 12748 68440 12788 68480
rect 13708 68440 13748 68480
rect 14956 68440 14996 68480
rect 15340 68440 15380 68480
rect 16588 68440 16628 68480
rect 16972 68440 17012 68480
rect 18220 68440 18260 68480
rect 18604 68440 18644 68480
rect 18700 68440 18740 68480
rect 18892 68440 18932 68480
rect 19084 68440 19124 68480
rect 19276 68440 19316 68480
rect 19372 68440 19412 68480
rect 5260 68356 5300 68396
rect 9100 68356 9140 68396
rect 19372 68272 19412 68312
rect 3820 68188 3860 68228
rect 4396 68188 4436 68228
rect 6700 68188 6740 68228
rect 12940 68188 12980 68228
rect 15148 68188 15188 68228
rect 16780 68188 16820 68228
rect 18412 68188 18452 68228
rect 3688 68020 3728 68060
rect 3770 68020 3810 68060
rect 3852 68020 3892 68060
rect 3934 68020 3974 68060
rect 4016 68020 4056 68060
rect 18808 68020 18848 68060
rect 18890 68020 18930 68060
rect 18972 68020 19012 68060
rect 19054 68020 19094 68060
rect 19136 68020 19176 68060
rect 7372 67852 7412 67892
rect 2860 67684 2900 67724
rect 10156 67684 10196 67724
rect 14188 67684 14228 67724
rect 15340 67684 15380 67724
rect 15436 67684 15476 67724
rect 18028 67684 18068 67724
rect 2380 67600 2420 67640
rect 2476 67600 2516 67640
rect 2956 67600 2996 67640
rect 3436 67600 3476 67640
rect 3964 67609 4004 67649
rect 4492 67600 4532 67640
rect 5740 67600 5780 67640
rect 5932 67600 5972 67640
rect 7180 67600 7220 67640
rect 7852 67600 7892 67640
rect 9100 67600 9140 67640
rect 9580 67600 9620 67640
rect 9676 67600 9716 67640
rect 10060 67600 10100 67640
rect 10636 67600 10676 67640
rect 11116 67605 11156 67645
rect 12076 67600 12116 67640
rect 13324 67600 13364 67640
rect 14092 67600 14132 67640
rect 14284 67600 14324 67640
rect 14860 67600 14900 67640
rect 14956 67600 14996 67640
rect 15916 67600 15956 67640
rect 16396 67605 16436 67645
rect 16780 67600 16820 67640
rect 16972 67600 17012 67640
rect 17068 67600 17108 67640
rect 17548 67600 17588 67640
rect 17644 67600 17684 67640
rect 18124 67600 18164 67640
rect 18604 67600 18644 67640
rect 19084 67605 19124 67645
rect 19468 67600 19508 67640
rect 19564 67600 19604 67640
rect 19660 67600 19700 67640
rect 19948 67600 19988 67640
rect 20236 67600 20276 67640
rect 9292 67516 9332 67556
rect 19276 67516 19316 67556
rect 19756 67516 19796 67556
rect 4108 67432 4148 67472
rect 4300 67432 4340 67472
rect 11308 67432 11348 67472
rect 13516 67432 13556 67472
rect 16588 67432 16628 67472
rect 16876 67432 16916 67472
rect 20044 67432 20084 67472
rect 4928 67264 4968 67304
rect 5010 67264 5050 67304
rect 5092 67264 5132 67304
rect 5174 67264 5214 67304
rect 5256 67264 5296 67304
rect 20048 67264 20088 67304
rect 20130 67264 20170 67304
rect 20212 67264 20252 67304
rect 20294 67264 20334 67304
rect 20376 67264 20416 67304
rect 9676 67096 9716 67136
rect 11692 67096 11732 67136
rect 13804 67096 13844 67136
rect 19468 67096 19508 67136
rect 8908 67012 8948 67052
rect 1708 66928 1748 66968
rect 2956 66928 2996 66968
rect 3532 66928 3572 66968
rect 4780 66928 4820 66968
rect 5356 66928 5396 66968
rect 6604 66928 6644 66968
rect 6796 66928 6836 66968
rect 8044 66928 8084 66968
rect 8620 66928 8660 66968
rect 8716 66928 8756 66968
rect 8812 66928 8852 66968
rect 9100 66928 9140 66968
rect 9292 66928 9332 66968
rect 9388 66928 9428 66968
rect 9580 66928 9620 66968
rect 9772 66928 9812 66968
rect 10252 66928 10292 66968
rect 11500 66928 11540 66968
rect 12076 66928 12116 66968
rect 12172 66928 12212 66968
rect 13132 66928 13172 66968
rect 13612 66923 13652 66963
rect 14188 66928 14228 66968
rect 15436 66928 15476 66968
rect 15628 66928 15668 66968
rect 16876 66928 16916 66968
rect 17260 66928 17300 66968
rect 17356 66928 17396 66968
rect 17548 66928 17588 66968
rect 18028 66928 18068 66968
rect 19276 66928 19316 66968
rect 19756 66928 19796 66968
rect 12556 66844 12596 66884
rect 12652 66844 12692 66884
rect 8236 66760 8276 66800
rect 9388 66760 9428 66800
rect 13996 66760 14036 66800
rect 17548 66760 17588 66800
rect 19756 66760 19796 66800
rect 19948 66760 19988 66800
rect 3148 66676 3188 66716
rect 4972 66676 5012 66716
rect 5164 66676 5204 66716
rect 17068 66676 17108 66716
rect 3688 66508 3728 66548
rect 3770 66508 3810 66548
rect 3852 66508 3892 66548
rect 3934 66508 3974 66548
rect 4016 66508 4056 66548
rect 18808 66508 18848 66548
rect 18890 66508 18930 66548
rect 18972 66508 19012 66548
rect 19054 66508 19094 66548
rect 19136 66508 19176 66548
rect 9100 66340 9140 66380
rect 9676 66340 9716 66380
rect 12364 66340 12404 66380
rect 16108 66340 16148 66380
rect 19852 66340 19892 66380
rect 7180 66256 7220 66296
rect 9964 66256 10004 66296
rect 5068 66172 5108 66212
rect 16876 66172 16916 66212
rect 1228 66088 1268 66128
rect 2476 66088 2516 66128
rect 3532 66088 3572 66128
rect 3628 66088 3668 66128
rect 3724 66088 3764 66128
rect 3916 66088 3956 66128
rect 4012 66088 4052 66128
rect 4108 66088 4148 66128
rect 4204 66088 4244 66128
rect 4492 66088 4532 66128
rect 4588 66088 4628 66128
rect 4972 66088 5012 66128
rect 5548 66088 5588 66128
rect 6028 66093 6068 66133
rect 6508 66088 6548 66128
rect 6796 66088 6836 66128
rect 6892 66088 6932 66128
rect 7660 66088 7700 66128
rect 8908 66088 8948 66128
rect 9388 66088 9428 66128
rect 9676 66081 9716 66121
rect 9964 66088 10004 66128
rect 12364 66088 12404 66128
rect 12556 66088 12596 66128
rect 12748 66088 12788 66128
rect 12844 66088 12884 66128
rect 13036 66088 13076 66128
rect 13132 66088 13172 66128
rect 13228 66088 13268 66128
rect 13516 66107 13556 66147
rect 13612 66088 13652 66128
rect 13804 66088 13844 66128
rect 14188 66088 14228 66128
rect 14284 66088 14324 66128
rect 14476 66088 14516 66128
rect 16012 66088 16052 66128
rect 16300 66088 16340 66128
rect 16396 66088 16436 66128
rect 16492 66088 16532 66128
rect 16588 66088 16628 66128
rect 16780 66088 16820 66128
rect 16972 66088 17012 66128
rect 18412 66088 18452 66128
rect 19660 66088 19700 66128
rect 13708 66004 13748 66044
rect 2668 65920 2708 65960
rect 3436 65920 3476 65960
rect 6220 65920 6260 65960
rect 9100 65920 9140 65960
rect 10156 65920 10196 65960
rect 13324 65920 13364 65960
rect 14380 65920 14420 65960
rect 4928 65752 4968 65792
rect 5010 65752 5050 65792
rect 5092 65752 5132 65792
rect 5174 65752 5214 65792
rect 5256 65752 5296 65792
rect 20048 65752 20088 65792
rect 20130 65752 20170 65792
rect 20212 65752 20252 65792
rect 20294 65752 20334 65792
rect 20376 65752 20416 65792
rect 5932 65584 5972 65624
rect 9292 65584 9332 65624
rect 9484 65584 9524 65624
rect 13036 65584 13076 65624
rect 3340 65500 3380 65540
rect 6508 65500 6548 65540
rect 13324 65500 13364 65540
rect 15916 65500 15956 65540
rect 17932 65500 17972 65540
rect 1612 65416 1652 65456
rect 1708 65416 1748 65456
rect 2092 65416 2132 65456
rect 2188 65416 2228 65456
rect 2668 65416 2708 65456
rect 3148 65411 3188 65451
rect 4300 65416 4340 65456
rect 5548 65416 5588 65456
rect 6124 65416 6164 65456
rect 6220 65416 6260 65456
rect 6412 65416 6452 65456
rect 6604 65416 6644 65456
rect 6700 65416 6740 65456
rect 6988 65416 7028 65456
rect 7276 65416 7316 65456
rect 7564 65416 7604 65456
rect 7660 65416 7700 65456
rect 8044 65416 8084 65456
rect 8140 65416 8180 65456
rect 8620 65416 8660 65456
rect 9100 65411 9140 65451
rect 9676 65416 9716 65456
rect 10924 65416 10964 65456
rect 11116 65416 11156 65456
rect 12364 65416 12404 65456
rect 12748 65416 12788 65456
rect 12844 65416 12884 65456
rect 12940 65437 12980 65477
rect 13228 65416 13268 65456
rect 13420 65416 13460 65456
rect 13516 65416 13556 65456
rect 14476 65416 14516 65456
rect 15724 65416 15764 65456
rect 16204 65416 16244 65456
rect 16300 65416 16340 65456
rect 16684 65416 16724 65456
rect 17260 65416 17300 65456
rect 17740 65402 17780 65442
rect 16780 65332 16820 65372
rect 6988 65248 7028 65288
rect 12556 65248 12596 65288
rect 5740 65164 5780 65204
rect 3688 64996 3728 65036
rect 3770 64996 3810 65036
rect 3852 64996 3892 65036
rect 3934 64996 3974 65036
rect 4016 64996 4056 65036
rect 18808 64996 18848 65036
rect 18890 64996 18930 65036
rect 18972 64996 19012 65036
rect 19054 64996 19094 65036
rect 19136 64996 19176 65036
rect 11020 64828 11060 64868
rect 13708 64828 13748 64868
rect 17644 64828 17684 64868
rect 5260 64660 5300 64700
rect 11788 64660 11828 64700
rect 11884 64660 11924 64700
rect 1228 64576 1268 64616
rect 2476 64576 2516 64616
rect 3532 64576 3572 64616
rect 4780 64576 4820 64616
rect 5164 64576 5204 64616
rect 5356 64576 5396 64616
rect 5548 64576 5588 64616
rect 6796 64576 6836 64616
rect 7372 64576 7412 64616
rect 8620 64576 8660 64616
rect 8908 64576 8948 64616
rect 9004 64576 9044 64616
rect 9580 64576 9620 64616
rect 10828 64576 10868 64616
rect 11308 64576 11348 64616
rect 11404 64576 11444 64616
rect 12364 64576 12404 64616
rect 12844 64581 12884 64621
rect 13228 64576 13268 64616
rect 13324 64576 13364 64616
rect 13420 64576 13460 64616
rect 13516 64576 13556 64616
rect 13708 64576 13748 64616
rect 13900 64576 13940 64616
rect 14092 64576 14132 64616
rect 15340 64576 15380 64616
rect 15724 64576 15764 64616
rect 16012 64576 16052 64616
rect 16204 64576 16244 64616
rect 17452 64576 17492 64616
rect 17836 64576 17876 64616
rect 7180 64492 7220 64532
rect 13036 64492 13076 64532
rect 2668 64408 2708 64448
rect 4972 64408 5012 64448
rect 6988 64408 7028 64448
rect 9196 64408 9236 64448
rect 15532 64408 15572 64448
rect 15916 64408 15956 64448
rect 17932 64408 17972 64448
rect 4928 64240 4968 64280
rect 5010 64240 5050 64280
rect 5092 64240 5132 64280
rect 5174 64240 5214 64280
rect 5256 64240 5296 64280
rect 20048 64240 20088 64280
rect 20130 64240 20170 64280
rect 20212 64240 20252 64280
rect 20294 64240 20334 64280
rect 20376 64240 20416 64280
rect 4012 64072 4052 64112
rect 7180 64072 7220 64112
rect 8332 64072 8372 64112
rect 12268 64072 12308 64112
rect 8140 64030 8180 64070
rect 17356 64072 17396 64112
rect 18028 64072 18068 64112
rect 12940 63988 12980 64028
rect 15532 64030 15572 64070
rect 2284 63904 2324 63944
rect 2380 63904 2420 63944
rect 2764 63904 2804 63944
rect 2860 63904 2900 63944
rect 3340 63904 3380 63944
rect 3820 63899 3860 63939
rect 5452 63904 5492 63944
rect 5548 63904 5588 63944
rect 6028 63904 6068 63944
rect 6508 63904 6548 63944
rect 6988 63899 7028 63939
rect 7852 63904 7892 63944
rect 7948 63904 7988 63944
rect 8428 63904 8468 63944
rect 8812 63904 8852 63944
rect 10060 63904 10100 63944
rect 10828 63904 10868 63944
rect 12076 63904 12116 63944
rect 12556 63904 12596 63944
rect 12844 63904 12884 63944
rect 13804 63904 13844 63944
rect 13900 63904 13940 63944
rect 14380 63904 14420 63944
rect 14860 63904 14900 63944
rect 15340 63890 15380 63930
rect 15724 63904 15764 63944
rect 15916 63904 15956 63944
rect 16012 63904 16052 63944
rect 16204 63904 16244 63944
rect 16396 63904 16436 63944
rect 16492 63904 16532 63944
rect 16780 63904 16820 63944
rect 17351 63904 17391 63944
rect 17452 63904 17492 63944
rect 17548 63904 17588 63944
rect 17740 63904 17780 63944
rect 17836 63904 17876 63944
rect 18220 63904 18260 63944
rect 18316 63904 18356 63944
rect 5932 63820 5972 63860
rect 14284 63820 14324 63860
rect 13228 63736 13268 63776
rect 16492 63736 16532 63776
rect 16780 63736 16820 63776
rect 8620 63652 8660 63692
rect 10252 63652 10292 63692
rect 16972 63652 17012 63692
rect 3688 63484 3728 63524
rect 3770 63484 3810 63524
rect 3852 63484 3892 63524
rect 3934 63484 3974 63524
rect 4016 63484 4056 63524
rect 18808 63484 18848 63524
rect 18890 63484 18930 63524
rect 18972 63484 19012 63524
rect 19054 63484 19094 63524
rect 19136 63484 19176 63524
rect 14668 63316 14708 63356
rect 14860 63316 14900 63356
rect 17932 63316 17972 63356
rect 18124 63232 18164 63272
rect 3244 63148 3284 63188
rect 3340 63148 3380 63188
rect 8140 63148 8180 63188
rect 8236 63148 8276 63188
rect 2764 63083 2804 63123
rect 2860 63064 2900 63104
rect 3820 63064 3860 63104
rect 4300 63078 4340 63118
rect 5932 63064 5972 63104
rect 7180 63064 7220 63104
rect 7660 63064 7700 63104
rect 7756 63064 7796 63104
rect 8716 63064 8756 63104
rect 9196 63078 9236 63118
rect 9772 63064 9812 63104
rect 9868 63064 9908 63104
rect 10060 63064 10100 63104
rect 10252 63106 10292 63146
rect 11212 63148 11252 63188
rect 10348 63064 10388 63104
rect 10444 63064 10484 63104
rect 10540 63064 10580 63104
rect 10732 63064 10772 63104
rect 10924 63064 10964 63104
rect 11116 63064 11156 63104
rect 12556 63064 12596 63104
rect 12652 63064 12692 63104
rect 13228 63064 13268 63104
rect 14476 63064 14516 63104
rect 15052 63064 15092 63104
rect 16300 63064 16340 63104
rect 16492 63064 16532 63104
rect 17740 63064 17780 63104
rect 18124 63064 18164 63104
rect 18220 63064 18260 63104
rect 18412 63064 18452 63104
rect 4492 62980 4532 63020
rect 7372 62980 7412 63020
rect 9388 62980 9428 63020
rect 9964 62980 10004 63020
rect 10828 62980 10868 63020
rect 12844 62896 12884 62936
rect 14668 62896 14708 62936
rect 14860 62896 14900 62936
rect 4928 62728 4968 62768
rect 5010 62728 5050 62768
rect 5092 62728 5132 62768
rect 5174 62728 5214 62768
rect 5256 62728 5296 62768
rect 20048 62728 20088 62768
rect 20130 62728 20170 62768
rect 20212 62728 20252 62768
rect 20294 62728 20334 62768
rect 20376 62728 20416 62768
rect 9388 62560 9428 62600
rect 9868 62560 9908 62600
rect 13708 62560 13748 62600
rect 15052 62560 15092 62600
rect 15724 62560 15764 62600
rect 17932 62560 17972 62600
rect 1708 62392 1748 62432
rect 2956 62392 2996 62432
rect 4204 62392 4244 62432
rect 5452 62392 5492 62432
rect 5836 62392 5876 62432
rect 7084 62392 7124 62432
rect 7468 62392 7508 62432
rect 8716 62392 8756 62432
rect 9100 62392 9140 62432
rect 9196 62392 9236 62432
rect 9292 62392 9332 62432
rect 9580 62392 9620 62432
rect 9676 62392 9716 62432
rect 9772 62392 9812 62432
rect 10252 62392 10292 62432
rect 11500 62392 11540 62432
rect 11980 62392 12020 62432
rect 12076 62392 12116 62432
rect 12460 62392 12500 62432
rect 13036 62392 13076 62432
rect 13516 62378 13556 62418
rect 14764 62392 14804 62432
rect 14860 62392 14900 62432
rect 14956 62392 14996 62432
rect 15244 62392 15284 62432
rect 15340 62392 15380 62432
rect 15436 62392 15476 62432
rect 15532 62392 15572 62432
rect 15820 62392 15860 62432
rect 16492 62392 16532 62432
rect 17740 62392 17780 62432
rect 12556 62308 12596 62348
rect 11692 62224 11732 62264
rect 3148 62140 3188 62180
rect 5644 62140 5684 62180
rect 7276 62140 7316 62180
rect 8908 62140 8948 62180
rect 16012 62140 16052 62180
rect 3688 61972 3728 62012
rect 3770 61972 3810 62012
rect 3852 61972 3892 62012
rect 3934 61972 3974 62012
rect 4016 61972 4056 62012
rect 18808 61972 18848 62012
rect 18890 61972 18930 62012
rect 18972 61972 19012 62012
rect 19054 61972 19094 62012
rect 19136 61972 19176 62012
rect 13612 61804 13652 61844
rect 2668 61636 2708 61676
rect 6220 61636 6260 61676
rect 2188 61552 2228 61592
rect 2284 61552 2324 61592
rect 2764 61552 2804 61592
rect 3244 61552 3284 61592
rect 3724 61566 3764 61606
rect 5644 61552 5684 61592
rect 5740 61552 5780 61592
rect 6124 61552 6164 61592
rect 6700 61552 6740 61592
rect 7180 61566 7220 61606
rect 7756 61552 7796 61592
rect 9004 61552 9044 61592
rect 9676 61552 9716 61592
rect 10924 61552 10964 61592
rect 12172 61552 12212 61592
rect 13420 61552 13460 61592
rect 14380 61552 14420 61592
rect 14572 61552 14612 61592
rect 14764 61552 14804 61592
rect 14860 61552 14900 61592
rect 15244 61531 15284 61571
rect 15340 61531 15380 61571
rect 15436 61531 15476 61571
rect 15916 61552 15956 61592
rect 17164 61552 17204 61592
rect 3916 61468 3956 61508
rect 7564 61468 7604 61508
rect 7372 61384 7412 61424
rect 11116 61384 11156 61424
rect 14476 61384 14516 61424
rect 15052 61384 15092 61424
rect 15532 61384 15572 61424
rect 15724 61384 15764 61424
rect 4928 61216 4968 61256
rect 5010 61216 5050 61256
rect 5092 61216 5132 61256
rect 5174 61216 5214 61256
rect 5256 61216 5296 61256
rect 20048 61216 20088 61256
rect 20130 61216 20170 61256
rect 20212 61216 20252 61256
rect 20294 61216 20334 61256
rect 20376 61216 20416 61256
rect 10924 61048 10964 61088
rect 15628 61048 15668 61088
rect 4588 60964 4628 61004
rect 6796 60964 6836 61004
rect 8908 60964 8948 61004
rect 2860 60880 2900 60920
rect 2956 60880 2996 60920
rect 3436 60880 3476 60920
rect 3916 60880 3956 60920
rect 4444 60870 4484 60910
rect 5068 60880 5108 60920
rect 5356 60880 5396 60920
rect 6604 60880 6644 60920
rect 6988 60880 7028 60920
rect 7180 60880 7220 60920
rect 7276 60880 7316 60920
rect 7468 60880 7508 60920
rect 8716 60880 8756 60920
rect 9196 60880 9236 60920
rect 9292 60880 9332 60920
rect 9676 60880 9716 60920
rect 10252 60880 10292 60920
rect 10780 60870 10820 60910
rect 11116 60880 11156 60920
rect 12364 60859 12404 60899
rect 12748 60880 12788 60920
rect 12844 60880 12884 60920
rect 13036 60880 13076 60920
rect 13900 60880 13940 60920
rect 13996 60880 14036 60920
rect 14380 60880 14420 60920
rect 14956 60880 14996 60920
rect 15436 60866 15476 60906
rect 15820 60880 15860 60920
rect 16012 60880 16052 60920
rect 16108 60880 16148 60920
rect 16396 60880 16436 60920
rect 17644 60880 17684 60920
rect 18220 60880 18260 60920
rect 19468 60880 19508 60920
rect 3340 60796 3380 60836
rect 9772 60796 9812 60836
rect 14476 60796 14516 60836
rect 7276 60712 7316 60752
rect 12940 60712 12980 60752
rect 5164 60628 5204 60668
rect 12556 60628 12596 60668
rect 15820 60628 15860 60668
rect 17836 60628 17876 60668
rect 19660 60628 19700 60668
rect 3688 60460 3728 60500
rect 3770 60460 3810 60500
rect 3852 60460 3892 60500
rect 3934 60460 3974 60500
rect 4016 60460 4056 60500
rect 18808 60460 18848 60500
rect 18890 60460 18930 60500
rect 18972 60460 19012 60500
rect 19054 60460 19094 60500
rect 19136 60460 19176 60500
rect 14188 60292 14228 60332
rect 9676 60124 9716 60164
rect 9772 60124 9812 60164
rect 1420 60040 1460 60080
rect 2668 60040 2708 60080
rect 4300 60040 4340 60080
rect 5356 60040 5396 60080
rect 6604 60040 6644 60080
rect 6988 60040 7028 60080
rect 3052 59998 3092 60038
rect 7084 60040 7124 60080
rect 7468 60040 7508 60080
rect 8716 60040 8756 60080
rect 9196 60040 9236 60080
rect 9292 60040 9332 60080
rect 10252 60040 10292 60080
rect 10732 60049 10772 60089
rect 11884 60040 11924 60080
rect 12268 60040 12308 60080
rect 12364 60040 12404 60080
rect 12748 60040 12788 60080
rect 12844 60040 12884 60080
rect 13324 60040 13364 60080
rect 13804 60045 13844 60085
rect 14380 60040 14420 60080
rect 15628 60040 15668 60080
rect 15820 60040 15860 60080
rect 17068 60040 17108 60080
rect 17548 60040 17588 60080
rect 17644 60040 17684 60080
rect 18028 60040 18068 60080
rect 18124 60040 18164 60080
rect 18604 60040 18644 60080
rect 19084 60054 19124 60094
rect 6796 59956 6836 59996
rect 8908 59956 8948 59996
rect 2860 59872 2900 59912
rect 4492 59872 4532 59912
rect 7276 59872 7316 59912
rect 10924 59872 10964 59912
rect 11980 59872 12020 59912
rect 13996 59872 14036 59912
rect 17260 59872 17300 59912
rect 19276 59872 19316 59912
rect 4928 59704 4968 59744
rect 5010 59704 5050 59744
rect 5092 59704 5132 59744
rect 5174 59704 5214 59744
rect 5256 59704 5296 59744
rect 20048 59704 20088 59744
rect 20130 59704 20170 59744
rect 20212 59704 20252 59744
rect 20294 59704 20334 59744
rect 20376 59704 20416 59744
rect 10924 59536 10964 59576
rect 12748 59536 12788 59576
rect 14380 59536 14420 59576
rect 14572 59536 14612 59576
rect 4300 59452 4340 59492
rect 17164 59452 17204 59492
rect 19276 59452 19316 59492
rect 2572 59368 2612 59408
rect 2668 59368 2708 59408
rect 3052 59368 3092 59408
rect 3148 59368 3188 59408
rect 3628 59368 3668 59408
rect 4156 59358 4196 59398
rect 5164 59368 5204 59408
rect 6412 59368 6452 59408
rect 6796 59368 6836 59408
rect 8044 59368 8084 59408
rect 8428 59368 8468 59408
rect 8524 59368 8564 59408
rect 8716 59368 8756 59408
rect 8812 59368 8852 59408
rect 8913 59368 8953 59408
rect 9484 59368 9524 59408
rect 10732 59368 10772 59408
rect 11308 59368 11348 59408
rect 12556 59368 12596 59408
rect 12940 59368 12980 59408
rect 14188 59368 14228 59408
rect 14764 59368 14804 59408
rect 16012 59368 16052 59408
rect 16300 59368 16340 59408
rect 17548 59368 17588 59408
rect 17644 59368 17684 59408
rect 18604 59368 18644 59408
rect 19084 59354 19124 59394
rect 2092 59284 2132 59324
rect 18028 59284 18068 59324
rect 18124 59284 18164 59324
rect 1900 59116 1940 59156
rect 6604 59116 6644 59156
rect 8236 59116 8276 59156
rect 8428 59116 8468 59156
rect 12748 59116 12788 59156
rect 16972 59116 17012 59156
rect 3688 58948 3728 58988
rect 3770 58948 3810 58988
rect 3852 58948 3892 58988
rect 3934 58948 3974 58988
rect 4016 58948 4056 58988
rect 18808 58948 18848 58988
rect 18890 58948 18930 58988
rect 18972 58948 19012 58988
rect 19054 58948 19094 58988
rect 19136 58948 19176 58988
rect 19852 58780 19892 58820
rect 12556 58696 12596 58736
rect 15532 58696 15572 58736
rect 1228 58528 1268 58568
rect 2476 58528 2516 58568
rect 3724 58528 3764 58568
rect 4972 58528 5012 58568
rect 5356 58528 5396 58568
rect 6604 58528 6644 58568
rect 7372 58528 7412 58568
rect 8620 58528 8660 58568
rect 9004 58528 9044 58568
rect 10252 58528 10292 58568
rect 11116 58528 11156 58568
rect 12364 58528 12404 58568
rect 12839 58528 12879 58568
rect 12940 58528 12980 58568
rect 13036 58528 13076 58568
rect 13228 58528 13268 58568
rect 13324 58528 13364 58568
rect 13516 58528 13556 58568
rect 13612 58528 13652 58568
rect 14092 58528 14132 58568
rect 15340 58528 15380 58568
rect 16012 58528 16052 58568
rect 16108 58528 16148 58568
rect 16300 58528 16340 58568
rect 16396 58528 16436 58568
rect 16492 58528 16532 58568
rect 16588 58528 16628 58568
rect 16780 58528 16820 58568
rect 18028 58528 18068 58568
rect 18412 58528 18452 58568
rect 19660 58528 19700 58568
rect 2668 58360 2708 58400
rect 5164 58360 5204 58400
rect 6796 58360 6836 58400
rect 8812 58360 8852 58400
rect 10444 58360 10484 58400
rect 13132 58360 13172 58400
rect 13804 58360 13844 58400
rect 15820 58360 15860 58400
rect 18220 58360 18260 58400
rect 4928 58192 4968 58232
rect 5010 58192 5050 58232
rect 5092 58192 5132 58232
rect 5174 58192 5214 58232
rect 5256 58192 5296 58232
rect 20048 58192 20088 58232
rect 20130 58192 20170 58232
rect 20212 58192 20252 58232
rect 20294 58192 20334 58232
rect 20376 58192 20416 58232
rect 5356 57940 5396 57980
rect 10156 57940 10196 57980
rect 2092 57856 2132 57896
rect 3340 57856 3380 57896
rect 3628 57856 3668 57896
rect 3724 57856 3764 57896
rect 4684 57856 4724 57896
rect 5212 57846 5252 57886
rect 6316 57856 6356 57896
rect 7564 57856 7604 57896
rect 8428 57856 8468 57896
rect 8524 57856 8564 57896
rect 8908 57856 8948 57896
rect 9484 57856 9524 57896
rect 9964 57851 10004 57891
rect 11692 57856 11732 57896
rect 12940 57856 12980 57896
rect 13516 57856 13556 57896
rect 14764 57856 14804 57896
rect 15916 57856 15956 57896
rect 17164 57856 17204 57896
rect 17548 57856 17588 57896
rect 17644 57856 17684 57896
rect 4108 57772 4148 57812
rect 4204 57772 4244 57812
rect 9004 57772 9044 57812
rect 11500 57772 11540 57812
rect 11308 57688 11348 57728
rect 13324 57688 13364 57728
rect 1900 57604 1940 57644
rect 7756 57604 7796 57644
rect 13132 57604 13172 57644
rect 17356 57604 17396 57644
rect 3688 57436 3728 57476
rect 3770 57436 3810 57476
rect 3852 57436 3892 57476
rect 3934 57436 3974 57476
rect 4016 57436 4056 57476
rect 18808 57436 18848 57476
rect 18890 57436 18930 57476
rect 18972 57436 19012 57476
rect 19054 57436 19094 57476
rect 19136 57436 19176 57476
rect 1804 57268 1844 57308
rect 16300 57268 16340 57308
rect 1996 57100 2036 57140
rect 7756 57100 7796 57140
rect 9676 57100 9716 57140
rect 12172 57100 12212 57140
rect 14284 57100 14324 57140
rect 14380 57100 14420 57140
rect 16012 57100 16052 57140
rect 16492 57100 16532 57140
rect 2188 57016 2228 57056
rect 3436 57016 3476 57056
rect 3820 57016 3860 57056
rect 5068 57016 5108 57056
rect 5452 57016 5492 57056
rect 6700 57016 6740 57056
rect 7180 57016 7220 57056
rect 7276 57016 7316 57056
rect 7660 57016 7700 57056
rect 8236 57016 8276 57056
rect 8716 57030 8756 57070
rect 9868 57016 9908 57056
rect 11116 57016 11156 57056
rect 11596 57016 11636 57056
rect 11692 57016 11732 57056
rect 12076 57016 12116 57056
rect 12652 57016 12692 57056
rect 13132 57030 13172 57070
rect 13804 57016 13844 57056
rect 13900 57016 13940 57056
rect 14860 57016 14900 57056
rect 15340 57030 15380 57070
rect 16780 57016 16820 57056
rect 16876 57016 16916 57056
rect 17260 57016 17300 57056
rect 17356 57016 17396 57056
rect 17836 57016 17876 57056
rect 18316 57030 18356 57070
rect 20140 57058 20180 57098
rect 18892 57016 18932 57056
rect 8908 56932 8948 56972
rect 11308 56932 11348 56972
rect 13324 56932 13364 56972
rect 18508 56932 18548 56972
rect 3628 56848 3668 56888
rect 5260 56848 5300 56888
rect 6892 56848 6932 56888
rect 9484 56848 9524 56888
rect 15532 56848 15572 56888
rect 15820 56848 15860 56888
rect 18700 56848 18740 56888
rect 4928 56680 4968 56720
rect 5010 56680 5050 56720
rect 5092 56680 5132 56720
rect 5174 56680 5214 56720
rect 5256 56680 5296 56720
rect 20048 56680 20088 56720
rect 20130 56680 20170 56720
rect 20212 56680 20252 56720
rect 20294 56680 20334 56720
rect 20376 56680 20416 56720
rect 12364 56512 12404 56552
rect 16684 56512 16724 56552
rect 16876 56512 16916 56552
rect 19564 56512 19604 56552
rect 3052 56428 3092 56468
rect 7180 56428 7220 56468
rect 9196 56428 9236 56468
rect 19180 56428 19220 56468
rect 1420 56344 1460 56384
rect 2668 56344 2708 56384
rect 3244 56339 3284 56379
rect 3724 56344 3764 56384
rect 4204 56344 4244 56384
rect 4684 56344 4724 56384
rect 4780 56344 4820 56384
rect 5740 56344 5780 56384
rect 6988 56344 7028 56384
rect 7468 56344 7508 56384
rect 7564 56344 7604 56384
rect 7948 56344 7988 56384
rect 8044 56344 8084 56384
rect 8524 56344 8564 56384
rect 9004 56339 9044 56379
rect 10732 56344 10772 56384
rect 13228 56344 13268 56384
rect 14476 56344 14516 56384
rect 15244 56344 15284 56384
rect 16492 56344 16532 56384
rect 17452 56344 17492 56384
rect 11980 56302 12020 56342
rect 17548 56344 17588 56384
rect 17932 56344 17972 56384
rect 18508 56344 18548 56384
rect 18988 56339 19028 56379
rect 4300 56260 4340 56300
rect 10348 56260 10388 56300
rect 12556 56260 12596 56300
rect 15052 56260 15092 56300
rect 17068 56260 17108 56300
rect 18028 56260 18068 56300
rect 19372 56260 19412 56300
rect 2860 56176 2900 56216
rect 10540 56092 10580 56132
rect 12172 56092 12212 56132
rect 14668 56092 14708 56132
rect 14860 56092 14900 56132
rect 3688 55924 3728 55964
rect 3770 55924 3810 55964
rect 3852 55924 3892 55964
rect 3934 55924 3974 55964
rect 4016 55924 4056 55964
rect 18808 55924 18848 55964
rect 18890 55924 18930 55964
rect 18972 55924 19012 55964
rect 19054 55924 19094 55964
rect 19136 55924 19176 55964
rect 2860 55672 2900 55712
rect 19564 55672 19604 55712
rect 3244 55588 3284 55628
rect 5644 55588 5684 55628
rect 5740 55588 5780 55628
rect 8428 55588 8468 55628
rect 8524 55588 8564 55628
rect 10060 55599 10100 55639
rect 11212 55588 11252 55628
rect 11308 55588 11348 55628
rect 19372 55588 19412 55628
rect 1420 55504 1460 55544
rect 2668 55504 2708 55544
rect 3436 55504 3476 55544
rect 4684 55504 4724 55544
rect 5164 55504 5204 55544
rect 5260 55504 5300 55544
rect 6220 55504 6260 55544
rect 6700 55518 6740 55558
rect 7948 55504 7988 55544
rect 8044 55504 8084 55544
rect 9004 55504 9044 55544
rect 9484 55509 9524 55549
rect 10732 55504 10772 55544
rect 10828 55504 10868 55544
rect 11788 55504 11828 55544
rect 12268 55518 12308 55558
rect 13132 55504 13172 55544
rect 14380 55504 14420 55544
rect 15052 55504 15092 55544
rect 16300 55504 16340 55544
rect 16876 55504 16916 55544
rect 18124 55504 18164 55544
rect 6892 55420 6932 55460
rect 9676 55420 9716 55460
rect 12460 55420 12500 55460
rect 3052 55336 3092 55376
rect 4876 55336 4916 55376
rect 9868 55336 9908 55376
rect 14572 55336 14612 55376
rect 16492 55336 16532 55376
rect 16684 55336 16724 55376
rect 4928 55168 4968 55208
rect 5010 55168 5050 55208
rect 5092 55168 5132 55208
rect 5174 55168 5214 55208
rect 5256 55168 5296 55208
rect 20048 55168 20088 55208
rect 20130 55168 20170 55208
rect 20212 55168 20252 55208
rect 20294 55168 20334 55208
rect 20376 55168 20416 55208
rect 9388 55000 9428 55040
rect 11020 55000 11060 55040
rect 16780 55000 16820 55040
rect 20236 55000 20276 55040
rect 2188 54916 2228 54956
rect 12748 54916 12788 54956
rect 14764 54916 14804 54956
rect 19084 54916 19124 54956
rect 2332 54822 2372 54862
rect 2860 54832 2900 54872
rect 3340 54832 3380 54872
rect 3820 54832 3860 54872
rect 3916 54832 3956 54872
rect 5452 54832 5492 54872
rect 6700 54832 6740 54872
rect 7948 54832 7988 54872
rect 9196 54832 9236 54872
rect 9580 54832 9620 54872
rect 10828 54832 10868 54872
rect 11308 54832 11348 54872
rect 12556 54811 12596 54851
rect 13036 54832 13076 54872
rect 13132 54832 13172 54872
rect 13612 54832 13652 54872
rect 14092 54832 14132 54872
rect 14572 54827 14612 54867
rect 15052 54832 15092 54872
rect 15148 54832 15188 54872
rect 15532 54832 15572 54872
rect 15628 54832 15668 54872
rect 16108 54832 16148 54872
rect 16588 54827 16628 54867
rect 17356 54832 17396 54872
rect 17452 54832 17492 54872
rect 17932 54832 17972 54872
rect 18412 54832 18452 54872
rect 1996 54748 2036 54788
rect 3436 54748 3476 54788
rect 13516 54748 13556 54788
rect 17836 54748 17876 54788
rect 18940 54790 18980 54830
rect 19468 54748 19508 54788
rect 19660 54748 19700 54788
rect 20044 54748 20084 54788
rect 1804 54580 1844 54620
rect 6892 54580 6932 54620
rect 19276 54580 19316 54620
rect 19852 54580 19892 54620
rect 3688 54412 3728 54452
rect 3770 54412 3810 54452
rect 3852 54412 3892 54452
rect 3934 54412 3974 54452
rect 4016 54412 4056 54452
rect 18808 54412 18848 54452
rect 18890 54412 18930 54452
rect 18972 54412 19012 54452
rect 19054 54412 19094 54452
rect 19136 54412 19176 54452
rect 19276 54244 19316 54284
rect 17164 54160 17204 54200
rect 9964 54076 10004 54116
rect 12172 54076 12212 54116
rect 17356 54076 17396 54116
rect 19468 54076 19508 54116
rect 19852 54076 19892 54116
rect 1228 53992 1268 54032
rect 2476 53992 2516 54032
rect 3340 53992 3380 54032
rect 3436 53992 3476 54032
rect 3820 53992 3860 54032
rect 3916 53992 3956 54032
rect 4396 53992 4436 54032
rect 4876 54006 4916 54046
rect 6700 53992 6740 54032
rect 7948 53992 7988 54032
rect 8332 53992 8372 54032
rect 9580 53992 9620 54032
rect 10348 53992 10388 54032
rect 11596 53992 11636 54032
rect 13804 53992 13844 54032
rect 15052 53992 15092 54032
rect 15532 53992 15572 54032
rect 16780 53992 16820 54032
rect 17836 53992 17876 54032
rect 19084 53992 19124 54032
rect 5068 53908 5108 53948
rect 2668 53824 2708 53864
rect 8140 53824 8180 53864
rect 9772 53824 9812 53864
rect 10156 53824 10196 53864
rect 11788 53824 11828 53864
rect 11980 53824 12020 53864
rect 15244 53824 15284 53864
rect 16972 53824 17012 53864
rect 19660 53824 19700 53864
rect 20044 53824 20084 53864
rect 4928 53656 4968 53696
rect 5010 53656 5050 53696
rect 5092 53656 5132 53696
rect 5174 53656 5214 53696
rect 5256 53656 5296 53696
rect 20048 53656 20088 53696
rect 20130 53656 20170 53696
rect 20212 53656 20252 53696
rect 20294 53656 20334 53696
rect 20376 53656 20416 53696
rect 3148 53488 3188 53528
rect 9292 53488 9332 53528
rect 16876 53488 16916 53528
rect 2956 53404 2996 53444
rect 7276 53404 7316 53444
rect 1516 53320 1556 53360
rect 2764 53320 2804 53360
rect 3292 53310 3332 53350
rect 3820 53320 3860 53360
rect 4780 53320 4820 53360
rect 4876 53320 4916 53360
rect 5836 53320 5876 53360
rect 7084 53320 7124 53360
rect 7564 53320 7604 53360
rect 7660 53320 7700 53360
rect 8620 53320 8660 53360
rect 9100 53315 9140 53355
rect 9484 53320 9524 53360
rect 10732 53320 10772 53360
rect 11116 53320 11156 53360
rect 12364 53320 12404 53360
rect 12748 53320 12788 53360
rect 13996 53320 14036 53360
rect 15148 53320 15188 53360
rect 15244 53320 15284 53360
rect 15724 53320 15764 53360
rect 16204 53320 16244 53360
rect 16684 53315 16724 53355
rect 18508 53320 18548 53360
rect 19756 53320 19796 53360
rect 4300 53236 4340 53276
rect 4396 53236 4436 53276
rect 8044 53236 8084 53276
rect 8140 53236 8180 53276
rect 15628 53236 15668 53276
rect 17260 53236 17300 53276
rect 14188 53152 14228 53192
rect 10924 53068 10964 53108
rect 12556 53068 12596 53108
rect 17068 53068 17108 53108
rect 19948 53068 19988 53108
rect 3688 52900 3728 52940
rect 3770 52900 3810 52940
rect 3852 52900 3892 52940
rect 3934 52900 3974 52940
rect 4016 52900 4056 52940
rect 18808 52900 18848 52940
rect 18890 52900 18930 52940
rect 18972 52900 19012 52940
rect 19054 52900 19094 52940
rect 19136 52900 19176 52940
rect 1804 52732 1844 52772
rect 1612 52564 1652 52604
rect 1996 52564 2036 52604
rect 10924 52564 10964 52604
rect 19564 52564 19604 52604
rect 19756 52564 19796 52604
rect 2380 52480 2420 52520
rect 3628 52480 3668 52520
rect 3820 52480 3860 52520
rect 5068 52480 5108 52520
rect 6892 52480 6932 52520
rect 6988 52480 7028 52520
rect 7372 52480 7412 52520
rect 7468 52480 7508 52520
rect 7948 52480 7988 52520
rect 8428 52494 8468 52534
rect 10348 52480 10388 52520
rect 10444 52480 10484 52520
rect 10828 52480 10868 52520
rect 11404 52480 11444 52520
rect 11884 52494 11924 52534
rect 12652 52480 12692 52520
rect 12748 52480 12788 52520
rect 13132 52480 13172 52520
rect 13228 52480 13268 52520
rect 13719 52479 13759 52519
rect 14188 52494 14228 52534
rect 14572 52480 14612 52520
rect 15820 52480 15860 52520
rect 17452 52480 17492 52520
rect 18700 52480 18740 52520
rect 8620 52396 8660 52436
rect 12076 52396 12116 52436
rect 14380 52396 14420 52436
rect 1420 52312 1460 52352
rect 2188 52312 2228 52352
rect 5260 52312 5300 52352
rect 16012 52312 16052 52352
rect 18892 52312 18932 52352
rect 19372 52312 19412 52352
rect 19948 52312 19988 52352
rect 4928 52144 4968 52184
rect 5010 52144 5050 52184
rect 5092 52144 5132 52184
rect 5174 52144 5214 52184
rect 5256 52144 5296 52184
rect 20048 52144 20088 52184
rect 20130 52144 20170 52184
rect 20212 52144 20252 52184
rect 20294 52144 20334 52184
rect 20376 52144 20416 52184
rect 17452 51976 17492 52016
rect 20044 51976 20084 52016
rect 2380 51892 2420 51932
rect 2572 51803 2612 51843
rect 3052 51808 3092 51848
rect 3532 51808 3572 51848
rect 4012 51808 4052 51848
rect 4108 51808 4148 51848
rect 5932 51808 5972 51848
rect 7180 51808 7220 51848
rect 8620 51808 8660 51848
rect 9868 51808 9908 51848
rect 10252 51808 10292 51848
rect 11500 51808 11540 51848
rect 11884 51808 11924 51848
rect 13132 51808 13172 51848
rect 13516 51808 13556 51848
rect 14764 51808 14804 51848
rect 15724 51808 15764 51848
rect 15820 51808 15860 51848
rect 16300 51808 16340 51848
rect 16780 51808 16820 51848
rect 17260 51794 17300 51834
rect 18316 51808 18356 51848
rect 18412 51808 18452 51848
rect 18892 51808 18932 51848
rect 19372 51808 19412 51848
rect 19852 51803 19892 51843
rect 1708 51724 1748 51764
rect 2092 51724 2132 51764
rect 3628 51724 3668 51764
rect 16204 51724 16244 51764
rect 18796 51724 18836 51764
rect 1516 51556 1556 51596
rect 1900 51556 1940 51596
rect 7372 51556 7412 51596
rect 10060 51556 10100 51596
rect 11692 51556 11732 51596
rect 13324 51556 13364 51596
rect 14956 51556 14996 51596
rect 3688 51388 3728 51428
rect 3770 51388 3810 51428
rect 3852 51388 3892 51428
rect 3934 51388 3974 51428
rect 4016 51388 4056 51428
rect 18808 51388 18848 51428
rect 18890 51388 18930 51428
rect 18972 51388 19012 51428
rect 19054 51388 19094 51428
rect 19136 51388 19176 51428
rect 2860 51220 2900 51260
rect 12364 51220 12404 51260
rect 17644 51220 17684 51260
rect 3052 51052 3092 51092
rect 5932 51052 5972 51092
rect 8044 51052 8084 51092
rect 12556 51052 12596 51092
rect 19756 51052 19796 51092
rect 19948 51052 19988 51092
rect 1228 50968 1268 51008
rect 2476 50968 2516 51008
rect 3340 50968 3380 51008
rect 4588 50968 4628 51008
rect 5356 50968 5396 51008
rect 5452 50968 5492 51008
rect 5836 50968 5876 51008
rect 6412 50968 6452 51008
rect 6892 50982 6932 51022
rect 7564 50968 7604 51008
rect 7660 50968 7700 51008
rect 8140 50968 8180 51008
rect 8620 50968 8660 51008
rect 9100 50973 9140 51013
rect 10444 50968 10484 51008
rect 10540 50968 10580 51008
rect 10924 50968 10964 51008
rect 11020 50968 11060 51008
rect 11500 50968 11540 51008
rect 11980 50982 12020 51022
rect 13228 50968 13268 51008
rect 13324 50968 13364 51008
rect 13708 50968 13748 51008
rect 14812 51010 14852 51050
rect 13804 50968 13844 51008
rect 14284 50968 14324 51008
rect 16204 50968 16244 51008
rect 17452 50968 17492 51008
rect 17932 50968 17972 51008
rect 19180 50968 19220 51008
rect 9292 50884 9332 50924
rect 12172 50884 12212 50924
rect 2668 50800 2708 50840
rect 4780 50800 4820 50840
rect 7084 50800 7124 50840
rect 14956 50800 14996 50840
rect 19372 50800 19412 50840
rect 19564 50800 19604 50840
rect 20140 50800 20180 50840
rect 4928 50632 4968 50672
rect 5010 50632 5050 50672
rect 5092 50632 5132 50672
rect 5174 50632 5214 50672
rect 5256 50632 5296 50672
rect 20048 50632 20088 50672
rect 20130 50632 20170 50672
rect 20212 50632 20252 50672
rect 20294 50632 20334 50672
rect 20376 50632 20416 50672
rect 9004 50464 9044 50504
rect 19276 50464 19316 50504
rect 4684 50380 4724 50420
rect 1420 50296 1460 50336
rect 2668 50296 2708 50336
rect 3052 50296 3092 50336
rect 4300 50296 4340 50336
rect 4876 50282 4916 50322
rect 5356 50296 5396 50336
rect 6316 50296 6356 50336
rect 6412 50296 6452 50336
rect 7564 50296 7604 50336
rect 8812 50296 8852 50336
rect 9196 50296 9236 50336
rect 10444 50296 10484 50336
rect 11596 50296 11636 50336
rect 12844 50296 12884 50336
rect 13996 50296 14036 50336
rect 15244 50296 15284 50336
rect 17164 50296 17204 50336
rect 17548 50296 17588 50336
rect 17644 50296 17684 50336
rect 18124 50296 18164 50336
rect 18604 50296 18644 50336
rect 19132 50286 19172 50326
rect 5836 50212 5876 50252
rect 5932 50212 5972 50252
rect 13420 50212 13460 50252
rect 16012 50212 16052 50252
rect 18028 50212 18068 50252
rect 19468 50212 19508 50252
rect 19852 50212 19892 50252
rect 13228 50128 13268 50168
rect 20044 50128 20084 50168
rect 2860 50044 2900 50084
rect 4492 50044 4532 50084
rect 10636 50044 10676 50084
rect 13036 50044 13076 50084
rect 15436 50044 15476 50084
rect 15820 50044 15860 50084
rect 16492 50044 16532 50084
rect 19660 50044 19700 50084
rect 3688 49876 3728 49916
rect 3770 49876 3810 49916
rect 3852 49876 3892 49916
rect 3934 49876 3974 49916
rect 4016 49876 4056 49916
rect 18808 49876 18848 49916
rect 18890 49876 18930 49916
rect 18972 49876 19012 49916
rect 19054 49876 19094 49916
rect 19136 49876 19176 49916
rect 1900 49708 1940 49748
rect 7276 49708 7316 49748
rect 17260 49708 17300 49748
rect 18988 49708 19028 49748
rect 11308 49624 11348 49664
rect 1708 49540 1748 49580
rect 2092 49540 2132 49580
rect 3436 49540 3476 49580
rect 3532 49540 3572 49580
rect 12076 49540 12116 49580
rect 12172 49540 12212 49580
rect 15916 49540 15956 49580
rect 19180 49540 19220 49580
rect 19372 49540 19412 49580
rect 19756 49540 19796 49580
rect 2476 49470 2516 49510
rect 2956 49456 2996 49496
rect 3916 49456 3956 49496
rect 4012 49456 4052 49496
rect 5836 49456 5876 49496
rect 7084 49456 7124 49496
rect 7468 49456 7508 49496
rect 8716 49456 8756 49496
rect 9868 49456 9908 49496
rect 11116 49456 11156 49496
rect 11596 49456 11636 49496
rect 11692 49456 11732 49496
rect 12652 49456 12692 49496
rect 13132 49470 13172 49510
rect 13516 49456 13556 49496
rect 14764 49456 14804 49496
rect 15340 49456 15380 49496
rect 15436 49436 15476 49476
rect 15820 49456 15860 49496
rect 16396 49456 16436 49496
rect 16924 49465 16964 49505
rect 17452 49456 17492 49496
rect 18700 49456 18740 49496
rect 2284 49372 2324 49412
rect 13324 49372 13364 49412
rect 17068 49372 17108 49412
rect 1516 49288 1556 49328
rect 8908 49288 8948 49328
rect 14956 49288 14996 49328
rect 19564 49288 19604 49328
rect 19948 49288 19988 49328
rect 4928 49120 4968 49160
rect 5010 49120 5050 49160
rect 5092 49120 5132 49160
rect 5174 49120 5214 49160
rect 5256 49120 5296 49160
rect 20048 49120 20088 49160
rect 20130 49120 20170 49160
rect 20212 49120 20252 49160
rect 20294 49120 20334 49160
rect 20376 49120 20416 49160
rect 2860 48952 2900 48992
rect 14956 48952 14996 48992
rect 17068 48952 17108 48992
rect 19756 48952 19796 48992
rect 10540 48868 10580 48908
rect 12940 48868 12980 48908
rect 1228 48784 1268 48824
rect 2476 48784 2516 48824
rect 3436 48784 3476 48824
rect 4684 48784 4724 48824
rect 5068 48784 5108 48824
rect 6316 48784 6356 48824
rect 6796 48784 6836 48824
rect 8044 48784 8084 48824
rect 8812 48784 8852 48824
rect 8908 48784 8948 48824
rect 9292 48784 9332 48824
rect 9388 48784 9428 48824
rect 9868 48784 9908 48824
rect 10396 48774 10436 48814
rect 11500 48784 11540 48824
rect 12748 48784 12788 48824
rect 13228 48784 13268 48824
rect 13324 48784 13364 48824
rect 14284 48784 14324 48824
rect 14812 48774 14852 48814
rect 15628 48784 15668 48824
rect 16876 48784 16916 48824
rect 18028 48784 18068 48824
rect 18124 48784 18164 48824
rect 18604 48784 18644 48824
rect 19084 48784 19124 48824
rect 3052 48700 3092 48740
rect 13708 48700 13748 48740
rect 13804 48700 13844 48740
rect 18508 48700 18548 48740
rect 19612 48742 19652 48782
rect 19948 48700 19988 48740
rect 2668 48532 2708 48572
rect 4876 48532 4916 48572
rect 6508 48532 6548 48572
rect 8236 48532 8276 48572
rect 20140 48532 20180 48572
rect 3688 48364 3728 48404
rect 3770 48364 3810 48404
rect 3852 48364 3892 48404
rect 3934 48364 3974 48404
rect 4016 48364 4056 48404
rect 18808 48364 18848 48404
rect 18890 48364 18930 48404
rect 18972 48364 19012 48404
rect 19054 48364 19094 48404
rect 19136 48364 19176 48404
rect 1612 48196 1652 48236
rect 16204 48196 16244 48236
rect 18028 48196 18068 48236
rect 19660 48196 19700 48236
rect 1804 48028 1844 48068
rect 6412 48028 6452 48068
rect 6508 48028 6548 48068
rect 8908 48028 8948 48068
rect 9004 48028 9044 48068
rect 16396 48028 16436 48068
rect 19852 48028 19892 48068
rect 1996 47944 2036 47984
rect 3244 47944 3284 47984
rect 3628 47944 3668 47984
rect 4876 47944 4916 47984
rect 5452 47949 5492 47989
rect 5932 47944 5972 47984
rect 6892 47944 6932 47984
rect 6988 47944 7028 47984
rect 7948 47949 7988 47989
rect 8428 47944 8468 47984
rect 9388 47944 9428 47984
rect 9484 47944 9524 47984
rect 10252 47944 10292 47984
rect 11500 47944 11540 47984
rect 13612 47944 13652 47984
rect 14860 47944 14900 47984
rect 16588 47944 16628 47984
rect 17836 47944 17876 47984
rect 18220 47944 18260 47984
rect 19468 47944 19508 47984
rect 5068 47860 5108 47900
rect 5260 47860 5300 47900
rect 7756 47860 7796 47900
rect 3436 47776 3476 47816
rect 11692 47776 11732 47816
rect 15052 47776 15092 47816
rect 20044 47776 20084 47816
rect 4928 47608 4968 47648
rect 5010 47608 5050 47648
rect 5092 47608 5132 47648
rect 5174 47608 5214 47648
rect 5256 47608 5296 47648
rect 20048 47608 20088 47648
rect 20130 47608 20170 47648
rect 20212 47608 20252 47648
rect 20294 47608 20334 47648
rect 20376 47608 20416 47648
rect 1804 47440 1844 47480
rect 6700 47440 6740 47480
rect 8044 47440 8084 47480
rect 10636 47440 10676 47480
rect 16780 47440 16820 47480
rect 4012 47356 4052 47396
rect 2284 47272 2324 47312
rect 2380 47272 2420 47312
rect 2860 47272 2900 47312
rect 3340 47272 3380 47312
rect 3820 47267 3860 47307
rect 4972 47272 5012 47312
rect 5068 47272 5108 47312
rect 5452 47272 5492 47312
rect 5548 47272 5588 47312
rect 6028 47272 6068 47312
rect 6556 47262 6596 47302
rect 8236 47272 8276 47312
rect 9484 47272 9524 47312
rect 11116 47272 11156 47312
rect 12364 47272 12404 47312
rect 12748 47272 12788 47312
rect 13996 47272 14036 47312
rect 15052 47272 15092 47312
rect 15148 47272 15188 47312
rect 15532 47272 15572 47312
rect 15628 47272 15668 47312
rect 16108 47272 16148 47312
rect 16972 47272 17012 47312
rect 18220 47272 18260 47312
rect 18604 47272 18644 47312
rect 19852 47272 19892 47312
rect 1996 47188 2036 47228
rect 16636 47230 16676 47270
rect 2764 47188 2804 47228
rect 10828 47188 10868 47228
rect 12556 47020 12596 47060
rect 14188 47020 14228 47060
rect 18412 47020 18452 47060
rect 20044 47020 20084 47060
rect 3688 46852 3728 46892
rect 3770 46852 3810 46892
rect 3852 46852 3892 46892
rect 3934 46852 3974 46892
rect 4016 46852 4056 46892
rect 18808 46852 18848 46892
rect 18890 46852 18930 46892
rect 18972 46852 19012 46892
rect 19054 46852 19094 46892
rect 19136 46852 19176 46892
rect 16684 46684 16724 46724
rect 5932 46600 5972 46640
rect 11884 46516 11924 46556
rect 13132 46516 13172 46556
rect 1228 46432 1268 46472
rect 2476 46432 2516 46472
rect 4492 46432 4532 46472
rect 5740 46432 5780 46472
rect 6124 46432 6164 46472
rect 7372 46432 7412 46472
rect 8140 46432 8180 46472
rect 9388 46432 9428 46472
rect 9868 46432 9908 46472
rect 9964 46432 10004 46472
rect 10348 46432 10388 46472
rect 10444 46432 10484 46472
rect 10924 46432 10964 46472
rect 11452 46441 11492 46481
rect 12556 46432 12596 46472
rect 12652 46432 12692 46472
rect 14140 46474 14180 46514
rect 18412 46516 18452 46556
rect 19852 46516 19892 46556
rect 13036 46432 13076 46472
rect 13612 46432 13652 46472
rect 15244 46432 15284 46472
rect 16492 46432 16532 46472
rect 17932 46432 17972 46472
rect 18028 46432 18068 46472
rect 19516 46474 19556 46514
rect 18508 46432 18548 46472
rect 18988 46432 19028 46472
rect 2668 46264 2708 46304
rect 7564 46264 7604 46304
rect 9580 46264 9620 46304
rect 11596 46264 11636 46304
rect 12076 46264 12116 46304
rect 14284 46264 14324 46304
rect 19660 46264 19700 46304
rect 20044 46264 20084 46304
rect 4928 46096 4968 46136
rect 5010 46096 5050 46136
rect 5092 46096 5132 46136
rect 5174 46096 5214 46136
rect 5256 46096 5296 46136
rect 20048 46096 20088 46136
rect 20130 46096 20170 46136
rect 20212 46096 20252 46136
rect 20294 46096 20334 46136
rect 20376 46096 20416 46136
rect 1516 45928 1556 45968
rect 1900 45928 1940 45968
rect 11212 45928 11252 45968
rect 12940 45928 12980 45968
rect 19180 45928 19220 45968
rect 14860 45844 14900 45884
rect 16876 45844 16916 45884
rect 2668 45760 2708 45800
rect 3916 45760 3956 45800
rect 4108 45760 4148 45800
rect 5356 45760 5396 45800
rect 6316 45760 6356 45800
rect 7564 45760 7604 45800
rect 9484 45760 9524 45800
rect 9580 45760 9620 45800
rect 10060 45760 10100 45800
rect 10540 45760 10580 45800
rect 11020 45746 11060 45786
rect 13420 45760 13460 45800
rect 14668 45760 14708 45800
rect 15148 45760 15188 45800
rect 15244 45760 15284 45800
rect 15724 45760 15764 45800
rect 16204 45760 16244 45800
rect 16684 45746 16724 45786
rect 17068 45760 17108 45800
rect 18316 45760 18356 45800
rect 1708 45676 1748 45716
rect 2092 45676 2132 45716
rect 9964 45676 10004 45716
rect 11596 45676 11636 45716
rect 13132 45676 13172 45716
rect 15628 45676 15668 45716
rect 18988 45676 19028 45716
rect 19372 45676 19412 45716
rect 19564 45676 19604 45716
rect 2476 45508 2516 45548
rect 5548 45508 5588 45548
rect 7756 45508 7796 45548
rect 11404 45508 11444 45548
rect 18508 45508 18548 45548
rect 18796 45508 18836 45548
rect 19756 45508 19796 45548
rect 3688 45340 3728 45380
rect 3770 45340 3810 45380
rect 3852 45340 3892 45380
rect 3934 45340 3974 45380
rect 4016 45340 4056 45380
rect 18808 45340 18848 45380
rect 18890 45340 18930 45380
rect 18972 45340 19012 45380
rect 19054 45340 19094 45380
rect 19136 45340 19176 45380
rect 1516 45172 1556 45212
rect 9388 45172 9428 45212
rect 11020 45172 11060 45212
rect 13708 45172 13748 45212
rect 16684 45172 16724 45212
rect 16876 45172 16916 45212
rect 1708 45004 1748 45044
rect 2092 45004 2132 45044
rect 2524 44962 2564 45002
rect 6124 45004 6164 45044
rect 13900 45004 13940 45044
rect 17068 45004 17108 45044
rect 18412 45004 18452 45044
rect 18508 45004 18548 45044
rect 19852 45004 19892 45044
rect 3052 44920 3092 44960
rect 3532 44920 3572 44960
rect 3628 44920 3668 44960
rect 4012 44920 4052 44960
rect 4108 44920 4148 44960
rect 5644 44920 5684 44960
rect 5740 44920 5780 44960
rect 6220 44920 6260 44960
rect 6700 44920 6740 44960
rect 7180 44934 7220 44974
rect 7948 44920 7988 44960
rect 9196 44920 9236 44960
rect 9580 44920 9620 44960
rect 10828 44920 10868 44960
rect 12076 44920 12116 44960
rect 13324 44920 13364 44960
rect 15244 44920 15284 44960
rect 16492 44920 16532 44960
rect 17932 44920 17972 44960
rect 18028 44920 18068 44960
rect 18988 44920 19028 44960
rect 19516 44929 19556 44969
rect 2380 44836 2420 44876
rect 7372 44836 7412 44876
rect 19660 44836 19700 44876
rect 1900 44752 1940 44792
rect 13516 44752 13556 44792
rect 20044 44752 20084 44792
rect 4928 44584 4968 44624
rect 5010 44584 5050 44624
rect 5092 44584 5132 44624
rect 5174 44584 5214 44624
rect 5256 44584 5296 44624
rect 20048 44584 20088 44624
rect 20130 44584 20170 44624
rect 20212 44584 20252 44624
rect 20294 44584 20334 44624
rect 20376 44584 20416 44624
rect 1804 44416 1844 44456
rect 7276 44416 7316 44456
rect 9676 44416 9716 44456
rect 13516 44416 13556 44456
rect 15436 44416 15476 44456
rect 19564 44416 19604 44456
rect 17452 44332 17492 44372
rect 2380 44248 2420 44288
rect 3628 44248 3668 44288
rect 3820 44248 3860 44288
rect 5068 44248 5108 44288
rect 5548 44248 5588 44288
rect 5644 44248 5684 44288
rect 6028 44248 6068 44288
rect 6124 44248 6164 44288
rect 6604 44248 6644 44288
rect 7084 44243 7124 44283
rect 10060 44248 10100 44288
rect 11308 44248 11348 44288
rect 11788 44248 11828 44288
rect 11884 44248 11924 44288
rect 13996 44290 14036 44330
rect 12364 44248 12404 44288
rect 12844 44248 12884 44288
rect 13324 44234 13364 44274
rect 15244 44248 15284 44288
rect 15724 44248 15764 44288
rect 15820 44248 15860 44288
rect 16204 44248 16244 44288
rect 16300 44248 16340 44288
rect 16780 44248 16820 44288
rect 17260 44234 17300 44274
rect 18124 44248 18164 44288
rect 19372 44248 19412 44288
rect 1996 44164 2036 44204
rect 9196 44164 9236 44204
rect 9868 44164 9908 44204
rect 12268 44164 12308 44204
rect 19756 44164 19796 44204
rect 5260 44080 5300 44120
rect 2188 43996 2228 44036
rect 9004 43996 9044 44036
rect 11500 43996 11540 44036
rect 19948 43996 19988 44036
rect 3688 43828 3728 43868
rect 3770 43828 3810 43868
rect 3852 43828 3892 43868
rect 3934 43828 3974 43868
rect 4016 43828 4056 43868
rect 18808 43828 18848 43868
rect 18890 43828 18930 43868
rect 18972 43828 19012 43868
rect 19054 43828 19094 43868
rect 19136 43828 19176 43868
rect 11404 43660 11444 43700
rect 15052 43660 15092 43700
rect 17260 43660 17300 43700
rect 17452 43660 17492 43700
rect 19180 43660 19220 43700
rect 3628 43492 3668 43532
rect 8524 43492 8564 43532
rect 12268 43492 12308 43532
rect 14092 43492 14132 43532
rect 14860 43492 14900 43532
rect 17644 43492 17684 43532
rect 17836 43492 17876 43532
rect 18988 43492 19028 43532
rect 19372 43492 19412 43532
rect 2668 43422 2708 43462
rect 3148 43408 3188 43448
rect 3724 43408 3764 43448
rect 4108 43408 4148 43448
rect 4204 43408 4244 43448
rect 6220 43408 6260 43448
rect 7468 43408 7508 43448
rect 7948 43408 7988 43448
rect 8044 43408 8084 43448
rect 8428 43408 8468 43448
rect 9004 43408 9044 43448
rect 9532 43417 9572 43457
rect 9964 43408 10004 43448
rect 11212 43408 11252 43448
rect 11692 43408 11732 43448
rect 11788 43408 11828 43448
rect 12172 43408 12212 43448
rect 12748 43408 12788 43448
rect 13276 43417 13316 43457
rect 15820 43408 15860 43448
rect 17068 43408 17108 43448
rect 2476 43324 2516 43364
rect 7660 43324 7700 43364
rect 9676 43324 9716 43364
rect 13420 43240 13460 43280
rect 13900 43240 13940 43280
rect 18028 43240 18068 43280
rect 19564 43240 19604 43280
rect 4928 43072 4968 43112
rect 5010 43072 5050 43112
rect 5092 43072 5132 43112
rect 5174 43072 5214 43112
rect 5256 43072 5296 43112
rect 20048 43072 20088 43112
rect 20130 43072 20170 43112
rect 20212 43072 20252 43112
rect 20294 43072 20334 43112
rect 20376 43072 20416 43112
rect 9580 42904 9620 42944
rect 2668 42820 2708 42860
rect 4684 42820 4724 42860
rect 6700 42820 6740 42860
rect 13804 42820 13844 42860
rect 1228 42736 1268 42776
rect 2476 42736 2516 42776
rect 3244 42736 3284 42776
rect 4492 42736 4532 42776
rect 4972 42736 5012 42776
rect 5068 42736 5108 42776
rect 6028 42736 6068 42776
rect 8140 42736 8180 42776
rect 9388 42736 9428 42776
rect 12364 42736 12404 42776
rect 13612 42736 13652 42776
rect 5452 42652 5492 42692
rect 5548 42652 5588 42692
rect 6556 42694 6596 42734
rect 18604 42652 18644 42692
rect 18988 42652 19028 42692
rect 19372 42652 19412 42692
rect 19756 42652 19796 42692
rect 19180 42568 19220 42608
rect 19564 42568 19604 42608
rect 18796 42484 18836 42524
rect 19948 42484 19988 42524
rect 3688 42316 3728 42356
rect 3770 42316 3810 42356
rect 3852 42316 3892 42356
rect 3934 42316 3974 42356
rect 4016 42316 4056 42356
rect 18808 42316 18848 42356
rect 18890 42316 18930 42356
rect 18972 42316 19012 42356
rect 19054 42316 19094 42356
rect 19136 42316 19176 42356
rect 1900 42148 1940 42188
rect 6700 42148 6740 42188
rect 17164 42148 17204 42188
rect 19276 42148 19316 42188
rect 20044 42148 20084 42188
rect 4876 42064 4916 42104
rect 18892 42064 18932 42104
rect 2092 41980 2132 42020
rect 3436 41980 3476 42020
rect 16972 41980 17012 42020
rect 18316 41980 18356 42020
rect 18700 41980 18740 42020
rect 19084 41980 19124 42020
rect 19468 41980 19508 42020
rect 19852 41980 19892 42020
rect 2476 41901 2516 41941
rect 2956 41896 2996 41936
rect 3532 41896 3572 41936
rect 3916 41896 3956 41936
rect 4012 41896 4052 41936
rect 5260 41896 5300 41936
rect 6508 41896 6548 41936
rect 7564 41896 7604 41936
rect 8812 41896 8852 41936
rect 9196 41896 9236 41936
rect 10444 41896 10484 41936
rect 10828 41896 10868 41936
rect 12076 41896 12116 41936
rect 2284 41812 2324 41852
rect 9004 41728 9044 41768
rect 10636 41728 10676 41768
rect 12268 41728 12308 41768
rect 18508 41728 18548 41768
rect 19660 41728 19700 41768
rect 4928 41560 4968 41600
rect 5010 41560 5050 41600
rect 5092 41560 5132 41600
rect 5174 41560 5214 41600
rect 5256 41560 5296 41600
rect 20048 41560 20088 41600
rect 20130 41560 20170 41600
rect 20212 41560 20252 41600
rect 20294 41560 20334 41600
rect 20376 41560 20416 41600
rect 3340 41392 3380 41432
rect 9292 41392 9332 41432
rect 12940 41392 12980 41432
rect 19084 41392 19124 41432
rect 5068 41308 5108 41348
rect 7084 41308 7124 41348
rect 9100 41308 9140 41348
rect 12172 41308 12212 41348
rect 1900 41224 1940 41264
rect 3148 41224 3188 41264
rect 3628 41224 3668 41264
rect 4876 41224 4916 41264
rect 5356 41224 5396 41264
rect 5452 41224 5492 41264
rect 6412 41224 6452 41264
rect 6940 41214 6980 41254
rect 7660 41224 7700 41264
rect 8908 41224 8948 41264
rect 10444 41224 10484 41264
rect 10540 41224 10580 41264
rect 11020 41224 11060 41264
rect 11500 41224 11540 41264
rect 12028 41214 12068 41254
rect 5836 41140 5876 41180
rect 5932 41140 5972 41180
rect 10924 41140 10964 41180
rect 12748 41140 12788 41180
rect 18892 41140 18932 41180
rect 19276 41140 19316 41180
rect 19660 41140 19700 41180
rect 19468 40972 19508 41012
rect 19852 40972 19892 41012
rect 3688 40804 3728 40844
rect 3770 40804 3810 40844
rect 3852 40804 3892 40844
rect 3934 40804 3974 40844
rect 4016 40804 4056 40844
rect 18808 40804 18848 40844
rect 18890 40804 18930 40844
rect 18972 40804 19012 40844
rect 19054 40804 19094 40844
rect 19136 40804 19176 40844
rect 2668 40636 2708 40676
rect 7372 40636 7412 40676
rect 13228 40636 13268 40676
rect 19084 40636 19124 40676
rect 19468 40636 19508 40676
rect 9964 40468 10004 40508
rect 2476 40426 2516 40466
rect 13036 40468 13076 40508
rect 18892 40468 18932 40508
rect 19276 40468 19316 40508
rect 19660 40468 19700 40508
rect 20044 40468 20084 40508
rect 1228 40384 1268 40424
rect 3916 40384 3956 40424
rect 5164 40384 5204 40424
rect 5932 40384 5972 40424
rect 7180 40384 7220 40424
rect 7756 40384 7796 40424
rect 9004 40384 9044 40424
rect 9388 40384 9428 40424
rect 9484 40384 9524 40424
rect 9868 40384 9908 40424
rect 10444 40384 10484 40424
rect 10924 40398 10964 40438
rect 7564 40300 7604 40340
rect 5356 40216 5396 40256
rect 11116 40216 11156 40256
rect 19852 40216 19892 40256
rect 20236 40216 20276 40256
rect 4928 40048 4968 40088
rect 5010 40048 5050 40088
rect 5092 40048 5132 40088
rect 5174 40048 5214 40088
rect 5256 40048 5296 40088
rect 20048 40048 20088 40088
rect 20130 40048 20170 40088
rect 20212 40048 20252 40088
rect 20294 40048 20334 40088
rect 20376 40048 20416 40088
rect 3724 39880 3764 39920
rect 5740 39880 5780 39920
rect 9388 39880 9428 39920
rect 19564 39880 19604 39920
rect 19948 39880 19988 39920
rect 1996 39712 2036 39752
rect 2092 39712 2132 39752
rect 3052 39712 3092 39752
rect 3532 39707 3572 39747
rect 4012 39712 4052 39752
rect 4108 39712 4148 39752
rect 5068 39712 5108 39752
rect 5548 39707 5588 39747
rect 5932 39712 5972 39752
rect 6124 39712 6164 39752
rect 6220 39712 6260 39752
rect 6412 39712 6452 39752
rect 6508 39712 6548 39752
rect 6700 39712 6740 39752
rect 6796 39712 6836 39752
rect 6897 39712 6937 39752
rect 7660 39712 7700 39752
rect 8908 39712 8948 39752
rect 10636 39712 10676 39752
rect 11884 39712 11924 39752
rect 12652 39712 12692 39752
rect 12844 39712 12884 39752
rect 12940 39712 12980 39752
rect 2476 39628 2516 39668
rect 2572 39628 2612 39668
rect 4492 39628 4532 39668
rect 4588 39628 4628 39668
rect 18988 39628 19028 39668
rect 19372 39628 19412 39668
rect 19756 39628 19796 39668
rect 6220 39544 6260 39584
rect 9292 39544 9332 39584
rect 12844 39544 12884 39584
rect 6412 39460 6452 39500
rect 9100 39460 9140 39500
rect 10444 39460 10484 39500
rect 19180 39460 19220 39500
rect 3688 39292 3728 39332
rect 3770 39292 3810 39332
rect 3852 39292 3892 39332
rect 3934 39292 3974 39332
rect 4016 39292 4056 39332
rect 18808 39292 18848 39332
rect 18890 39292 18930 39332
rect 18972 39292 19012 39332
rect 19054 39292 19094 39332
rect 19136 39292 19176 39332
rect 3436 39124 3476 39164
rect 6700 39124 6740 39164
rect 12940 39124 12980 39164
rect 9196 38956 9236 38996
rect 14476 38956 14516 38996
rect 19372 38956 19412 38996
rect 1996 38872 2036 38912
rect 3244 38872 3284 38912
rect 3628 38872 3668 38912
rect 4876 38872 4916 38912
rect 5260 38872 5300 38912
rect 6508 38872 6548 38912
rect 6892 38872 6932 38912
rect 8140 38872 8180 38912
rect 8620 38872 8660 38912
rect 8716 38872 8756 38912
rect 9100 38872 9140 38912
rect 9676 38872 9716 38912
rect 10156 38886 10196 38926
rect 12748 38914 12788 38954
rect 11500 38872 11540 38912
rect 13132 38872 13172 38912
rect 13420 38872 13460 38912
rect 8332 38788 8372 38828
rect 5068 38704 5108 38744
rect 10348 38704 10388 38744
rect 13324 38704 13364 38744
rect 14668 38704 14708 38744
rect 19564 38704 19604 38744
rect 4928 38536 4968 38576
rect 5010 38536 5050 38576
rect 5092 38536 5132 38576
rect 5174 38536 5214 38576
rect 5256 38536 5296 38576
rect 20048 38536 20088 38576
rect 20130 38536 20170 38576
rect 20212 38536 20252 38576
rect 20294 38536 20334 38576
rect 20376 38536 20416 38576
rect 3052 38368 3092 38408
rect 7180 38368 7220 38408
rect 7468 38368 7508 38408
rect 8044 38368 8084 38408
rect 12940 38368 12980 38408
rect 14572 38368 14612 38408
rect 5164 38284 5204 38324
rect 10252 38284 10292 38324
rect 13804 38284 13844 38324
rect 1612 38200 1652 38240
rect 2860 38200 2900 38240
rect 3724 38200 3764 38240
rect 4972 38200 5012 38240
rect 5452 38200 5492 38240
rect 5548 38200 5588 38240
rect 6508 38200 6548 38240
rect 6988 38195 7028 38235
rect 7660 38200 7700 38240
rect 7756 38200 7796 38240
rect 7948 38200 7988 38240
rect 8524 38200 8564 38240
rect 8620 38200 8660 38240
rect 9004 38200 9044 38240
rect 9100 38200 9140 38240
rect 9580 38200 9620 38240
rect 10060 38186 10100 38226
rect 11500 38200 11540 38240
rect 12748 38200 12788 38240
rect 13132 38200 13172 38240
rect 13324 38200 13364 38240
rect 13420 38200 13460 38240
rect 13612 38200 13652 38240
rect 13708 38200 13748 38240
rect 13900 38200 13940 38240
rect 14092 38200 14132 38240
rect 14188 38200 14228 38240
rect 5932 38116 5972 38156
rect 6028 38116 6068 38156
rect 14380 38116 14420 38156
rect 15340 38105 15380 38145
rect 18604 38116 18644 38156
rect 19372 38116 19412 38156
rect 13420 38032 13460 38072
rect 15532 38032 15572 38072
rect 19564 38032 19604 38072
rect 12940 37948 12980 37988
rect 18796 37948 18836 37988
rect 3688 37780 3728 37820
rect 3770 37780 3810 37820
rect 3852 37780 3892 37820
rect 3934 37780 3974 37820
rect 4016 37780 4056 37820
rect 18808 37780 18848 37820
rect 18890 37780 18930 37820
rect 18972 37780 19012 37820
rect 19054 37780 19094 37820
rect 19136 37780 19176 37820
rect 15052 37612 15092 37652
rect 19948 37612 19988 37652
rect 10444 37528 10484 37568
rect 11884 37528 11924 37568
rect 12556 37528 12596 37568
rect 19564 37528 19604 37568
rect 18988 37444 19028 37484
rect 19372 37444 19412 37484
rect 19756 37444 19796 37484
rect 2380 37360 2420 37400
rect 2476 37360 2516 37400
rect 2860 37360 2900 37400
rect 2956 37360 2996 37400
rect 3436 37360 3476 37400
rect 3964 37369 4004 37409
rect 4300 37360 4340 37400
rect 5548 37360 5588 37400
rect 6028 37360 6068 37400
rect 6124 37360 6164 37400
rect 6508 37360 6548 37400
rect 6604 37360 6644 37400
rect 7084 37360 7124 37400
rect 7564 37365 7604 37405
rect 9004 37360 9044 37400
rect 10252 37360 10292 37400
rect 11116 37360 11156 37400
rect 11308 37360 11348 37400
rect 11404 37360 11444 37400
rect 11596 37360 11636 37400
rect 11788 37360 11828 37400
rect 11884 37360 11924 37400
rect 12076 37360 12116 37400
rect 12268 37360 12308 37400
rect 12364 37360 12404 37400
rect 12556 37360 12596 37400
rect 12844 37360 12884 37400
rect 13036 37360 13076 37400
rect 13132 37360 13172 37400
rect 13324 37360 13364 37400
rect 13612 37360 13652 37400
rect 14860 37360 14900 37400
rect 5740 37276 5780 37316
rect 12172 37276 12212 37316
rect 4108 37192 4148 37232
rect 7756 37192 7796 37232
rect 11212 37192 11252 37232
rect 13324 37192 13364 37232
rect 19180 37192 19220 37232
rect 4928 37024 4968 37064
rect 5010 37024 5050 37064
rect 5092 37024 5132 37064
rect 5174 37024 5214 37064
rect 5256 37024 5296 37064
rect 20048 37024 20088 37064
rect 20130 37024 20170 37064
rect 20212 37024 20252 37064
rect 20294 37024 20334 37064
rect 20376 37024 20416 37064
rect 2668 36856 2708 36896
rect 4300 36856 4340 36896
rect 8908 36856 8948 36896
rect 10828 36856 10868 36896
rect 12364 36856 12404 36896
rect 13036 36856 13076 36896
rect 13804 36856 13844 36896
rect 19564 36856 19604 36896
rect 1228 36688 1268 36728
rect 2476 36688 2516 36728
rect 2860 36688 2900 36728
rect 4108 36688 4148 36728
rect 4492 36688 4532 36728
rect 4684 36688 4724 36728
rect 4780 36688 4820 36728
rect 4972 36688 5012 36728
rect 5164 36688 5204 36728
rect 5836 36688 5876 36728
rect 7084 36688 7124 36728
rect 7468 36688 7508 36728
rect 8716 36688 8756 36728
rect 10252 36688 10292 36728
rect 10348 36688 10388 36728
rect 10540 36688 10580 36728
rect 10732 36688 10772 36728
rect 10924 36688 10964 36728
rect 11020 36688 11060 36728
rect 11308 36703 11348 36743
rect 11596 36688 11636 36728
rect 11692 36688 11732 36728
rect 12172 36688 12212 36728
rect 12268 36688 12308 36728
rect 12460 36688 12500 36728
rect 12556 36688 12596 36728
rect 12657 36688 12697 36728
rect 12940 36688 12980 36728
rect 13228 36688 13268 36728
rect 13612 36688 13652 36728
rect 13900 36688 13940 36728
rect 13996 36688 14036 36728
rect 14092 36688 14132 36728
rect 14284 36688 14324 36728
rect 13324 36604 13364 36644
rect 13516 36604 13556 36644
rect 18988 36604 19028 36644
rect 19372 36604 19412 36644
rect 5068 36520 5108 36560
rect 7276 36520 7316 36560
rect 10540 36520 10580 36560
rect 11980 36520 12020 36560
rect 13420 36520 13460 36560
rect 14380 36520 14420 36560
rect 4492 36436 4532 36476
rect 19180 36436 19220 36476
rect 3688 36268 3728 36308
rect 3770 36268 3810 36308
rect 3852 36268 3892 36308
rect 3934 36268 3974 36308
rect 4016 36268 4056 36308
rect 18808 36268 18848 36308
rect 18890 36268 18930 36308
rect 18972 36268 19012 36308
rect 19054 36268 19094 36308
rect 19136 36268 19176 36308
rect 2668 36100 2708 36140
rect 4300 36100 4340 36140
rect 11020 36100 11060 36140
rect 12268 36100 12308 36140
rect 19564 36100 19604 36140
rect 13324 36016 13364 36056
rect 19180 36016 19220 36056
rect 10444 35932 10484 35972
rect 18988 35932 19028 35972
rect 19372 35932 19412 35972
rect 19756 35932 19796 35972
rect 1228 35848 1268 35888
rect 2476 35848 2516 35888
rect 2860 35848 2900 35888
rect 4108 35848 4148 35888
rect 4492 35848 4532 35888
rect 4588 35848 4628 35888
rect 4972 35848 5012 35888
rect 6220 35848 6260 35888
rect 6604 35848 6644 35888
rect 7852 35848 7892 35888
rect 8332 35848 8372 35888
rect 8428 35848 8468 35888
rect 8812 35848 8852 35888
rect 8908 35848 8948 35888
rect 9388 35848 9428 35888
rect 9916 35857 9956 35897
rect 10252 35848 10292 35888
rect 10540 35848 10580 35888
rect 10732 35848 10772 35888
rect 11020 35848 11060 35888
rect 11308 35848 11348 35888
rect 11596 35848 11636 35888
rect 11788 35848 11828 35888
rect 11884 35848 11924 35888
rect 12076 35848 12116 35888
rect 12268 35848 12308 35888
rect 12556 35848 12596 35888
rect 12748 35848 12788 35888
rect 12844 35848 12884 35888
rect 13228 35848 13268 35888
rect 13324 35848 13364 35888
rect 13516 35848 13556 35888
rect 13708 35848 13748 35888
rect 13804 35848 13844 35888
rect 13900 35848 13940 35888
rect 13996 35848 14036 35888
rect 14188 35848 14228 35888
rect 14284 35848 14324 35888
rect 14380 35848 14420 35888
rect 8044 35764 8084 35804
rect 4300 35680 4340 35720
rect 4780 35680 4820 35720
rect 6412 35680 6452 35720
rect 10060 35680 10100 35720
rect 11500 35680 11540 35720
rect 12076 35680 12116 35720
rect 13036 35680 13076 35720
rect 14476 35680 14516 35720
rect 19948 35680 19988 35720
rect 4928 35512 4968 35552
rect 5010 35512 5050 35552
rect 5092 35512 5132 35552
rect 5174 35512 5214 35552
rect 5256 35512 5296 35552
rect 20048 35512 20088 35552
rect 20130 35512 20170 35552
rect 20212 35512 20252 35552
rect 20294 35512 20334 35552
rect 20376 35512 20416 35552
rect 9964 35344 10004 35384
rect 13228 35344 13268 35384
rect 13708 35344 13748 35384
rect 2860 35260 2900 35300
rect 6604 35260 6644 35300
rect 10540 35260 10580 35300
rect 1420 35176 1460 35216
rect 2668 35176 2708 35216
rect 3052 35176 3092 35216
rect 3244 35176 3284 35216
rect 3724 35176 3764 35216
rect 3820 35176 3860 35216
rect 4108 35176 4148 35216
rect 4492 35176 4532 35216
rect 5740 35176 5780 35216
rect 6412 35176 6452 35216
rect 6508 35176 6548 35216
rect 6892 35218 6932 35258
rect 12556 35260 12596 35300
rect 6700 35176 6740 35216
rect 8140 35176 8180 35216
rect 8524 35176 8564 35216
rect 9772 35176 9812 35216
rect 10444 35176 10484 35216
rect 10636 35176 10676 35216
rect 10828 35176 10868 35216
rect 11116 35176 11156 35216
rect 11404 35176 11444 35216
rect 11692 35176 11732 35216
rect 11788 35176 11828 35216
rect 12268 35176 12308 35216
rect 12364 35176 12404 35216
rect 12460 35176 12500 35216
rect 12940 35176 12980 35216
rect 13036 35176 13076 35216
rect 13132 35176 13172 35216
rect 13420 35176 13460 35216
rect 13516 35176 13556 35216
rect 14284 35176 14324 35216
rect 15532 35176 15572 35216
rect 16396 35092 16436 35132
rect 18988 35092 19028 35132
rect 19372 35092 19412 35132
rect 3436 35008 3476 35048
rect 12076 35008 12116 35048
rect 14092 35008 14132 35048
rect 19180 35008 19220 35048
rect 19564 35008 19604 35048
rect 3244 34924 3284 34964
rect 5932 34924 5972 34964
rect 8332 34924 8372 34964
rect 11116 34924 11156 34964
rect 16588 34924 16628 34964
rect 3688 34756 3728 34796
rect 3770 34756 3810 34796
rect 3852 34756 3892 34796
rect 3934 34756 3974 34796
rect 4016 34756 4056 34796
rect 18808 34756 18848 34796
rect 18890 34756 18930 34796
rect 18972 34756 19012 34796
rect 19054 34756 19094 34796
rect 19136 34756 19176 34796
rect 7468 34588 7508 34628
rect 7948 34588 7988 34628
rect 13420 34588 13460 34628
rect 19564 34588 19604 34628
rect 13228 34504 13268 34544
rect 14188 34504 14228 34544
rect 2668 34420 2708 34460
rect 6028 34420 6068 34460
rect 11116 34420 11156 34460
rect 19372 34420 19412 34460
rect 2188 34336 2228 34376
rect 2284 34336 2324 34376
rect 2764 34336 2804 34376
rect 3244 34336 3284 34376
rect 3724 34341 3764 34381
rect 4108 34336 4148 34376
rect 4204 34336 4244 34376
rect 5068 34336 5108 34376
rect 5164 34336 5204 34376
rect 5260 34336 5300 34376
rect 5548 34336 5588 34376
rect 5644 34336 5684 34376
rect 6124 34336 6164 34376
rect 6604 34336 6644 34376
rect 7084 34341 7124 34381
rect 7468 34336 7508 34376
rect 7756 34336 7796 34376
rect 7948 34336 7988 34376
rect 8140 34336 8180 34376
rect 8428 34336 8468 34376
rect 8524 34336 8564 34376
rect 8908 34336 8948 34376
rect 9004 34336 9044 34376
rect 9484 34336 9524 34376
rect 9964 34341 10004 34381
rect 10540 34336 10580 34376
rect 10636 34336 10676 34376
rect 11020 34336 11060 34376
rect 11596 34336 11636 34376
rect 12076 34341 12116 34381
rect 12556 34336 12596 34376
rect 12844 34336 12884 34376
rect 12940 34336 12980 34376
rect 13420 34336 13460 34376
rect 13516 34336 13556 34376
rect 13708 34336 13748 34376
rect 13804 34336 13844 34376
rect 13959 34336 13999 34376
rect 14188 34336 14228 34376
rect 14380 34333 14420 34373
rect 14764 34336 14804 34376
rect 16012 34336 16052 34376
rect 19756 34336 19796 34376
rect 3916 34252 3956 34292
rect 7276 34252 7316 34292
rect 4396 34168 4436 34208
rect 4972 34168 5012 34208
rect 10156 34168 10196 34208
rect 12268 34168 12308 34208
rect 14572 34168 14612 34208
rect 19852 34168 19892 34208
rect 4928 34000 4968 34040
rect 5010 34000 5050 34040
rect 5092 34000 5132 34040
rect 5174 34000 5214 34040
rect 5256 34000 5296 34040
rect 20048 34000 20088 34040
rect 20130 34000 20170 34040
rect 20212 34000 20252 34040
rect 20294 34000 20334 34040
rect 20376 34000 20416 34040
rect 3148 33832 3188 33872
rect 6220 33832 6260 33872
rect 7756 33832 7796 33872
rect 9772 33832 9812 33872
rect 11404 33832 11444 33872
rect 11692 33832 11732 33872
rect 12460 33832 12500 33872
rect 12748 33832 12788 33872
rect 14284 33832 14324 33872
rect 14668 33832 14708 33872
rect 5644 33748 5684 33788
rect 6988 33748 7028 33788
rect 1708 33664 1748 33704
rect 2956 33664 2996 33704
rect 3532 33664 3572 33704
rect 3820 33664 3860 33704
rect 4204 33664 4244 33704
rect 5452 33664 5492 33704
rect 6028 33664 6068 33704
rect 6124 33664 6164 33704
rect 6316 33664 6356 33704
rect 6604 33664 6644 33704
rect 6892 33664 6932 33704
rect 7468 33664 7508 33704
rect 7564 33664 7604 33704
rect 8332 33664 8372 33704
rect 9580 33664 9620 33704
rect 9964 33664 10004 33704
rect 11212 33664 11252 33704
rect 11596 33664 11636 33704
rect 11788 33664 11828 33704
rect 11884 33664 11924 33704
rect 12364 33664 12404 33704
rect 12652 33664 12692 33704
rect 12844 33664 12884 33704
rect 12940 33664 12980 33704
rect 13132 33664 13172 33704
rect 13516 33664 13556 33704
rect 13708 33664 13748 33704
rect 13900 33664 13940 33704
rect 13996 33664 14036 33704
rect 14188 33664 14228 33704
rect 14476 33664 14516 33704
rect 14860 33664 14900 33704
rect 16108 33664 16148 33704
rect 13228 33580 13268 33620
rect 13420 33580 13460 33620
rect 13324 33496 13364 33536
rect 13996 33496 14036 33536
rect 3532 33412 3572 33452
rect 7276 33412 7316 33452
rect 3688 33244 3728 33284
rect 3770 33244 3810 33284
rect 3852 33244 3892 33284
rect 3934 33244 3974 33284
rect 4016 33244 4056 33284
rect 18808 33244 18848 33284
rect 18890 33244 18930 33284
rect 18972 33244 19012 33284
rect 19054 33244 19094 33284
rect 19136 33244 19176 33284
rect 13708 33076 13748 33116
rect 7948 32992 7988 33032
rect 13420 32992 13460 33032
rect 3148 32908 3188 32948
rect 8428 32908 8468 32948
rect 2668 32804 2708 32844
rect 2764 32824 2804 32864
rect 3244 32824 3284 32864
rect 3724 32824 3764 32864
rect 4204 32829 4244 32869
rect 6124 32824 6164 32864
rect 7372 32824 7412 32864
rect 7756 32824 7796 32864
rect 7948 32820 7988 32860
rect 8044 32824 8084 32864
rect 8236 32817 8276 32857
rect 8524 32824 8564 32864
rect 12268 32824 12308 32864
rect 12460 32824 12500 32864
rect 13228 32824 13268 32864
rect 13420 32824 13460 32864
rect 13516 32824 13556 32864
rect 13804 32824 13844 32864
rect 13996 32824 14036 32864
rect 15244 32824 15284 32864
rect 16204 32824 16244 32864
rect 17452 32824 17492 32864
rect 4396 32740 4436 32780
rect 12364 32740 12404 32780
rect 7564 32656 7604 32696
rect 15436 32656 15476 32696
rect 17644 32656 17684 32696
rect 4928 32488 4968 32528
rect 5010 32488 5050 32528
rect 5092 32488 5132 32528
rect 5174 32488 5214 32528
rect 5256 32488 5296 32528
rect 20048 32488 20088 32528
rect 20130 32488 20170 32528
rect 20212 32488 20252 32528
rect 20294 32488 20334 32528
rect 20376 32488 20416 32528
rect 3916 32320 3956 32360
rect 5548 32320 5588 32360
rect 10732 32320 10772 32360
rect 11212 32320 11252 32360
rect 13708 32320 13748 32360
rect 7564 32236 7604 32276
rect 8428 32236 8468 32276
rect 2476 32152 2516 32192
rect 3724 32152 3764 32192
rect 4108 32152 4148 32192
rect 5356 32152 5396 32192
rect 5836 32152 5876 32192
rect 5932 32172 5972 32212
rect 6892 32152 6932 32192
rect 7372 32138 7412 32178
rect 8044 32152 8084 32192
rect 8332 32152 8372 32192
rect 9292 32152 9332 32192
rect 10540 32152 10580 32192
rect 10924 32152 10964 32192
rect 11020 32152 11060 32192
rect 11404 32152 11444 32192
rect 12652 32152 12692 32192
rect 12844 32152 12884 32192
rect 12940 32152 12980 32192
rect 13132 32152 13172 32192
rect 13804 32152 13844 32192
rect 14380 32152 14420 32192
rect 14476 32152 14516 32192
rect 14668 32152 14708 32192
rect 14860 32152 14900 32192
rect 15148 32152 15188 32192
rect 15340 32152 15380 32192
rect 16588 32152 16628 32192
rect 6316 32068 6356 32108
rect 6412 32068 6452 32108
rect 14956 32068 14996 32108
rect 14668 31984 14708 32024
rect 8716 31900 8756 31940
rect 9100 31900 9140 31940
rect 11212 31900 11252 31940
rect 12940 31900 12980 31940
rect 16780 31900 16820 31940
rect 3688 31732 3728 31772
rect 3770 31732 3810 31772
rect 3852 31732 3892 31772
rect 3934 31732 3974 31772
rect 4016 31732 4056 31772
rect 18808 31732 18848 31772
rect 18890 31732 18930 31772
rect 18972 31732 19012 31772
rect 19054 31732 19094 31772
rect 19136 31732 19176 31772
rect 8332 31564 8372 31604
rect 10828 31564 10868 31604
rect 12940 31564 12980 31604
rect 2668 31480 2708 31520
rect 6700 31480 6740 31520
rect 14956 31480 14996 31520
rect 15628 31480 15668 31520
rect 5068 31396 5108 31436
rect 1228 31312 1268 31352
rect 2476 31312 2516 31352
rect 2860 31312 2900 31352
rect 2956 31312 2996 31352
rect 3148 31312 3188 31352
rect 3244 31312 3284 31352
rect 3345 31312 3385 31352
rect 3628 31312 3668 31352
rect 3729 31322 3769 31362
rect 4492 31312 4532 31352
rect 4588 31312 4628 31352
rect 4972 31312 5012 31352
rect 5548 31312 5588 31352
rect 6028 31317 6068 31357
rect 6508 31312 6548 31352
rect 6700 31312 6740 31352
rect 6892 31312 6932 31352
rect 8140 31312 8180 31352
rect 9100 31312 9140 31352
rect 9388 31312 9428 31352
rect 10636 31312 10676 31352
rect 11212 31312 11252 31352
rect 11308 31312 11348 31352
rect 11500 31312 11540 31352
rect 12748 31312 12788 31352
rect 13132 31312 13172 31352
rect 13324 31312 13364 31352
rect 13516 31312 13556 31352
rect 14764 31312 14804 31352
rect 15148 31312 15188 31352
rect 15244 31312 15284 31352
rect 15436 31312 15476 31352
rect 15628 31312 15668 31352
rect 15820 31312 15860 31352
rect 16108 31312 16148 31352
rect 16204 31292 16244 31332
rect 16588 31312 16628 31352
rect 16684 31312 16724 31352
rect 17164 31312 17204 31352
rect 17644 31326 17684 31366
rect 18220 31312 18260 31352
rect 19468 31312 19508 31352
rect 19852 31312 19892 31352
rect 20044 31312 20084 31352
rect 6220 31228 6260 31268
rect 15340 31228 15380 31268
rect 17836 31228 17876 31268
rect 3052 31144 3092 31184
rect 3916 31144 3956 31184
rect 9196 31144 9236 31184
rect 10828 31144 10868 31184
rect 11020 31144 11060 31184
rect 13228 31144 13268 31184
rect 19660 31144 19700 31184
rect 19948 31144 19988 31184
rect 4928 30976 4968 31016
rect 5010 30976 5050 31016
rect 5092 30976 5132 31016
rect 5174 30976 5214 31016
rect 5256 30976 5296 31016
rect 20048 30976 20088 31016
rect 20130 30976 20170 31016
rect 20212 30976 20252 31016
rect 20294 30976 20334 31016
rect 20376 30976 20416 31016
rect 1708 30808 1748 30848
rect 1996 30808 2036 30848
rect 3820 30808 3860 30848
rect 13228 30808 13268 30848
rect 15436 30808 15476 30848
rect 15916 30808 15956 30848
rect 19756 30808 19796 30848
rect 5836 30724 5876 30764
rect 8524 30724 8564 30764
rect 10540 30724 10580 30764
rect 11212 30724 11252 30764
rect 12460 30724 12500 30764
rect 18796 30724 18836 30764
rect 1612 30640 1652 30680
rect 1900 30640 1940 30680
rect 2092 30640 2132 30680
rect 2188 30640 2228 30680
rect 2380 30640 2420 30680
rect 3628 30640 3668 30680
rect 4108 30640 4148 30680
rect 4204 30640 4244 30680
rect 4684 30640 4724 30680
rect 5164 30640 5204 30680
rect 5644 30626 5684 30666
rect 7084 30640 7124 30680
rect 8332 30640 8372 30680
rect 8812 30640 8852 30680
rect 8908 30640 8948 30680
rect 9292 30640 9332 30680
rect 9868 30640 9908 30680
rect 4588 30556 4628 30596
rect 9388 30598 9428 30638
rect 10348 30626 10388 30666
rect 10828 30640 10868 30680
rect 11116 30640 11156 30680
rect 12076 30640 12116 30680
rect 12364 30640 12404 30680
rect 12940 30640 12980 30680
rect 13036 30640 13076 30680
rect 13708 30640 13748 30680
rect 13804 30640 13844 30680
rect 14188 30640 14228 30680
rect 14764 30640 14804 30680
rect 15244 30635 15284 30675
rect 14284 30556 14324 30596
rect 15628 30595 15668 30635
rect 15724 30640 15764 30680
rect 15820 30640 15860 30680
rect 16492 30640 16532 30680
rect 17740 30640 17780 30680
rect 18412 30640 18452 30680
rect 18700 30640 18740 30680
rect 19276 30640 19316 30680
rect 19468 30640 19508 30680
rect 19564 30640 19604 30680
rect 19948 30640 19988 30680
rect 20044 30640 20084 30680
rect 11500 30472 11540 30512
rect 12748 30472 12788 30512
rect 19276 30472 19316 30512
rect 17932 30388 17972 30428
rect 19084 30388 19124 30428
rect 3688 30220 3728 30260
rect 3770 30220 3810 30260
rect 3852 30220 3892 30260
rect 3934 30220 3974 30260
rect 4016 30220 4056 30260
rect 18808 30220 18848 30260
rect 18890 30220 18930 30260
rect 18972 30220 19012 30260
rect 19054 30220 19094 30260
rect 19136 30220 19176 30260
rect 2668 30052 2708 30092
rect 4396 30052 4436 30092
rect 6028 30052 6068 30092
rect 14668 30052 14708 30092
rect 20236 30052 20276 30092
rect 9196 29968 9236 30008
rect 10156 29968 10196 30008
rect 15628 29968 15668 30008
rect 18124 29884 18164 29924
rect 1228 29800 1268 29840
rect 2476 29800 2516 29840
rect 2956 29800 2996 29840
rect 4204 29800 4244 29840
rect 4588 29800 4628 29840
rect 5836 29800 5876 29840
rect 7084 29800 7124 29840
rect 8332 29800 8372 29840
rect 9004 29800 9044 29840
rect 9196 29800 9236 29840
rect 9484 29800 9524 29840
rect 9772 29800 9812 29840
rect 10444 29800 10484 29840
rect 10636 29800 10676 29840
rect 10732 29800 10772 29840
rect 10924 29800 10964 29840
rect 12172 29800 12212 29840
rect 12652 29800 12692 29840
rect 12940 29800 12980 29840
rect 13228 29800 13268 29840
rect 14476 29800 14516 29840
rect 14956 29800 14996 29840
rect 15244 29800 15284 29840
rect 15820 29800 15860 29840
rect 15916 29800 15956 29840
rect 17548 29800 17588 29840
rect 17644 29800 17684 29840
rect 18028 29800 18068 29840
rect 18604 29800 18644 29840
rect 19084 29805 19124 29845
rect 19564 29800 19604 29840
rect 19852 29800 19892 29840
rect 9868 29716 9908 29756
rect 15340 29716 15380 29756
rect 19276 29716 19316 29756
rect 19948 29716 19988 29756
rect 8524 29632 8564 29672
rect 10540 29632 10580 29672
rect 12364 29632 12404 29672
rect 12748 29632 12788 29672
rect 16108 29632 16148 29672
rect 4928 29464 4968 29504
rect 5010 29464 5050 29504
rect 5092 29464 5132 29504
rect 5174 29464 5214 29504
rect 5256 29464 5296 29504
rect 20048 29464 20088 29504
rect 20130 29464 20170 29504
rect 20212 29464 20252 29504
rect 20294 29464 20334 29504
rect 20376 29464 20416 29504
rect 1900 29296 1940 29336
rect 3820 29296 3860 29336
rect 10732 29296 10772 29336
rect 11404 29296 11444 29336
rect 13612 29296 13652 29336
rect 16300 29296 16340 29336
rect 17740 29296 17780 29336
rect 20044 29296 20084 29336
rect 6604 29212 6644 29252
rect 8620 29212 8660 29252
rect 2380 29128 2420 29168
rect 3628 29128 3668 29168
rect 4012 29128 4052 29168
rect 4204 29128 4244 29168
rect 5164 29128 5204 29168
rect 6412 29128 6452 29168
rect 6892 29128 6932 29168
rect 6988 29128 7028 29168
rect 7372 29128 7412 29168
rect 7948 29128 7988 29168
rect 8476 29118 8516 29158
rect 9004 29128 9044 29168
rect 10252 29128 10292 29168
rect 10636 29128 10676 29168
rect 10828 29128 10868 29168
rect 10924 29128 10964 29168
rect 11116 29128 11156 29168
rect 11212 29128 11252 29168
rect 11884 29148 11924 29188
rect 11980 29128 12020 29168
rect 12364 29128 12404 29168
rect 12460 29128 12500 29168
rect 12940 29128 12980 29168
rect 14476 29128 14516 29168
rect 15724 29128 15764 29168
rect 16204 29128 16244 29168
rect 2092 29044 2132 29084
rect 7468 29044 7508 29084
rect 13468 29086 13508 29126
rect 16396 29128 16436 29168
rect 16492 29128 16532 29168
rect 16684 29128 16724 29168
rect 16780 29128 16820 29168
rect 16972 29128 17012 29168
rect 17068 29128 17108 29168
rect 17220 29128 17260 29168
rect 17452 29128 17492 29168
rect 17548 29128 17588 29168
rect 18028 29128 18068 29168
rect 18124 29128 18164 29168
rect 18316 29128 18356 29168
rect 19564 29128 19604 29168
rect 19948 29128 19988 29168
rect 20140 29128 20180 29168
rect 20236 29128 20276 29168
rect 19756 28960 19796 29000
rect 4108 28876 4148 28916
rect 10444 28876 10484 28916
rect 15916 28876 15956 28916
rect 16684 28876 16724 28916
rect 3688 28708 3728 28748
rect 3770 28708 3810 28748
rect 3852 28708 3892 28748
rect 3934 28708 3974 28748
rect 4016 28708 4056 28748
rect 18808 28708 18848 28748
rect 18890 28708 18930 28748
rect 18972 28708 19012 28748
rect 19054 28708 19094 28748
rect 19136 28708 19176 28748
rect 2668 28540 2708 28580
rect 13516 28540 13556 28580
rect 16396 28540 16436 28580
rect 5548 28456 5588 28496
rect 6412 28372 6452 28412
rect 15052 28372 15092 28412
rect 1228 28288 1268 28328
rect 2476 28288 2516 28328
rect 3148 28288 3188 28328
rect 3244 28288 3284 28328
rect 3628 28288 3668 28328
rect 3724 28288 3764 28328
rect 3916 28288 3956 28328
rect 4108 28288 4148 28328
rect 5356 28288 5396 28328
rect 5836 28288 5876 28328
rect 5932 28288 5972 28328
rect 6316 28288 6356 28328
rect 6892 28288 6932 28328
rect 7372 28293 7412 28333
rect 8044 28288 8084 28328
rect 9292 28288 9332 28328
rect 9868 28288 9908 28328
rect 11116 28288 11156 28328
rect 11500 28288 11540 28328
rect 11596 28288 11636 28328
rect 11692 28288 11732 28328
rect 12076 28288 12116 28328
rect 13324 28288 13364 28328
rect 14476 28288 14516 28328
rect 14572 28288 14612 28328
rect 14956 28288 14996 28328
rect 15532 28288 15572 28328
rect 16012 28302 16052 28342
rect 16588 28288 16628 28328
rect 17836 28288 17876 28328
rect 18220 28288 18260 28328
rect 19468 28288 19508 28328
rect 19852 28288 19892 28328
rect 19948 28288 19988 28328
rect 20044 28288 20084 28328
rect 3436 28120 3476 28160
rect 3916 28120 3956 28160
rect 7564 28120 7604 28160
rect 9484 28120 9524 28160
rect 11308 28120 11348 28160
rect 11788 28120 11828 28160
rect 16204 28120 16244 28160
rect 19660 28120 19700 28160
rect 20140 28120 20180 28160
rect 4928 27952 4968 27992
rect 5010 27952 5050 27992
rect 5092 27952 5132 27992
rect 5174 27952 5214 27992
rect 5256 27952 5296 27992
rect 20048 27952 20088 27992
rect 20130 27952 20170 27992
rect 20212 27952 20252 27992
rect 20294 27952 20334 27992
rect 20376 27952 20416 27992
rect 4492 27784 4532 27824
rect 7372 27784 7412 27824
rect 14476 27784 14516 27824
rect 17356 27784 17396 27824
rect 20044 27784 20084 27824
rect 2668 27700 2708 27740
rect 4300 27700 4340 27740
rect 10348 27700 10388 27740
rect 1228 27616 1268 27656
rect 2476 27616 2516 27656
rect 2860 27616 2900 27656
rect 4108 27616 4148 27656
rect 4684 27616 4724 27656
rect 4780 27616 4820 27656
rect 4972 27616 5012 27656
rect 5260 27616 5300 27656
rect 5452 27616 5492 27656
rect 5644 27616 5684 27656
rect 5932 27616 5972 27656
rect 7180 27616 7220 27656
rect 8620 27616 8660 27656
rect 8716 27616 8756 27656
rect 9100 27616 9140 27656
rect 9676 27616 9716 27656
rect 10204 27606 10244 27646
rect 10924 27616 10964 27656
rect 12172 27616 12212 27656
rect 13036 27616 13076 27656
rect 14284 27616 14324 27656
rect 15628 27616 15668 27656
rect 15724 27616 15764 27656
rect 15916 27616 15956 27656
rect 17164 27616 17204 27656
rect 18124 27616 18164 27656
rect 19372 27595 19412 27635
rect 19756 27617 19796 27657
rect 19852 27616 19892 27656
rect 9196 27532 9236 27572
rect 5452 27448 5492 27488
rect 5260 27364 5300 27404
rect 12364 27364 12404 27404
rect 19564 27364 19604 27404
rect 3688 27196 3728 27236
rect 3770 27196 3810 27236
rect 3852 27196 3892 27236
rect 3934 27196 3974 27236
rect 4016 27196 4056 27236
rect 18808 27196 18848 27236
rect 18890 27196 18930 27236
rect 18972 27196 19012 27236
rect 19054 27196 19094 27236
rect 19136 27196 19176 27236
rect 4108 27028 4148 27068
rect 1996 26860 2036 26900
rect 6796 26860 6836 26900
rect 17836 26860 17876 26900
rect 1420 26776 1460 26816
rect 1516 26776 1556 26816
rect 1900 26776 1940 26816
rect 2476 26776 2516 26816
rect 3004 26785 3044 26825
rect 3436 26776 3476 26816
rect 3724 26776 3764 26816
rect 4492 26776 4532 26816
rect 5740 26776 5780 26816
rect 6220 26776 6260 26816
rect 6316 26776 6356 26816
rect 6700 26776 6740 26816
rect 7276 26776 7316 26816
rect 7756 26781 7796 26821
rect 8332 26776 8372 26816
rect 9580 26776 9620 26816
rect 10060 26776 10100 26816
rect 10156 26776 10196 26816
rect 10252 26776 10292 26816
rect 10540 26776 10580 26816
rect 10636 26776 10676 26816
rect 11020 26776 11060 26816
rect 11116 26776 11156 26816
rect 11788 26776 11828 26816
rect 11884 26776 11924 26816
rect 12268 26776 12308 26816
rect 12364 26776 12404 26816
rect 12844 26776 12884 26816
rect 13372 26785 13412 26825
rect 14188 26776 14228 26816
rect 15436 26776 15476 26816
rect 15820 26776 15860 26816
rect 16012 26776 16052 26816
rect 16108 26776 16148 26816
rect 17356 26776 17396 26816
rect 17452 26776 17492 26816
rect 17932 26776 17972 26816
rect 18412 26776 18452 26816
rect 18940 26785 18980 26825
rect 19276 26776 19316 26816
rect 19372 26776 19412 26816
rect 19468 26776 19508 26816
rect 19756 26776 19796 26816
rect 19852 26776 19892 26816
rect 3148 26692 3188 26732
rect 3820 26692 3860 26732
rect 5932 26692 5972 26732
rect 7948 26692 7988 26732
rect 8140 26692 8180 26732
rect 10348 26692 10388 26732
rect 15628 26692 15668 26732
rect 10828 26608 10868 26648
rect 11308 26608 11348 26648
rect 13516 26608 13556 26648
rect 15916 26608 15956 26648
rect 19084 26608 19124 26648
rect 19564 26608 19604 26648
rect 20044 26608 20084 26648
rect 4928 26440 4968 26480
rect 5010 26440 5050 26480
rect 5092 26440 5132 26480
rect 5174 26440 5214 26480
rect 5256 26440 5296 26480
rect 20048 26440 20088 26480
rect 20130 26440 20170 26480
rect 20212 26440 20252 26480
rect 20294 26440 20334 26480
rect 20376 26440 20416 26480
rect 2956 26272 2996 26312
rect 5452 26272 5492 26312
rect 11212 26272 11252 26312
rect 13420 26272 13460 26312
rect 17644 26272 17684 26312
rect 19276 26272 19316 26312
rect 15820 26188 15860 26228
rect 1516 26104 1556 26144
rect 2764 26104 2804 26144
rect 3532 26104 3572 26144
rect 4780 26104 4820 26144
rect 5164 26104 5204 26144
rect 5260 26104 5300 26144
rect 6124 26104 6164 26144
rect 7372 26104 7412 26144
rect 7756 26104 7796 26144
rect 9004 26104 9044 26144
rect 9484 26104 9524 26144
rect 9580 26104 9620 26144
rect 10540 26104 10580 26144
rect 11068 26094 11108 26134
rect 11980 26104 12020 26144
rect 13228 26104 13268 26144
rect 14092 26104 14132 26144
rect 14188 26104 14228 26144
rect 14668 26104 14708 26144
rect 15148 26104 15188 26144
rect 15628 26099 15668 26139
rect 16204 26104 16244 26144
rect 17452 26104 17492 26144
rect 17836 26104 17876 26144
rect 19084 26104 19124 26144
rect 19468 26104 19508 26144
rect 19564 26104 19604 26144
rect 9964 26020 10004 26060
rect 10060 26020 10100 26060
rect 14572 26020 14612 26060
rect 4972 25852 5012 25892
rect 7564 25852 7604 25892
rect 9196 25852 9236 25892
rect 16012 25852 16052 25892
rect 3688 25684 3728 25724
rect 3770 25684 3810 25724
rect 3852 25684 3892 25724
rect 3934 25684 3974 25724
rect 4016 25684 4056 25724
rect 18808 25684 18848 25724
rect 18890 25684 18930 25724
rect 18972 25684 19012 25724
rect 19054 25684 19094 25724
rect 19136 25684 19176 25724
rect 11212 25516 11252 25556
rect 14572 25516 14612 25556
rect 15148 25516 15188 25556
rect 15628 25516 15668 25556
rect 16300 25432 16340 25472
rect 17356 25432 17396 25472
rect 2380 25264 2420 25304
rect 2476 25264 2516 25304
rect 2764 25264 2804 25304
rect 2860 25264 2900 25304
rect 3244 25264 3284 25304
rect 3340 25264 3380 25304
rect 3820 25264 3860 25304
rect 4300 25269 4340 25309
rect 4684 25264 4724 25304
rect 4780 25264 4820 25304
rect 4876 25264 4916 25304
rect 5164 25264 5204 25304
rect 5260 25264 5300 25304
rect 5356 25264 5396 25304
rect 5452 25243 5492 25283
rect 5836 25264 5876 25304
rect 5932 25264 5972 25304
rect 6220 25264 6260 25304
rect 6316 25264 6356 25304
rect 6700 25264 6740 25304
rect 6796 25264 6836 25304
rect 7276 25264 7316 25304
rect 7756 25278 7796 25318
rect 8140 25264 8180 25304
rect 8236 25264 8276 25304
rect 9772 25264 9812 25304
rect 11020 25264 11060 25304
rect 13132 25264 13172 25304
rect 14380 25264 14420 25304
rect 14956 25264 14996 25304
rect 15148 25264 15188 25304
rect 15340 25264 15380 25304
rect 15628 25264 15668 25304
rect 15916 25264 15956 25304
rect 16012 25264 16052 25304
rect 16108 25264 16148 25304
rect 16684 25264 16724 25304
rect 16972 25264 17012 25304
rect 17068 25264 17108 25304
rect 4492 25180 4532 25220
rect 7948 25180 7988 25220
rect 2188 25096 2228 25136
rect 4972 25096 5012 25136
rect 5644 25096 5684 25136
rect 8428 25096 8468 25136
rect 4928 24928 4968 24968
rect 5010 24928 5050 24968
rect 5092 24928 5132 24968
rect 5174 24928 5214 24968
rect 5256 24928 5296 24968
rect 20048 24928 20088 24968
rect 20130 24928 20170 24968
rect 20212 24928 20252 24968
rect 20294 24928 20334 24968
rect 20376 24928 20416 24968
rect 2764 24760 2804 24800
rect 2956 24760 2996 24800
rect 6316 24760 6356 24800
rect 11020 24802 11060 24842
rect 16780 24760 16820 24800
rect 9004 24676 9044 24716
rect 1324 24592 1364 24632
rect 2572 24592 2612 24632
rect 3148 24592 3188 24632
rect 4396 24592 4436 24632
rect 4876 24592 4916 24632
rect 6124 24592 6164 24632
rect 6700 24592 6740 24632
rect 6988 24592 7028 24632
rect 7084 24592 7124 24632
rect 7564 24592 7604 24632
rect 8812 24592 8852 24632
rect 9292 24573 9332 24613
rect 9388 24573 9428 24613
rect 9868 24592 9908 24632
rect 10348 24592 10388 24632
rect 10828 24578 10868 24618
rect 11404 24592 11444 24632
rect 12652 24592 12692 24632
rect 13132 24592 13172 24632
rect 14380 24592 14420 24632
rect 15340 24592 15380 24632
rect 16588 24592 16628 24632
rect 16972 24592 17012 24632
rect 17068 24592 17108 24632
rect 17164 24592 17204 24632
rect 17260 24592 17300 24632
rect 18220 24592 18260 24632
rect 19468 24592 19508 24632
rect 9772 24508 9812 24548
rect 7372 24424 7412 24464
rect 11212 24340 11252 24380
rect 14572 24340 14612 24380
rect 18028 24340 18068 24380
rect 3688 24172 3728 24212
rect 3770 24172 3810 24212
rect 3852 24172 3892 24212
rect 3934 24172 3974 24212
rect 4016 24172 4056 24212
rect 18808 24172 18848 24212
rect 18890 24172 18930 24212
rect 18972 24172 19012 24212
rect 19054 24172 19094 24212
rect 19136 24172 19176 24212
rect 1228 24004 1268 24044
rect 3820 24004 3860 24044
rect 10924 24004 10964 24044
rect 12364 24004 12404 24044
rect 15628 24004 15668 24044
rect 8428 23920 8468 23960
rect 9100 23920 9140 23960
rect 11692 23920 11732 23960
rect 6220 23836 6260 23876
rect 6316 23836 6356 23876
rect 16492 23836 16532 23876
rect 1420 23752 1460 23792
rect 2668 23752 2708 23792
rect 3148 23752 3188 23792
rect 3436 23752 3476 23792
rect 4012 23752 4052 23792
rect 5260 23752 5300 23792
rect 5740 23752 5780 23792
rect 5836 23752 5876 23792
rect 6796 23752 6836 23792
rect 7276 23766 7316 23806
rect 7756 23752 7796 23792
rect 8044 23752 8084 23792
rect 8620 23752 8660 23792
rect 8716 23752 8756 23792
rect 8908 23752 8948 23792
rect 9100 23752 9140 23792
rect 9292 23752 9332 23792
rect 9484 23752 9524 23792
rect 10732 23752 10772 23792
rect 11500 23752 11540 23792
rect 11692 23752 11732 23792
rect 11884 23752 11924 23792
rect 12076 23752 12116 23792
rect 12172 23752 12212 23792
rect 12364 23752 12404 23792
rect 12556 23752 12596 23792
rect 12652 23752 12692 23792
rect 13036 23752 13076 23792
rect 13132 23752 13172 23792
rect 13516 23752 13556 23792
rect 13612 23752 13652 23792
rect 13996 23752 14036 23792
rect 14092 23752 14132 23792
rect 14572 23752 14612 23792
rect 15052 23757 15092 23797
rect 15532 23741 15572 23781
rect 15916 23752 15956 23792
rect 16012 23752 16052 23792
rect 16396 23752 16436 23792
rect 16972 23752 17012 23792
rect 17452 23757 17492 23797
rect 18124 23752 18164 23792
rect 19372 23752 19412 23792
rect 19756 23752 19796 23792
rect 19852 23752 19892 23792
rect 3532 23668 3572 23708
rect 5452 23668 5492 23708
rect 7468 23668 7508 23708
rect 8140 23668 8180 23708
rect 15244 23668 15284 23708
rect 17644 23668 17684 23708
rect 8812 23584 8852 23624
rect 12844 23584 12884 23624
rect 19564 23584 19604 23624
rect 20044 23584 20084 23624
rect 4928 23416 4968 23456
rect 5010 23416 5050 23456
rect 5092 23416 5132 23456
rect 5174 23416 5214 23456
rect 5256 23416 5296 23456
rect 20048 23416 20088 23456
rect 20130 23416 20170 23456
rect 20212 23416 20252 23456
rect 20294 23416 20334 23456
rect 20376 23416 20416 23456
rect 3724 23248 3764 23288
rect 7084 23248 7124 23288
rect 11692 23248 11732 23288
rect 15436 23248 15476 23288
rect 18220 23248 18260 23288
rect 19468 23248 19508 23288
rect 19948 23248 19988 23288
rect 8716 23164 8756 23204
rect 11500 23164 11540 23204
rect 1420 23080 1460 23120
rect 1708 23080 1748 23120
rect 1996 23080 2036 23120
rect 2092 23080 2132 23120
rect 2476 23080 2516 23120
rect 2572 23080 2612 23120
rect 3052 23080 3092 23120
rect 3532 23066 3572 23106
rect 3916 23080 3956 23120
rect 5164 23080 5204 23120
rect 5644 23080 5684 23120
rect 6892 23080 6932 23120
rect 7276 23080 7316 23120
rect 8524 23080 8564 23120
rect 9004 23080 9044 23120
rect 10060 23080 10100 23120
rect 11308 23080 11348 23120
rect 11884 23066 11924 23106
rect 12364 23080 12404 23120
rect 12844 23080 12884 23120
rect 13324 23080 13364 23120
rect 13420 23080 13460 23120
rect 13996 23080 14036 23120
rect 15244 23080 15284 23120
rect 15724 23080 15764 23120
rect 16012 23107 16052 23147
rect 16780 23080 16820 23120
rect 18028 23080 18068 23120
rect 18412 23080 18452 23120
rect 16108 23038 16148 23078
rect 18508 23080 18548 23120
rect 18604 23080 18644 23120
rect 18700 23080 18740 23120
rect 19180 23080 19220 23120
rect 19276 23080 19316 23120
rect 19660 23080 19700 23120
rect 19756 23080 19796 23120
rect 19852 23080 19892 23120
rect 12940 22996 12980 23036
rect 16396 22912 16436 22952
rect 1708 22828 1748 22868
rect 5356 22828 5396 22868
rect 7084 22828 7124 22868
rect 8908 22828 8948 22868
rect 3688 22660 3728 22700
rect 3770 22660 3810 22700
rect 3852 22660 3892 22700
rect 3934 22660 3974 22700
rect 4016 22660 4056 22700
rect 18808 22660 18848 22700
rect 18890 22660 18930 22700
rect 18972 22660 19012 22700
rect 19054 22660 19094 22700
rect 19136 22660 19176 22700
rect 2668 22492 2708 22532
rect 2860 22492 2900 22532
rect 8332 22492 8372 22532
rect 12844 22492 12884 22532
rect 6124 22408 6164 22448
rect 1228 22240 1268 22280
rect 2476 22240 2516 22280
rect 3052 22240 3092 22280
rect 4300 22240 4340 22280
rect 4492 22240 4532 22280
rect 5740 22240 5780 22280
rect 6124 22240 6164 22280
rect 6220 22240 6260 22280
rect 6412 22240 6452 22280
rect 6604 22240 6644 22280
rect 6796 22240 6836 22280
rect 8044 22240 8084 22280
rect 8140 22240 8180 22280
rect 8332 22240 8372 22280
rect 11596 22240 11636 22280
rect 11692 22240 11732 22280
rect 11788 22240 11828 22280
rect 11884 22240 11924 22280
rect 12172 22240 12212 22280
rect 12460 22240 12500 22280
rect 13036 22240 13076 22280
rect 13228 22240 13268 22280
rect 13324 22240 13364 22280
rect 13708 22240 13748 22280
rect 14956 22240 14996 22280
rect 16972 22240 17012 22280
rect 17452 22240 17492 22280
rect 17548 22240 17588 22280
rect 6700 22156 6740 22196
rect 12556 22156 12596 22196
rect 13132 22156 13172 22196
rect 5932 22072 5972 22112
rect 15148 22072 15188 22112
rect 17068 22072 17108 22112
rect 17740 22072 17780 22112
rect 4928 21904 4968 21944
rect 5010 21904 5050 21944
rect 5092 21904 5132 21944
rect 5174 21904 5214 21944
rect 5256 21904 5296 21944
rect 20048 21904 20088 21944
rect 20130 21904 20170 21944
rect 20212 21904 20252 21944
rect 20294 21904 20334 21944
rect 20376 21904 20416 21944
rect 3148 21736 3188 21776
rect 6988 21736 7028 21776
rect 12844 21736 12884 21776
rect 15244 21736 15284 21776
rect 5356 21652 5396 21692
rect 5932 21652 5972 21692
rect 9004 21652 9044 21692
rect 11020 21652 11060 21692
rect 17356 21652 17396 21692
rect 1708 21568 1748 21608
rect 2956 21568 2996 21608
rect 3628 21568 3668 21608
rect 3724 21568 3764 21608
rect 4108 21568 4148 21608
rect 4204 21568 4244 21608
rect 4684 21568 4724 21608
rect 5164 21563 5204 21603
rect 5740 21568 5780 21608
rect 5836 21568 5876 21608
rect 6028 21568 6068 21608
rect 6220 21568 6260 21608
rect 6316 21568 6356 21608
rect 6508 21568 6548 21608
rect 6700 21568 6740 21608
rect 6796 21568 6836 21608
rect 6892 21568 6932 21608
rect 7180 21568 7220 21608
rect 7372 21568 7412 21608
rect 7564 21568 7604 21608
rect 8812 21568 8852 21608
rect 9292 21568 9332 21608
rect 9388 21568 9428 21608
rect 9772 21568 9812 21608
rect 9868 21568 9908 21608
rect 10348 21568 10388 21608
rect 10876 21558 10916 21598
rect 11404 21568 11444 21608
rect 12652 21568 12692 21608
rect 13516 21568 13556 21608
rect 13612 21568 13652 21608
rect 13996 21568 14036 21608
rect 14092 21568 14132 21608
rect 14572 21568 14612 21608
rect 15100 21558 15140 21598
rect 15628 21568 15668 21608
rect 15724 21568 15764 21608
rect 16108 21568 16148 21608
rect 16204 21568 16244 21608
rect 16684 21568 16724 21608
rect 17164 21554 17204 21594
rect 17740 21568 17780 21608
rect 18988 21568 19028 21608
rect 7180 21400 7220 21440
rect 17548 21400 17588 21440
rect 3688 21148 3728 21188
rect 3770 21148 3810 21188
rect 3852 21148 3892 21188
rect 3934 21148 3974 21188
rect 4016 21148 4056 21188
rect 18808 21148 18848 21188
rect 18890 21148 18930 21188
rect 18972 21148 19012 21188
rect 19054 21148 19094 21188
rect 19136 21148 19176 21188
rect 4876 20980 4916 21020
rect 11020 20980 11060 21020
rect 13708 20980 13748 21020
rect 15820 20980 15860 21020
rect 16876 20896 16916 20936
rect 17836 20896 17876 20936
rect 1996 20812 2036 20852
rect 2092 20812 2132 20852
rect 7756 20812 7796 20852
rect 7852 20812 7892 20852
rect 1516 20728 1556 20768
rect 1612 20728 1652 20768
rect 2572 20728 2612 20768
rect 3052 20733 3092 20773
rect 3436 20728 3476 20768
rect 4684 20728 4724 20768
rect 5068 20728 5108 20768
rect 5164 20728 5204 20768
rect 5548 20728 5588 20768
rect 6796 20728 6836 20768
rect 7276 20728 7316 20768
rect 7372 20728 7412 20768
rect 8332 20728 8372 20768
rect 8860 20737 8900 20777
rect 9580 20728 9620 20768
rect 10828 20728 10868 20768
rect 12268 20728 12308 20768
rect 13516 20728 13556 20768
rect 14380 20728 14420 20768
rect 15628 20728 15668 20768
rect 16204 20728 16244 20768
rect 16492 20728 16532 20768
rect 16588 20728 16628 20768
rect 17164 20728 17204 20768
rect 17452 20728 17492 20768
rect 18028 20728 18068 20768
rect 18124 20728 18164 20768
rect 18508 20728 18548 20768
rect 18700 20728 18740 20768
rect 17548 20644 17588 20684
rect 5356 20602 5396 20642
rect 3244 20560 3284 20600
rect 6988 20560 7028 20600
rect 9004 20560 9044 20600
rect 18316 20560 18356 20600
rect 18604 20560 18644 20600
rect 4928 20392 4968 20432
rect 5010 20392 5050 20432
rect 5092 20392 5132 20432
rect 5174 20392 5214 20432
rect 5256 20392 5296 20432
rect 20048 20392 20088 20432
rect 20130 20392 20170 20432
rect 20212 20392 20252 20432
rect 20294 20392 20334 20432
rect 20376 20392 20416 20432
rect 8908 20224 8948 20264
rect 3916 20140 3956 20180
rect 5164 20140 5204 20180
rect 10540 20140 10580 20180
rect 12556 20140 12596 20180
rect 2476 20056 2516 20096
rect 3724 20056 3764 20096
rect 4396 20056 4436 20096
rect 4492 20056 4532 20096
rect 4684 20056 4724 20096
rect 5260 20056 5300 20096
rect 5548 20056 5588 20096
rect 5836 20056 5876 20096
rect 7084 20056 7124 20096
rect 7468 20056 7508 20096
rect 8716 20056 8756 20096
rect 9100 20056 9140 20096
rect 10348 20056 10388 20096
rect 10828 20056 10868 20096
rect 10924 20056 10964 20096
rect 11404 20056 11444 20096
rect 11884 20014 11924 20054
rect 12364 20046 12404 20086
rect 12748 20056 12788 20096
rect 13996 20056 14036 20096
rect 14380 20056 14420 20096
rect 15628 20056 15668 20096
rect 16876 20056 16916 20096
rect 17260 20056 17300 20096
rect 17452 20042 17492 20082
rect 17552 20037 17592 20077
rect 17740 20056 17780 20096
rect 17932 20056 17972 20096
rect 18028 20056 18068 20096
rect 11308 19972 11348 20012
rect 4684 19888 4724 19928
rect 4876 19888 4916 19928
rect 17068 19888 17108 19928
rect 7276 19804 7316 19844
rect 14188 19804 14228 19844
rect 14476 19804 14516 19844
rect 17260 19804 17300 19844
rect 17740 19804 17780 19844
rect 3688 19636 3728 19676
rect 3770 19636 3810 19676
rect 3852 19636 3892 19676
rect 3934 19636 3974 19676
rect 4016 19636 4056 19676
rect 18808 19636 18848 19676
rect 18890 19636 18930 19676
rect 18972 19636 19012 19676
rect 19054 19636 19094 19676
rect 19136 19636 19176 19676
rect 2764 19468 2804 19508
rect 12652 19468 12692 19508
rect 6508 19300 6548 19340
rect 9100 19300 9140 19340
rect 13996 19300 14036 19340
rect 1324 19216 1364 19256
rect 2572 19216 2612 19256
rect 4204 19216 4244 19256
rect 5452 19216 5492 19256
rect 5932 19216 5972 19256
rect 6028 19216 6068 19256
rect 6412 19216 6452 19256
rect 6988 19216 7028 19256
rect 7468 19230 7508 19270
rect 8620 19216 8660 19256
rect 8716 19216 8756 19256
rect 9196 19216 9236 19256
rect 9676 19216 9716 19256
rect 10204 19225 10244 19265
rect 11212 19216 11252 19256
rect 12460 19216 12500 19256
rect 13516 19216 13556 19256
rect 13612 19216 13652 19256
rect 14092 19216 14132 19256
rect 14572 19216 14612 19256
rect 15100 19225 15140 19265
rect 17452 19216 17492 19256
rect 18700 19216 18740 19256
rect 5644 19048 5684 19088
rect 7660 19048 7700 19088
rect 10348 19048 10388 19088
rect 15244 19048 15284 19088
rect 18892 19048 18932 19088
rect 4928 18880 4968 18920
rect 5010 18880 5050 18920
rect 5092 18880 5132 18920
rect 5174 18880 5214 18920
rect 5256 18880 5296 18920
rect 20048 18880 20088 18920
rect 20130 18880 20170 18920
rect 20212 18880 20252 18920
rect 20294 18880 20334 18920
rect 20376 18880 20416 18920
rect 2668 18712 2708 18752
rect 3148 18712 3188 18752
rect 15244 18712 15284 18752
rect 15724 18712 15764 18752
rect 7756 18628 7796 18668
rect 10732 18628 10772 18668
rect 12748 18628 12788 18668
rect 18700 18628 18740 18668
rect 1228 18544 1268 18584
rect 2476 18544 2516 18584
rect 2860 18544 2900 18584
rect 2956 18544 2996 18584
rect 4300 18544 4340 18584
rect 5548 18544 5588 18584
rect 6028 18544 6068 18584
rect 6124 18544 6164 18584
rect 6508 18544 6548 18584
rect 6604 18544 6644 18584
rect 7084 18544 7124 18584
rect 7564 18530 7604 18570
rect 9292 18544 9332 18584
rect 10540 18544 10580 18584
rect 11020 18544 11060 18584
rect 11116 18544 11156 18584
rect 11500 18544 11540 18584
rect 12076 18544 12116 18584
rect 12556 18530 12596 18570
rect 13804 18544 13844 18584
rect 15052 18544 15092 18584
rect 15436 18544 15476 18584
rect 15532 18529 15572 18569
rect 15724 18544 15764 18584
rect 15820 18544 15860 18584
rect 15921 18544 15961 18584
rect 16972 18544 17012 18584
rect 17068 18544 17108 18584
rect 17548 18544 17588 18584
rect 18028 18544 18068 18584
rect 18556 18534 18596 18574
rect 11596 18460 11636 18500
rect 17452 18460 17492 18500
rect 5740 18376 5780 18416
rect 3688 18124 3728 18164
rect 3770 18124 3810 18164
rect 3852 18124 3892 18164
rect 3934 18124 3974 18164
rect 4016 18124 4056 18164
rect 18808 18124 18848 18164
rect 18890 18124 18930 18164
rect 18972 18124 19012 18164
rect 19054 18124 19094 18164
rect 19136 18124 19176 18164
rect 7084 17956 7124 17996
rect 8716 17956 8756 17996
rect 10348 17956 10388 17996
rect 12940 17956 12980 17996
rect 14956 17956 14996 17996
rect 17068 17956 17108 17996
rect 4108 17788 4148 17828
rect 1324 17704 1364 17744
rect 1516 17704 1556 17744
rect 1612 17704 1652 17744
rect 1804 17704 1844 17744
rect 3052 17704 3092 17744
rect 3532 17704 3572 17744
rect 3628 17704 3668 17744
rect 4588 17746 4628 17786
rect 4012 17704 4052 17744
rect 5068 17709 5108 17749
rect 5644 17704 5684 17744
rect 6892 17704 6932 17744
rect 7276 17704 7316 17744
rect 8524 17704 8564 17744
rect 8908 17704 8948 17744
rect 10156 17704 10196 17744
rect 11500 17704 11540 17744
rect 12748 17704 12788 17744
rect 13516 17704 13556 17744
rect 14764 17704 14804 17744
rect 15148 17704 15188 17744
rect 15244 17704 15284 17744
rect 15628 17704 15668 17744
rect 16876 17704 16916 17744
rect 17644 17704 17684 17744
rect 18892 17704 18932 17744
rect 3244 17620 3284 17660
rect 19084 17620 19124 17660
rect 1420 17536 1460 17576
rect 5260 17536 5300 17576
rect 14956 17536 14996 17576
rect 15436 17536 15476 17576
rect 4928 17368 4968 17408
rect 5010 17368 5050 17408
rect 5092 17368 5132 17408
rect 5174 17368 5214 17408
rect 5256 17368 5296 17408
rect 20048 17368 20088 17408
rect 20130 17368 20170 17408
rect 20212 17368 20252 17408
rect 20294 17368 20334 17408
rect 20376 17368 20416 17408
rect 2668 17200 2708 17240
rect 15052 17200 15092 17240
rect 5164 17116 5204 17156
rect 9100 17116 9140 17156
rect 11116 17116 11156 17156
rect 11308 17116 11348 17156
rect 18700 17116 18740 17156
rect 1228 17032 1268 17072
rect 2476 17032 2516 17072
rect 2860 17032 2900 17072
rect 2956 17032 2996 17072
rect 3148 17032 3188 17072
rect 3244 17032 3284 17072
rect 3345 17032 3385 17072
rect 3724 17032 3764 17072
rect 4972 17032 5012 17072
rect 6028 17032 6068 17072
rect 7276 17032 7316 17072
rect 7660 17032 7700 17072
rect 8908 17032 8948 17072
rect 9388 17032 9428 17072
rect 9484 17032 9524 17072
rect 9868 17032 9908 17072
rect 9964 17032 10004 17072
rect 10444 17032 10484 17072
rect 10924 17027 10964 17067
rect 11500 17032 11540 17072
rect 12748 17032 12788 17072
rect 13612 17032 13652 17072
rect 14860 17032 14900 17072
rect 15244 17032 15284 17072
rect 16492 17032 16532 17072
rect 16972 17032 17012 17072
rect 17068 17032 17108 17072
rect 18028 17032 18068 17072
rect 18508 17027 18548 17067
rect 17452 16948 17492 16988
rect 17548 16948 17588 16988
rect 16684 16864 16724 16904
rect 2860 16780 2900 16820
rect 7468 16780 7508 16820
rect 15052 16780 15092 16820
rect 3688 16612 3728 16652
rect 3770 16612 3810 16652
rect 3852 16612 3892 16652
rect 3934 16612 3974 16652
rect 4016 16612 4056 16652
rect 18808 16612 18848 16652
rect 18890 16612 18930 16652
rect 18972 16612 19012 16652
rect 19054 16612 19094 16652
rect 19136 16612 19176 16652
rect 2668 16444 2708 16484
rect 5548 16360 5588 16400
rect 14668 16360 14708 16400
rect 3052 16263 3092 16303
rect 6412 16276 6452 16316
rect 1228 16192 1268 16232
rect 2476 16192 2516 16232
rect 3244 16192 3284 16232
rect 3340 16192 3380 16232
rect 3532 16192 3572 16232
rect 4108 16192 4148 16232
rect 5356 16192 5396 16232
rect 5836 16211 5876 16251
rect 5932 16192 5972 16232
rect 7420 16234 7460 16274
rect 9868 16276 9908 16316
rect 6316 16192 6356 16232
rect 6892 16192 6932 16232
rect 9292 16192 9332 16232
rect 9388 16192 9428 16232
rect 9772 16192 9812 16232
rect 10348 16192 10388 16232
rect 10876 16201 10916 16241
rect 12460 16192 12500 16232
rect 13708 16192 13748 16232
rect 14476 16192 14516 16232
rect 14668 16192 14708 16232
rect 14764 16192 14804 16232
rect 14956 16192 14996 16232
rect 16204 16192 16244 16232
rect 16684 16192 16724 16232
rect 16780 16192 16820 16232
rect 17164 16192 17204 16232
rect 17260 16192 17300 16232
rect 17740 16192 17780 16232
rect 18220 16197 18260 16237
rect 16396 16108 16436 16148
rect 18412 16108 18452 16148
rect 2860 16024 2900 16064
rect 3436 16024 3476 16064
rect 7564 16024 7604 16064
rect 11020 16024 11060 16064
rect 13900 16024 13940 16064
rect 4928 15856 4968 15896
rect 5010 15856 5050 15896
rect 5092 15856 5132 15896
rect 5174 15856 5214 15896
rect 5256 15856 5296 15896
rect 20048 15856 20088 15896
rect 20130 15856 20170 15896
rect 20212 15856 20252 15896
rect 20294 15856 20334 15896
rect 20376 15856 20416 15896
rect 14092 15688 14132 15728
rect 18028 15688 18068 15728
rect 8716 15604 8756 15644
rect 1804 15562 1844 15602
rect 12076 15604 12116 15644
rect 3052 15520 3092 15560
rect 3436 15516 3476 15556
rect 3532 15520 3572 15560
rect 3724 15520 3764 15560
rect 3820 15520 3860 15560
rect 3975 15520 4015 15560
rect 5260 15520 5300 15560
rect 6508 15520 6548 15560
rect 6988 15520 7028 15560
rect 7084 15520 7124 15560
rect 7468 15520 7508 15560
rect 8044 15520 8084 15560
rect 10636 15520 10676 15560
rect 11884 15520 11924 15560
rect 12364 15520 12404 15560
rect 1612 15436 1652 15476
rect 4396 15436 4436 15476
rect 7564 15436 7604 15476
rect 8572 15478 8612 15518
rect 12460 15520 12500 15560
rect 13420 15520 13460 15560
rect 13900 15515 13940 15555
rect 14284 15520 14324 15560
rect 15532 15520 15572 15560
rect 16588 15520 16628 15560
rect 17836 15520 17876 15560
rect 12844 15436 12884 15476
rect 12940 15436 12980 15476
rect 1420 15352 1460 15392
rect 6700 15352 6740 15392
rect 3244 15268 3284 15308
rect 3436 15268 3476 15308
rect 4204 15268 4244 15308
rect 15724 15268 15764 15308
rect 3688 15100 3728 15140
rect 3770 15100 3810 15140
rect 3852 15100 3892 15140
rect 3934 15100 3974 15140
rect 4016 15100 4056 15140
rect 18808 15100 18848 15140
rect 18890 15100 18930 15140
rect 18972 15100 19012 15140
rect 19054 15100 19094 15140
rect 19136 15100 19176 15140
rect 1420 14932 1460 14972
rect 3244 14932 3284 14972
rect 9484 14932 9524 14972
rect 11212 14932 11252 14972
rect 7660 14848 7700 14888
rect 1612 14764 1652 14804
rect 4588 14764 4628 14804
rect 4684 14764 4724 14804
rect 7852 14764 7892 14804
rect 13996 14764 14036 14804
rect 17548 14764 17588 14804
rect 1804 14680 1844 14720
rect 3052 14680 3092 14720
rect 3436 14680 3476 14720
rect 3532 14680 3572 14720
rect 4108 14680 4148 14720
rect 4204 14680 4244 14720
rect 5164 14680 5204 14720
rect 5644 14685 5684 14725
rect 8044 14680 8084 14720
rect 9292 14680 9332 14720
rect 9772 14680 9812 14720
rect 11020 14680 11060 14720
rect 11788 14680 11828 14720
rect 13036 14680 13076 14720
rect 13516 14680 13556 14720
rect 13612 14680 13652 14720
rect 14092 14680 14132 14720
rect 14572 14680 14612 14720
rect 15052 14694 15092 14734
rect 17068 14680 17108 14720
rect 17164 14680 17204 14720
rect 17644 14680 17684 14720
rect 18124 14680 18164 14720
rect 18604 14685 18644 14725
rect 5836 14596 5876 14636
rect 13228 14596 13268 14636
rect 15244 14596 15284 14636
rect 3724 14512 3764 14552
rect 18796 14512 18836 14552
rect 4928 14344 4968 14384
rect 5010 14344 5050 14384
rect 5092 14344 5132 14384
rect 5174 14344 5214 14384
rect 5256 14344 5296 14384
rect 20048 14344 20088 14384
rect 20130 14344 20170 14384
rect 20212 14344 20252 14384
rect 20294 14344 20334 14384
rect 20376 14344 20416 14384
rect 1324 14176 1364 14216
rect 4012 14176 4052 14216
rect 5644 14176 5684 14216
rect 8812 14176 8852 14216
rect 17356 14176 17396 14216
rect 19180 14176 19220 14216
rect 11116 14092 11156 14132
rect 15340 14092 15380 14132
rect 2092 14008 2132 14048
rect 2284 14008 2324 14048
rect 2380 14008 2420 14048
rect 2572 14008 2612 14048
rect 3820 14008 3860 14048
rect 5452 14008 5492 14048
rect 7372 14008 7412 14048
rect 8620 14008 8660 14048
rect 9388 14008 9428 14048
rect 4204 13966 4244 14006
rect 9484 14008 9524 14048
rect 9868 14008 9908 14048
rect 9964 14008 10004 14048
rect 10444 14008 10484 14048
rect 11884 14008 11924 14048
rect 13132 14008 13172 14048
rect 13900 14008 13940 14048
rect 15148 14008 15188 14048
rect 15628 14008 15668 14048
rect 10972 13966 11012 14006
rect 15724 14008 15764 14048
rect 16108 14008 16148 14048
rect 16684 14008 16724 14048
rect 17212 13998 17252 14038
rect 17740 14008 17780 14048
rect 18988 14008 19028 14048
rect 1516 13924 1556 13964
rect 1900 13924 1940 13964
rect 16204 13924 16244 13964
rect 2188 13840 2228 13880
rect 1708 13756 1748 13796
rect 13324 13756 13364 13796
rect 3688 13588 3728 13628
rect 3770 13588 3810 13628
rect 3852 13588 3892 13628
rect 3934 13588 3974 13628
rect 4016 13588 4056 13628
rect 18808 13588 18848 13628
rect 18890 13588 18930 13628
rect 18972 13588 19012 13628
rect 19054 13588 19094 13628
rect 19136 13588 19176 13628
rect 2668 13420 2708 13460
rect 11212 13420 11252 13460
rect 17356 13420 17396 13460
rect 5068 13252 5108 13292
rect 8044 13252 8084 13292
rect 13804 13252 13844 13292
rect 13900 13252 13940 13292
rect 1228 13168 1268 13208
rect 2476 13168 2516 13208
rect 2860 13168 2900 13208
rect 4108 13168 4148 13208
rect 4588 13168 4628 13208
rect 4684 13168 4724 13208
rect 5164 13168 5204 13208
rect 5644 13168 5684 13208
rect 6124 13173 6164 13213
rect 6988 13173 7028 13213
rect 7468 13168 7508 13208
rect 7948 13168 7988 13208
rect 8428 13168 8468 13208
rect 8524 13168 8564 13208
rect 9772 13168 9812 13208
rect 11020 13189 11060 13229
rect 13324 13168 13364 13208
rect 13420 13168 13460 13208
rect 14380 13168 14420 13208
rect 14908 13177 14948 13217
rect 15916 13168 15956 13208
rect 17164 13168 17204 13208
rect 4300 13084 4340 13124
rect 6796 13084 6836 13124
rect 6316 13000 6356 13040
rect 15052 13000 15092 13040
rect 4928 12832 4968 12872
rect 5010 12832 5050 12872
rect 5092 12832 5132 12872
rect 5174 12832 5214 12872
rect 5256 12832 5296 12872
rect 20048 12832 20088 12872
rect 20130 12832 20170 12872
rect 20212 12832 20252 12872
rect 20294 12832 20334 12872
rect 20376 12832 20416 12872
rect 2668 12664 2708 12704
rect 3916 12664 3956 12704
rect 6028 12664 6068 12704
rect 7660 12580 7700 12620
rect 9292 12580 9332 12620
rect 12940 12580 12980 12620
rect 15148 12580 15188 12620
rect 17452 12580 17492 12620
rect 1228 12496 1268 12536
rect 2476 12496 2516 12536
rect 2860 12496 2900 12536
rect 2956 12496 2996 12536
rect 3148 12496 3188 12536
rect 3244 12496 3284 12536
rect 3345 12496 3385 12536
rect 3628 12496 3668 12536
rect 3724 12496 3764 12536
rect 4588 12496 4628 12536
rect 5836 12496 5876 12536
rect 6220 12496 6260 12536
rect 7468 12496 7508 12536
rect 7852 12496 7892 12536
rect 9100 12496 9140 12536
rect 9484 12496 9524 12536
rect 10732 12496 10772 12536
rect 11212 12496 11252 12536
rect 11308 12496 11348 12536
rect 12268 12496 12308 12536
rect 12748 12482 12788 12522
rect 13708 12496 13748 12536
rect 14956 12496 14996 12536
rect 16012 12496 16052 12536
rect 17260 12496 17300 12536
rect 18316 12496 18356 12536
rect 19564 12496 19604 12536
rect 11692 12412 11732 12452
rect 11788 12412 11828 12452
rect 17836 12412 17876 12452
rect 17644 12328 17684 12368
rect 2860 12244 2900 12284
rect 10924 12244 10964 12284
rect 18124 12244 18164 12284
rect 3688 12076 3728 12116
rect 3770 12076 3810 12116
rect 3852 12076 3892 12116
rect 3934 12076 3974 12116
rect 4016 12076 4056 12116
rect 18808 12076 18848 12116
rect 18890 12076 18930 12116
rect 18972 12076 19012 12116
rect 19054 12076 19094 12116
rect 19136 12076 19176 12116
rect 1804 11908 1844 11948
rect 7276 11908 7316 11948
rect 7468 11908 7508 11948
rect 12652 11908 12692 11948
rect 1612 11740 1652 11780
rect 1996 11740 2036 11780
rect 4396 11740 4436 11780
rect 4492 11740 4532 11780
rect 7660 11740 7700 11780
rect 8812 11740 8852 11780
rect 2188 11656 2228 11696
rect 3436 11656 3476 11696
rect 3916 11656 3956 11696
rect 4012 11656 4052 11696
rect 4972 11656 5012 11696
rect 5500 11665 5540 11705
rect 5836 11698 5876 11738
rect 8908 11740 8948 11780
rect 10732 11740 10772 11780
rect 13612 11740 13652 11780
rect 13708 11740 13748 11780
rect 16396 11740 16436 11780
rect 16492 11740 16532 11780
rect 7084 11656 7124 11696
rect 8332 11656 8372 11696
rect 8428 11656 8468 11696
rect 9388 11656 9428 11696
rect 9868 11661 9908 11701
rect 11212 11656 11252 11696
rect 12460 11656 12500 11696
rect 13132 11656 13172 11696
rect 13228 11656 13268 11696
rect 14188 11656 14228 11696
rect 14716 11665 14756 11705
rect 15916 11656 15956 11696
rect 16012 11656 16052 11696
rect 16972 11656 17012 11696
rect 17452 11661 17492 11701
rect 18028 11656 18068 11696
rect 19276 11656 19316 11696
rect 3628 11572 3668 11612
rect 1420 11488 1460 11528
rect 5644 11530 5684 11570
rect 17836 11572 17876 11612
rect 10060 11488 10100 11528
rect 10540 11488 10580 11528
rect 14860 11488 14900 11528
rect 17644 11488 17684 11528
rect 4928 11320 4968 11360
rect 5010 11320 5050 11360
rect 5092 11320 5132 11360
rect 5174 11320 5214 11360
rect 5256 11320 5296 11360
rect 20048 11320 20088 11360
rect 20130 11320 20170 11360
rect 20212 11320 20252 11360
rect 20294 11320 20334 11360
rect 20376 11320 20416 11360
rect 1708 11152 1748 11192
rect 5740 11152 5780 11192
rect 10156 11152 10196 11192
rect 10636 11152 10676 11192
rect 13132 11152 13172 11192
rect 14860 11152 14900 11192
rect 16492 11152 16532 11192
rect 7756 11068 7796 11108
rect 17740 11068 17780 11108
rect 2092 10984 2132 11024
rect 3340 10984 3380 11024
rect 4300 10984 4340 11024
rect 5548 10984 5588 11024
rect 6028 10984 6068 11024
rect 6124 10984 6164 11024
rect 6508 10984 6548 11024
rect 7084 10984 7124 11024
rect 8716 10984 8756 11024
rect 9964 10984 10004 11024
rect 10348 10984 10388 11024
rect 1526 10889 1566 10929
rect 1900 10900 1940 10940
rect 6604 10900 6644 10940
rect 7612 10942 7652 10982
rect 10444 10984 10484 11024
rect 11692 10984 11732 11024
rect 12940 10984 12980 11024
rect 13420 10984 13460 11024
rect 14668 10984 14708 11024
rect 15052 10984 15092 11024
rect 16300 10984 16340 11024
rect 17932 10979 17972 11019
rect 18412 10984 18452 11024
rect 18988 10984 19028 11024
rect 19372 10984 19412 11024
rect 19468 10984 19508 11024
rect 8140 10900 8180 10940
rect 18892 10900 18932 10940
rect 1324 10732 1364 10772
rect 3532 10732 3572 10772
rect 7948 10732 7988 10772
rect 3688 10564 3728 10604
rect 3770 10564 3810 10604
rect 3852 10564 3892 10604
rect 3934 10564 3974 10604
rect 4016 10564 4056 10604
rect 18808 10564 18848 10604
rect 18890 10564 18930 10604
rect 18972 10564 19012 10604
rect 19054 10564 19094 10604
rect 19136 10564 19176 10604
rect 1420 10396 1460 10436
rect 6124 10396 6164 10436
rect 8524 10396 8564 10436
rect 18700 10396 18740 10436
rect 3244 10312 3284 10352
rect 10540 10312 10580 10352
rect 1612 10228 1652 10268
rect 11884 10228 11924 10268
rect 13708 10228 13748 10268
rect 15820 10228 15860 10268
rect 1804 10144 1844 10184
rect 3052 10144 3092 10184
rect 3436 10144 3476 10184
rect 3532 10144 3572 10184
rect 3724 10144 3764 10184
rect 3820 10144 3860 10184
rect 3977 10159 4017 10199
rect 4204 10144 4244 10184
rect 4300 10144 4340 10184
rect 4684 10144 4724 10184
rect 5932 10144 5972 10184
rect 7084 10144 7124 10184
rect 8332 10144 8372 10184
rect 9100 10144 9140 10184
rect 10348 10144 10388 10184
rect 10876 10153 10916 10193
rect 11404 10144 11444 10184
rect 11980 10144 12020 10184
rect 12364 10144 12404 10184
rect 12460 10144 12500 10184
rect 13228 10144 13268 10184
rect 13324 10144 13364 10184
rect 13804 10144 13844 10184
rect 14284 10144 14324 10184
rect 14812 10153 14852 10193
rect 15340 10144 15380 10184
rect 15436 10144 15476 10184
rect 15916 10144 15956 10184
rect 16396 10144 16436 10184
rect 16924 10153 16964 10193
rect 17260 10144 17300 10184
rect 18508 10144 18548 10184
rect 3628 9976 3668 10016
rect 4492 9976 4532 10016
rect 10732 9976 10772 10016
rect 14956 9976 14996 10016
rect 17068 10018 17108 10058
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 1900 9640 1940 9680
rect 2284 9640 2324 9680
rect 3340 9640 3380 9680
rect 7756 9640 7796 9680
rect 10348 9640 10388 9680
rect 13420 9640 13460 9680
rect 15052 9640 15092 9680
rect 17260 9640 17300 9680
rect 2764 9472 2804 9512
rect 2860 9472 2900 9512
rect 3052 9472 3092 9512
rect 3244 9472 3284 9512
rect 3436 9472 3476 9512
rect 3532 9472 3572 9512
rect 4108 9472 4148 9512
rect 4300 9472 4340 9512
rect 4396 9472 4436 9512
rect 4588 9472 4628 9512
rect 4684 9472 4724 9512
rect 4876 9472 4916 9512
rect 4972 9472 5012 9512
rect 5073 9472 5113 9512
rect 6316 9472 6356 9512
rect 7564 9472 7604 9512
rect 7948 9472 7988 9512
rect 8140 9472 8180 9512
rect 8236 9472 8276 9512
rect 8620 9472 8660 9512
rect 9868 9472 9908 9512
rect 10540 9472 10580 9512
rect 11788 9472 11828 9512
rect 13228 9472 13268 9512
rect 13612 9472 13652 9512
rect 14860 9472 14900 9512
rect 15820 9472 15860 9512
rect 17068 9472 17108 9512
rect 17740 9472 17780 9512
rect 18988 9472 19028 9512
rect 11980 9430 12020 9470
rect 1708 9388 1748 9428
rect 2092 9388 2132 9428
rect 2476 9388 2516 9428
rect 2956 9304 2996 9344
rect 4396 9304 4436 9344
rect 8236 9304 8276 9344
rect 1516 9220 1556 9260
rect 4588 9220 4628 9260
rect 8428 9220 8468 9260
rect 19180 9220 19220 9260
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 3724 8800 3764 8840
rect 8332 8800 8372 8840
rect 15628 8800 15668 8840
rect 1708 8716 1748 8756
rect 2092 8716 2132 8756
rect 3916 8716 3956 8756
rect 6988 8716 7028 8756
rect 17932 8716 17972 8756
rect 18028 8716 18068 8756
rect 2668 8632 2708 8672
rect 2764 8632 2804 8672
rect 2956 8632 2996 8672
rect 3052 8632 3092 8672
rect 3244 8632 3284 8672
rect 3340 8632 3380 8672
rect 3468 8632 3508 8672
rect 4108 8632 4148 8672
rect 5356 8632 5396 8672
rect 5932 8637 5972 8677
rect 6412 8632 6452 8672
rect 6892 8632 6932 8672
rect 7372 8632 7412 8672
rect 7468 8632 7508 8672
rect 8524 8632 8564 8672
rect 9772 8632 9812 8672
rect 9964 8632 10004 8672
rect 10060 8632 10100 8672
rect 10252 8632 10292 8672
rect 10348 8632 10388 8672
rect 10505 8647 10545 8687
rect 10828 8632 10868 8672
rect 10924 8632 10964 8672
rect 11308 8632 11348 8672
rect 11404 8632 11444 8672
rect 11884 8632 11924 8672
rect 12412 8641 12452 8681
rect 14188 8632 14228 8672
rect 15436 8632 15476 8672
rect 17452 8632 17492 8672
rect 17548 8632 17588 8672
rect 18508 8632 18548 8672
rect 19036 8641 19076 8681
rect 5548 8548 5588 8588
rect 12556 8548 12596 8588
rect 1516 8464 1556 8504
rect 1900 8464 1940 8504
rect 2476 8464 2516 8504
rect 3436 8464 3476 8504
rect 5740 8464 5780 8504
rect 10156 8464 10196 8504
rect 19180 8464 19220 8504
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 1228 8128 1268 8168
rect 3052 8128 3092 8168
rect 5068 8128 5108 8168
rect 6700 8128 6740 8168
rect 10636 8128 10676 8168
rect 12460 8128 12500 8168
rect 14572 8128 14612 8168
rect 16780 8128 16820 8168
rect 16972 8128 17012 8168
rect 8716 8044 8756 8084
rect 1612 7960 1652 8000
rect 2860 7960 2900 8000
rect 3628 7960 3668 8000
rect 4876 7960 4916 8000
rect 5260 7960 5300 8000
rect 6508 7960 6548 8000
rect 6988 7960 7028 8000
rect 7084 7960 7124 8000
rect 7468 7960 7508 8000
rect 7564 7960 7604 8000
rect 8044 7960 8084 8000
rect 9196 7960 9236 8000
rect 10444 7960 10484 8000
rect 11020 7960 11060 8000
rect 12268 7960 12308 8000
rect 12844 7960 12884 8000
rect 8572 7918 8612 7958
rect 12940 7960 12980 8000
rect 13900 7960 13940 8000
rect 1420 7876 1460 7916
rect 3436 7876 3476 7916
rect 13324 7876 13364 7916
rect 13420 7876 13460 7916
rect 14428 7918 14468 7958
rect 15052 7960 15092 8000
rect 15148 7960 15188 8000
rect 16108 7960 16148 8000
rect 17164 7960 17204 8000
rect 18412 7960 18452 8000
rect 15532 7876 15572 7916
rect 15628 7876 15668 7916
rect 16636 7918 16676 7958
rect 18796 7876 18836 7916
rect 3244 7792 3284 7832
rect 18604 7708 18644 7748
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 2956 7372 2996 7412
rect 7180 7372 7220 7412
rect 8812 7372 8852 7412
rect 12940 7372 12980 7412
rect 14572 7372 14612 7412
rect 14764 7372 14804 7412
rect 10636 7288 10676 7328
rect 3340 7204 3380 7244
rect 1516 7120 1556 7160
rect 2764 7120 2804 7160
rect 3532 7120 3572 7160
rect 4780 7120 4820 7160
rect 5164 7120 5204 7160
rect 5260 7120 5300 7160
rect 5740 7120 5780 7160
rect 6988 7120 7028 7160
rect 7372 7120 7412 7160
rect 8620 7120 8660 7160
rect 9196 7120 9236 7160
rect 10444 7120 10484 7160
rect 10835 7125 10875 7165
rect 10931 7116 10971 7156
rect 11123 7125 11163 7165
rect 11500 7120 11540 7160
rect 12748 7120 12788 7160
rect 13132 7120 13172 7160
rect 14380 7120 14420 7160
rect 14956 7120 14996 7160
rect 16204 7120 16244 7160
rect 3148 6952 3188 6992
rect 4972 6952 5012 6992
rect 5452 6952 5492 6992
rect 11020 6952 11060 6992
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 1324 6616 1364 6656
rect 1708 6616 1748 6656
rect 4300 6616 4340 6656
rect 6796 6616 6836 6656
rect 8716 6616 8756 6656
rect 11692 6616 11732 6656
rect 14284 6616 14324 6656
rect 16876 6616 16916 6656
rect 2188 6532 2228 6572
rect 9196 6532 9236 6572
rect 2092 6448 2132 6488
rect 2284 6448 2324 6488
rect 2380 6448 2420 6488
rect 2572 6448 2612 6488
rect 2668 6448 2708 6488
rect 2860 6448 2900 6488
rect 2956 6448 2996 6488
rect 3057 6448 3097 6488
rect 3628 6448 3668 6488
rect 3820 6448 3860 6488
rect 3916 6448 3956 6488
rect 4108 6448 4148 6488
rect 4204 6448 4244 6488
rect 4396 6448 4436 6488
rect 4492 6448 4532 6488
rect 4593 6448 4633 6488
rect 4876 6448 4916 6488
rect 6124 6448 6164 6488
rect 6508 6448 6548 6488
rect 6604 6448 6644 6488
rect 6988 6448 7028 6488
rect 8236 6448 8276 6488
rect 8908 6448 8948 6488
rect 9004 6448 9044 6488
rect 9388 6448 9428 6488
rect 10636 6448 10676 6488
rect 10828 6448 10868 6488
rect 10924 6448 10964 6488
rect 11116 6448 11156 6488
rect 11212 6448 11252 6488
rect 11369 6441 11409 6481
rect 11630 6433 11670 6473
rect 11788 6448 11828 6488
rect 11884 6448 11924 6488
rect 12076 6448 12116 6488
rect 12172 6448 12212 6488
rect 12556 6448 12596 6488
rect 12652 6448 12692 6488
rect 13132 6448 13172 6488
rect 13612 6448 13652 6488
rect 14140 6438 14180 6478
rect 15436 6448 15476 6488
rect 16684 6448 16724 6488
rect 17164 6448 17204 6488
rect 18412 6448 18452 6488
rect 1516 6364 1556 6404
rect 1900 6364 1940 6404
rect 13036 6364 13076 6404
rect 3916 6280 3956 6320
rect 2572 6196 2612 6236
rect 6316 6196 6356 6236
rect 8428 6196 8468 6236
rect 10828 6196 10868 6236
rect 18604 6196 18644 6236
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 4588 5860 4628 5900
rect 6220 5860 6260 5900
rect 12748 5860 12788 5900
rect 14380 5860 14420 5900
rect 2860 5776 2900 5816
rect 6988 5692 7028 5732
rect 7084 5692 7124 5732
rect 17644 5692 17684 5732
rect 17740 5692 17780 5732
rect 1420 5608 1460 5648
rect 2668 5608 2708 5648
rect 3148 5608 3188 5648
rect 4396 5608 4436 5648
rect 4780 5608 4820 5648
rect 6028 5608 6068 5648
rect 6508 5608 6548 5648
rect 6604 5608 6644 5648
rect 7564 5608 7604 5648
rect 8044 5622 8084 5662
rect 8524 5608 8564 5648
rect 9772 5608 9812 5648
rect 10156 5608 10196 5648
rect 10252 5608 10292 5648
rect 10444 5608 10484 5648
rect 10540 5608 10580 5648
rect 10697 5623 10737 5663
rect 11308 5608 11348 5648
rect 12556 5608 12596 5648
rect 12940 5608 12980 5648
rect 14188 5608 14228 5648
rect 15148 5608 15188 5648
rect 15244 5608 15284 5648
rect 15628 5608 15668 5648
rect 15724 5608 15764 5648
rect 16204 5608 16244 5648
rect 16732 5617 16772 5657
rect 17164 5608 17204 5648
rect 17260 5608 17300 5648
rect 18220 5608 18260 5648
rect 18700 5622 18740 5662
rect 16876 5524 16916 5564
rect 6220 5440 6260 5480
rect 8236 5440 8276 5480
rect 9964 5440 10004 5480
rect 10636 5440 10676 5480
rect 18892 5440 18932 5480
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 2860 5104 2900 5144
rect 5356 5104 5396 5144
rect 10348 5104 10388 5144
rect 12268 5104 12308 5144
rect 15244 5104 15284 5144
rect 16972 5104 17012 5144
rect 4876 5020 4916 5060
rect 7180 5020 7220 5060
rect 9868 5020 9908 5060
rect 12940 5020 12980 5060
rect 1420 4936 1460 4976
rect 2668 4936 2708 4976
rect 3436 4936 3476 4976
rect 5068 4936 5108 4976
rect 4684 4894 4724 4934
rect 5164 4936 5204 4976
rect 5740 4936 5780 4976
rect 6988 4936 7028 4976
rect 7372 4936 7412 4976
rect 7468 4936 7508 4976
rect 7660 4936 7700 4976
rect 7756 4936 7796 4976
rect 7857 4936 7897 4976
rect 8428 4936 8468 4976
rect 9676 4936 9716 4976
rect 10060 4936 10100 4976
rect 10156 4936 10196 4976
rect 10636 4936 10676 4976
rect 11884 4936 11924 4976
rect 12460 4936 12500 4976
rect 12556 4936 12596 4976
rect 12748 4936 12788 4976
rect 12844 4936 12884 4976
rect 13036 4936 13076 4976
rect 13804 4936 13844 4976
rect 15052 4936 15092 4976
rect 15532 4936 15572 4976
rect 16780 4936 16820 4976
rect 3244 4852 3284 4892
rect 3052 4768 3092 4808
rect 12076 4768 12116 4808
rect 7372 4684 7412 4724
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 1516 4348 1556 4388
rect 1900 4348 1940 4388
rect 2284 4348 2324 4388
rect 12172 4348 12212 4388
rect 9772 4264 9812 4304
rect 1708 4180 1748 4220
rect 2092 4180 2132 4220
rect 2476 4180 2516 4220
rect 3052 4096 3092 4136
rect 3148 4096 3188 4136
rect 3628 4096 3668 4136
rect 4876 4096 4916 4136
rect 5740 4096 5780 4136
rect 5836 4096 5876 4136
rect 6892 4096 6932 4136
rect 7084 4096 7124 4136
rect 7180 4096 7220 4136
rect 7372 4096 7412 4136
rect 7468 4096 7508 4136
rect 7660 4096 7700 4136
rect 7756 4096 7796 4136
rect 7884 4096 7924 4136
rect 9580 4096 9620 4136
rect 9772 4096 9812 4136
rect 9868 4096 9908 4136
rect 10348 4096 10388 4136
rect 10444 4096 10484 4136
rect 10732 4096 10772 4136
rect 11980 4096 12020 4136
rect 12940 4096 12980 4136
rect 14188 4096 14228 4136
rect 14668 4096 14708 4136
rect 14764 4096 14804 4136
rect 15148 4096 15188 4136
rect 15244 4096 15284 4136
rect 15724 4096 15764 4136
rect 16252 4105 16292 4145
rect 14380 4012 14420 4052
rect 16396 4012 16436 4052
rect 2860 3928 2900 3968
rect 5068 3928 5108 3968
rect 5548 3928 5588 3968
rect 6988 3928 7028 3968
rect 7564 3928 7604 3968
rect 10156 3928 10196 3968
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 1516 3592 1556 3632
rect 1900 3592 1940 3632
rect 2284 3592 2324 3632
rect 2668 3592 2708 3632
rect 7852 3592 7892 3632
rect 8332 3592 8372 3632
rect 16876 3592 16916 3632
rect 5260 3508 5300 3548
rect 12556 3508 12596 3548
rect 14572 3508 14612 3548
rect 3628 3424 3668 3464
rect 4876 3424 4916 3464
rect 5260 3401 5300 3441
rect 5356 3424 5396 3464
rect 5548 3424 5588 3464
rect 5644 3424 5684 3464
rect 5772 3421 5812 3461
rect 6412 3424 6452 3464
rect 7660 3424 7700 3464
rect 8044 3424 8084 3464
rect 8140 3424 8180 3464
rect 8620 3424 8660 3464
rect 9868 3424 9908 3464
rect 10252 3424 10292 3464
rect 10540 3424 10580 3464
rect 10732 3424 10772 3464
rect 10924 3424 10964 3464
rect 11116 3424 11156 3464
rect 12364 3424 12404 3464
rect 12844 3424 12884 3464
rect 12940 3424 12980 3464
rect 13324 3424 13364 3464
rect 13420 3424 13460 3464
rect 13900 3424 13940 3464
rect 14380 3410 14420 3450
rect 15436 3424 15476 3464
rect 16684 3424 16724 3464
rect 1708 3340 1748 3380
rect 2092 3340 2132 3380
rect 2476 3340 2516 3380
rect 2860 3340 2900 3380
rect 3244 3340 3284 3380
rect 10540 3256 10580 3296
rect 10828 3256 10868 3296
rect 3052 3172 3092 3212
rect 5068 3172 5108 3212
rect 7852 3172 7892 3212
rect 10060 3172 10100 3212
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 1516 2836 1556 2876
rect 1900 2836 1940 2876
rect 4972 2836 5012 2876
rect 5164 2836 5204 2876
rect 7756 2836 7796 2876
rect 14380 2836 14420 2876
rect 16300 2836 16340 2876
rect 9580 2752 9620 2792
rect 10540 2752 10580 2792
rect 1708 2668 1748 2708
rect 2092 2668 2132 2708
rect 2572 2668 2612 2708
rect 10828 2668 10868 2708
rect 11308 2668 11348 2708
rect 3532 2584 3572 2624
rect 4780 2584 4820 2624
rect 5164 2607 5204 2647
rect 5260 2584 5300 2624
rect 5452 2584 5492 2624
rect 5548 2584 5588 2624
rect 5705 2599 5745 2639
rect 6316 2584 6356 2624
rect 7564 2584 7604 2624
rect 8140 2584 8180 2624
rect 9388 2584 9428 2624
rect 9868 2584 9908 2624
rect 10156 2584 10196 2624
rect 10732 2584 10772 2624
rect 10924 2597 10964 2637
rect 12940 2584 12980 2624
rect 14188 2584 14228 2624
rect 14860 2584 14900 2624
rect 16108 2584 16148 2624
rect 10252 2500 10292 2540
rect 2380 2416 2420 2456
rect 11116 2416 11156 2456
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 1900 2080 1940 2120
rect 5356 2080 5396 2120
rect 5932 2080 5972 2120
rect 6604 2080 6644 2120
rect 6988 2080 7028 2120
rect 7468 2080 7508 2120
rect 9676 2080 9716 2120
rect 10156 2080 10196 2120
rect 3532 1912 3572 1952
rect 4780 1912 4820 1952
rect 5164 1912 5204 1952
rect 5260 1912 5300 1952
rect 5452 1912 5492 1952
rect 5644 1912 5684 1952
rect 5740 1912 5780 1952
rect 7372 1912 7412 1952
rect 7564 1912 7604 1952
rect 7660 1912 7700 1952
rect 9388 1912 9428 1952
rect 9484 1912 9524 1952
rect 9868 1912 9908 1952
rect 9964 1912 10004 1952
rect 10156 1912 10196 1952
rect 1708 1828 1748 1868
rect 2092 1828 2132 1868
rect 2476 1828 2516 1868
rect 2860 1828 2900 1868
rect 3148 1828 3188 1868
rect 6412 1828 6452 1868
rect 6796 1817 6836 1857
rect 7180 1828 7220 1868
rect 7852 1828 7892 1868
rect 8236 1828 8276 1868
rect 8620 1828 8660 1868
rect 9004 1828 9044 1868
rect 10540 1828 10580 1868
rect 10924 1828 10964 1868
rect 11308 1828 11348 1868
rect 11884 1828 11924 1868
rect 12268 1828 12308 1868
rect 12940 1828 12980 1868
rect 13228 1828 13268 1868
rect 13900 1828 13940 1868
rect 14284 1828 14324 1868
rect 14668 1828 14708 1868
rect 15244 1828 15284 1868
rect 15628 1828 15668 1868
rect 16012 1828 16052 1868
rect 16396 1828 16436 1868
rect 1516 1744 1556 1784
rect 4972 1744 5012 1784
rect 2284 1660 2324 1700
rect 2668 1660 2708 1700
rect 3340 1660 3380 1700
rect 6220 1660 6260 1700
rect 8044 1660 8084 1700
rect 8428 1660 8468 1700
rect 8812 1660 8852 1700
rect 9196 1660 9236 1700
rect 10732 1660 10772 1700
rect 11116 1660 11156 1700
rect 11500 1660 11540 1700
rect 11692 1660 11732 1700
rect 12076 1660 12116 1700
rect 12748 1660 12788 1700
rect 13420 1660 13460 1700
rect 14092 1660 14132 1700
rect 14476 1660 14516 1700
rect 14860 1660 14900 1700
rect 15052 1660 15092 1700
rect 15436 1660 15476 1700
rect 15820 1660 15860 1700
rect 16204 1660 16244 1700
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 5356 1240 5396 1280
rect 6700 1240 6740 1280
rect 7372 1240 7412 1280
rect 7756 1240 7796 1280
rect 1708 1156 1748 1196
rect 2092 1156 2132 1196
rect 2476 1156 2516 1196
rect 6124 1156 6164 1196
rect 6508 1156 6548 1196
rect 6892 1156 6932 1196
rect 7564 1156 7604 1196
rect 7948 1156 7988 1196
rect 9004 1156 9044 1196
rect 9388 1156 9428 1196
rect 9772 1156 9812 1196
rect 10156 1156 10196 1196
rect 10540 1156 10580 1196
rect 10924 1156 10964 1196
rect 15148 1156 15188 1196
rect 16012 1156 16052 1196
rect 5164 1072 5204 1112
rect 5260 1072 5300 1112
rect 5452 1072 5492 1112
rect 1516 904 1556 944
rect 1900 904 1940 944
rect 2284 904 2324 944
rect 5932 904 5972 944
rect 6316 904 6356 944
rect 9196 904 9236 944
rect 9580 904 9620 944
rect 9964 904 10004 944
rect 10348 904 10388 944
rect 10732 904 10772 944
rect 11116 904 11156 944
rect 14956 904 14996 944
rect 15820 904 15860 944
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
<< metal2 >>
rect 1784 85936 1864 86016
rect 1976 85936 2056 86016
rect 2168 85952 2248 86016
rect 2168 85936 2188 85952
rect 267 85784 309 85793
rect 267 85744 268 85784
rect 308 85744 309 85784
rect 267 85735 309 85744
rect 75 83768 117 83777
rect 75 83728 76 83768
rect 116 83728 117 83768
rect 75 83719 117 83728
rect 76 77552 116 83719
rect 268 81920 308 85735
rect 1323 84104 1365 84113
rect 1323 84064 1324 84104
rect 1364 84064 1365 84104
rect 1323 84055 1365 84064
rect 1131 82088 1173 82097
rect 1131 82048 1132 82088
rect 1172 82048 1173 82088
rect 1131 82039 1173 82048
rect 1228 82088 1268 82099
rect 268 81880 500 81920
rect 363 79736 405 79745
rect 363 79696 364 79736
rect 404 79696 405 79736
rect 363 79687 405 79696
rect 76 77512 308 77552
rect 171 76376 213 76385
rect 171 76336 172 76376
rect 212 76336 213 76376
rect 171 76327 213 76336
rect 172 65213 212 76327
rect 268 72941 308 77512
rect 267 72932 309 72941
rect 267 72892 268 72932
rect 308 72892 309 72932
rect 267 72883 309 72892
rect 364 72773 404 79687
rect 460 75125 500 81880
rect 459 75116 501 75125
rect 459 75076 460 75116
rect 500 75076 501 75116
rect 459 75067 501 75076
rect 939 75116 981 75125
rect 939 75076 940 75116
rect 980 75076 981 75116
rect 939 75067 981 75076
rect 555 74360 597 74369
rect 555 74320 556 74360
rect 596 74320 597 74360
rect 555 74311 597 74320
rect 363 72764 405 72773
rect 363 72724 364 72764
rect 404 72724 405 72764
rect 363 72715 405 72724
rect 556 67397 596 74311
rect 555 67388 597 67397
rect 555 67348 556 67388
rect 596 67348 597 67388
rect 555 67339 597 67348
rect 940 66977 980 75067
rect 1132 74108 1172 82039
rect 1228 82013 1268 82048
rect 1227 82004 1269 82013
rect 1227 81964 1228 82004
rect 1268 81964 1269 82004
rect 1227 81955 1269 81964
rect 1228 81173 1268 81258
rect 1227 81164 1269 81173
rect 1227 81124 1228 81164
rect 1268 81124 1269 81164
rect 1227 81115 1269 81124
rect 1228 79568 1268 79577
rect 1228 79409 1268 79528
rect 1227 79400 1269 79409
rect 1227 79360 1228 79400
rect 1268 79360 1269 79400
rect 1227 79351 1269 79360
rect 1228 78224 1268 78233
rect 1324 78224 1364 84055
rect 1804 84029 1844 85936
rect 1803 84020 1845 84029
rect 1803 83980 1804 84020
rect 1844 83980 1845 84020
rect 1803 83971 1845 83980
rect 1900 83768 1940 83777
rect 1996 83768 2036 85936
rect 2187 85912 2188 85936
rect 2228 85936 2248 85952
rect 2360 85936 2440 86016
rect 2552 85936 2632 86016
rect 2744 85936 2824 86016
rect 2936 85936 3016 86016
rect 3128 85936 3208 86016
rect 3320 85936 3400 86016
rect 3512 85936 3592 86016
rect 3704 85936 3784 86016
rect 3896 85936 3976 86016
rect 4088 85936 4168 86016
rect 4280 85936 4360 86016
rect 4472 85936 4552 86016
rect 4664 85936 4744 86016
rect 4856 85936 4936 86016
rect 5048 85936 5128 86016
rect 5240 85936 5320 86016
rect 5432 85936 5512 86016
rect 5624 85936 5704 86016
rect 5816 85936 5896 86016
rect 6008 85936 6088 86016
rect 6200 85936 6280 86016
rect 6392 85936 6472 86016
rect 6584 85936 6664 86016
rect 6776 85936 6856 86016
rect 6968 85936 7048 86016
rect 7160 85936 7240 86016
rect 7352 85936 7432 86016
rect 7544 85936 7624 86016
rect 7736 85936 7816 86016
rect 7928 85936 8008 86016
rect 8120 85936 8200 86016
rect 8312 85936 8392 86016
rect 8504 85936 8584 86016
rect 8696 85936 8776 86016
rect 8888 85936 8968 86016
rect 9080 85936 9160 86016
rect 9272 85936 9352 86016
rect 9464 85936 9544 86016
rect 9656 85936 9736 86016
rect 9848 85936 9928 86016
rect 10040 85936 10120 86016
rect 10232 85936 10312 86016
rect 10424 85936 10504 86016
rect 10616 85936 10696 86016
rect 10808 85936 10888 86016
rect 11000 85936 11080 86016
rect 11192 85936 11272 86016
rect 11384 85936 11464 86016
rect 11576 85936 11656 86016
rect 11768 85936 11848 86016
rect 11960 85936 12040 86016
rect 12152 85936 12232 86016
rect 12344 85936 12424 86016
rect 12536 85936 12616 86016
rect 12728 85936 12808 86016
rect 12920 85936 13000 86016
rect 13112 85936 13192 86016
rect 13304 85936 13384 86016
rect 13496 85936 13576 86016
rect 13688 85936 13768 86016
rect 13880 85936 13960 86016
rect 14072 85936 14152 86016
rect 14264 85936 14344 86016
rect 14456 85936 14536 86016
rect 14648 85936 14728 86016
rect 14840 85936 14920 86016
rect 15032 85936 15112 86016
rect 15224 85936 15304 86016
rect 15416 85936 15496 86016
rect 15608 85936 15688 86016
rect 15800 85936 15880 86016
rect 15992 85936 16072 86016
rect 16184 85936 16264 86016
rect 16376 85936 16456 86016
rect 16568 85936 16648 86016
rect 16760 85936 16840 86016
rect 16952 85936 17032 86016
rect 17144 85936 17224 86016
rect 17336 85936 17416 86016
rect 17528 85936 17608 86016
rect 17720 85936 17800 86016
rect 17912 85936 17992 86016
rect 18104 85936 18184 86016
rect 18296 85936 18376 86016
rect 18488 85936 18568 86016
rect 18680 85936 18760 86016
rect 18872 85936 18952 86016
rect 19064 85936 19144 86016
rect 19256 85936 19336 86016
rect 19448 85936 19528 86016
rect 2228 85912 2229 85936
rect 2187 85903 2229 85912
rect 2380 84692 2420 85936
rect 2188 84652 2420 84692
rect 2091 84440 2133 84449
rect 2091 84400 2092 84440
rect 2132 84400 2133 84440
rect 2091 84391 2133 84400
rect 1940 83728 2036 83768
rect 1900 83719 1940 83728
rect 2092 83684 2132 84391
rect 2188 83861 2228 84652
rect 2572 84440 2612 85936
rect 2667 85280 2709 85289
rect 2667 85240 2668 85280
rect 2708 85240 2709 85280
rect 2667 85231 2709 85240
rect 2284 84400 2612 84440
rect 2187 83852 2229 83861
rect 2187 83812 2188 83852
rect 2228 83812 2229 83852
rect 2187 83803 2229 83812
rect 2284 83768 2324 84400
rect 2284 83719 2324 83728
rect 2668 83768 2708 85231
rect 2764 84440 2804 85936
rect 2956 84617 2996 85936
rect 3148 85289 3188 85936
rect 3147 85280 3189 85289
rect 3147 85240 3148 85280
rect 3188 85240 3189 85280
rect 3147 85231 3189 85240
rect 2955 84608 2997 84617
rect 2955 84568 2956 84608
rect 2996 84568 2997 84608
rect 2955 84559 2997 84568
rect 3052 84440 3092 84449
rect 2764 84400 3052 84440
rect 3052 84391 3092 84400
rect 3243 84356 3285 84365
rect 3243 84316 3244 84356
rect 3284 84316 3285 84356
rect 3243 84307 3285 84316
rect 3244 84222 3284 84307
rect 2668 83719 2708 83728
rect 3051 83768 3093 83777
rect 3051 83728 3052 83768
rect 3092 83728 3093 83768
rect 3051 83719 3093 83728
rect 1996 83644 2132 83684
rect 1707 83516 1749 83525
rect 1707 83476 1708 83516
rect 1748 83476 1749 83516
rect 1707 83467 1749 83476
rect 1708 83382 1748 83467
rect 1900 82760 1940 82769
rect 1707 82256 1749 82265
rect 1707 82216 1708 82256
rect 1748 82216 1749 82256
rect 1707 82207 1749 82216
rect 1420 81248 1460 81257
rect 1420 80669 1460 81208
rect 1515 81164 1557 81173
rect 1515 81124 1516 81164
rect 1556 81124 1557 81164
rect 1515 81115 1557 81124
rect 1419 80660 1461 80669
rect 1419 80620 1420 80660
rect 1460 80620 1461 80660
rect 1419 80611 1461 80620
rect 1420 79736 1460 80611
rect 1420 79687 1460 79696
rect 1419 79400 1461 79409
rect 1419 79360 1420 79400
rect 1460 79360 1461 79400
rect 1419 79351 1461 79360
rect 1268 78184 1364 78224
rect 1228 78175 1268 78184
rect 1228 75200 1268 75209
rect 1324 75200 1364 78184
rect 1268 75160 1364 75200
rect 1228 75151 1268 75160
rect 1324 74696 1364 75160
rect 1420 74873 1460 79351
rect 1516 76040 1556 81115
rect 1611 80576 1653 80585
rect 1611 80536 1612 80576
rect 1652 80536 1653 80576
rect 1611 80527 1653 80536
rect 1612 80442 1652 80527
rect 1516 75991 1556 76000
rect 1611 76040 1653 76049
rect 1611 76000 1612 76040
rect 1652 76000 1653 76040
rect 1611 75991 1653 76000
rect 1612 75906 1652 75991
rect 1708 75788 1748 82207
rect 1803 82004 1845 82013
rect 1803 81964 1804 82004
rect 1844 81964 1845 82004
rect 1803 81955 1845 81964
rect 1804 80417 1844 81955
rect 1900 80501 1940 82720
rect 1996 81920 2036 83644
rect 3052 83634 3092 83719
rect 2092 83516 2132 83525
rect 2476 83516 2516 83525
rect 2132 83476 2228 83516
rect 2092 83467 2132 83476
rect 1996 81880 2132 81920
rect 1899 80492 1941 80501
rect 1899 80452 1900 80492
rect 1940 80452 1941 80492
rect 1899 80443 1941 80452
rect 1803 80408 1845 80417
rect 1803 80368 1804 80408
rect 1844 80368 1845 80408
rect 1803 80359 1845 80368
rect 1900 79064 1940 79075
rect 1900 78989 1940 79024
rect 1899 78980 1941 78989
rect 1899 78940 1900 78980
rect 1940 78940 1941 78980
rect 1899 78931 1941 78940
rect 1803 78140 1845 78149
rect 1803 78100 1804 78140
rect 1844 78100 1845 78140
rect 1803 78091 1845 78100
rect 1804 75965 1844 78091
rect 2092 76712 2132 81880
rect 2092 76628 2132 76672
rect 1900 76588 2132 76628
rect 1803 75956 1845 75965
rect 1803 75916 1804 75956
rect 1844 75916 1845 75956
rect 1803 75907 1845 75916
rect 1612 75748 1748 75788
rect 1419 74864 1461 74873
rect 1419 74824 1420 74864
rect 1460 74824 1461 74864
rect 1419 74815 1461 74824
rect 1324 74656 1556 74696
rect 1419 74528 1461 74537
rect 1419 74488 1420 74528
rect 1460 74488 1461 74528
rect 1419 74479 1461 74488
rect 1420 74394 1460 74479
rect 1228 74285 1268 74370
rect 1227 74276 1269 74285
rect 1227 74236 1228 74276
rect 1268 74236 1269 74276
rect 1227 74227 1269 74236
rect 1132 74068 1268 74108
rect 1131 73352 1173 73361
rect 1131 73312 1132 73352
rect 1172 73312 1173 73352
rect 1131 73303 1173 73312
rect 1035 72932 1077 72941
rect 1035 72892 1036 72932
rect 1076 72892 1077 72932
rect 1035 72883 1077 72892
rect 1036 68489 1076 72883
rect 1132 72353 1172 73303
rect 1228 73268 1268 74068
rect 1323 74024 1365 74033
rect 1323 73984 1324 74024
rect 1364 73984 1365 74024
rect 1323 73975 1365 73984
rect 1324 73529 1364 73975
rect 1323 73520 1365 73529
rect 1323 73480 1324 73520
rect 1364 73480 1365 73520
rect 1323 73471 1365 73480
rect 1516 73445 1556 74656
rect 1612 74369 1652 75748
rect 1900 75620 1940 76588
rect 2188 76301 2228 83476
rect 2476 82265 2516 83476
rect 2859 83516 2901 83525
rect 2859 83476 2860 83516
rect 2900 83476 2901 83516
rect 2859 83467 2901 83476
rect 3244 83516 3284 83525
rect 2860 83382 2900 83467
rect 3148 82760 3188 82769
rect 3148 82601 3188 82720
rect 2571 82592 2613 82601
rect 2571 82552 2572 82592
rect 2612 82552 2613 82592
rect 2571 82543 2613 82552
rect 3147 82592 3189 82601
rect 3147 82552 3148 82592
rect 3188 82552 3189 82592
rect 3147 82543 3189 82552
rect 2475 82256 2517 82265
rect 2475 82216 2476 82256
rect 2516 82216 2517 82256
rect 2475 82207 2517 82216
rect 2476 82088 2516 82097
rect 2572 82088 2612 82543
rect 2516 82048 2612 82088
rect 2476 82039 2516 82048
rect 2668 81836 2708 81845
rect 2708 81796 2804 81836
rect 2668 81787 2708 81796
rect 2668 81248 2708 81257
rect 2668 80753 2708 81208
rect 2667 80744 2709 80753
rect 2667 80704 2668 80744
rect 2708 80704 2709 80744
rect 2667 80695 2709 80704
rect 2571 80408 2613 80417
rect 2571 80368 2572 80408
rect 2612 80368 2613 80408
rect 2571 80359 2613 80368
rect 2379 79148 2421 79157
rect 2379 79108 2380 79148
rect 2420 79108 2421 79148
rect 2379 79099 2421 79108
rect 2283 76796 2325 76805
rect 2283 76756 2284 76796
rect 2324 76756 2325 76796
rect 2283 76747 2325 76756
rect 2187 76292 2229 76301
rect 2187 76252 2188 76292
rect 2228 76252 2229 76292
rect 2187 76243 2229 76252
rect 1708 75580 1940 75620
rect 1996 75956 2036 75965
rect 1708 74789 1748 75580
rect 1899 75452 1941 75461
rect 1899 75412 1900 75452
rect 1940 75412 1941 75452
rect 1899 75403 1941 75412
rect 1803 74864 1845 74873
rect 1803 74824 1804 74864
rect 1844 74824 1845 74864
rect 1803 74815 1845 74824
rect 1707 74780 1749 74789
rect 1707 74740 1708 74780
rect 1748 74740 1749 74780
rect 1707 74731 1749 74740
rect 1611 74360 1653 74369
rect 1611 74320 1612 74360
rect 1652 74320 1653 74360
rect 1611 74311 1653 74320
rect 1707 74276 1749 74285
rect 1707 74236 1708 74276
rect 1748 74236 1749 74276
rect 1707 74227 1749 74236
rect 1611 73688 1653 73697
rect 1611 73648 1612 73688
rect 1652 73648 1653 73688
rect 1611 73639 1653 73648
rect 1515 73436 1557 73445
rect 1515 73396 1516 73436
rect 1556 73396 1557 73436
rect 1515 73387 1557 73396
rect 1228 73228 1364 73268
rect 1228 73025 1268 73110
rect 1227 73016 1269 73025
rect 1227 72976 1228 73016
rect 1268 72976 1269 73016
rect 1227 72967 1269 72976
rect 1324 72848 1364 73228
rect 1228 72808 1364 72848
rect 1131 72344 1173 72353
rect 1131 72304 1132 72344
rect 1172 72304 1173 72344
rect 1131 72295 1173 72304
rect 1132 69245 1172 72295
rect 1228 71504 1268 72808
rect 1612 72689 1652 73639
rect 1611 72680 1653 72689
rect 1611 72640 1612 72680
rect 1652 72640 1653 72680
rect 1611 72631 1653 72640
rect 1419 72176 1461 72185
rect 1419 72136 1420 72176
rect 1460 72136 1461 72176
rect 1419 72127 1461 72136
rect 1228 70589 1268 71464
rect 1227 70580 1269 70589
rect 1227 70540 1228 70580
rect 1268 70540 1269 70580
rect 1227 70531 1269 70540
rect 1228 69992 1268 70001
rect 1323 69992 1365 70001
rect 1268 69952 1324 69992
rect 1364 69952 1365 69992
rect 1228 69943 1268 69952
rect 1323 69943 1365 69952
rect 1131 69236 1173 69245
rect 1131 69196 1132 69236
rect 1172 69196 1173 69236
rect 1131 69187 1173 69196
rect 1035 68480 1077 68489
rect 1035 68440 1036 68480
rect 1076 68440 1077 68480
rect 1035 68431 1077 68440
rect 1131 67640 1173 67649
rect 1131 67600 1132 67640
rect 1172 67600 1173 67640
rect 1131 67591 1173 67600
rect 939 66968 981 66977
rect 939 66928 940 66968
rect 980 66928 981 66968
rect 939 66919 981 66928
rect 171 65204 213 65213
rect 171 65164 172 65204
rect 212 65164 213 65204
rect 171 65155 213 65164
rect 1132 63785 1172 67591
rect 1227 66884 1269 66893
rect 1227 66844 1228 66884
rect 1268 66844 1269 66884
rect 1227 66835 1269 66844
rect 1228 66128 1268 66835
rect 1228 66079 1268 66088
rect 1323 65036 1365 65045
rect 1323 64996 1324 65036
rect 1364 64996 1365 65036
rect 1323 64987 1365 64996
rect 1324 64625 1364 64987
rect 1420 64700 1460 72127
rect 1515 72092 1557 72101
rect 1515 72052 1516 72092
rect 1556 72052 1557 72092
rect 1515 72043 1557 72052
rect 1516 65045 1556 72043
rect 1612 68060 1652 72631
rect 1708 69152 1748 74227
rect 1804 73688 1844 74815
rect 1900 73865 1940 75403
rect 1996 73949 2036 75916
rect 2092 75956 2132 75965
rect 2092 75461 2132 75916
rect 2187 75956 2229 75965
rect 2187 75916 2188 75956
rect 2228 75916 2229 75956
rect 2187 75907 2229 75916
rect 2091 75452 2133 75461
rect 2091 75412 2092 75452
rect 2132 75412 2133 75452
rect 2091 75403 2133 75412
rect 2188 74192 2228 75907
rect 2092 74152 2228 74192
rect 1995 73940 2037 73949
rect 1995 73900 1996 73940
rect 2036 73900 2037 73940
rect 1995 73891 2037 73900
rect 1899 73856 1941 73865
rect 1899 73816 1900 73856
rect 1940 73816 1941 73856
rect 1899 73807 1941 73816
rect 1804 73639 1844 73648
rect 1900 73688 1940 73697
rect 1803 73520 1845 73529
rect 1803 73480 1804 73520
rect 1844 73480 1845 73520
rect 1803 73471 1845 73480
rect 1804 71588 1844 73471
rect 1900 72185 1940 73648
rect 2092 73100 2132 74152
rect 2187 73940 2229 73949
rect 2187 73900 2188 73940
rect 2228 73900 2229 73940
rect 2187 73891 2229 73900
rect 1996 73060 2132 73100
rect 1899 72176 1941 72185
rect 1899 72136 1900 72176
rect 1940 72136 1941 72176
rect 1899 72127 1941 72136
rect 1996 72176 2036 73060
rect 1996 72127 2036 72136
rect 2091 72176 2133 72185
rect 2091 72136 2092 72176
rect 2132 72136 2133 72176
rect 2091 72127 2133 72136
rect 2092 72042 2132 72127
rect 2188 71924 2228 73891
rect 2284 73865 2324 76747
rect 2380 75209 2420 79099
rect 2572 78401 2612 80359
rect 2667 79736 2709 79745
rect 2667 79696 2668 79736
rect 2708 79696 2709 79736
rect 2667 79687 2709 79696
rect 2668 79602 2708 79687
rect 2667 79064 2709 79073
rect 2667 79024 2668 79064
rect 2708 79024 2709 79064
rect 2667 79015 2709 79024
rect 2668 78905 2708 79015
rect 2667 78896 2709 78905
rect 2667 78856 2668 78896
rect 2708 78856 2709 78896
rect 2667 78847 2709 78856
rect 2571 78392 2613 78401
rect 2571 78352 2572 78392
rect 2612 78352 2613 78392
rect 2571 78343 2613 78352
rect 2476 78224 2516 78233
rect 2476 76805 2516 78184
rect 2572 77300 2612 78343
rect 2667 78140 2709 78149
rect 2667 78100 2668 78140
rect 2708 78100 2709 78140
rect 2667 78091 2709 78100
rect 2668 78006 2708 78091
rect 2764 77552 2804 81796
rect 3147 81416 3189 81425
rect 3147 81376 3148 81416
rect 3188 81376 3189 81416
rect 3147 81367 3189 81376
rect 2860 81248 2900 81257
rect 2900 81208 2996 81248
rect 2860 81199 2900 81208
rect 2860 80669 2900 80700
rect 2859 80660 2901 80669
rect 2859 80620 2860 80660
rect 2900 80620 2901 80660
rect 2859 80611 2901 80620
rect 2860 80576 2900 80611
rect 2860 79157 2900 80536
rect 2859 79148 2901 79157
rect 2859 79108 2860 79148
rect 2900 79108 2901 79148
rect 2859 79099 2901 79108
rect 2956 78065 2996 81208
rect 3052 80324 3092 80333
rect 2955 78056 2997 78065
rect 2955 78016 2956 78056
rect 2996 78016 2997 78056
rect 2955 78007 2997 78016
rect 2860 77552 2900 77561
rect 2764 77512 2860 77552
rect 2860 77503 2900 77512
rect 2955 77552 2997 77561
rect 2955 77512 2956 77552
rect 2996 77512 2997 77552
rect 2955 77503 2997 77512
rect 2956 77418 2996 77503
rect 2572 77260 2996 77300
rect 2475 76796 2517 76805
rect 2475 76756 2476 76796
rect 2516 76756 2517 76796
rect 2475 76747 2517 76756
rect 2572 76040 2612 76051
rect 2572 75965 2612 76000
rect 2571 75956 2613 75965
rect 2571 75916 2572 75956
rect 2612 75916 2613 75956
rect 2571 75907 2613 75916
rect 2379 75200 2421 75209
rect 2476 75200 2516 75228
rect 2379 75160 2380 75200
rect 2420 75160 2476 75200
rect 2379 75151 2421 75160
rect 2476 75151 2516 75160
rect 2763 75200 2805 75209
rect 2763 75160 2764 75200
rect 2804 75160 2805 75200
rect 2763 75151 2805 75160
rect 2668 75032 2708 75041
rect 2476 74992 2668 75032
rect 2283 73856 2325 73865
rect 2283 73816 2284 73856
rect 2324 73816 2325 73856
rect 2283 73807 2325 73816
rect 2380 73697 2420 73782
rect 2284 73688 2324 73697
rect 2284 72101 2324 73648
rect 2379 73688 2421 73697
rect 2379 73648 2380 73688
rect 2420 73648 2421 73688
rect 2379 73639 2421 73648
rect 2476 73520 2516 74992
rect 2668 74983 2708 74992
rect 2571 74864 2613 74873
rect 2571 74824 2572 74864
rect 2612 74824 2613 74864
rect 2571 74815 2613 74824
rect 2572 73781 2612 74815
rect 2667 74612 2709 74621
rect 2667 74572 2668 74612
rect 2708 74572 2709 74612
rect 2667 74563 2709 74572
rect 2668 74528 2708 74563
rect 2668 74477 2708 74488
rect 2764 74453 2804 75151
rect 2859 74780 2901 74789
rect 2859 74740 2860 74780
rect 2900 74740 2901 74780
rect 2859 74731 2901 74740
rect 2860 74537 2900 74731
rect 2859 74528 2901 74537
rect 2859 74488 2860 74528
rect 2900 74488 2901 74528
rect 2859 74479 2901 74488
rect 2763 74444 2805 74453
rect 2763 74404 2764 74444
rect 2804 74404 2805 74444
rect 2763 74395 2805 74404
rect 2860 74394 2900 74479
rect 2763 74276 2805 74285
rect 2763 74236 2764 74276
rect 2804 74236 2805 74276
rect 2763 74227 2805 74236
rect 2571 73772 2613 73781
rect 2571 73732 2572 73772
rect 2612 73732 2613 73772
rect 2571 73723 2613 73732
rect 2380 73480 2516 73520
rect 2283 72092 2325 72101
rect 2283 72052 2284 72092
rect 2324 72052 2325 72092
rect 2283 72043 2325 72052
rect 2188 71884 2324 71924
rect 1804 71548 2132 71588
rect 1900 69152 1940 69161
rect 1708 69112 1900 69152
rect 1900 69103 1940 69112
rect 1996 69152 2036 69161
rect 1612 68020 1940 68060
rect 1803 67808 1845 67817
rect 1803 67768 1804 67808
rect 1844 67768 1845 67808
rect 1803 67759 1845 67768
rect 1707 66968 1749 66977
rect 1707 66928 1708 66968
rect 1748 66928 1749 66968
rect 1707 66919 1749 66928
rect 1708 66834 1748 66919
rect 1611 65456 1653 65465
rect 1611 65416 1612 65456
rect 1652 65416 1653 65456
rect 1611 65407 1653 65416
rect 1708 65456 1748 65467
rect 1612 65322 1652 65407
rect 1708 65381 1748 65416
rect 1707 65372 1749 65381
rect 1707 65332 1708 65372
rect 1748 65332 1749 65372
rect 1707 65323 1749 65332
rect 1804 65297 1844 67759
rect 1803 65288 1845 65297
rect 1803 65248 1804 65288
rect 1844 65248 1845 65288
rect 1803 65239 1845 65248
rect 1515 65036 1557 65045
rect 1515 64996 1516 65036
rect 1556 64996 1557 65036
rect 1515 64987 1557 64996
rect 1803 65036 1845 65045
rect 1803 64996 1804 65036
rect 1844 64996 1845 65036
rect 1803 64987 1845 64996
rect 1420 64660 1652 64700
rect 1228 64616 1268 64625
rect 1131 63776 1173 63785
rect 1131 63736 1132 63776
rect 1172 63736 1173 63776
rect 1131 63727 1173 63736
rect 1228 63188 1268 64576
rect 1323 64616 1365 64625
rect 1323 64576 1324 64616
rect 1364 64576 1365 64616
rect 1323 64567 1365 64576
rect 1228 63148 1556 63188
rect 1419 63020 1461 63029
rect 1419 62980 1420 63020
rect 1460 62980 1461 63020
rect 1419 62971 1461 62980
rect 1420 60080 1460 62971
rect 1420 59240 1460 60040
rect 1516 59753 1556 63148
rect 1612 61937 1652 64660
rect 1707 62432 1749 62441
rect 1707 62392 1708 62432
rect 1748 62392 1749 62432
rect 1707 62383 1749 62392
rect 1708 62298 1748 62383
rect 1611 61928 1653 61937
rect 1611 61888 1612 61928
rect 1652 61888 1653 61928
rect 1611 61879 1653 61888
rect 1611 59996 1653 60005
rect 1611 59956 1612 59996
rect 1652 59956 1653 59996
rect 1611 59947 1653 59956
rect 1515 59744 1557 59753
rect 1515 59704 1516 59744
rect 1556 59704 1557 59744
rect 1515 59695 1557 59704
rect 1324 59200 1460 59240
rect 1324 58736 1364 59200
rect 1132 58696 1364 58736
rect 1132 58400 1172 58696
rect 1228 58568 1268 58577
rect 1516 58568 1556 59695
rect 1268 58528 1556 58568
rect 1228 58519 1268 58528
rect 1612 58484 1652 59947
rect 1804 59240 1844 64987
rect 1900 64205 1940 68020
rect 1996 67649 2036 69112
rect 1995 67640 2037 67649
rect 1995 67600 1996 67640
rect 2036 67600 2037 67640
rect 1995 67591 2037 67600
rect 1899 64196 1941 64205
rect 1899 64156 1900 64196
rect 1940 64156 1941 64196
rect 1899 64147 1941 64156
rect 1996 62609 2036 67591
rect 2092 66557 2132 71548
rect 2187 71420 2229 71429
rect 2187 71380 2188 71420
rect 2228 71380 2229 71420
rect 2187 71371 2229 71380
rect 2188 68237 2228 71371
rect 2187 68228 2229 68237
rect 2187 68188 2188 68228
rect 2228 68188 2229 68228
rect 2187 68179 2229 68188
rect 2284 68060 2324 71884
rect 2380 70678 2420 73480
rect 2475 73016 2517 73025
rect 2475 72976 2476 73016
rect 2516 72976 2517 73016
rect 2475 72967 2517 72976
rect 2476 72882 2516 72967
rect 2572 72260 2612 73723
rect 2572 72211 2612 72220
rect 2668 72764 2708 72773
rect 2476 72176 2516 72187
rect 2476 72101 2516 72136
rect 2475 72092 2517 72101
rect 2475 72052 2476 72092
rect 2516 72052 2517 72092
rect 2475 72043 2517 72052
rect 2475 71924 2517 71933
rect 2475 71884 2476 71924
rect 2516 71884 2517 71924
rect 2475 71875 2517 71884
rect 2476 71504 2516 71875
rect 2476 70832 2516 71464
rect 2668 71429 2708 72724
rect 2667 71420 2709 71429
rect 2667 71380 2668 71420
rect 2708 71380 2709 71420
rect 2667 71371 2709 71380
rect 2667 71252 2709 71261
rect 2667 71212 2668 71252
rect 2708 71212 2709 71252
rect 2667 71203 2709 71212
rect 2668 71118 2708 71203
rect 2476 70792 2708 70832
rect 2380 70664 2516 70678
rect 2380 70638 2476 70664
rect 2476 70615 2516 70624
rect 2571 70664 2613 70673
rect 2571 70624 2572 70664
rect 2612 70624 2613 70664
rect 2571 70615 2613 70624
rect 2379 70580 2421 70589
rect 2379 70540 2380 70580
rect 2420 70540 2421 70580
rect 2379 70531 2421 70540
rect 2380 69404 2420 70531
rect 2572 70530 2612 70615
rect 2668 70001 2708 70792
rect 2475 69992 2517 70001
rect 2475 69952 2476 69992
rect 2516 69952 2517 69992
rect 2475 69943 2517 69952
rect 2667 69992 2709 70001
rect 2667 69952 2668 69992
rect 2708 69952 2709 69992
rect 2667 69943 2709 69952
rect 2476 69858 2516 69943
rect 2667 69740 2709 69749
rect 2667 69700 2668 69740
rect 2708 69700 2709 69740
rect 2667 69691 2709 69700
rect 2668 69606 2708 69691
rect 2764 69488 2804 74227
rect 2859 74192 2901 74201
rect 2859 74152 2860 74192
rect 2900 74152 2901 74192
rect 2859 74143 2901 74152
rect 2860 73688 2900 74143
rect 2860 73100 2900 73648
rect 2956 73445 2996 77260
rect 3052 76035 3092 80284
rect 3148 79409 3188 81367
rect 3147 79400 3189 79409
rect 3147 79360 3148 79400
rect 3188 79360 3189 79400
rect 3147 79351 3189 79360
rect 3147 79064 3189 79073
rect 3147 79024 3148 79064
rect 3188 79024 3189 79064
rect 3147 79015 3189 79024
rect 3148 78930 3188 79015
rect 3244 78980 3284 83476
rect 3340 83096 3380 85936
rect 3435 84608 3477 84617
rect 3435 84568 3436 84608
rect 3476 84568 3477 84608
rect 3435 84559 3477 84568
rect 3436 84440 3476 84559
rect 3436 84391 3476 84400
rect 3436 83768 3476 83777
rect 3532 83768 3572 85936
rect 3724 85877 3764 85936
rect 3723 85868 3765 85877
rect 3723 85828 3724 85868
rect 3764 85828 3765 85868
rect 3723 85819 3765 85828
rect 3916 84860 3956 85936
rect 4108 85028 4148 85936
rect 4300 85793 4340 85936
rect 4299 85784 4341 85793
rect 4299 85744 4300 85784
rect 4340 85744 4341 85784
rect 4299 85735 4341 85744
rect 4108 84988 4340 85028
rect 4203 84860 4245 84869
rect 3916 84820 4148 84860
rect 3688 84692 4056 84701
rect 3728 84652 3770 84692
rect 3810 84652 3852 84692
rect 3892 84652 3934 84692
rect 3974 84652 4016 84692
rect 3688 84643 4056 84652
rect 3628 84356 3668 84365
rect 3628 84197 3668 84316
rect 3627 84188 3669 84197
rect 3627 84148 3628 84188
rect 3668 84148 3669 84188
rect 3627 84139 3669 84148
rect 3476 83728 3572 83768
rect 3820 83768 3860 83777
rect 4108 83768 4148 84820
rect 4203 84820 4204 84860
rect 4244 84820 4245 84860
rect 4203 84811 4245 84820
rect 3860 83728 4148 83768
rect 4204 83768 4244 84811
rect 4300 83777 4340 84988
rect 3436 83719 3476 83728
rect 3820 83719 3860 83728
rect 4204 83719 4244 83728
rect 4299 83768 4341 83777
rect 4299 83728 4300 83768
rect 4340 83728 4341 83768
rect 4299 83719 4341 83728
rect 3628 83516 3668 83525
rect 3628 83357 3668 83476
rect 4012 83516 4052 83525
rect 4395 83516 4437 83525
rect 4052 83476 4244 83516
rect 4012 83467 4052 83476
rect 3627 83348 3669 83357
rect 3627 83308 3628 83348
rect 3668 83308 3669 83348
rect 3627 83299 3669 83308
rect 3688 83180 4056 83189
rect 3728 83140 3770 83180
rect 3810 83140 3852 83180
rect 3892 83140 3934 83180
rect 3974 83140 4016 83180
rect 3688 83131 4056 83140
rect 3340 83056 3572 83096
rect 3532 83012 3572 83056
rect 3628 83012 3668 83021
rect 3532 82972 3628 83012
rect 3628 82963 3668 82972
rect 3820 82844 3860 82853
rect 3340 82592 3380 82601
rect 3380 82552 3572 82592
rect 3340 82543 3380 82552
rect 3435 82088 3477 82097
rect 3435 82048 3436 82088
rect 3476 82048 3477 82088
rect 3435 82039 3477 82048
rect 3436 81920 3476 82039
rect 3340 81880 3476 81920
rect 3340 80081 3380 81880
rect 3435 81752 3477 81761
rect 3435 81712 3436 81752
rect 3476 81712 3477 81752
rect 3435 81703 3477 81712
rect 3339 80072 3381 80081
rect 3339 80032 3340 80072
rect 3380 80032 3381 80072
rect 3339 80023 3381 80032
rect 3436 79064 3476 81703
rect 3532 79736 3572 82552
rect 3723 82088 3765 82097
rect 3723 82048 3724 82088
rect 3764 82048 3765 82088
rect 3723 82039 3765 82048
rect 3724 81954 3764 82039
rect 3820 81929 3860 82804
rect 4108 82769 4148 82854
rect 4107 82760 4149 82769
rect 4107 82720 4108 82760
rect 4148 82720 4149 82760
rect 4107 82711 4149 82720
rect 4107 82592 4149 82601
rect 4107 82552 4108 82592
rect 4148 82552 4149 82592
rect 4107 82543 4149 82552
rect 3819 81920 3861 81929
rect 3819 81880 3820 81920
rect 3860 81880 3861 81920
rect 3819 81871 3861 81880
rect 4108 81845 4148 82543
rect 4107 81836 4149 81845
rect 4107 81796 4108 81836
rect 4148 81796 4149 81836
rect 4107 81787 4149 81796
rect 3688 81668 4056 81677
rect 3728 81628 3770 81668
rect 3810 81628 3852 81668
rect 3892 81628 3934 81668
rect 3974 81628 4016 81668
rect 3688 81619 4056 81628
rect 4011 81500 4053 81509
rect 4011 81460 4012 81500
rect 4052 81460 4053 81500
rect 4011 81451 4053 81460
rect 3724 80576 3764 80585
rect 3724 80417 3764 80536
rect 3723 80408 3765 80417
rect 3723 80368 3724 80408
rect 3764 80368 3765 80408
rect 3723 80359 3765 80368
rect 4012 80324 4052 81451
rect 4108 81248 4148 81787
rect 4108 81199 4148 81208
rect 4204 80576 4244 83476
rect 4395 83476 4396 83516
rect 4436 83476 4437 83516
rect 4395 83467 4437 83476
rect 4396 83382 4436 83467
rect 4492 83264 4532 85936
rect 4684 84869 4724 85936
rect 4683 84860 4725 84869
rect 4683 84820 4684 84860
rect 4724 84820 4725 84860
rect 4683 84811 4725 84820
rect 4876 84692 4916 85936
rect 4588 84652 4916 84692
rect 4588 83432 4628 84652
rect 5068 84113 5108 85936
rect 5260 84449 5300 85936
rect 5259 84440 5301 84449
rect 5259 84400 5260 84440
rect 5300 84400 5301 84440
rect 5259 84391 5301 84400
rect 5067 84104 5109 84113
rect 5067 84064 5068 84104
rect 5108 84064 5109 84104
rect 5067 84055 5109 84064
rect 4928 83936 5296 83945
rect 4968 83896 5010 83936
rect 5050 83896 5092 83936
rect 5132 83896 5174 83936
rect 5214 83896 5256 83936
rect 4928 83887 5296 83896
rect 5356 83768 5396 83777
rect 5452 83768 5492 85936
rect 5644 84608 5684 85936
rect 5548 84568 5684 84608
rect 5548 84281 5588 84568
rect 5836 84449 5876 85936
rect 6028 84533 6068 85936
rect 6027 84524 6069 84533
rect 6027 84484 6028 84524
rect 6068 84484 6069 84524
rect 6027 84475 6069 84484
rect 6220 84449 6260 85936
rect 6412 84449 6452 85936
rect 6604 84533 6644 85936
rect 6603 84524 6645 84533
rect 6603 84484 6604 84524
rect 6644 84484 6645 84524
rect 6603 84475 6645 84484
rect 6796 84449 6836 85936
rect 6988 84449 7028 85936
rect 5643 84440 5685 84449
rect 5643 84400 5644 84440
rect 5684 84400 5685 84440
rect 5643 84391 5685 84400
rect 5835 84440 5877 84449
rect 5835 84400 5836 84440
rect 5876 84400 5877 84440
rect 5835 84391 5877 84400
rect 6219 84440 6261 84449
rect 6219 84400 6220 84440
rect 6260 84400 6261 84440
rect 6219 84391 6261 84400
rect 6411 84440 6453 84449
rect 6411 84400 6412 84440
rect 6452 84400 6453 84440
rect 6411 84391 6453 84400
rect 6795 84440 6837 84449
rect 6795 84400 6796 84440
rect 6836 84400 6837 84440
rect 6795 84391 6837 84400
rect 6987 84440 7029 84449
rect 6987 84400 6988 84440
rect 7028 84400 7029 84440
rect 6987 84391 7029 84400
rect 5547 84272 5589 84281
rect 5547 84232 5548 84272
rect 5588 84232 5589 84272
rect 5547 84223 5589 84232
rect 5547 83852 5589 83861
rect 5547 83812 5548 83852
rect 5588 83812 5589 83852
rect 5547 83803 5589 83812
rect 5396 83728 5492 83768
rect 5548 83768 5588 83803
rect 5356 83719 5396 83728
rect 5548 83717 5588 83728
rect 5644 83693 5684 84391
rect 6411 84020 6453 84029
rect 6411 83980 6412 84020
rect 6452 83980 6453 84020
rect 6411 83971 6453 83980
rect 6219 83852 6261 83861
rect 6219 83812 6220 83852
rect 6260 83812 6261 83852
rect 6219 83803 6261 83812
rect 6220 83768 6260 83803
rect 6220 83717 6260 83728
rect 6412 83768 6452 83971
rect 7180 83861 7220 85936
rect 7179 83852 7221 83861
rect 7179 83812 7180 83852
rect 7220 83812 7221 83852
rect 7372 83852 7412 85936
rect 7564 84440 7604 85936
rect 7564 84400 7700 84440
rect 7372 83812 7604 83852
rect 7179 83803 7221 83812
rect 6412 83719 6452 83728
rect 6987 83768 7029 83777
rect 6987 83728 6988 83768
rect 7028 83728 7029 83768
rect 6987 83719 7029 83728
rect 7564 83768 7604 83812
rect 7564 83719 7604 83728
rect 5643 83684 5685 83693
rect 5643 83644 5644 83684
rect 5684 83644 5685 83684
rect 5643 83635 5685 83644
rect 6988 83634 7028 83719
rect 4588 83383 4628 83392
rect 4972 83516 5012 83525
rect 4972 83357 5012 83476
rect 5164 83516 5204 83525
rect 5739 83516 5781 83525
rect 5204 83476 5684 83516
rect 5164 83467 5204 83476
rect 4780 83348 4820 83357
rect 4780 83264 4820 83308
rect 4971 83348 5013 83357
rect 4971 83308 4972 83348
rect 5012 83308 5013 83348
rect 4971 83299 5013 83308
rect 4492 83224 4820 83264
rect 5356 82760 5396 82769
rect 4683 82508 4725 82517
rect 4683 82468 4684 82508
rect 4724 82468 4725 82508
rect 4683 82459 4725 82468
rect 4492 81248 4532 81257
rect 4300 81080 4340 81089
rect 4340 81040 4436 81080
rect 4300 81031 4340 81040
rect 4204 80536 4340 80576
rect 4012 80284 4148 80324
rect 3688 80156 4056 80165
rect 3728 80116 3770 80156
rect 3810 80116 3852 80156
rect 3892 80116 3934 80156
rect 3974 80116 4016 80156
rect 3688 80107 4056 80116
rect 4108 79988 4148 80284
rect 4012 79948 4148 79988
rect 3628 79736 3668 79745
rect 3532 79696 3628 79736
rect 3628 79687 3668 79696
rect 3724 79736 3764 79747
rect 3724 79661 3764 79696
rect 3723 79652 3765 79661
rect 3723 79612 3724 79652
rect 3764 79612 3765 79652
rect 3723 79603 3765 79612
rect 3436 79024 3572 79064
rect 3244 78940 3476 78980
rect 3340 78812 3380 78821
rect 3244 78772 3340 78812
rect 3147 78056 3189 78065
rect 3147 78016 3148 78056
rect 3188 78016 3189 78056
rect 3147 78007 3189 78016
rect 3052 75986 3092 75995
rect 3051 75284 3093 75293
rect 3051 75244 3052 75284
rect 3092 75244 3093 75284
rect 3051 75235 3093 75244
rect 3052 74621 3092 75235
rect 3051 74612 3093 74621
rect 3051 74572 3052 74612
rect 3092 74572 3093 74612
rect 3051 74563 3093 74572
rect 3051 74444 3093 74453
rect 3051 74404 3052 74444
rect 3092 74404 3093 74444
rect 3051 74395 3093 74404
rect 2955 73436 2997 73445
rect 2955 73396 2956 73436
rect 2996 73396 2997 73436
rect 2955 73387 2997 73396
rect 3052 73193 3092 74395
rect 3148 73613 3188 78007
rect 3244 76460 3284 78772
rect 3340 78763 3380 78772
rect 3340 78233 3380 78318
rect 3339 78224 3381 78233
rect 3339 78184 3340 78224
rect 3380 78184 3381 78224
rect 3339 78175 3381 78184
rect 3339 77972 3381 77981
rect 3339 77932 3340 77972
rect 3380 77932 3381 77972
rect 3339 77923 3381 77932
rect 3340 77552 3380 77923
rect 3436 77645 3476 78940
rect 3435 77636 3477 77645
rect 3435 77596 3436 77636
rect 3476 77596 3477 77636
rect 3435 77587 3477 77596
rect 3340 77503 3380 77512
rect 3435 77468 3477 77477
rect 3435 77428 3436 77468
rect 3476 77428 3477 77468
rect 3435 77419 3477 77428
rect 3436 77334 3476 77419
rect 3339 76796 3381 76805
rect 3339 76756 3340 76796
rect 3380 76756 3381 76796
rect 3339 76747 3381 76756
rect 3340 76712 3380 76747
rect 3532 76712 3572 79024
rect 4012 78812 4052 79948
rect 4107 79820 4149 79829
rect 4107 79780 4108 79820
rect 4148 79780 4149 79820
rect 4107 79771 4149 79780
rect 4108 79686 4148 79771
rect 4203 79736 4245 79745
rect 4203 79696 4204 79736
rect 4244 79696 4245 79736
rect 4203 79687 4245 79696
rect 4204 79602 4244 79687
rect 4300 79661 4340 80536
rect 4299 79652 4341 79661
rect 4299 79612 4300 79652
rect 4340 79612 4341 79652
rect 4299 79603 4341 79612
rect 4204 79064 4244 79075
rect 4204 78989 4244 79024
rect 4203 78980 4245 78989
rect 4203 78940 4204 78980
rect 4244 78940 4245 78980
rect 4203 78931 4245 78940
rect 4012 78772 4148 78812
rect 3688 78644 4056 78653
rect 3728 78604 3770 78644
rect 3810 78604 3852 78644
rect 3892 78604 3934 78644
rect 3974 78604 4016 78644
rect 3688 78595 4056 78604
rect 3915 78476 3957 78485
rect 3915 78436 3916 78476
rect 3956 78436 3957 78476
rect 3915 78427 3957 78436
rect 3916 77552 3956 78427
rect 3916 77503 3956 77512
rect 3688 77132 4056 77141
rect 3728 77092 3770 77132
rect 3810 77092 3852 77132
rect 3892 77092 3934 77132
rect 3974 77092 4016 77132
rect 3688 77083 4056 77092
rect 4108 76721 4148 78772
rect 4299 78056 4341 78065
rect 4299 78016 4300 78056
rect 4340 78016 4341 78056
rect 4299 78007 4341 78016
rect 4203 77636 4245 77645
rect 4203 77596 4204 77636
rect 4244 77596 4245 77636
rect 4203 77587 4245 77596
rect 3340 76661 3380 76672
rect 3436 76672 3572 76712
rect 4107 76712 4149 76721
rect 4107 76672 4108 76712
rect 4148 76672 4149 76712
rect 3244 76420 3380 76460
rect 3243 76292 3285 76301
rect 3243 76252 3244 76292
rect 3284 76252 3285 76292
rect 3243 76243 3285 76252
rect 3244 76208 3284 76243
rect 3244 76157 3284 76168
rect 3243 74528 3285 74537
rect 3243 74488 3244 74528
rect 3284 74488 3285 74528
rect 3243 74479 3285 74488
rect 3147 73604 3189 73613
rect 3147 73564 3148 73604
rect 3188 73564 3189 73604
rect 3147 73555 3189 73564
rect 3147 73436 3189 73445
rect 3147 73396 3148 73436
rect 3188 73396 3189 73436
rect 3147 73387 3189 73396
rect 3051 73184 3093 73193
rect 3051 73144 3052 73184
rect 3092 73144 3093 73184
rect 3051 73135 3093 73144
rect 2860 73060 2996 73100
rect 2859 72764 2901 72773
rect 2859 72724 2860 72764
rect 2900 72724 2901 72764
rect 2859 72715 2901 72724
rect 2860 72630 2900 72715
rect 2956 72596 2996 73060
rect 3052 73016 3092 73135
rect 3052 72967 3092 72976
rect 2956 72556 3092 72596
rect 2955 72428 2997 72437
rect 2955 72388 2956 72428
rect 2996 72388 2997 72428
rect 2955 72379 2997 72388
rect 2956 72101 2996 72379
rect 3052 72176 3092 72556
rect 3148 72260 3188 73387
rect 3244 72437 3284 74479
rect 3340 73702 3380 76420
rect 3436 74285 3476 76672
rect 4107 76663 4149 76672
rect 3531 76544 3573 76553
rect 3531 76504 3532 76544
rect 3572 76504 3573 76544
rect 3531 76495 3573 76504
rect 3532 76410 3572 76495
rect 3688 75620 4056 75629
rect 3728 75580 3770 75620
rect 3810 75580 3852 75620
rect 3892 75580 3934 75620
rect 3974 75580 4016 75620
rect 3688 75571 4056 75580
rect 3723 75452 3765 75461
rect 3723 75412 3724 75452
rect 3764 75412 3765 75452
rect 3723 75403 3765 75412
rect 3724 74369 3764 75403
rect 4108 75041 4148 76663
rect 4107 75032 4149 75041
rect 4107 74992 4108 75032
rect 4148 74992 4149 75032
rect 4107 74983 4149 74992
rect 4107 74528 4149 74537
rect 4107 74488 4108 74528
rect 4148 74488 4149 74528
rect 4107 74479 4149 74488
rect 4108 74394 4148 74479
rect 3531 74360 3573 74369
rect 3531 74320 3532 74360
rect 3572 74320 3573 74360
rect 3531 74311 3573 74320
rect 3723 74360 3765 74369
rect 3723 74320 3724 74360
rect 3764 74320 3765 74360
rect 3723 74311 3765 74320
rect 3435 74276 3477 74285
rect 3435 74236 3436 74276
rect 3476 74236 3477 74276
rect 3435 74227 3477 74236
rect 3340 73653 3380 73662
rect 3532 73604 3572 74311
rect 3688 74108 4056 74117
rect 3728 74068 3770 74108
rect 3810 74068 3852 74108
rect 3892 74068 3934 74108
rect 3974 74068 4016 74108
rect 3688 74059 4056 74068
rect 3532 73555 3572 73564
rect 3339 73520 3381 73529
rect 3339 73480 3340 73520
rect 3380 73480 3381 73520
rect 3339 73471 3381 73480
rect 3340 72605 3380 73471
rect 3531 73100 3573 73109
rect 3531 73060 3532 73100
rect 3572 73060 3573 73100
rect 3531 73051 3573 73060
rect 3435 72764 3477 72773
rect 3435 72724 3436 72764
rect 3476 72724 3477 72764
rect 3435 72715 3477 72724
rect 3339 72596 3381 72605
rect 3339 72556 3340 72596
rect 3380 72556 3381 72596
rect 3339 72547 3381 72556
rect 3243 72428 3285 72437
rect 3243 72388 3244 72428
rect 3284 72388 3285 72428
rect 3243 72379 3285 72388
rect 3148 72220 3380 72260
rect 3092 72136 3188 72176
rect 3052 72127 3092 72136
rect 2955 72092 2997 72101
rect 2955 72052 2956 72092
rect 2996 72052 2997 72092
rect 2955 72043 2997 72052
rect 2859 71504 2901 71513
rect 2859 71464 2860 71504
rect 2900 71464 2901 71504
rect 2859 71455 2901 71464
rect 2860 71370 2900 71455
rect 3051 71252 3093 71261
rect 3051 71212 3052 71252
rect 3092 71212 3093 71252
rect 3051 71203 3093 71212
rect 2859 71168 2901 71177
rect 2859 71128 2860 71168
rect 2900 71128 2901 71168
rect 2859 71119 2901 71128
rect 2860 70673 2900 71119
rect 2955 70748 2997 70757
rect 2955 70708 2956 70748
rect 2996 70708 2997 70748
rect 2955 70699 2997 70708
rect 3052 70748 3092 71203
rect 3052 70699 3092 70708
rect 2859 70664 2901 70673
rect 2859 70624 2860 70664
rect 2900 70624 2901 70664
rect 2859 70615 2901 70624
rect 2860 70085 2900 70615
rect 2956 70614 2996 70699
rect 2859 70076 2901 70085
rect 2859 70036 2860 70076
rect 2900 70036 2901 70076
rect 2859 70027 2901 70036
rect 3052 70001 3092 70086
rect 3051 69992 3093 70001
rect 3051 69952 3052 69992
rect 3092 69952 3093 69992
rect 3051 69943 3093 69952
rect 3148 69824 3188 72136
rect 3243 72092 3285 72101
rect 3243 72052 3244 72092
rect 3284 72052 3285 72092
rect 3243 72043 3285 72052
rect 3052 69784 3188 69824
rect 2859 69740 2901 69749
rect 2859 69700 2860 69740
rect 2900 69700 2901 69740
rect 2859 69691 2901 69700
rect 2860 69606 2900 69691
rect 2668 69448 2804 69488
rect 2668 69404 2708 69448
rect 2380 69364 2612 69404
rect 2475 69236 2517 69245
rect 2475 69196 2476 69236
rect 2516 69196 2517 69236
rect 2475 69187 2517 69196
rect 2380 69152 2420 69161
rect 2380 68732 2420 69112
rect 2476 69102 2516 69187
rect 2572 68909 2612 69364
rect 2667 69364 2708 69404
rect 2667 69320 2707 69364
rect 2667 69280 2708 69320
rect 2571 68900 2613 68909
rect 2571 68860 2572 68900
rect 2612 68860 2613 68900
rect 2571 68851 2613 68860
rect 2380 68692 2516 68732
rect 2380 68489 2420 68574
rect 2379 68480 2421 68489
rect 2379 68440 2380 68480
rect 2420 68440 2421 68480
rect 2379 68431 2421 68440
rect 2379 68228 2421 68237
rect 2379 68188 2380 68228
rect 2420 68188 2421 68228
rect 2379 68179 2421 68188
rect 2188 68020 2324 68060
rect 2091 66548 2133 66557
rect 2091 66508 2092 66548
rect 2132 66508 2133 66548
rect 2091 66499 2133 66508
rect 2188 66380 2228 68020
rect 2380 67640 2420 68179
rect 2476 67817 2516 68692
rect 2475 67808 2517 67817
rect 2475 67768 2476 67808
rect 2516 67768 2517 67808
rect 2475 67759 2517 67768
rect 2380 67591 2420 67600
rect 2475 67640 2517 67649
rect 2475 67600 2476 67640
rect 2516 67600 2517 67640
rect 2475 67591 2517 67600
rect 2476 67506 2516 67591
rect 2571 67556 2613 67565
rect 2571 67516 2572 67556
rect 2612 67516 2613 67556
rect 2571 67507 2613 67516
rect 2572 67145 2612 67507
rect 2571 67136 2613 67145
rect 2571 67096 2572 67136
rect 2612 67096 2613 67136
rect 2571 67087 2613 67096
rect 2283 66548 2325 66557
rect 2283 66508 2284 66548
rect 2324 66508 2325 66548
rect 2283 66499 2325 66508
rect 2092 66340 2228 66380
rect 2092 65633 2132 66340
rect 2187 65792 2229 65801
rect 2284 65792 2324 66499
rect 2571 66212 2613 66221
rect 2571 66172 2572 66212
rect 2612 66172 2613 66212
rect 2571 66163 2613 66172
rect 2187 65752 2188 65792
rect 2228 65752 2324 65792
rect 2476 66128 2516 66137
rect 2187 65743 2229 65752
rect 2091 65624 2133 65633
rect 2091 65584 2092 65624
rect 2132 65584 2133 65624
rect 2091 65575 2133 65584
rect 2092 65456 2132 65575
rect 2092 65407 2132 65416
rect 2188 65456 2228 65743
rect 2188 65407 2228 65416
rect 2476 65129 2516 66088
rect 2572 65456 2612 66163
rect 2668 66128 2708 69280
rect 2956 69152 2996 69161
rect 2956 68993 2996 69112
rect 2955 68984 2997 68993
rect 2955 68944 2956 68984
rect 2996 68944 2997 68984
rect 2955 68935 2997 68944
rect 2859 67808 2901 67817
rect 2859 67768 2860 67808
rect 2900 67768 2901 67808
rect 2859 67759 2901 67768
rect 2860 67724 2900 67759
rect 2860 67673 2900 67684
rect 2956 67640 2996 67649
rect 2859 67556 2901 67565
rect 2859 67516 2860 67556
rect 2900 67516 2901 67556
rect 2859 67507 2901 67516
rect 2668 66088 2804 66128
rect 2667 65960 2709 65969
rect 2667 65920 2668 65960
rect 2708 65920 2709 65960
rect 2667 65911 2709 65920
rect 2668 65826 2708 65911
rect 2668 65456 2708 65465
rect 2572 65416 2668 65456
rect 2571 65288 2613 65297
rect 2571 65248 2572 65288
rect 2612 65248 2613 65288
rect 2571 65239 2613 65248
rect 2091 65120 2133 65129
rect 2091 65080 2092 65120
rect 2132 65080 2133 65120
rect 2091 65071 2133 65080
rect 2475 65120 2517 65129
rect 2475 65080 2476 65120
rect 2516 65080 2517 65120
rect 2475 65071 2517 65080
rect 1995 62600 2037 62609
rect 1995 62560 1996 62600
rect 2036 62560 2037 62600
rect 1995 62551 2037 62560
rect 2092 62432 2132 65071
rect 2572 65045 2612 65239
rect 2571 65036 2613 65045
rect 2571 64996 2572 65036
rect 2612 64996 2613 65036
rect 2571 64987 2613 64996
rect 2668 64709 2708 65416
rect 2667 64700 2709 64709
rect 2667 64660 2668 64700
rect 2708 64660 2709 64700
rect 2667 64651 2709 64660
rect 2764 64625 2804 66088
rect 2476 64616 2516 64625
rect 2283 64532 2325 64541
rect 2283 64492 2284 64532
rect 2324 64492 2325 64532
rect 2283 64483 2325 64492
rect 2284 63944 2324 64483
rect 2284 63895 2324 63904
rect 2380 63944 2420 63953
rect 2380 63197 2420 63904
rect 2379 63188 2421 63197
rect 2379 63148 2380 63188
rect 2420 63148 2421 63188
rect 2379 63139 2421 63148
rect 1420 58444 1652 58484
rect 1708 59200 1844 59240
rect 1996 62392 2132 62432
rect 1132 58360 1364 58400
rect 555 57896 597 57905
rect 555 57856 556 57896
rect 596 57856 597 57896
rect 555 57847 597 57856
rect 556 53789 596 57847
rect 747 56888 789 56897
rect 747 56848 748 56888
rect 788 56848 789 56888
rect 747 56839 789 56848
rect 555 53780 597 53789
rect 555 53740 556 53780
rect 596 53740 597 53780
rect 555 53731 597 53740
rect 748 52949 788 56839
rect 1324 56468 1364 58360
rect 1132 56428 1364 56468
rect 1132 53780 1172 56428
rect 1420 56384 1460 58444
rect 1515 58316 1557 58325
rect 1515 58276 1516 58316
rect 1556 58276 1557 58316
rect 1515 58267 1557 58276
rect 1324 56344 1420 56384
rect 1228 54032 1268 54041
rect 1228 53948 1268 53992
rect 1324 53957 1364 56344
rect 1420 56335 1460 56344
rect 1420 55544 1460 55553
rect 1516 55544 1556 58267
rect 1708 57140 1748 59200
rect 1900 59156 1940 59165
rect 1900 58913 1940 59116
rect 1899 58904 1941 58913
rect 1899 58864 1900 58904
rect 1940 58864 1941 58904
rect 1899 58855 1941 58864
rect 1996 58652 2036 62392
rect 2380 61685 2420 63139
rect 2476 62693 2516 64576
rect 2763 64616 2805 64625
rect 2763 64576 2764 64616
rect 2804 64576 2805 64616
rect 2763 64567 2805 64576
rect 2668 64448 2708 64457
rect 2572 64408 2668 64448
rect 2475 62684 2517 62693
rect 2475 62644 2476 62684
rect 2516 62644 2517 62684
rect 2475 62635 2517 62644
rect 2379 61676 2421 61685
rect 2379 61636 2380 61676
rect 2420 61636 2421 61676
rect 2379 61627 2421 61636
rect 2187 61592 2229 61601
rect 2187 61552 2188 61592
rect 2228 61552 2229 61592
rect 2187 61543 2229 61552
rect 2284 61592 2324 61601
rect 2188 61458 2228 61543
rect 2284 60593 2324 61552
rect 2283 60584 2325 60593
rect 2283 60544 2284 60584
rect 2324 60544 2325 60584
rect 2283 60535 2325 60544
rect 2092 59333 2132 59418
rect 2572 59408 2612 64408
rect 2668 64399 2708 64408
rect 2763 64364 2805 64373
rect 2763 64324 2764 64364
rect 2804 64324 2805 64364
rect 2763 64315 2805 64324
rect 2667 64280 2709 64289
rect 2667 64240 2668 64280
rect 2708 64240 2709 64280
rect 2667 64231 2709 64240
rect 2668 63692 2708 64231
rect 2764 63944 2804 64315
rect 2764 63895 2804 63904
rect 2860 63944 2900 67507
rect 2956 67397 2996 67600
rect 2955 67388 2997 67397
rect 2955 67348 2956 67388
rect 2996 67348 2997 67388
rect 2955 67339 2997 67348
rect 2955 67052 2997 67061
rect 2955 67012 2956 67052
rect 2996 67012 2997 67052
rect 2955 67003 2997 67012
rect 2956 66968 2996 67003
rect 2956 66917 2996 66928
rect 2955 66716 2997 66725
rect 2955 66676 2956 66716
rect 2996 66676 2997 66716
rect 2955 66667 2997 66676
rect 2956 65381 2996 66667
rect 2955 65372 2997 65381
rect 2955 65332 2956 65372
rect 2996 65332 2997 65372
rect 2955 65323 2997 65332
rect 2955 64700 2997 64709
rect 2955 64660 2956 64700
rect 2996 64660 2997 64700
rect 2955 64651 2997 64660
rect 2860 63895 2900 63904
rect 2668 63652 2804 63692
rect 2764 63123 2804 63652
rect 2956 63281 2996 64651
rect 2955 63272 2997 63281
rect 2955 63232 2956 63272
rect 2996 63232 2997 63272
rect 2955 63223 2997 63232
rect 2764 63074 2804 63083
rect 2860 63104 2900 63113
rect 2860 63020 2900 63064
rect 2955 63104 2997 63113
rect 2955 63064 2956 63104
rect 2996 63064 2997 63104
rect 2955 63055 2997 63064
rect 2764 62980 2900 63020
rect 2667 62936 2709 62945
rect 2667 62896 2668 62936
rect 2708 62896 2709 62936
rect 2667 62887 2709 62896
rect 2668 61676 2708 62887
rect 2764 62777 2804 62980
rect 2956 62936 2996 63055
rect 3052 63029 3092 69784
rect 3147 68564 3189 68573
rect 3147 68524 3148 68564
rect 3188 68524 3189 68564
rect 3147 68515 3189 68524
rect 3148 67061 3188 68515
rect 3244 67565 3284 72043
rect 3243 67556 3285 67565
rect 3243 67516 3244 67556
rect 3284 67516 3285 67556
rect 3243 67507 3285 67516
rect 3147 67052 3189 67061
rect 3147 67012 3148 67052
rect 3188 67012 3189 67052
rect 3147 67003 3189 67012
rect 3148 66716 3188 66725
rect 3188 66676 3284 66716
rect 3148 66667 3188 66676
rect 3147 65624 3189 65633
rect 3147 65584 3148 65624
rect 3188 65584 3189 65624
rect 3147 65575 3189 65584
rect 3148 65451 3188 65575
rect 3148 65402 3188 65411
rect 3244 64532 3284 66676
rect 3340 65717 3380 72220
rect 3436 69166 3476 72715
rect 3532 72190 3572 73051
rect 3688 72596 4056 72605
rect 3728 72556 3770 72596
rect 3810 72556 3852 72596
rect 3892 72556 3934 72596
rect 3974 72556 4016 72596
rect 3688 72547 4056 72556
rect 3532 72141 3572 72150
rect 3723 72008 3765 72017
rect 3723 71968 3724 72008
rect 3764 71968 3765 72008
rect 3723 71959 3765 71968
rect 3724 71874 3764 71959
rect 3915 71924 3957 71933
rect 3915 71884 3916 71924
rect 3956 71884 3957 71924
rect 3915 71875 3957 71884
rect 3627 71840 3669 71849
rect 3627 71800 3628 71840
rect 3668 71800 3669 71840
rect 3627 71791 3669 71800
rect 3531 71504 3573 71513
rect 3531 71464 3532 71504
rect 3572 71464 3573 71504
rect 3531 71455 3573 71464
rect 3532 70916 3572 71455
rect 3628 71261 3668 71791
rect 3916 71513 3956 71875
rect 4108 71513 4148 71598
rect 3915 71504 3957 71513
rect 3915 71464 3916 71504
rect 3956 71464 3957 71504
rect 3915 71455 3957 71464
rect 4107 71504 4149 71513
rect 4107 71464 4108 71504
rect 4148 71464 4149 71504
rect 4107 71455 4149 71464
rect 3627 71252 3669 71261
rect 3627 71212 3628 71252
rect 3668 71212 3669 71252
rect 3627 71203 3669 71212
rect 3688 71084 4056 71093
rect 3728 71044 3770 71084
rect 3810 71044 3852 71084
rect 3892 71044 3934 71084
rect 3974 71044 4016 71084
rect 3688 71035 4056 71044
rect 3532 70876 3668 70916
rect 3532 70673 3572 70758
rect 3531 70664 3573 70673
rect 3531 70624 3532 70664
rect 3572 70624 3573 70664
rect 3531 70615 3573 70624
rect 3628 70496 3668 70876
rect 3723 70832 3765 70841
rect 3723 70792 3724 70832
rect 3764 70792 3765 70832
rect 3723 70783 3765 70792
rect 3436 69117 3476 69126
rect 3532 70456 3668 70496
rect 3435 68984 3477 68993
rect 3435 68944 3436 68984
rect 3476 68944 3477 68984
rect 3435 68935 3477 68944
rect 3436 67640 3476 68935
rect 3436 67591 3476 67600
rect 3532 67565 3572 70456
rect 3724 69749 3764 70783
rect 4011 70748 4053 70757
rect 4011 70708 4012 70748
rect 4052 70708 4053 70748
rect 4011 70699 4053 70708
rect 4012 70678 4052 70699
rect 4012 70613 4052 70638
rect 4204 70580 4244 77587
rect 4300 75200 4340 78007
rect 4396 77547 4436 81040
rect 4492 78905 4532 81208
rect 4587 80492 4629 80501
rect 4587 80452 4588 80492
rect 4628 80452 4629 80492
rect 4587 80443 4629 80452
rect 4491 78896 4533 78905
rect 4491 78856 4492 78896
rect 4532 78856 4533 78896
rect 4491 78847 4533 78856
rect 4588 78224 4628 80443
rect 4684 79736 4724 82459
rect 4928 82424 5296 82433
rect 4968 82384 5010 82424
rect 5050 82384 5092 82424
rect 5132 82384 5174 82424
rect 5214 82384 5256 82424
rect 4928 82375 5296 82384
rect 4972 82088 5012 82097
rect 5356 82088 5396 82720
rect 5548 82592 5588 82601
rect 5012 82048 5396 82088
rect 5452 82552 5548 82592
rect 4972 81845 5012 82048
rect 4971 81836 5013 81845
rect 4971 81796 4972 81836
rect 5012 81796 5013 81836
rect 4971 81787 5013 81796
rect 5164 81836 5204 81845
rect 5204 81796 5396 81836
rect 5164 81787 5204 81796
rect 4928 80912 5296 80921
rect 4968 80872 5010 80912
rect 5050 80872 5092 80912
rect 5132 80872 5174 80912
rect 5214 80872 5256 80912
rect 4928 80863 5296 80872
rect 4972 80669 5012 80700
rect 4971 80660 5013 80669
rect 4971 80620 4972 80660
rect 5012 80620 5013 80660
rect 4971 80611 5013 80620
rect 4972 80576 5012 80611
rect 4972 80501 5012 80536
rect 4971 80492 5013 80501
rect 4971 80452 4972 80492
rect 5012 80452 5013 80492
rect 4971 80443 5013 80452
rect 5163 80324 5205 80333
rect 5163 80284 5164 80324
rect 5204 80284 5205 80324
rect 5163 80275 5205 80284
rect 5164 80190 5204 80275
rect 5212 79745 5252 79754
rect 5356 79736 5396 81796
rect 5452 80576 5492 82552
rect 5548 82543 5588 82552
rect 5644 81920 5684 83476
rect 5739 83476 5740 83516
rect 5780 83476 5781 83516
rect 5739 83467 5781 83476
rect 6028 83516 6068 83525
rect 5740 83382 5780 83467
rect 5452 80527 5492 80536
rect 5548 81880 5684 81920
rect 5548 80576 5588 81880
rect 5740 81248 5780 81257
rect 5740 80669 5780 81208
rect 5932 81080 5972 81089
rect 5836 81040 5932 81080
rect 5739 80660 5781 80669
rect 5739 80620 5740 80660
rect 5780 80620 5781 80660
rect 5739 80611 5781 80620
rect 5451 80324 5493 80333
rect 5451 80284 5452 80324
rect 5492 80284 5493 80324
rect 5451 80275 5493 80284
rect 5252 79705 5396 79736
rect 5212 79696 5396 79705
rect 4684 79687 4724 79696
rect 5356 79568 5396 79577
rect 4928 79400 5296 79409
rect 4968 79360 5010 79400
rect 5050 79360 5092 79400
rect 5132 79360 5174 79400
rect 5214 79360 5256 79400
rect 4928 79351 5296 79360
rect 5259 79148 5301 79157
rect 5259 79108 5260 79148
rect 5300 79108 5301 79148
rect 5259 79099 5301 79108
rect 4875 78896 4917 78905
rect 4875 78856 4876 78896
rect 4916 78856 4917 78896
rect 4875 78847 4917 78856
rect 4396 77498 4436 77507
rect 4492 78184 4588 78224
rect 4492 76805 4532 78184
rect 4588 78175 4628 78184
rect 4876 78149 4916 78847
rect 5260 78569 5300 79099
rect 5259 78560 5301 78569
rect 5259 78520 5260 78560
rect 5300 78520 5301 78560
rect 5259 78511 5301 78520
rect 5356 78401 5396 79528
rect 5452 79325 5492 80275
rect 5548 79997 5588 80536
rect 5547 79988 5589 79997
rect 5547 79948 5548 79988
rect 5588 79948 5589 79988
rect 5547 79939 5589 79948
rect 5548 79736 5588 79745
rect 5548 79409 5588 79696
rect 5547 79400 5589 79409
rect 5547 79360 5548 79400
rect 5588 79360 5589 79400
rect 5547 79351 5589 79360
rect 5451 79316 5493 79325
rect 5451 79276 5452 79316
rect 5492 79276 5493 79316
rect 5451 79267 5493 79276
rect 5548 79157 5588 79351
rect 5836 79316 5876 81040
rect 5932 81031 5972 81040
rect 6028 80660 6068 83476
rect 6604 83516 6644 83525
rect 6507 83096 6549 83105
rect 6507 83056 6508 83096
rect 6548 83056 6549 83096
rect 6507 83047 6549 83056
rect 6315 81752 6357 81761
rect 6315 81712 6316 81752
rect 6356 81712 6357 81752
rect 6315 81703 6357 81712
rect 6124 81248 6164 81257
rect 6164 81208 6260 81248
rect 6124 81199 6164 81208
rect 6028 80620 6164 80660
rect 5932 80492 5972 80503
rect 5932 80417 5972 80452
rect 6027 80492 6069 80501
rect 6027 80452 6028 80492
rect 6068 80452 6069 80492
rect 6027 80443 6069 80452
rect 5931 80408 5973 80417
rect 5931 80368 5932 80408
rect 5972 80368 5973 80408
rect 5931 80359 5973 80368
rect 6028 80358 6068 80443
rect 5644 79276 5876 79316
rect 5547 79148 5589 79157
rect 5547 79108 5548 79148
rect 5588 79108 5589 79148
rect 5547 79099 5589 79108
rect 5451 79064 5493 79073
rect 5451 79024 5452 79064
rect 5492 79024 5493 79064
rect 5451 79015 5493 79024
rect 5355 78392 5397 78401
rect 5355 78352 5356 78392
rect 5396 78352 5397 78392
rect 5355 78343 5397 78352
rect 5164 78224 5204 78233
rect 5452 78224 5492 79015
rect 5644 78980 5684 79276
rect 5931 79232 5973 79241
rect 5931 79192 5932 79232
rect 5972 79192 5973 79232
rect 5931 79183 5973 79192
rect 5836 79073 5876 79158
rect 5932 79098 5972 79183
rect 5835 79064 5877 79073
rect 5835 79024 5836 79064
rect 5876 79024 5877 79064
rect 5835 79015 5877 79024
rect 6028 79064 6068 79073
rect 5204 78184 5492 78224
rect 5548 78940 5684 78980
rect 5164 78175 5204 78184
rect 4875 78140 4917 78149
rect 4875 78100 4876 78140
rect 4916 78100 4917 78140
rect 4875 78091 4917 78100
rect 4972 78065 5012 78150
rect 4780 78056 4820 78065
rect 4684 78016 4780 78056
rect 4588 77636 4628 77645
rect 4588 76889 4628 77596
rect 4587 76880 4629 76889
rect 4587 76840 4588 76880
rect 4628 76840 4629 76880
rect 4587 76831 4629 76840
rect 4491 76796 4533 76805
rect 4491 76756 4492 76796
rect 4532 76756 4533 76796
rect 4491 76747 4533 76756
rect 4395 76712 4437 76721
rect 4395 76672 4396 76712
rect 4436 76672 4437 76712
rect 4395 76663 4437 76672
rect 4396 76578 4436 76663
rect 4395 76040 4437 76049
rect 4395 76000 4396 76040
rect 4436 76000 4437 76040
rect 4395 75991 4437 76000
rect 4300 75151 4340 75160
rect 4396 75200 4436 75991
rect 4436 75160 4628 75200
rect 4396 75151 4436 75160
rect 4395 75032 4437 75041
rect 4395 74992 4396 75032
rect 4436 74992 4437 75032
rect 4395 74983 4437 74992
rect 4299 74276 4341 74285
rect 4299 74236 4300 74276
rect 4340 74236 4341 74276
rect 4299 74227 4341 74236
rect 4300 74142 4340 74227
rect 4396 73100 4436 74983
rect 4588 73520 4628 75160
rect 4684 73688 4724 78016
rect 4780 78007 4820 78016
rect 4971 78056 5013 78065
rect 4971 78016 4972 78056
rect 5012 78016 5013 78056
rect 4971 78007 5013 78016
rect 4928 77888 5296 77897
rect 4968 77848 5010 77888
rect 5050 77848 5092 77888
rect 5132 77848 5174 77888
rect 5214 77848 5256 77888
rect 4928 77839 5296 77848
rect 5548 77720 5588 78940
rect 5835 78896 5877 78905
rect 5835 78856 5836 78896
rect 5876 78856 5877 78896
rect 5835 78847 5877 78856
rect 5644 78812 5684 78821
rect 5684 78772 5780 78812
rect 5644 78763 5684 78772
rect 5643 78392 5685 78401
rect 5643 78352 5644 78392
rect 5684 78352 5685 78392
rect 5643 78343 5685 78352
rect 5164 77680 5588 77720
rect 5164 77552 5204 77680
rect 5164 77503 5204 77512
rect 5259 77552 5301 77561
rect 5259 77512 5260 77552
rect 5300 77512 5301 77552
rect 5259 77503 5301 77512
rect 5260 76544 5300 77503
rect 5356 76721 5396 77680
rect 5452 77552 5492 77561
rect 5355 76712 5397 76721
rect 5355 76672 5356 76712
rect 5396 76672 5397 76712
rect 5355 76663 5397 76672
rect 5260 76504 5396 76544
rect 4928 76376 5296 76385
rect 4968 76336 5010 76376
rect 5050 76336 5092 76376
rect 5132 76336 5174 76376
rect 5214 76336 5256 76376
rect 4928 76327 5296 76336
rect 5356 76208 5396 76504
rect 5452 76301 5492 77512
rect 5548 77552 5588 77561
rect 5644 77552 5684 78343
rect 5588 77512 5684 77552
rect 5451 76292 5493 76301
rect 5451 76252 5452 76292
rect 5492 76252 5493 76292
rect 5451 76243 5493 76252
rect 5260 76168 5396 76208
rect 4972 76040 5012 76049
rect 4972 75881 5012 76000
rect 5067 76040 5109 76049
rect 5067 76000 5068 76040
rect 5108 76000 5109 76040
rect 5067 75991 5109 76000
rect 5068 75906 5108 75991
rect 4971 75872 5013 75881
rect 4971 75832 4972 75872
rect 5012 75832 5013 75872
rect 4971 75823 5013 75832
rect 4875 75620 4917 75629
rect 4875 75580 4876 75620
rect 4916 75580 4917 75620
rect 4875 75571 4917 75580
rect 4779 75536 4821 75545
rect 4779 75496 4780 75536
rect 4820 75496 4821 75536
rect 4779 75487 4821 75496
rect 4780 75284 4820 75487
rect 4780 74957 4820 75244
rect 4876 75200 4916 75571
rect 5260 75209 5300 76168
rect 5548 76124 5588 77512
rect 5643 76796 5685 76805
rect 5643 76756 5644 76796
rect 5684 76756 5685 76796
rect 5643 76747 5685 76756
rect 5644 76712 5684 76747
rect 5644 76661 5684 76672
rect 5643 76544 5685 76553
rect 5643 76504 5644 76544
rect 5684 76504 5685 76544
rect 5643 76495 5685 76504
rect 5356 76084 5588 76124
rect 5356 75461 5396 76084
rect 5451 75956 5493 75965
rect 5451 75916 5452 75956
rect 5492 75916 5493 75956
rect 5451 75907 5493 75916
rect 5548 75956 5588 75965
rect 5452 75822 5492 75907
rect 5548 75797 5588 75916
rect 5547 75788 5589 75797
rect 5547 75748 5548 75788
rect 5588 75748 5589 75788
rect 5547 75739 5589 75748
rect 5644 75629 5684 76495
rect 5740 76376 5780 78772
rect 5836 77384 5876 78847
rect 6028 77729 6068 79024
rect 6027 77720 6069 77729
rect 6027 77680 6028 77720
rect 6068 77680 6069 77720
rect 6027 77671 6069 77680
rect 6027 77552 6069 77561
rect 6027 77512 6028 77552
rect 6068 77512 6069 77552
rect 6027 77503 6069 77512
rect 6028 77418 6068 77503
rect 5836 77335 5876 77344
rect 6124 77300 6164 80620
rect 6220 80585 6260 81208
rect 6219 80576 6261 80585
rect 6219 80536 6220 80576
rect 6260 80536 6261 80576
rect 6219 80527 6261 80536
rect 6220 79064 6260 80527
rect 6220 79015 6260 79024
rect 5932 77260 6164 77300
rect 5836 76553 5876 76638
rect 5835 76544 5877 76553
rect 5835 76504 5836 76544
rect 5876 76504 5877 76544
rect 5835 76495 5877 76504
rect 5740 76336 5876 76376
rect 5739 76208 5781 76217
rect 5739 76168 5740 76208
rect 5780 76168 5781 76208
rect 5739 76159 5781 76168
rect 5643 75620 5685 75629
rect 5548 75580 5644 75620
rect 5684 75580 5685 75620
rect 5451 75536 5493 75545
rect 5451 75496 5452 75536
rect 5492 75496 5493 75536
rect 5451 75487 5493 75496
rect 5355 75452 5397 75461
rect 5355 75412 5356 75452
rect 5396 75412 5397 75452
rect 5355 75403 5397 75412
rect 4876 75151 4916 75160
rect 5259 75200 5301 75209
rect 5259 75160 5260 75200
rect 5300 75160 5301 75200
rect 5259 75151 5301 75160
rect 5356 75200 5396 75209
rect 4779 74948 4821 74957
rect 4779 74908 4780 74948
rect 4820 74908 4821 74948
rect 4779 74899 4821 74908
rect 4928 74864 5296 74873
rect 4968 74824 5010 74864
rect 5050 74824 5092 74864
rect 5132 74824 5174 74864
rect 5214 74824 5256 74864
rect 4928 74815 5296 74824
rect 5356 73949 5396 75160
rect 5452 74789 5492 75487
rect 5451 74780 5493 74789
rect 5451 74740 5452 74780
rect 5492 74740 5493 74780
rect 5451 74731 5493 74740
rect 5548 74621 5588 75580
rect 5643 75571 5685 75580
rect 5643 75368 5685 75377
rect 5643 75328 5644 75368
rect 5684 75328 5685 75368
rect 5643 75319 5685 75328
rect 5547 74612 5589 74621
rect 5547 74572 5548 74612
rect 5588 74572 5589 74612
rect 5547 74563 5589 74572
rect 5451 74528 5493 74537
rect 5451 74488 5452 74528
rect 5492 74488 5493 74528
rect 5451 74479 5493 74488
rect 5452 74394 5492 74479
rect 5547 74360 5589 74369
rect 5547 74320 5548 74360
rect 5588 74320 5589 74360
rect 5547 74311 5589 74320
rect 5451 74276 5493 74285
rect 5451 74236 5452 74276
rect 5492 74236 5493 74276
rect 5451 74227 5493 74236
rect 5355 73940 5397 73949
rect 5355 73900 5356 73940
rect 5396 73900 5397 73940
rect 5355 73891 5397 73900
rect 5259 73772 5301 73781
rect 5259 73732 5260 73772
rect 5300 73732 5301 73772
rect 5259 73723 5301 73732
rect 5356 73772 5396 73781
rect 5452 73772 5492 74227
rect 5548 74226 5588 74311
rect 5644 74108 5684 75319
rect 5740 75116 5780 76159
rect 5836 75214 5876 76336
rect 5836 75165 5876 75174
rect 5740 75076 5876 75116
rect 5836 74873 5876 75076
rect 5835 74864 5877 74873
rect 5835 74824 5836 74864
rect 5876 74824 5877 74864
rect 5835 74815 5877 74824
rect 5739 74780 5781 74789
rect 5739 74740 5740 74780
rect 5780 74740 5781 74780
rect 5739 74731 5781 74740
rect 5740 74528 5780 74731
rect 5740 74479 5780 74488
rect 5836 74360 5876 74815
rect 5396 73732 5492 73772
rect 5548 74068 5684 74108
rect 5740 74320 5876 74360
rect 5356 73723 5396 73732
rect 4780 73688 4820 73697
rect 4684 73648 4780 73688
rect 4780 73639 4820 73648
rect 4876 73688 4916 73697
rect 4876 73520 4916 73648
rect 5260 73638 5300 73723
rect 4588 73480 4916 73520
rect 4683 73352 4725 73361
rect 4683 73312 4684 73352
rect 4724 73312 4725 73352
rect 4683 73303 4725 73312
rect 4300 73060 4436 73100
rect 4300 73016 4340 73060
rect 4300 72967 4340 72976
rect 4491 73016 4533 73025
rect 4491 72976 4492 73016
rect 4532 72976 4533 73016
rect 4491 72967 4533 72976
rect 4492 72882 4532 72967
rect 4587 72428 4629 72437
rect 4587 72388 4588 72428
rect 4628 72388 4629 72428
rect 4587 72379 4629 72388
rect 4588 72176 4628 72379
rect 4588 72017 4628 72136
rect 4587 72008 4629 72017
rect 4587 71968 4588 72008
rect 4628 71968 4629 72008
rect 4587 71959 4629 71968
rect 4684 71597 4724 73303
rect 4780 71933 4820 73480
rect 4928 73352 5296 73361
rect 4968 73312 5010 73352
rect 5050 73312 5092 73352
rect 5132 73312 5174 73352
rect 5214 73312 5256 73352
rect 4928 73303 5296 73312
rect 5548 73100 5588 74068
rect 5740 74024 5780 74320
rect 5356 73060 5588 73100
rect 5644 73984 5780 74024
rect 4779 71924 4821 71933
rect 4779 71884 4780 71924
rect 4820 71884 4821 71924
rect 4779 71875 4821 71884
rect 4683 71588 4725 71597
rect 4683 71548 4684 71588
rect 4724 71548 4725 71588
rect 4683 71539 4725 71548
rect 4300 71252 4340 71261
rect 4340 71212 4436 71252
rect 4300 71203 4340 71212
rect 4204 70531 4244 70540
rect 4107 69992 4149 70001
rect 4107 69952 4108 69992
rect 4148 69952 4149 69992
rect 4107 69943 4149 69952
rect 4299 69992 4341 70001
rect 4299 69952 4300 69992
rect 4340 69952 4341 69992
rect 4299 69943 4341 69952
rect 3723 69740 3765 69749
rect 3723 69700 3724 69740
rect 3764 69700 3765 69740
rect 3723 69691 3765 69700
rect 3688 69572 4056 69581
rect 3728 69532 3770 69572
rect 3810 69532 3852 69572
rect 3892 69532 3934 69572
rect 3974 69532 4016 69572
rect 3688 69523 4056 69532
rect 3627 69404 3669 69413
rect 3627 69364 3628 69404
rect 3668 69364 3669 69404
rect 3627 69355 3669 69364
rect 3628 69068 3668 69355
rect 3628 69019 3668 69028
rect 4012 69152 4052 69161
rect 4108 69152 4148 69943
rect 4300 69858 4340 69943
rect 4052 69112 4148 69152
rect 3820 68984 3860 68993
rect 3860 68944 3956 68984
rect 3820 68935 3860 68944
rect 3819 68732 3861 68741
rect 3819 68692 3820 68732
rect 3860 68692 3861 68732
rect 3819 68683 3861 68692
rect 3627 68564 3669 68573
rect 3627 68524 3628 68564
rect 3668 68524 3669 68564
rect 3627 68515 3669 68524
rect 3628 68480 3668 68515
rect 3820 68489 3860 68683
rect 3628 68429 3668 68440
rect 3819 68480 3861 68489
rect 3819 68440 3820 68480
rect 3860 68440 3861 68480
rect 3819 68431 3861 68440
rect 3820 68237 3860 68322
rect 3819 68228 3861 68237
rect 3819 68188 3820 68228
rect 3860 68188 3861 68228
rect 3916 68228 3956 68944
rect 4012 68312 4052 69112
rect 4396 68648 4436 71212
rect 4683 70076 4725 70085
rect 4683 70036 4684 70076
rect 4724 70036 4725 70076
rect 4683 70027 4725 70036
rect 4587 69992 4629 70001
rect 4587 69952 4588 69992
rect 4628 69952 4629 69992
rect 4587 69943 4629 69952
rect 4684 69992 4724 70027
rect 4300 68608 4436 68648
rect 4492 69740 4532 69749
rect 4107 68564 4149 68573
rect 4107 68524 4108 68564
rect 4148 68524 4149 68564
rect 4107 68515 4149 68524
rect 4108 68480 4148 68515
rect 4204 68489 4244 68574
rect 4108 68429 4148 68440
rect 4203 68480 4245 68489
rect 4203 68440 4204 68480
rect 4244 68440 4245 68480
rect 4203 68431 4245 68440
rect 4012 68272 4244 68312
rect 3916 68188 4148 68228
rect 3819 68179 3861 68188
rect 3688 68060 4056 68069
rect 3728 68020 3770 68060
rect 3810 68020 3852 68060
rect 3892 68020 3934 68060
rect 3974 68020 4016 68060
rect 3688 68011 4056 68020
rect 4108 67808 4148 68188
rect 4204 68069 4244 68272
rect 4203 68060 4245 68069
rect 4203 68020 4204 68060
rect 4244 68020 4245 68060
rect 4203 68011 4245 68020
rect 3820 67768 4148 67808
rect 3627 67640 3669 67649
rect 3627 67600 3628 67640
rect 3668 67600 3669 67640
rect 3627 67591 3669 67600
rect 3531 67556 3573 67565
rect 3531 67516 3532 67556
rect 3572 67516 3573 67556
rect 3531 67507 3573 67516
rect 3435 67472 3477 67481
rect 3435 67432 3436 67472
rect 3476 67432 3477 67472
rect 3435 67423 3477 67432
rect 3436 66809 3476 67423
rect 3531 67052 3573 67061
rect 3628 67052 3668 67591
rect 3531 67012 3532 67052
rect 3572 67012 3668 67052
rect 3531 67003 3573 67012
rect 3532 66968 3572 67003
rect 3532 66917 3572 66928
rect 3435 66800 3477 66809
rect 3435 66760 3436 66800
rect 3476 66760 3477 66800
rect 3435 66751 3477 66760
rect 3820 66716 3860 67768
rect 3964 67649 4004 67658
rect 4300 67640 4340 68608
rect 4492 68489 4532 69700
rect 4396 68480 4436 68489
rect 4491 68480 4533 68489
rect 4436 68440 4492 68480
rect 4532 68440 4533 68480
rect 4396 68431 4436 68440
rect 4491 68431 4533 68440
rect 4492 68346 4532 68431
rect 4396 68228 4436 68237
rect 4588 68228 4628 69943
rect 4684 69941 4724 69952
rect 4683 69320 4725 69329
rect 4683 69280 4684 69320
rect 4724 69280 4725 69320
rect 4683 69271 4725 69280
rect 4684 68573 4724 69271
rect 4780 68648 4820 71875
rect 4928 71840 5296 71849
rect 4968 71800 5010 71840
rect 5050 71800 5092 71840
rect 5132 71800 5174 71840
rect 5214 71800 5256 71840
rect 4928 71791 5296 71800
rect 5067 71504 5109 71513
rect 5067 71464 5068 71504
rect 5108 71464 5109 71504
rect 5067 71455 5109 71464
rect 5068 70664 5108 71455
rect 5259 71420 5301 71429
rect 5259 71380 5260 71420
rect 5300 71380 5301 71420
rect 5259 71371 5301 71380
rect 5260 70841 5300 71371
rect 5356 71336 5396 73060
rect 5644 72344 5684 73984
rect 5835 73940 5877 73949
rect 5835 73900 5836 73940
rect 5876 73900 5877 73940
rect 5835 73891 5877 73900
rect 5836 73688 5876 73891
rect 5836 73639 5876 73648
rect 5932 73100 5972 77260
rect 6316 77048 6356 81703
rect 6508 80576 6548 83047
rect 6604 81929 6644 83476
rect 6796 83516 6836 83525
rect 6796 83273 6836 83476
rect 7180 83516 7220 83525
rect 6795 83264 6837 83273
rect 6795 83224 6796 83264
rect 6836 83224 6837 83264
rect 6795 83215 6837 83224
rect 6891 82844 6933 82853
rect 6891 82804 6892 82844
rect 6932 82804 6933 82844
rect 6891 82795 6933 82804
rect 6603 81920 6645 81929
rect 6603 81880 6604 81920
rect 6644 81880 6645 81920
rect 6603 81871 6645 81880
rect 6795 80660 6837 80669
rect 6795 80620 6796 80660
rect 6836 80620 6837 80660
rect 6795 80611 6837 80620
rect 6508 80527 6548 80536
rect 6411 80072 6453 80081
rect 6411 80032 6412 80072
rect 6452 80032 6453 80072
rect 6411 80023 6453 80032
rect 6412 78224 6452 80023
rect 6796 79736 6836 80611
rect 6796 79687 6836 79696
rect 6700 78224 6740 78233
rect 6452 78184 6700 78224
rect 6412 78175 6452 78184
rect 6411 77552 6453 77561
rect 6411 77512 6412 77552
rect 6452 77512 6453 77552
rect 6411 77503 6453 77512
rect 6220 77008 6356 77048
rect 6220 76805 6260 77008
rect 6315 76880 6357 76889
rect 6315 76840 6316 76880
rect 6356 76840 6357 76880
rect 6315 76831 6357 76840
rect 6219 76796 6261 76805
rect 6219 76756 6220 76796
rect 6260 76756 6261 76796
rect 6219 76747 6261 76756
rect 6028 76712 6068 76723
rect 6028 76637 6068 76672
rect 6123 76712 6165 76721
rect 6123 76672 6124 76712
rect 6164 76672 6165 76712
rect 6123 76663 6165 76672
rect 6027 76628 6069 76637
rect 6027 76588 6028 76628
rect 6068 76588 6069 76628
rect 6027 76579 6069 76588
rect 6124 76578 6164 76663
rect 6219 76544 6261 76553
rect 6219 76504 6220 76544
rect 6260 76504 6261 76544
rect 6219 76495 6261 76504
rect 6316 76544 6356 76831
rect 6316 76495 6356 76504
rect 6028 76040 6068 76049
rect 6068 76000 6164 76040
rect 6028 75991 6068 76000
rect 6027 75116 6069 75125
rect 6027 75076 6028 75116
rect 6068 75076 6069 75116
rect 6027 75067 6069 75076
rect 6028 74982 6068 75067
rect 5836 73060 5972 73100
rect 5740 73016 5780 73025
rect 5740 72605 5780 72976
rect 5739 72596 5781 72605
rect 5739 72556 5740 72596
rect 5780 72556 5781 72596
rect 5739 72547 5781 72556
rect 5836 72521 5876 73060
rect 5931 72764 5973 72773
rect 5931 72724 5932 72764
rect 5972 72724 5973 72764
rect 5931 72715 5973 72724
rect 5932 72630 5972 72715
rect 6124 72521 6164 76000
rect 6220 75620 6260 76495
rect 6220 75580 6356 75620
rect 6219 75200 6261 75209
rect 6219 75160 6220 75200
rect 6260 75160 6261 75200
rect 6219 75151 6261 75160
rect 5835 72512 5877 72521
rect 5835 72472 5836 72512
rect 5876 72472 5877 72512
rect 5835 72463 5877 72472
rect 6123 72512 6165 72521
rect 6123 72472 6124 72512
rect 6164 72472 6165 72512
rect 6123 72463 6165 72472
rect 5931 72428 5973 72437
rect 5931 72388 5932 72428
rect 5972 72388 5973 72428
rect 5931 72379 5973 72388
rect 5644 72304 5780 72344
rect 5643 72176 5685 72185
rect 5643 72136 5644 72176
rect 5684 72136 5685 72176
rect 5643 72127 5685 72136
rect 5451 72092 5493 72101
rect 5451 72052 5452 72092
rect 5492 72052 5493 72092
rect 5451 72043 5493 72052
rect 5452 71513 5492 72043
rect 5644 71672 5684 72127
rect 5740 72008 5780 72304
rect 5836 72176 5876 72185
rect 5932 72176 5972 72379
rect 6220 72344 6260 75151
rect 6316 73702 6356 75580
rect 6412 74453 6452 77503
rect 6508 76973 6548 78184
rect 6700 78175 6740 78184
rect 6603 77720 6645 77729
rect 6603 77680 6604 77720
rect 6644 77680 6645 77720
rect 6603 77671 6645 77680
rect 6507 76964 6549 76973
rect 6507 76924 6508 76964
rect 6548 76924 6549 76964
rect 6507 76915 6549 76924
rect 6507 76712 6549 76721
rect 6507 76672 6508 76712
rect 6548 76672 6549 76712
rect 6507 76663 6549 76672
rect 6508 76049 6548 76663
rect 6604 76553 6644 77671
rect 6892 77561 6932 82795
rect 7180 81920 7220 83476
rect 7371 83432 7413 83441
rect 7371 83392 7372 83432
rect 7412 83392 7413 83432
rect 7371 83383 7413 83392
rect 7372 83298 7412 83383
rect 7660 83264 7700 84400
rect 7756 83777 7796 85936
rect 7948 84776 7988 85936
rect 7948 84736 8084 84776
rect 7755 83768 7797 83777
rect 7755 83728 7756 83768
rect 7796 83728 7797 83768
rect 7755 83719 7797 83728
rect 7755 83516 7797 83525
rect 7755 83476 7756 83516
rect 7796 83476 7797 83516
rect 7755 83467 7797 83476
rect 7756 83382 7796 83467
rect 7948 83348 7988 83357
rect 7948 83264 7988 83308
rect 7660 83224 7988 83264
rect 8044 83189 8084 84736
rect 8140 83777 8180 85936
rect 8332 84365 8372 85936
rect 8331 84356 8373 84365
rect 8331 84316 8332 84356
rect 8372 84316 8373 84356
rect 8331 84307 8373 84316
rect 8331 84188 8373 84197
rect 8331 84148 8332 84188
rect 8372 84148 8373 84188
rect 8331 84139 8373 84148
rect 8139 83768 8181 83777
rect 8139 83728 8140 83768
rect 8180 83728 8181 83768
rect 8139 83719 8181 83728
rect 8140 83516 8180 83525
rect 8140 83273 8180 83476
rect 8139 83264 8181 83273
rect 8139 83224 8140 83264
rect 8180 83224 8181 83264
rect 8139 83215 8181 83224
rect 7467 83180 7509 83189
rect 7467 83140 7468 83180
rect 7508 83140 7509 83180
rect 7467 83131 7509 83140
rect 8043 83180 8085 83189
rect 8043 83140 8044 83180
rect 8084 83140 8085 83180
rect 8043 83131 8085 83140
rect 7468 83012 7508 83131
rect 7468 82963 7508 82972
rect 7275 82844 7317 82853
rect 7275 82804 7276 82844
rect 7316 82804 7317 82844
rect 7275 82795 7317 82804
rect 7276 82710 7316 82795
rect 7947 82760 7989 82769
rect 7947 82720 7948 82760
rect 7988 82720 7989 82760
rect 7947 82711 7989 82720
rect 7180 81880 7316 81920
rect 6987 81080 7029 81089
rect 6987 81040 6988 81080
rect 7028 81040 7029 81080
rect 6987 81031 7029 81040
rect 6988 80571 7028 81031
rect 7180 80660 7220 80669
rect 6988 80522 7028 80531
rect 7084 80620 7180 80660
rect 6988 79568 7028 79577
rect 6988 79073 7028 79528
rect 6987 79064 7029 79073
rect 6987 79024 6988 79064
rect 7028 79024 7029 79064
rect 6987 79015 7029 79024
rect 6988 78821 7028 79015
rect 6987 78812 7029 78821
rect 6987 78772 6988 78812
rect 7028 78772 7029 78812
rect 6987 78763 7029 78772
rect 6891 77552 6933 77561
rect 6891 77512 6892 77552
rect 6932 77512 6933 77552
rect 6891 77503 6933 77512
rect 6699 77216 6741 77225
rect 6699 77176 6700 77216
rect 6740 77176 6741 77216
rect 6699 77167 6741 77176
rect 6700 76712 6740 77167
rect 7084 77048 7124 80620
rect 7180 80611 7220 80620
rect 7276 79820 7316 81880
rect 7371 81752 7413 81761
rect 7371 81712 7372 81752
rect 7412 81712 7413 81752
rect 7371 81703 7413 81712
rect 7372 81341 7412 81703
rect 7371 81332 7413 81341
rect 7371 81292 7372 81332
rect 7412 81292 7413 81332
rect 7371 81283 7413 81292
rect 7372 81248 7412 81283
rect 7372 81198 7412 81208
rect 7563 81080 7605 81089
rect 7563 81040 7564 81080
rect 7604 81040 7605 81080
rect 7563 81031 7605 81040
rect 7564 80946 7604 81031
rect 7276 79771 7316 79780
rect 7180 79736 7220 79745
rect 7180 79241 7220 79696
rect 7372 79736 7412 79745
rect 7275 79316 7317 79325
rect 7275 79276 7276 79316
rect 7316 79276 7317 79316
rect 7275 79267 7317 79276
rect 7179 79232 7221 79241
rect 7179 79192 7180 79232
rect 7220 79192 7221 79232
rect 7179 79183 7221 79192
rect 7179 78224 7221 78233
rect 7179 78184 7180 78224
rect 7220 78184 7221 78224
rect 7179 78175 7221 78184
rect 7180 77552 7220 78175
rect 7276 77888 7316 79267
rect 7372 79241 7412 79696
rect 7948 79736 7988 82711
rect 7948 79687 7988 79696
rect 8043 79316 8085 79325
rect 8043 79276 8044 79316
rect 8084 79276 8085 79316
rect 8043 79267 8085 79276
rect 7371 79232 7413 79241
rect 7371 79192 7372 79232
rect 7412 79192 7413 79232
rect 7371 79183 7413 79192
rect 7947 79232 7989 79241
rect 7947 79192 7948 79232
rect 7988 79192 7989 79232
rect 7947 79183 7989 79192
rect 7948 79098 7988 79183
rect 7467 79064 7509 79073
rect 7852 79064 7892 79073
rect 7467 79024 7468 79064
rect 7508 79024 7509 79064
rect 7467 79015 7509 79024
rect 7564 79024 7852 79064
rect 7468 78233 7508 79015
rect 7467 78224 7509 78233
rect 7467 78184 7468 78224
rect 7508 78184 7509 78224
rect 7467 78175 7509 78184
rect 7276 77848 7412 77888
rect 7276 77552 7316 77561
rect 7180 77512 7276 77552
rect 7276 77225 7316 77512
rect 7275 77216 7317 77225
rect 7275 77176 7276 77216
rect 7316 77176 7317 77216
rect 7275 77167 7317 77176
rect 6603 76544 6645 76553
rect 6603 76504 6604 76544
rect 6644 76504 6645 76544
rect 6603 76495 6645 76504
rect 6700 76469 6740 76672
rect 6796 77008 7124 77048
rect 7275 77048 7317 77057
rect 7275 77008 7276 77048
rect 7316 77008 7317 77048
rect 6699 76460 6741 76469
rect 6699 76420 6700 76460
rect 6740 76420 6741 76460
rect 6699 76411 6741 76420
rect 6699 76208 6741 76217
rect 6699 76168 6700 76208
rect 6740 76168 6741 76208
rect 6699 76159 6741 76168
rect 6603 76124 6645 76133
rect 6603 76084 6604 76124
rect 6644 76084 6645 76124
rect 6603 76075 6645 76084
rect 6507 76040 6549 76049
rect 6507 75995 6508 76040
rect 6548 75995 6549 76040
rect 6507 75991 6549 75995
rect 6508 75906 6548 75991
rect 6507 75620 6549 75629
rect 6507 75580 6508 75620
rect 6548 75580 6549 75620
rect 6507 75571 6549 75580
rect 6411 74444 6453 74453
rect 6411 74404 6412 74444
rect 6452 74404 6453 74444
rect 6411 74395 6453 74404
rect 6411 74276 6453 74285
rect 6411 74236 6412 74276
rect 6452 74236 6453 74276
rect 6411 74227 6453 74236
rect 6412 73781 6452 74227
rect 6411 73772 6453 73781
rect 6411 73732 6412 73772
rect 6452 73732 6453 73772
rect 6411 73723 6453 73732
rect 6316 73653 6356 73662
rect 6315 73436 6357 73445
rect 6315 73396 6316 73436
rect 6356 73396 6357 73436
rect 6315 73387 6357 73396
rect 6316 73016 6356 73387
rect 6316 72967 6356 72976
rect 6315 72764 6357 72773
rect 6315 72724 6316 72764
rect 6356 72724 6357 72764
rect 6315 72715 6357 72724
rect 5876 72136 5972 72176
rect 6124 72304 6260 72344
rect 5836 72127 5876 72136
rect 6028 72008 6068 72017
rect 5740 71968 5876 72008
rect 5644 71623 5684 71632
rect 5446 71504 5492 71513
rect 5446 71464 5447 71504
rect 5446 71455 5492 71464
rect 5547 71504 5589 71513
rect 5547 71464 5548 71504
rect 5588 71464 5589 71504
rect 5547 71455 5589 71464
rect 5740 71504 5780 71515
rect 5548 71370 5588 71455
rect 5740 71429 5780 71464
rect 5739 71420 5781 71429
rect 5739 71380 5740 71420
rect 5780 71380 5781 71420
rect 5739 71371 5781 71380
rect 5356 71296 5492 71336
rect 5259 70832 5301 70841
rect 5259 70792 5260 70832
rect 5300 70792 5301 70832
rect 5259 70783 5301 70792
rect 5164 70673 5204 70758
rect 5068 70615 5108 70624
rect 5163 70664 5205 70673
rect 5163 70624 5164 70664
rect 5204 70624 5205 70664
rect 5163 70615 5205 70624
rect 5355 70664 5397 70673
rect 5355 70624 5356 70664
rect 5396 70624 5397 70664
rect 5355 70615 5397 70624
rect 4928 70328 5296 70337
rect 4968 70288 5010 70328
rect 5050 70288 5092 70328
rect 5132 70288 5174 70328
rect 5214 70288 5256 70328
rect 4928 70279 5296 70288
rect 5260 69152 5300 69163
rect 5260 69077 5300 69112
rect 5259 69068 5301 69077
rect 5259 69028 5260 69068
rect 5300 69028 5301 69068
rect 5259 69019 5301 69028
rect 4928 68816 5296 68825
rect 4968 68776 5010 68816
rect 5050 68776 5092 68816
rect 5132 68776 5174 68816
rect 5214 68776 5256 68816
rect 4928 68767 5296 68776
rect 5163 68648 5205 68657
rect 4780 68608 4916 68648
rect 4683 68564 4725 68573
rect 4683 68524 4684 68564
rect 4724 68524 4725 68564
rect 4683 68515 4725 68524
rect 4684 68480 4724 68515
rect 4684 68430 4724 68440
rect 4780 68480 4820 68489
rect 4436 68188 4628 68228
rect 4396 68179 4436 68188
rect 4491 68060 4533 68069
rect 4491 68020 4492 68060
rect 4532 68020 4533 68060
rect 4491 68011 4533 68020
rect 4492 67649 4532 68011
rect 4587 67892 4629 67901
rect 4587 67852 4588 67892
rect 4628 67852 4629 67892
rect 4587 67843 4629 67852
rect 4004 67609 4340 67640
rect 3964 67600 4340 67609
rect 4491 67640 4533 67649
rect 4491 67600 4492 67640
rect 4532 67600 4533 67640
rect 4491 67591 4533 67600
rect 4107 67472 4149 67481
rect 4300 67472 4340 67481
rect 4107 67432 4108 67472
rect 4148 67432 4149 67472
rect 4107 67423 4149 67432
rect 4204 67432 4300 67472
rect 4108 67338 4148 67423
rect 3532 66676 3860 66716
rect 3532 66380 3572 66676
rect 3688 66548 4056 66557
rect 3728 66508 3770 66548
rect 3810 66508 3852 66548
rect 3892 66508 3934 66548
rect 3974 66508 4016 66548
rect 3688 66499 4056 66508
rect 3532 66340 3764 66380
rect 3724 66221 3764 66340
rect 4204 66296 4244 67432
rect 4300 67423 4340 67432
rect 4492 66809 4532 67591
rect 4588 66884 4628 67843
rect 4780 67136 4820 68440
rect 4876 67901 4916 68608
rect 5163 68608 5164 68648
rect 5204 68608 5205 68648
rect 5163 68599 5205 68608
rect 5164 68480 5204 68599
rect 5164 68431 5204 68440
rect 5260 68396 5300 68405
rect 5260 67901 5300 68356
rect 4875 67892 4917 67901
rect 4875 67852 4876 67892
rect 4916 67852 4917 67892
rect 4875 67843 4917 67852
rect 5259 67892 5301 67901
rect 5259 67852 5260 67892
rect 5300 67852 5301 67892
rect 5259 67843 5301 67852
rect 4928 67304 5296 67313
rect 4968 67264 5010 67304
rect 5050 67264 5092 67304
rect 5132 67264 5174 67304
rect 5214 67264 5256 67304
rect 4928 67255 5296 67264
rect 5356 67229 5396 70615
rect 5452 69488 5492 71296
rect 5836 71000 5876 71968
rect 5931 71588 5973 71597
rect 5931 71548 5932 71588
rect 5972 71548 5973 71588
rect 5931 71539 5973 71548
rect 5932 71504 5972 71539
rect 5932 71453 5972 71464
rect 6028 71429 6068 71968
rect 6027 71420 6069 71429
rect 6027 71380 6028 71420
rect 6068 71380 6069 71420
rect 6027 71371 6069 71380
rect 5644 70960 5876 71000
rect 5644 70748 5684 70960
rect 5739 70832 5781 70841
rect 5739 70792 5740 70832
rect 5780 70792 5781 70832
rect 5739 70783 5781 70792
rect 5644 70699 5684 70708
rect 5548 70664 5588 70673
rect 5548 69665 5588 70624
rect 5643 70076 5685 70085
rect 5643 70036 5644 70076
rect 5684 70036 5685 70076
rect 5643 70027 5685 70036
rect 5547 69656 5589 69665
rect 5547 69616 5548 69656
rect 5588 69616 5589 69656
rect 5547 69607 5589 69616
rect 5452 69448 5588 69488
rect 5451 69320 5493 69329
rect 5451 69280 5452 69320
rect 5492 69280 5493 69320
rect 5451 69271 5493 69280
rect 5452 69186 5492 69271
rect 5451 69068 5493 69077
rect 5548 69068 5588 69448
rect 5451 69028 5452 69068
rect 5492 69028 5588 69068
rect 5644 69152 5684 70027
rect 5451 69019 5493 69028
rect 5355 67220 5397 67229
rect 5355 67180 5356 67220
rect 5396 67180 5397 67220
rect 5355 67171 5397 67180
rect 4780 67096 4916 67136
rect 4780 66968 4820 66977
rect 4588 66844 4724 66884
rect 4491 66800 4533 66809
rect 4491 66760 4492 66800
rect 4532 66760 4533 66800
rect 4491 66751 4533 66760
rect 4395 66716 4437 66725
rect 4395 66676 4396 66716
rect 4436 66676 4437 66716
rect 4395 66667 4437 66676
rect 4299 66380 4341 66389
rect 4299 66340 4300 66380
rect 4340 66340 4341 66380
rect 4299 66331 4341 66340
rect 4108 66256 4244 66296
rect 3723 66212 3765 66221
rect 3723 66172 3724 66212
rect 3764 66172 3765 66212
rect 3723 66163 3765 66172
rect 3532 66128 3572 66139
rect 3532 66053 3572 66088
rect 3627 66128 3669 66137
rect 3627 66088 3628 66128
rect 3668 66088 3669 66128
rect 3627 66079 3669 66088
rect 3724 66128 3764 66163
rect 4108 66137 4148 66256
rect 3531 66044 3573 66053
rect 3531 66004 3532 66044
rect 3572 66004 3573 66044
rect 3531 65995 3573 66004
rect 3628 65994 3668 66079
rect 3724 66078 3764 66088
rect 3915 66128 3957 66137
rect 3915 66088 3916 66128
rect 3956 66088 3957 66128
rect 3915 66079 3957 66088
rect 4012 66128 4052 66137
rect 3916 65994 3956 66079
rect 3436 65960 3476 65969
rect 3339 65708 3381 65717
rect 3339 65668 3340 65708
rect 3380 65668 3381 65708
rect 3339 65659 3381 65668
rect 3339 65540 3381 65549
rect 3339 65500 3340 65540
rect 3380 65500 3381 65540
rect 3339 65491 3381 65500
rect 3340 65406 3380 65491
rect 3436 65465 3476 65920
rect 4012 65717 4052 66088
rect 4107 66128 4149 66137
rect 4107 66088 4108 66128
rect 4148 66088 4149 66128
rect 4107 66079 4149 66088
rect 4204 66128 4244 66137
rect 4300 66128 4340 66331
rect 4244 66088 4340 66128
rect 4108 65994 4148 66079
rect 4204 65801 4244 66088
rect 4203 65792 4245 65801
rect 4203 65752 4204 65792
rect 4244 65752 4245 65792
rect 4203 65743 4245 65752
rect 3531 65708 3573 65717
rect 3531 65668 3532 65708
rect 3572 65668 3573 65708
rect 3531 65659 3573 65668
rect 4011 65708 4053 65717
rect 4011 65668 4012 65708
rect 4052 65668 4053 65708
rect 4011 65659 4053 65668
rect 3435 65456 3477 65465
rect 3435 65416 3436 65456
rect 3476 65416 3477 65456
rect 3435 65407 3477 65416
rect 3532 65381 3572 65659
rect 4300 65456 4340 65467
rect 4300 65381 4340 65416
rect 3531 65372 3573 65381
rect 4299 65372 4341 65381
rect 3531 65332 3532 65372
rect 3572 65332 3573 65372
rect 3531 65323 3573 65332
rect 4204 65332 4300 65372
rect 4340 65332 4341 65372
rect 3531 65204 3573 65213
rect 3531 65164 3532 65204
rect 3572 65164 3573 65204
rect 3531 65155 3573 65164
rect 3532 64625 3572 65155
rect 3688 65036 4056 65045
rect 3728 64996 3770 65036
rect 3810 64996 3852 65036
rect 3892 64996 3934 65036
rect 3974 64996 4016 65036
rect 3688 64987 4056 64996
rect 4011 64700 4053 64709
rect 4011 64660 4012 64700
rect 4052 64660 4053 64700
rect 4011 64651 4053 64660
rect 3531 64616 3573 64625
rect 3531 64576 3532 64616
rect 3572 64576 3573 64616
rect 3531 64567 3573 64576
rect 3244 64492 3476 64532
rect 3243 64364 3285 64373
rect 3243 64324 3244 64364
rect 3284 64324 3285 64364
rect 3243 64315 3285 64324
rect 3147 63944 3189 63953
rect 3147 63904 3148 63944
rect 3188 63904 3189 63944
rect 3147 63895 3189 63904
rect 3051 63020 3093 63029
rect 3051 62980 3052 63020
rect 3092 62980 3093 63020
rect 3051 62971 3093 62980
rect 2860 62896 2996 62936
rect 2763 62768 2805 62777
rect 2763 62728 2764 62768
rect 2804 62728 2805 62768
rect 2763 62719 2805 62728
rect 2668 60929 2708 61636
rect 2764 61592 2804 61601
rect 2764 61013 2804 61552
rect 2763 61004 2805 61013
rect 2763 60964 2764 61004
rect 2804 60964 2805 61004
rect 2763 60955 2805 60964
rect 2667 60920 2709 60929
rect 2667 60880 2668 60920
rect 2708 60880 2709 60920
rect 2667 60871 2709 60880
rect 2860 60920 2900 62896
rect 3051 62768 3093 62777
rect 3051 62728 3052 62768
rect 3092 62728 3093 62768
rect 3051 62719 3093 62728
rect 2956 62432 2996 62441
rect 2956 61097 2996 62392
rect 2955 61088 2997 61097
rect 2955 61048 2956 61088
rect 2996 61048 2997 61088
rect 2955 61039 2997 61048
rect 2860 60871 2900 60880
rect 2956 60920 2996 60929
rect 2956 60425 2996 60880
rect 2955 60416 2997 60425
rect 2955 60376 2956 60416
rect 2996 60376 2997 60416
rect 2955 60367 2997 60376
rect 3052 60248 3092 62719
rect 3148 62348 3188 63895
rect 3244 63188 3284 64315
rect 3340 63944 3380 63953
rect 3340 63365 3380 63904
rect 3339 63356 3381 63365
rect 3339 63316 3340 63356
rect 3380 63316 3381 63356
rect 3339 63307 3381 63316
rect 3244 63139 3284 63148
rect 3339 63188 3381 63197
rect 3339 63148 3340 63188
rect 3380 63148 3381 63188
rect 3339 63139 3381 63148
rect 3340 63054 3380 63139
rect 3148 62308 3380 62348
rect 3147 62180 3189 62189
rect 3147 62140 3148 62180
rect 3188 62140 3189 62180
rect 3147 62131 3189 62140
rect 3148 62046 3188 62131
rect 3243 61676 3285 61685
rect 3243 61636 3244 61676
rect 3284 61636 3285 61676
rect 3243 61627 3285 61636
rect 3244 61592 3284 61627
rect 3244 61541 3284 61552
rect 3147 61256 3189 61265
rect 3147 61216 3148 61256
rect 3188 61216 3189 61256
rect 3147 61207 3189 61216
rect 2764 60208 3092 60248
rect 2668 60080 2708 60089
rect 2668 59837 2708 60040
rect 2667 59828 2709 59837
rect 2667 59788 2668 59828
rect 2708 59788 2709 59828
rect 2667 59779 2709 59788
rect 2764 59660 2804 60208
rect 3052 60038 3092 60047
rect 2955 59996 2997 60005
rect 3052 59996 3092 59998
rect 2955 59956 2956 59996
rect 2996 59956 3092 59996
rect 2955 59947 2997 59956
rect 2859 59912 2901 59921
rect 3148 59912 3188 61207
rect 3340 61004 3380 62308
rect 3436 61853 3476 64492
rect 3532 64482 3572 64567
rect 3819 64112 3861 64121
rect 3819 64072 3820 64112
rect 3860 64072 3861 64112
rect 3819 64063 3861 64072
rect 4012 64112 4052 64651
rect 4204 64280 4244 65332
rect 4299 65323 4341 65332
rect 4396 64952 4436 66667
rect 4491 66212 4533 66221
rect 4491 66172 4492 66212
rect 4532 66172 4533 66212
rect 4491 66163 4533 66172
rect 4492 66128 4532 66163
rect 4492 65381 4532 66088
rect 4588 66128 4628 66137
rect 4491 65372 4533 65381
rect 4491 65332 4492 65372
rect 4532 65332 4533 65372
rect 4491 65323 4533 65332
rect 4012 64063 4052 64072
rect 4108 64240 4244 64280
rect 4300 64912 4436 64952
rect 3820 63939 3860 64063
rect 3820 63890 3860 63899
rect 3688 63524 4056 63533
rect 3728 63484 3770 63524
rect 3810 63484 3852 63524
rect 3892 63484 3934 63524
rect 3974 63484 4016 63524
rect 3688 63475 4056 63484
rect 3723 63356 3765 63365
rect 3723 63316 3724 63356
rect 3764 63316 3765 63356
rect 3723 63307 3765 63316
rect 3531 63272 3573 63281
rect 3531 63232 3532 63272
rect 3572 63232 3573 63272
rect 3531 63223 3573 63232
rect 3435 61844 3477 61853
rect 3435 61804 3436 61844
rect 3476 61804 3477 61844
rect 3435 61795 3477 61804
rect 2859 59872 2860 59912
rect 2900 59872 2901 59912
rect 2859 59863 2901 59872
rect 3052 59872 3188 59912
rect 3244 60964 3380 61004
rect 2860 59778 2900 59863
rect 2955 59828 2997 59837
rect 2955 59788 2956 59828
rect 2996 59788 2997 59828
rect 2955 59779 2997 59788
rect 2764 59620 2900 59660
rect 2667 59492 2709 59501
rect 2667 59452 2668 59492
rect 2708 59452 2709 59492
rect 2667 59443 2709 59452
rect 2572 59359 2612 59368
rect 2668 59408 2708 59443
rect 2668 59357 2708 59368
rect 2091 59324 2133 59333
rect 2091 59284 2092 59324
rect 2132 59284 2133 59324
rect 2091 59275 2133 59284
rect 2571 58736 2613 58745
rect 2571 58696 2572 58736
rect 2612 58696 2613 58736
rect 2571 58687 2613 58696
rect 1996 58612 2516 58652
rect 2092 57896 2132 58612
rect 2476 58568 2516 58612
rect 2476 58519 2516 58528
rect 2092 57847 2132 57856
rect 1900 57644 1940 57653
rect 1940 57604 2324 57644
rect 1900 57595 1940 57604
rect 1803 57560 1845 57569
rect 1803 57520 1804 57560
rect 1844 57520 1845 57560
rect 1803 57511 1845 57520
rect 1804 57308 1844 57511
rect 1804 57259 1844 57268
rect 1900 57268 2228 57308
rect 1900 57140 1940 57268
rect 1708 57100 1940 57140
rect 1611 56552 1653 56561
rect 1611 56512 1612 56552
rect 1652 56512 1653 56552
rect 1611 56503 1653 56512
rect 1460 55504 1556 55544
rect 1323 53948 1365 53957
rect 1228 53908 1324 53948
rect 1364 53908 1365 53948
rect 1323 53899 1365 53908
rect 1132 53740 1364 53780
rect 747 52940 789 52949
rect 747 52900 748 52940
rect 788 52900 789 52940
rect 747 52891 789 52900
rect 1324 52856 1364 53740
rect 1228 52816 1364 52856
rect 1228 51353 1268 52816
rect 1323 52688 1365 52697
rect 1323 52648 1324 52688
rect 1364 52648 1365 52688
rect 1323 52639 1365 52648
rect 1227 51344 1269 51353
rect 1227 51304 1228 51344
rect 1268 51304 1269 51344
rect 1227 51295 1269 51304
rect 1228 51008 1268 51295
rect 1228 50959 1268 50968
rect 1228 48824 1268 48833
rect 1228 48665 1268 48784
rect 1227 48656 1269 48665
rect 1227 48616 1228 48656
rect 1268 48616 1269 48656
rect 1227 48607 1269 48616
rect 1228 46472 1268 46481
rect 1228 46313 1268 46432
rect 1227 46304 1269 46313
rect 1227 46264 1228 46304
rect 1268 46264 1269 46304
rect 1227 46255 1269 46264
rect 1227 45800 1269 45809
rect 1227 45760 1228 45800
rect 1268 45760 1269 45800
rect 1227 45751 1269 45760
rect 1228 44960 1268 45751
rect 1324 45044 1364 52639
rect 1420 52613 1460 55504
rect 1516 53369 1556 53454
rect 1515 53360 1557 53369
rect 1515 53320 1516 53360
rect 1556 53320 1557 53360
rect 1515 53311 1557 53320
rect 1612 53192 1652 56503
rect 1804 54620 1844 54629
rect 1707 53864 1749 53873
rect 1707 53824 1708 53864
rect 1748 53824 1749 53864
rect 1707 53815 1749 53824
rect 1516 53152 1652 53192
rect 1419 52604 1461 52613
rect 1419 52564 1420 52604
rect 1460 52564 1461 52604
rect 1419 52555 1461 52564
rect 1420 52352 1460 52361
rect 1516 52352 1556 53152
rect 1708 52772 1748 53815
rect 1804 53537 1844 54580
rect 1803 53528 1845 53537
rect 1803 53488 1804 53528
rect 1844 53488 1845 53528
rect 1803 53479 1845 53488
rect 1900 52781 1940 57100
rect 1996 57140 2036 57149
rect 1996 55133 2036 57100
rect 2188 57056 2228 57268
rect 2188 57007 2228 57016
rect 2091 55712 2133 55721
rect 2091 55672 2092 55712
rect 2132 55672 2133 55712
rect 2091 55663 2133 55672
rect 1995 55124 2037 55133
rect 1995 55084 1996 55124
rect 2036 55084 2037 55124
rect 1995 55075 2037 55084
rect 1995 54788 2037 54797
rect 1995 54748 1996 54788
rect 2036 54748 2037 54788
rect 1995 54739 2037 54748
rect 1996 54654 2036 54739
rect 1804 52772 1844 52781
rect 1708 52732 1804 52772
rect 1804 52723 1844 52732
rect 1899 52772 1941 52781
rect 1899 52732 1900 52772
rect 1940 52732 1941 52772
rect 1899 52723 1941 52732
rect 1612 52648 1748 52688
rect 1612 52604 1652 52648
rect 1708 52604 1748 52648
rect 1995 52604 2037 52613
rect 1708 52564 1940 52604
rect 1612 52555 1652 52564
rect 1803 52436 1845 52445
rect 1803 52396 1804 52436
rect 1844 52396 1845 52436
rect 1803 52387 1845 52396
rect 1707 52352 1749 52361
rect 1516 52312 1652 52352
rect 1420 52193 1460 52312
rect 1419 52184 1461 52193
rect 1419 52144 1420 52184
rect 1460 52144 1461 52184
rect 1419 52135 1461 52144
rect 1419 51932 1461 51941
rect 1419 51892 1420 51932
rect 1460 51892 1461 51932
rect 1419 51883 1461 51892
rect 1420 50336 1460 51883
rect 1516 51596 1556 51605
rect 1516 50849 1556 51556
rect 1515 50840 1557 50849
rect 1515 50800 1516 50840
rect 1556 50800 1557 50840
rect 1515 50791 1557 50800
rect 1515 50420 1557 50429
rect 1515 50380 1516 50420
rect 1556 50380 1557 50420
rect 1515 50371 1557 50380
rect 1420 50287 1460 50296
rect 1516 49664 1556 50371
rect 1420 49624 1556 49664
rect 1420 47993 1460 49624
rect 1515 49496 1557 49505
rect 1515 49456 1516 49496
rect 1556 49456 1557 49496
rect 1515 49447 1557 49456
rect 1516 49328 1556 49447
rect 1516 49279 1556 49288
rect 1515 48488 1557 48497
rect 1515 48448 1516 48488
rect 1556 48448 1557 48488
rect 1515 48439 1557 48448
rect 1419 47984 1461 47993
rect 1419 47944 1420 47984
rect 1460 47944 1461 47984
rect 1419 47935 1461 47944
rect 1516 46976 1556 48439
rect 1612 48236 1652 52312
rect 1707 52312 1708 52352
rect 1748 52312 1749 52352
rect 1707 52303 1749 52312
rect 1708 51764 1748 52303
rect 1708 51715 1748 51724
rect 1804 49748 1844 52387
rect 1900 51773 1940 52564
rect 1995 52564 1996 52604
rect 2036 52564 2037 52604
rect 1995 52555 2037 52564
rect 1996 52470 2036 52555
rect 2092 52361 2132 55663
rect 2188 54956 2228 54965
rect 2188 52697 2228 54916
rect 2284 54872 2324 57604
rect 2572 56384 2612 58687
rect 2668 58400 2708 58409
rect 2708 58360 2804 58400
rect 2668 58351 2708 58360
rect 2764 56393 2804 58360
rect 2860 56561 2900 59620
rect 2956 57065 2996 59779
rect 3052 59408 3092 59872
rect 3052 59359 3092 59368
rect 3148 59408 3188 59417
rect 3244 59408 3284 60964
rect 3435 60920 3477 60929
rect 3435 60880 3436 60920
rect 3476 60880 3477 60920
rect 3435 60871 3477 60880
rect 3340 60836 3380 60845
rect 3340 60593 3380 60796
rect 3436 60786 3476 60871
rect 3339 60584 3381 60593
rect 3339 60544 3340 60584
rect 3380 60544 3381 60584
rect 3339 60535 3381 60544
rect 3339 59996 3381 60005
rect 3339 59956 3340 59996
rect 3380 59956 3381 59996
rect 3339 59947 3381 59956
rect 3188 59368 3284 59408
rect 3148 59359 3188 59368
rect 3340 58661 3380 59947
rect 3339 58652 3381 58661
rect 3339 58612 3340 58652
rect 3380 58612 3381 58652
rect 3339 58603 3381 58612
rect 3340 57896 3380 58603
rect 3340 57847 3380 57856
rect 3532 57728 3572 63223
rect 3724 63104 3764 63307
rect 3820 63104 3860 63113
rect 3724 63064 3820 63104
rect 3724 62777 3764 63064
rect 3820 63055 3860 63064
rect 3723 62768 3765 62777
rect 3723 62728 3724 62768
rect 3764 62728 3765 62768
rect 3723 62719 3765 62728
rect 3688 62012 4056 62021
rect 3728 61972 3770 62012
rect 3810 61972 3852 62012
rect 3892 61972 3934 62012
rect 3974 61972 4016 62012
rect 3688 61963 4056 61972
rect 3723 61844 3765 61853
rect 3723 61804 3724 61844
rect 3764 61804 3765 61844
rect 3723 61795 3765 61804
rect 3724 61606 3764 61795
rect 3915 61760 3957 61769
rect 3915 61720 3916 61760
rect 3956 61720 3957 61760
rect 3915 61711 3957 61720
rect 3819 61676 3861 61685
rect 3819 61636 3820 61676
rect 3860 61636 3861 61676
rect 3819 61627 3861 61636
rect 3724 61557 3764 61566
rect 3820 60920 3860 61627
rect 3916 61508 3956 61711
rect 3916 61459 3956 61468
rect 3916 60920 3956 60929
rect 3820 60880 3916 60920
rect 3916 60871 3956 60880
rect 4108 60761 4148 64240
rect 4300 63118 4340 64912
rect 4588 63953 4628 66088
rect 4587 63944 4629 63953
rect 4587 63904 4588 63944
rect 4628 63904 4629 63944
rect 4587 63895 4629 63904
rect 4300 63069 4340 63078
rect 4491 63020 4533 63029
rect 4491 62980 4492 63020
rect 4532 62980 4533 63020
rect 4491 62971 4533 62980
rect 4492 62886 4532 62971
rect 4299 62684 4341 62693
rect 4299 62644 4300 62684
rect 4340 62644 4341 62684
rect 4299 62635 4341 62644
rect 4203 62432 4245 62441
rect 4203 62392 4204 62432
rect 4244 62392 4245 62432
rect 4203 62383 4245 62392
rect 4204 62298 4244 62383
rect 4107 60752 4149 60761
rect 4107 60712 4108 60752
rect 4148 60712 4149 60752
rect 4107 60703 4149 60712
rect 3688 60500 4056 60509
rect 3728 60460 3770 60500
rect 3810 60460 3852 60500
rect 3892 60460 3934 60500
rect 3974 60460 4016 60500
rect 3688 60451 4056 60460
rect 3627 60332 3669 60341
rect 3627 60292 3628 60332
rect 3668 60292 3669 60332
rect 3627 60283 3669 60292
rect 3628 59408 3668 60283
rect 4300 60080 4340 62635
rect 4491 62600 4533 62609
rect 4491 62560 4492 62600
rect 4532 62560 4533 62600
rect 4491 62551 4533 62560
rect 4492 60920 4532 62551
rect 4587 61004 4629 61013
rect 4587 60964 4588 61004
rect 4628 60964 4629 61004
rect 4587 60955 4629 60964
rect 4444 60910 4532 60920
rect 4484 60880 4532 60910
rect 4588 60870 4628 60955
rect 4444 60861 4484 60870
rect 4684 60425 4724 66844
rect 4780 66809 4820 66928
rect 4779 66800 4821 66809
rect 4779 66760 4780 66800
rect 4820 66760 4821 66800
rect 4779 66751 4821 66760
rect 4876 66128 4916 67096
rect 5356 66968 5396 66977
rect 5356 66809 5396 66928
rect 5355 66800 5397 66809
rect 5355 66760 5356 66800
rect 5396 66760 5397 66800
rect 5355 66751 5397 66760
rect 5452 66725 5492 69019
rect 5644 68564 5684 69112
rect 5740 68825 5780 70783
rect 5739 68816 5781 68825
rect 5739 68776 5740 68816
rect 5780 68776 5781 68816
rect 5739 68767 5781 68776
rect 5740 68657 5780 68767
rect 5739 68648 5781 68657
rect 5739 68608 5740 68648
rect 5780 68608 5781 68648
rect 5739 68599 5781 68608
rect 5548 68524 5684 68564
rect 5548 68069 5588 68524
rect 5740 68480 5780 68489
rect 5644 68440 5740 68480
rect 5547 68060 5589 68069
rect 5547 68020 5548 68060
rect 5588 68020 5589 68060
rect 5547 68011 5589 68020
rect 4971 66716 5013 66725
rect 4971 66676 4972 66716
rect 5012 66676 5013 66716
rect 4971 66667 5013 66676
rect 5164 66716 5204 66725
rect 4972 66582 5012 66667
rect 5067 66212 5109 66221
rect 5067 66172 5068 66212
rect 5108 66172 5109 66212
rect 5067 66163 5109 66172
rect 4972 66128 5012 66137
rect 4876 66088 4972 66128
rect 4779 66044 4821 66053
rect 4779 66004 4780 66044
rect 4820 66004 4821 66044
rect 4779 65995 4821 66004
rect 4780 65297 4820 65995
rect 4972 65969 5012 66088
rect 5068 66078 5108 66163
rect 5164 66053 5204 66676
rect 5451 66716 5493 66725
rect 5451 66676 5452 66716
rect 5492 66676 5493 66716
rect 5451 66667 5493 66676
rect 5547 66296 5589 66305
rect 5644 66296 5684 68440
rect 5740 68431 5780 68440
rect 5739 67640 5781 67649
rect 5739 67600 5740 67640
rect 5780 67600 5781 67640
rect 5739 67591 5781 67600
rect 5740 66893 5780 67591
rect 5739 66884 5781 66893
rect 5739 66844 5740 66884
rect 5780 66844 5781 66884
rect 5739 66835 5781 66844
rect 5547 66256 5548 66296
rect 5588 66256 5684 66296
rect 5547 66247 5589 66256
rect 5548 66128 5588 66247
rect 5548 66079 5588 66088
rect 5163 66044 5205 66053
rect 5163 66004 5164 66044
rect 5204 66004 5205 66044
rect 5163 65995 5205 66004
rect 5451 66044 5493 66053
rect 5451 66004 5452 66044
rect 5492 66004 5493 66044
rect 5451 65995 5493 66004
rect 4971 65960 5013 65969
rect 4971 65920 4972 65960
rect 5012 65920 5013 65960
rect 4971 65911 5013 65920
rect 5355 65876 5397 65885
rect 5355 65836 5356 65876
rect 5396 65836 5397 65876
rect 5355 65827 5397 65836
rect 4928 65792 5296 65801
rect 4968 65752 5010 65792
rect 5050 65752 5092 65792
rect 5132 65752 5174 65792
rect 5214 65752 5256 65792
rect 4928 65743 5296 65752
rect 4779 65288 4821 65297
rect 4779 65248 4780 65288
rect 4820 65248 4821 65288
rect 4779 65239 4821 65248
rect 5163 65288 5205 65297
rect 5163 65248 5164 65288
rect 5204 65248 5205 65288
rect 5163 65239 5205 65248
rect 4779 65120 4821 65129
rect 4779 65080 4780 65120
rect 4820 65080 4821 65120
rect 4779 65071 4821 65080
rect 4780 64709 4820 65071
rect 4779 64700 4821 64709
rect 4779 64660 4780 64700
rect 4820 64660 4821 64700
rect 4779 64651 4821 64660
rect 4780 64616 4820 64651
rect 4780 64566 4820 64576
rect 5164 64616 5204 65239
rect 5259 64952 5301 64961
rect 5259 64912 5260 64952
rect 5300 64912 5301 64952
rect 5259 64903 5301 64912
rect 5260 64700 5300 64903
rect 5260 64651 5300 64660
rect 5164 64567 5204 64576
rect 5356 64616 5396 65827
rect 5452 64616 5492 65995
rect 5548 65456 5588 65465
rect 5548 65129 5588 65416
rect 5836 65451 5876 70960
rect 6124 70832 6164 72304
rect 6220 72176 6260 72185
rect 6220 72017 6260 72136
rect 6316 72176 6356 72715
rect 6412 72680 6452 73723
rect 6508 73697 6548 75571
rect 6507 73688 6549 73697
rect 6507 73648 6508 73688
rect 6548 73648 6549 73688
rect 6507 73639 6549 73648
rect 6507 73520 6549 73529
rect 6507 73480 6508 73520
rect 6548 73480 6549 73520
rect 6507 73471 6549 73480
rect 6508 73386 6548 73471
rect 6604 73361 6644 76075
rect 6700 76074 6740 76159
rect 6796 74201 6836 77008
rect 7275 76999 7317 77008
rect 7083 76880 7125 76889
rect 7083 76840 7084 76880
rect 7124 76840 7125 76880
rect 7083 76831 7125 76840
rect 6892 76040 6932 76049
rect 6892 74285 6932 76000
rect 6987 76040 7029 76049
rect 6987 76000 6988 76040
rect 7028 76000 7029 76040
rect 6987 75991 7029 76000
rect 7084 76040 7124 76831
rect 7084 75991 7124 76000
rect 7179 76040 7221 76049
rect 7179 76000 7180 76040
rect 7220 76000 7221 76040
rect 7179 75991 7221 76000
rect 6988 75906 7028 75991
rect 7180 75906 7220 75991
rect 7276 75788 7316 76999
rect 7372 76040 7412 77848
rect 7467 77300 7509 77309
rect 7467 77260 7468 77300
rect 7508 77260 7509 77300
rect 7467 77251 7509 77260
rect 7468 77166 7508 77251
rect 7564 76208 7604 79024
rect 7852 79015 7892 79024
rect 8044 79064 8084 79267
rect 8044 79015 8084 79024
rect 8140 79064 8180 79073
rect 8140 78905 8180 79024
rect 8139 78896 8181 78905
rect 8139 78856 8140 78896
rect 8180 78856 8181 78896
rect 8139 78847 8181 78856
rect 7660 78812 7700 78821
rect 7660 77552 7700 78772
rect 7851 78812 7893 78821
rect 7851 78772 7852 78812
rect 7892 78772 7893 78812
rect 7851 78763 7893 78772
rect 7852 78056 7892 78763
rect 8332 78569 8372 84139
rect 8427 83768 8469 83777
rect 8427 83728 8428 83768
rect 8468 83728 8469 83768
rect 8427 83719 8469 83728
rect 8428 83634 8468 83719
rect 8524 83441 8564 85936
rect 8716 84953 8756 85936
rect 8715 84944 8757 84953
rect 8715 84904 8716 84944
rect 8756 84904 8757 84944
rect 8715 84895 8757 84904
rect 8811 84356 8853 84365
rect 8811 84316 8812 84356
rect 8852 84316 8853 84356
rect 8811 84307 8853 84316
rect 8812 83768 8852 84307
rect 8908 83768 8948 85936
rect 9100 84953 9140 85936
rect 9099 84944 9141 84953
rect 9099 84904 9100 84944
rect 9140 84904 9141 84944
rect 9099 84895 9141 84904
rect 8908 83728 9236 83768
rect 8812 83719 8852 83728
rect 8620 83516 8660 83525
rect 8523 83432 8565 83441
rect 8523 83392 8524 83432
rect 8564 83392 8565 83432
rect 8523 83383 8565 83392
rect 8331 78560 8373 78569
rect 8331 78520 8332 78560
rect 8372 78520 8373 78560
rect 8331 78511 8373 78520
rect 8620 78392 8660 83476
rect 9004 83516 9044 83525
rect 9044 83476 9140 83516
rect 9004 83467 9044 83476
rect 9003 83348 9045 83357
rect 9003 83308 9004 83348
rect 9044 83308 9045 83348
rect 9003 83299 9045 83308
rect 8907 82256 8949 82265
rect 8907 82216 8908 82256
rect 8948 82216 8949 82256
rect 8907 82207 8949 82216
rect 8908 79232 8948 82207
rect 9004 80585 9044 83299
rect 9003 80576 9045 80585
rect 9003 80536 9004 80576
rect 9044 80536 9045 80576
rect 9003 80527 9045 80536
rect 8908 79192 9044 79232
rect 8908 79064 8948 79073
rect 8908 78989 8948 79024
rect 8907 78980 8949 78989
rect 8907 78940 8908 78980
rect 8948 78940 8949 78980
rect 8907 78931 8949 78940
rect 8908 78392 8948 78931
rect 8044 78352 8660 78392
rect 8716 78352 8948 78392
rect 7948 78233 7988 78318
rect 7947 78224 7989 78233
rect 7947 78184 7948 78224
rect 7988 78184 7989 78224
rect 7947 78175 7989 78184
rect 7852 78016 7988 78056
rect 7852 77561 7892 77646
rect 7756 77552 7796 77561
rect 7660 77512 7756 77552
rect 7756 77503 7796 77512
rect 7851 77552 7893 77561
rect 7851 77512 7852 77552
rect 7892 77512 7893 77552
rect 7851 77503 7893 77512
rect 7948 77384 7988 78016
rect 7852 77344 7988 77384
rect 7755 76796 7797 76805
rect 7755 76756 7756 76796
rect 7796 76756 7797 76796
rect 7755 76747 7797 76756
rect 7756 76217 7796 76747
rect 7660 76208 7700 76217
rect 7564 76168 7660 76208
rect 7660 76159 7700 76168
rect 7755 76208 7797 76217
rect 7755 76168 7756 76208
rect 7796 76168 7797 76208
rect 7755 76159 7797 76168
rect 7468 76049 7508 76134
rect 7372 75881 7412 76000
rect 7467 76040 7509 76049
rect 7467 76000 7468 76040
rect 7508 76000 7509 76040
rect 7467 75991 7509 76000
rect 7564 76040 7604 76049
rect 7852 76040 7892 77344
rect 7947 76796 7989 76805
rect 7947 76756 7948 76796
rect 7988 76756 7989 76796
rect 7947 76747 7989 76756
rect 7948 76712 7988 76747
rect 7948 76661 7988 76672
rect 8044 76544 8084 78352
rect 8716 78308 8756 78352
rect 8620 78268 8756 78308
rect 9004 78308 9044 79192
rect 8428 78224 8468 78233
rect 8140 78140 8180 78149
rect 8428 78140 8468 78184
rect 8180 78100 8468 78140
rect 8524 78224 8564 78233
rect 8140 78091 8180 78100
rect 8524 77561 8564 78184
rect 8523 77552 8565 77561
rect 8523 77512 8524 77552
rect 8564 77512 8565 77552
rect 8523 77503 8565 77512
rect 8236 77468 8276 77477
rect 8236 76721 8276 77428
rect 8331 77468 8373 77477
rect 8331 77428 8332 77468
rect 8372 77428 8373 77468
rect 8331 77419 8373 77428
rect 8332 77334 8372 77419
rect 8427 77300 8469 77309
rect 8427 77260 8428 77300
rect 8468 77260 8469 77300
rect 8427 77251 8469 77260
rect 8331 77216 8373 77225
rect 8331 77176 8332 77216
rect 8372 77176 8373 77216
rect 8331 77167 8373 77176
rect 8235 76712 8277 76721
rect 8235 76672 8236 76712
rect 8276 76672 8277 76712
rect 8235 76663 8277 76672
rect 7604 76000 7892 76040
rect 7948 76504 8084 76544
rect 8140 76544 8180 76553
rect 7564 75991 7604 76000
rect 7371 75872 7413 75881
rect 7563 75872 7605 75881
rect 7371 75832 7372 75872
rect 7412 75832 7413 75872
rect 7371 75823 7413 75832
rect 7468 75832 7564 75872
rect 7604 75832 7605 75872
rect 7084 75748 7316 75788
rect 6987 75620 7029 75629
rect 6987 75580 6988 75620
rect 7028 75580 7029 75620
rect 6987 75571 7029 75580
rect 6988 74528 7028 75571
rect 6988 74479 7028 74488
rect 6891 74276 6933 74285
rect 6891 74236 6892 74276
rect 6932 74236 6933 74276
rect 6891 74227 6933 74236
rect 6795 74192 6837 74201
rect 6795 74152 6796 74192
rect 6836 74152 6837 74192
rect 6795 74143 6837 74152
rect 6891 74108 6933 74117
rect 7084 74108 7124 75748
rect 7360 75704 7402 75713
rect 7276 75664 7361 75704
rect 7401 75664 7402 75704
rect 6891 74068 6892 74108
rect 6932 74068 6933 74108
rect 6891 74059 6933 74068
rect 7058 74068 7124 74108
rect 7180 74276 7220 74285
rect 6796 73949 6836 74034
rect 6795 73940 6837 73949
rect 6795 73900 6796 73940
rect 6836 73900 6837 73940
rect 6795 73891 6837 73900
rect 6796 73688 6836 73697
rect 6700 73648 6796 73688
rect 6603 73352 6645 73361
rect 6603 73312 6604 73352
rect 6644 73312 6645 73352
rect 6603 73303 6645 73312
rect 6507 73268 6549 73277
rect 6507 73228 6508 73268
rect 6548 73228 6549 73268
rect 6507 73219 6549 73228
rect 6508 73016 6548 73219
rect 6603 73184 6645 73193
rect 6603 73144 6604 73184
rect 6644 73144 6645 73184
rect 6603 73135 6645 73144
rect 6508 72967 6548 72976
rect 6604 73020 6644 73135
rect 6604 72965 6644 72980
rect 6508 72848 6548 72857
rect 6508 72764 6548 72808
rect 6700 72764 6740 73648
rect 6796 73639 6836 73648
rect 6892 73688 6932 74059
rect 7058 73940 7098 74068
rect 7180 74024 7220 74236
rect 7180 73984 7225 74024
rect 6892 73639 6932 73648
rect 6988 73900 7098 73940
rect 6796 73016 6836 73025
rect 6836 72976 6932 73016
rect 6796 72967 6836 72976
rect 6508 72724 6740 72764
rect 6892 72689 6932 72976
rect 6891 72680 6933 72689
rect 6412 72640 6548 72680
rect 6316 72101 6356 72136
rect 6411 72176 6453 72185
rect 6411 72136 6412 72176
rect 6452 72136 6453 72176
rect 6508 72176 6548 72640
rect 6891 72640 6892 72680
rect 6932 72640 6933 72680
rect 6891 72631 6933 72640
rect 6796 72176 6836 72185
rect 6508 72136 6796 72176
rect 6411 72127 6453 72136
rect 6796 72127 6836 72136
rect 6315 72092 6357 72101
rect 6315 72052 6316 72092
rect 6356 72052 6357 72092
rect 6315 72043 6357 72052
rect 6412 72042 6452 72127
rect 6219 72008 6261 72017
rect 6219 71968 6220 72008
rect 6260 71968 6261 72008
rect 6219 71959 6261 71968
rect 6508 72008 6548 72017
rect 6700 72008 6740 72017
rect 6548 71968 6644 72008
rect 6508 71959 6548 71968
rect 6411 71840 6453 71849
rect 6411 71800 6412 71840
rect 6452 71800 6453 71840
rect 6411 71791 6453 71800
rect 6219 71336 6261 71345
rect 6219 71296 6220 71336
rect 6260 71296 6261 71336
rect 6219 71287 6261 71296
rect 5932 70792 6164 70832
rect 5932 70169 5972 70792
rect 6124 70655 6164 70664
rect 6027 70580 6069 70589
rect 6124 70580 6164 70615
rect 6027 70540 6028 70580
rect 6068 70540 6164 70580
rect 6027 70531 6069 70540
rect 6220 70496 6260 71287
rect 6412 70580 6452 71791
rect 6507 71420 6549 71429
rect 6507 71380 6508 71420
rect 6548 71380 6549 71420
rect 6507 71371 6549 71380
rect 6508 70664 6548 71371
rect 6604 71345 6644 71968
rect 6700 71513 6740 71968
rect 6795 72008 6837 72017
rect 6892 72008 6932 72631
rect 6988 72176 7028 73900
rect 7185 73856 7225 73984
rect 7276 73940 7316 75664
rect 7360 75655 7402 75664
rect 7468 75629 7508 75832
rect 7563 75823 7605 75832
rect 7563 75704 7605 75713
rect 7563 75664 7564 75704
rect 7604 75664 7605 75704
rect 7563 75655 7605 75664
rect 7467 75620 7509 75629
rect 7467 75580 7468 75620
rect 7508 75580 7509 75620
rect 7467 75571 7509 75580
rect 7468 75200 7508 75571
rect 7468 75151 7508 75160
rect 7564 74864 7604 75655
rect 7468 74824 7604 74864
rect 7660 75032 7700 75041
rect 7372 74696 7412 74705
rect 7372 74117 7412 74656
rect 7468 74360 7508 74824
rect 7563 74696 7605 74705
rect 7563 74656 7564 74696
rect 7604 74656 7605 74696
rect 7563 74647 7605 74656
rect 7564 74528 7604 74647
rect 7564 74479 7604 74488
rect 7660 74528 7700 74992
rect 7468 74320 7604 74360
rect 7467 74192 7509 74201
rect 7467 74152 7468 74192
rect 7508 74152 7509 74192
rect 7467 74143 7509 74152
rect 7371 74108 7413 74117
rect 7371 74068 7372 74108
rect 7412 74068 7413 74108
rect 7371 74059 7413 74068
rect 7276 73900 7412 73940
rect 7084 73816 7225 73856
rect 7084 73688 7124 73816
rect 7084 73277 7124 73648
rect 7179 73688 7221 73697
rect 7179 73648 7180 73688
rect 7220 73648 7221 73688
rect 7179 73639 7221 73648
rect 7281 73688 7321 73697
rect 7180 73554 7220 73639
rect 7281 73445 7321 73648
rect 7280 73436 7322 73445
rect 7280 73396 7281 73436
rect 7321 73396 7322 73436
rect 7280 73387 7322 73396
rect 7179 73352 7221 73361
rect 7179 73312 7180 73352
rect 7220 73312 7221 73352
rect 7179 73303 7221 73312
rect 7083 73268 7125 73277
rect 7083 73228 7084 73268
rect 7124 73228 7125 73268
rect 7083 73219 7125 73228
rect 7180 73100 7220 73303
rect 7372 73100 7412 73900
rect 6988 72101 7028 72136
rect 7084 73060 7220 73100
rect 7276 73060 7412 73100
rect 6987 72092 7029 72101
rect 6987 72052 6988 72092
rect 7028 72052 7029 72092
rect 6987 72043 7029 72052
rect 6795 71968 6796 72008
rect 6836 71968 6932 72008
rect 6795 71959 6837 71968
rect 7084 71597 7124 73060
rect 7179 72428 7221 72437
rect 7179 72388 7180 72428
rect 7220 72388 7221 72428
rect 7179 72379 7221 72388
rect 7083 71588 7125 71597
rect 7083 71548 7084 71588
rect 7124 71548 7125 71588
rect 7083 71539 7125 71548
rect 6699 71504 6741 71513
rect 6699 71464 6700 71504
rect 6740 71464 6741 71504
rect 6699 71455 6741 71464
rect 6603 71336 6645 71345
rect 6603 71296 6604 71336
rect 6644 71296 6645 71336
rect 6603 71287 6645 71296
rect 6987 71336 7029 71345
rect 6987 71296 6988 71336
rect 7028 71296 7029 71336
rect 6987 71287 7029 71296
rect 6891 71168 6933 71177
rect 6891 71128 6892 71168
rect 6932 71128 6933 71168
rect 6891 71119 6933 71128
rect 6699 70832 6741 70841
rect 6699 70792 6700 70832
rect 6740 70792 6741 70832
rect 6699 70783 6741 70792
rect 6604 70678 6644 70687
rect 6601 70664 6604 70678
rect 6508 70638 6604 70664
rect 6508 70629 6644 70638
rect 6508 70624 6641 70629
rect 6412 70540 6644 70580
rect 6124 70456 6260 70496
rect 5931 70160 5973 70169
rect 5931 70120 5932 70160
rect 5972 70120 5973 70160
rect 5931 70111 5973 70120
rect 5932 69992 5972 70001
rect 5932 69413 5972 69952
rect 6124 69992 6164 70456
rect 6124 69917 6164 69952
rect 6220 69992 6260 70001
rect 6123 69908 6165 69917
rect 6123 69868 6124 69908
rect 6164 69868 6165 69908
rect 6123 69859 6165 69868
rect 5931 69404 5973 69413
rect 5931 69364 5932 69404
rect 5972 69364 5973 69404
rect 5931 69355 5973 69364
rect 6220 69329 6260 69952
rect 6315 69992 6357 70001
rect 6315 69952 6316 69992
rect 6356 69952 6357 69992
rect 6315 69943 6357 69952
rect 6412 69992 6452 70001
rect 6316 69858 6356 69943
rect 6315 69656 6357 69665
rect 6315 69616 6316 69656
rect 6356 69616 6357 69656
rect 6315 69607 6357 69616
rect 6219 69320 6261 69329
rect 6219 69280 6220 69320
rect 6260 69280 6261 69320
rect 6219 69271 6261 69280
rect 6123 68732 6165 68741
rect 6123 68692 6124 68732
rect 6164 68692 6165 68732
rect 6123 68683 6165 68692
rect 5931 67808 5973 67817
rect 5931 67768 5932 67808
rect 5972 67768 5973 67808
rect 5931 67759 5973 67768
rect 5932 67640 5972 67759
rect 5932 66641 5972 67600
rect 6027 67556 6069 67565
rect 6027 67516 6028 67556
rect 6068 67516 6069 67556
rect 6027 67507 6069 67516
rect 6028 67313 6068 67507
rect 6027 67304 6069 67313
rect 6027 67264 6028 67304
rect 6068 67264 6069 67304
rect 6027 67255 6069 67264
rect 6124 67229 6164 68683
rect 6219 68480 6261 68489
rect 6219 68435 6220 68480
rect 6260 68435 6261 68480
rect 6219 68431 6261 68435
rect 6220 68345 6260 68431
rect 6123 67220 6165 67229
rect 6123 67180 6124 67220
rect 6164 67180 6165 67220
rect 6123 67171 6165 67180
rect 5931 66632 5973 66641
rect 5931 66592 5932 66632
rect 5972 66592 5973 66632
rect 5931 66583 5973 66592
rect 6028 66137 6068 66223
rect 6027 66133 6069 66137
rect 6027 66088 6028 66133
rect 6068 66088 6069 66133
rect 6027 66079 6069 66088
rect 6124 65876 6164 67171
rect 6316 66641 6356 69607
rect 6412 69161 6452 69952
rect 6507 69992 6549 70001
rect 6507 69952 6508 69992
rect 6548 69952 6549 69992
rect 6507 69943 6549 69952
rect 6411 69152 6453 69161
rect 6411 69112 6412 69152
rect 6452 69112 6453 69152
rect 6411 69103 6453 69112
rect 6412 68648 6452 68657
rect 6508 68648 6548 69943
rect 6604 69665 6644 70540
rect 6700 69824 6740 70783
rect 6795 70580 6837 70589
rect 6795 70540 6796 70580
rect 6836 70540 6837 70580
rect 6795 70531 6837 70540
rect 6796 70446 6836 70531
rect 6796 70001 6836 70086
rect 6892 70085 6932 71119
rect 6988 70664 7028 71287
rect 7084 70841 7124 71539
rect 7180 71504 7220 72379
rect 7180 71177 7220 71464
rect 7179 71168 7221 71177
rect 7179 71128 7180 71168
rect 7220 71128 7221 71168
rect 7179 71119 7221 71128
rect 7276 71000 7316 73060
rect 7371 71336 7413 71345
rect 7371 71296 7372 71336
rect 7412 71296 7413 71336
rect 7371 71287 7413 71296
rect 7372 71202 7412 71287
rect 7468 71084 7508 74143
rect 7564 73100 7604 74320
rect 7660 73445 7700 74488
rect 7851 74276 7893 74285
rect 7851 74236 7852 74276
rect 7892 74236 7893 74276
rect 7851 74227 7893 74236
rect 7755 74192 7797 74201
rect 7755 74152 7756 74192
rect 7796 74152 7797 74192
rect 7755 74143 7797 74152
rect 7756 73688 7796 74143
rect 7756 73639 7796 73648
rect 7852 73688 7892 74227
rect 7852 73639 7892 73648
rect 7659 73436 7701 73445
rect 7659 73396 7660 73436
rect 7700 73396 7701 73436
rect 7659 73387 7701 73396
rect 7564 73060 7892 73100
rect 7755 71756 7797 71765
rect 7755 71716 7756 71756
rect 7796 71716 7797 71756
rect 7755 71707 7797 71716
rect 7756 71504 7796 71707
rect 7756 71455 7796 71464
rect 7659 71336 7701 71345
rect 7659 71296 7660 71336
rect 7700 71296 7701 71336
rect 7659 71287 7701 71296
rect 7468 71044 7604 71084
rect 7276 70960 7412 71000
rect 7083 70832 7125 70841
rect 7083 70792 7084 70832
rect 7124 70792 7125 70832
rect 7083 70783 7125 70792
rect 7275 70832 7317 70841
rect 7275 70792 7276 70832
rect 7316 70792 7317 70832
rect 7275 70783 7317 70792
rect 7179 70748 7221 70757
rect 7179 70708 7180 70748
rect 7220 70708 7221 70748
rect 7179 70699 7221 70708
rect 6988 70615 7028 70624
rect 7083 70664 7125 70673
rect 7083 70624 7084 70664
rect 7124 70624 7125 70664
rect 7083 70615 7125 70624
rect 7084 70530 7124 70615
rect 7180 70580 7220 70699
rect 7276 70664 7316 70783
rect 7276 70615 7316 70624
rect 7180 70531 7220 70540
rect 6891 70076 6933 70085
rect 6891 70036 6892 70076
rect 6932 70036 6933 70076
rect 6891 70027 6933 70036
rect 6795 69992 6837 70001
rect 6795 69952 6796 69992
rect 6836 69952 6837 69992
rect 6795 69943 6837 69952
rect 6988 69992 7028 70001
rect 6891 69908 6933 69917
rect 6891 69868 6892 69908
rect 6932 69868 6933 69908
rect 6891 69859 6933 69868
rect 6700 69784 6836 69824
rect 6603 69656 6645 69665
rect 6603 69616 6604 69656
rect 6644 69616 6645 69656
rect 6603 69607 6645 69616
rect 6699 69320 6741 69329
rect 6699 69280 6700 69320
rect 6740 69280 6741 69320
rect 6699 69271 6741 69280
rect 6452 68608 6548 68648
rect 6412 68599 6452 68608
rect 6591 68491 6631 68500
rect 6508 68451 6591 68480
rect 6508 68440 6631 68451
rect 6700 68480 6740 69271
rect 6700 68440 6744 68480
rect 6315 66632 6357 66641
rect 6315 66592 6316 66632
rect 6356 66592 6357 66632
rect 6315 66583 6357 66592
rect 6508 66389 6548 68440
rect 6704 68396 6744 68440
rect 6604 68356 6744 68396
rect 6604 67145 6644 68356
rect 6699 68228 6741 68237
rect 6699 68188 6700 68228
rect 6740 68188 6741 68228
rect 6699 68179 6741 68188
rect 6700 68094 6740 68179
rect 6699 67892 6741 67901
rect 6699 67852 6700 67892
rect 6740 67852 6741 67892
rect 6699 67843 6741 67852
rect 6603 67136 6645 67145
rect 6603 67096 6604 67136
rect 6644 67096 6645 67136
rect 6603 67087 6645 67096
rect 6604 66968 6644 67087
rect 6604 66919 6644 66928
rect 6603 66800 6645 66809
rect 6603 66760 6604 66800
rect 6644 66760 6645 66800
rect 6603 66751 6645 66760
rect 6507 66380 6549 66389
rect 6412 66340 6508 66380
rect 6548 66340 6549 66380
rect 6315 66128 6357 66137
rect 6315 66088 6316 66128
rect 6356 66088 6357 66128
rect 6315 66079 6357 66088
rect 6220 65969 6260 66054
rect 6219 65960 6261 65969
rect 6219 65920 6220 65960
rect 6260 65920 6261 65960
rect 6219 65911 6261 65920
rect 6028 65836 6164 65876
rect 5931 65792 5973 65801
rect 5931 65752 5932 65792
rect 5972 65752 5973 65792
rect 5931 65743 5973 65752
rect 5932 65624 5972 65743
rect 5932 65575 5972 65584
rect 5836 65411 5972 65451
rect 5739 65204 5781 65213
rect 5739 65164 5740 65204
rect 5780 65164 5781 65204
rect 5739 65155 5781 65164
rect 5547 65120 5589 65129
rect 5547 65080 5548 65120
rect 5588 65080 5589 65120
rect 5547 65071 5589 65080
rect 5740 65070 5780 65155
rect 5548 64616 5588 64625
rect 5452 64576 5548 64616
rect 5588 64576 5684 64616
rect 5356 64567 5396 64576
rect 5548 64567 5588 64576
rect 4972 64448 5012 64457
rect 4780 64408 4972 64448
rect 4780 62609 4820 64408
rect 4972 64399 5012 64408
rect 5355 64448 5397 64457
rect 5355 64408 5356 64448
rect 5396 64408 5397 64448
rect 5355 64399 5397 64408
rect 4928 64280 5296 64289
rect 4968 64240 5010 64280
rect 5050 64240 5092 64280
rect 5132 64240 5174 64280
rect 5214 64240 5256 64280
rect 4928 64231 5296 64240
rect 4928 62768 5296 62777
rect 4968 62728 5010 62768
rect 5050 62728 5092 62768
rect 5132 62728 5174 62768
rect 5214 62728 5256 62768
rect 4928 62719 5296 62728
rect 4779 62600 4821 62609
rect 4779 62560 4780 62600
rect 4820 62560 4821 62600
rect 4779 62551 4821 62560
rect 4779 61676 4821 61685
rect 4779 61636 4780 61676
rect 4820 61636 4821 61676
rect 4779 61627 4821 61636
rect 4683 60416 4725 60425
rect 4683 60376 4684 60416
rect 4724 60376 4725 60416
rect 4683 60367 4725 60376
rect 4780 60080 4820 61627
rect 4928 61256 5296 61265
rect 4968 61216 5010 61256
rect 5050 61216 5092 61256
rect 5132 61216 5174 61256
rect 5214 61216 5256 61256
rect 4928 61207 5296 61216
rect 5067 60920 5109 60929
rect 5067 60880 5068 60920
rect 5108 60880 5109 60920
rect 5067 60871 5109 60880
rect 5356 60920 5396 64399
rect 5451 64112 5493 64121
rect 5451 64072 5452 64112
rect 5492 64072 5493 64112
rect 5451 64063 5493 64072
rect 5452 63944 5492 64063
rect 5452 63895 5492 63904
rect 5547 63944 5589 63953
rect 5547 63904 5548 63944
rect 5588 63904 5589 63944
rect 5547 63895 5589 63904
rect 5548 63810 5588 63895
rect 5644 63692 5684 64576
rect 5932 64373 5972 65411
rect 6028 64457 6068 65836
rect 6316 65792 6356 66079
rect 6124 65752 6356 65792
rect 6124 65456 6164 65752
rect 6412 65708 6452 66340
rect 6507 66331 6549 66340
rect 6507 66128 6549 66137
rect 6507 66088 6508 66128
rect 6548 66088 6549 66128
rect 6507 66079 6549 66088
rect 6508 65994 6548 66079
rect 6316 65668 6452 65708
rect 6220 65549 6260 65580
rect 6219 65540 6261 65549
rect 6219 65500 6220 65540
rect 6260 65500 6261 65540
rect 6219 65491 6261 65500
rect 6124 65407 6164 65416
rect 6220 65456 6260 65491
rect 6220 64952 6260 65416
rect 6124 64912 6260 64952
rect 6027 64448 6069 64457
rect 6027 64408 6028 64448
rect 6068 64408 6069 64448
rect 6027 64399 6069 64408
rect 5931 64364 5973 64373
rect 5931 64324 5932 64364
rect 5972 64324 5973 64364
rect 5931 64315 5973 64324
rect 5835 64112 5877 64121
rect 5835 64072 5836 64112
rect 5876 64072 5877 64112
rect 5835 64063 5877 64072
rect 5739 63944 5781 63953
rect 5739 63904 5740 63944
rect 5780 63904 5781 63944
rect 5739 63895 5781 63904
rect 5548 63652 5684 63692
rect 5451 62684 5493 62693
rect 5451 62644 5452 62684
rect 5492 62644 5493 62684
rect 5451 62635 5493 62644
rect 5452 62432 5492 62635
rect 5452 62383 5492 62392
rect 5068 60786 5108 60871
rect 5163 60668 5205 60677
rect 5163 60628 5164 60668
rect 5204 60628 5205 60668
rect 5163 60619 5205 60628
rect 5164 60534 5204 60619
rect 5356 60593 5396 60880
rect 5355 60584 5397 60593
rect 5355 60544 5356 60584
rect 5396 60544 5397 60584
rect 5355 60535 5397 60544
rect 5259 60500 5301 60509
rect 5259 60460 5260 60500
rect 5300 60460 5301 60500
rect 5259 60451 5301 60460
rect 5163 60416 5205 60425
rect 5163 60376 5164 60416
rect 5204 60376 5205 60416
rect 5163 60367 5205 60376
rect 4300 60031 4340 60040
rect 4684 60040 4820 60080
rect 4492 59912 4532 59921
rect 4204 59872 4492 59912
rect 4204 59408 4244 59872
rect 4492 59863 4532 59872
rect 4395 59744 4437 59753
rect 4395 59704 4396 59744
rect 4436 59704 4437 59744
rect 4395 59695 4437 59704
rect 4396 59585 4436 59695
rect 4395 59576 4437 59585
rect 4395 59536 4396 59576
rect 4436 59536 4437 59576
rect 4395 59527 4437 59536
rect 3628 59359 3668 59368
rect 4156 59398 4244 59408
rect 4196 59368 4244 59398
rect 4300 59492 4340 59501
rect 4156 59349 4196 59358
rect 3688 58988 4056 58997
rect 3728 58948 3770 58988
rect 3810 58948 3852 58988
rect 3892 58948 3934 58988
rect 3974 58948 4016 58988
rect 3688 58939 4056 58948
rect 3723 58820 3765 58829
rect 3723 58780 3724 58820
rect 3764 58780 3765 58820
rect 3723 58771 3765 58780
rect 3724 58568 3764 58771
rect 3724 58325 3764 58528
rect 3723 58316 3765 58325
rect 3723 58276 3724 58316
rect 3764 58276 3765 58316
rect 3723 58267 3765 58276
rect 4300 58073 4340 59452
rect 4299 58064 4341 58073
rect 4299 58024 4300 58064
rect 4340 58024 4341 58064
rect 4299 58015 4341 58024
rect 3627 57896 3669 57905
rect 3627 57856 3628 57896
rect 3668 57856 3669 57896
rect 3627 57847 3669 57856
rect 3724 57896 3764 57905
rect 3628 57762 3668 57847
rect 3436 57688 3572 57728
rect 3436 57224 3476 57688
rect 3724 57644 3764 57856
rect 4107 57812 4149 57821
rect 4107 57772 4108 57812
rect 4148 57772 4149 57812
rect 4107 57763 4149 57772
rect 4204 57812 4244 57821
rect 4108 57678 4148 57763
rect 3343 57184 3476 57224
rect 3532 57604 3764 57644
rect 2955 57056 2997 57065
rect 3343 57056 3383 57184
rect 2955 57016 2956 57056
rect 2996 57016 2997 57056
rect 2955 57007 2997 57016
rect 3340 57016 3383 57056
rect 3435 57056 3477 57065
rect 3435 57016 3436 57056
rect 3476 57016 3477 57056
rect 3532 57056 3572 57604
rect 3688 57476 4056 57485
rect 3728 57436 3770 57476
rect 3810 57436 3852 57476
rect 3892 57436 3934 57476
rect 3974 57436 4016 57476
rect 3688 57427 4056 57436
rect 3819 57056 3861 57065
rect 3532 57016 3764 57056
rect 2859 56552 2901 56561
rect 2859 56512 2860 56552
rect 2900 56512 2901 56552
rect 2859 56503 2901 56512
rect 2668 56384 2708 56393
rect 2572 56344 2668 56384
rect 2572 55469 2612 56344
rect 2668 56335 2708 56344
rect 2763 56384 2805 56393
rect 2763 56344 2764 56384
rect 2804 56344 2805 56384
rect 2763 56335 2805 56344
rect 2860 56216 2900 56225
rect 2667 56048 2709 56057
rect 2667 56008 2668 56048
rect 2708 56008 2709 56048
rect 2667 55999 2709 56008
rect 2668 55544 2708 55999
rect 2860 55880 2900 56176
rect 2956 56057 2996 57007
rect 3340 56972 3380 57016
rect 3435 57007 3477 57016
rect 3339 56932 3380 56972
rect 3243 56888 3285 56897
rect 3243 56848 3244 56888
rect 3284 56848 3285 56888
rect 3339 56888 3379 56932
rect 3436 56922 3476 57007
rect 3627 56888 3669 56897
rect 3339 56848 3380 56888
rect 3243 56839 3285 56848
rect 3052 56468 3092 56477
rect 3092 56428 3188 56468
rect 3052 56419 3092 56428
rect 2955 56048 2997 56057
rect 2955 56008 2956 56048
rect 2996 56008 2997 56048
rect 2955 55999 2997 56008
rect 2860 55840 3092 55880
rect 2860 55712 2900 55721
rect 2860 55628 2900 55672
rect 2860 55588 2901 55628
rect 2861 55544 2901 55588
rect 3052 55544 3092 55840
rect 3148 55628 3188 56428
rect 3244 56379 3284 56839
rect 3340 56804 3380 56848
rect 3627 56848 3628 56888
rect 3668 56848 3669 56888
rect 3627 56839 3669 56848
rect 3340 56764 3572 56804
rect 3339 56552 3381 56561
rect 3339 56512 3340 56552
rect 3380 56512 3381 56552
rect 3339 56503 3381 56512
rect 3244 56330 3284 56339
rect 3244 55628 3284 55637
rect 3148 55588 3244 55628
rect 3244 55579 3284 55588
rect 2861 55504 2996 55544
rect 3052 55504 3188 55544
rect 2571 55460 2613 55469
rect 2571 55420 2572 55460
rect 2612 55420 2613 55460
rect 2571 55411 2613 55420
rect 2284 54862 2372 54872
rect 2284 54832 2332 54862
rect 2332 54813 2372 54822
rect 2668 54704 2708 55504
rect 2859 55124 2901 55133
rect 2859 55084 2860 55124
rect 2900 55084 2901 55124
rect 2859 55075 2901 55084
rect 2476 54664 2708 54704
rect 2860 54872 2900 55075
rect 2476 54116 2516 54664
rect 2860 54200 2900 54832
rect 2956 54377 2996 55504
rect 3052 55376 3092 55385
rect 3052 54881 3092 55336
rect 3051 54872 3093 54881
rect 3051 54832 3052 54872
rect 3092 54832 3093 54872
rect 3051 54823 3093 54832
rect 3051 54704 3093 54713
rect 3051 54664 3052 54704
rect 3092 54664 3093 54704
rect 3051 54655 3093 54664
rect 2955 54368 2997 54377
rect 2955 54328 2956 54368
rect 2996 54328 2997 54368
rect 2955 54319 2997 54328
rect 2955 54200 2997 54209
rect 2860 54160 2956 54200
rect 2996 54160 2997 54200
rect 2955 54151 2997 54160
rect 2476 54076 2804 54116
rect 2476 54032 2516 54076
rect 2187 52688 2229 52697
rect 2187 52648 2188 52688
rect 2228 52648 2229 52688
rect 2187 52639 2229 52648
rect 2380 52520 2420 52529
rect 2476 52520 2516 53992
rect 2668 53864 2708 53873
rect 2571 53780 2613 53789
rect 2571 53740 2572 53780
rect 2612 53740 2613 53780
rect 2571 53731 2613 53740
rect 2420 52480 2516 52520
rect 2380 52471 2420 52480
rect 2572 52361 2612 53731
rect 2091 52352 2133 52361
rect 2091 52312 2092 52352
rect 2132 52312 2133 52352
rect 2091 52303 2133 52312
rect 2188 52352 2228 52361
rect 2091 52184 2133 52193
rect 2188 52184 2228 52312
rect 2379 52352 2421 52361
rect 2379 52312 2380 52352
rect 2420 52312 2421 52352
rect 2379 52303 2421 52312
rect 2571 52352 2613 52361
rect 2571 52312 2572 52352
rect 2612 52312 2613 52352
rect 2571 52303 2613 52312
rect 2091 52144 2092 52184
rect 2132 52144 2228 52184
rect 2091 52135 2133 52144
rect 2380 52100 2420 52303
rect 2571 52184 2613 52193
rect 2571 52144 2572 52184
rect 2612 52144 2613 52184
rect 2571 52135 2613 52144
rect 2284 52060 2420 52100
rect 1899 51764 1941 51773
rect 1899 51724 1900 51764
rect 1940 51724 1941 51764
rect 1899 51715 1941 51724
rect 2092 51764 2132 51773
rect 1900 51596 1940 51605
rect 1900 49925 1940 51556
rect 2092 50597 2132 51724
rect 2091 50588 2133 50597
rect 2091 50548 2092 50588
rect 2132 50548 2133 50588
rect 2091 50539 2133 50548
rect 2284 50420 2324 52060
rect 2380 51932 2420 51941
rect 2380 51773 2420 51892
rect 2572 51843 2612 52135
rect 2668 52109 2708 53824
rect 2764 53360 2804 54076
rect 3052 53528 3092 54655
rect 3148 54032 3188 55504
rect 3340 55133 3380 56503
rect 3532 56384 3572 56764
rect 3628 56754 3668 56839
rect 3724 56561 3764 57016
rect 3819 57016 3820 57056
rect 3860 57016 3861 57056
rect 3819 57007 3861 57016
rect 3820 56922 3860 57007
rect 4204 56981 4244 57772
rect 4396 57065 4436 59527
rect 4587 59072 4629 59081
rect 4587 59032 4588 59072
rect 4628 59032 4629 59072
rect 4587 59023 4629 59032
rect 4588 58241 4628 59023
rect 4587 58232 4629 58241
rect 4587 58192 4588 58232
rect 4628 58192 4629 58232
rect 4587 58183 4629 58192
rect 4684 57896 4724 60040
rect 4779 59912 4821 59921
rect 4779 59872 4780 59912
rect 4820 59872 4821 59912
rect 5164 59912 5204 60367
rect 5260 60080 5300 60451
rect 5548 60425 5588 63652
rect 5740 63029 5780 63895
rect 5739 63020 5781 63029
rect 5739 62980 5740 63020
rect 5780 62980 5781 63020
rect 5739 62971 5781 62980
rect 5644 62180 5684 62189
rect 5644 61592 5684 62140
rect 5740 61937 5780 62971
rect 5836 62600 5876 64063
rect 6027 63944 6069 63953
rect 6027 63904 6028 63944
rect 6068 63904 6069 63944
rect 6027 63895 6069 63904
rect 5932 63860 5972 63869
rect 5932 63356 5972 63820
rect 6028 63810 6068 63895
rect 6124 63356 6164 64912
rect 6316 64868 6356 65668
rect 6604 65624 6644 66751
rect 6700 66128 6740 67843
rect 6796 67565 6836 69784
rect 6892 69774 6932 69859
rect 6988 69404 7028 69952
rect 7275 69908 7317 69917
rect 7275 69868 7276 69908
rect 7316 69868 7317 69908
rect 7275 69859 7317 69868
rect 6988 69364 7220 69404
rect 6892 69245 6932 69247
rect 6891 69236 6933 69245
rect 6891 69196 6892 69236
rect 6932 69196 6933 69236
rect 6891 69187 6933 69196
rect 6892 69152 6932 69187
rect 6892 69103 6932 69112
rect 7083 69152 7125 69161
rect 7083 69112 7084 69152
rect 7124 69112 7125 69152
rect 7083 69103 7125 69112
rect 7180 69152 7220 69364
rect 7276 69152 7316 69859
rect 7372 69329 7412 70960
rect 7468 70841 7508 70926
rect 7467 70832 7509 70841
rect 7467 70792 7468 70832
rect 7508 70792 7509 70832
rect 7467 70783 7509 70792
rect 7468 70664 7508 70675
rect 7468 70589 7508 70624
rect 7467 70580 7509 70589
rect 7467 70540 7468 70580
rect 7508 70540 7509 70580
rect 7467 70531 7509 70540
rect 7564 70412 7604 71044
rect 7660 70673 7700 71287
rect 7659 70664 7701 70673
rect 7659 70624 7660 70664
rect 7700 70624 7701 70664
rect 7659 70615 7701 70624
rect 7660 70530 7700 70615
rect 7468 70372 7604 70412
rect 7371 69320 7413 69329
rect 7371 69280 7372 69320
rect 7412 69280 7413 69320
rect 7371 69271 7413 69280
rect 7372 69152 7412 69161
rect 7276 69112 7372 69152
rect 7084 69018 7124 69103
rect 6891 68900 6933 68909
rect 6891 68860 6892 68900
rect 6932 68860 6933 68900
rect 6891 68851 6933 68860
rect 6892 68489 6932 68851
rect 6891 68480 6933 68489
rect 6891 68440 6892 68480
rect 6932 68440 6933 68480
rect 6891 68431 6933 68440
rect 6892 68346 6932 68431
rect 7083 68060 7125 68069
rect 7083 68020 7084 68060
rect 7124 68020 7125 68060
rect 7083 68011 7125 68020
rect 7084 67640 7124 68011
rect 7180 67892 7220 69112
rect 7372 69103 7412 69112
rect 7275 68984 7317 68993
rect 7275 68944 7276 68984
rect 7316 68944 7317 68984
rect 7275 68935 7317 68944
rect 7276 68850 7316 68935
rect 7372 67892 7412 67901
rect 7180 67852 7372 67892
rect 7372 67843 7412 67852
rect 7180 67640 7220 67649
rect 7084 67600 7180 67640
rect 6795 67556 6837 67565
rect 6795 67516 6796 67556
rect 6836 67516 6837 67556
rect 6795 67507 6837 67516
rect 7083 67136 7125 67145
rect 7083 67096 7084 67136
rect 7124 67096 7125 67136
rect 6796 67061 6836 67092
rect 7083 67087 7125 67096
rect 6795 67052 6837 67061
rect 6795 67012 6796 67052
rect 6836 67012 6837 67052
rect 6795 67003 6837 67012
rect 6796 66968 6836 67003
rect 6796 66389 6836 66928
rect 6891 66548 6933 66557
rect 6891 66508 6892 66548
rect 6932 66508 6933 66548
rect 6891 66499 6933 66508
rect 6795 66380 6837 66389
rect 6795 66340 6796 66380
rect 6836 66340 6837 66380
rect 6795 66331 6837 66340
rect 6796 66128 6836 66137
rect 6700 66088 6796 66128
rect 6699 65792 6741 65801
rect 6699 65752 6700 65792
rect 6740 65752 6741 65792
rect 6699 65743 6741 65752
rect 6508 65584 6644 65624
rect 6412 65465 6452 65550
rect 6508 65540 6548 65584
rect 6508 65491 6548 65500
rect 6411 65456 6453 65465
rect 6411 65416 6412 65456
rect 6452 65416 6453 65456
rect 6411 65407 6453 65416
rect 6604 65456 6644 65467
rect 6604 65381 6644 65416
rect 6700 65456 6740 65743
rect 6796 65708 6836 66088
rect 6892 66128 6932 66499
rect 6892 66079 6932 66088
rect 6796 65668 6932 65708
rect 6700 65407 6740 65416
rect 6603 65372 6645 65381
rect 6603 65332 6604 65372
rect 6644 65332 6645 65372
rect 6603 65323 6645 65332
rect 6411 65288 6453 65297
rect 6411 65248 6412 65288
rect 6452 65248 6453 65288
rect 6411 65239 6453 65248
rect 5932 63316 6164 63356
rect 5931 63104 5973 63113
rect 5931 63064 5932 63104
rect 5972 63064 5973 63104
rect 5931 63055 5973 63064
rect 5932 62970 5972 63055
rect 6027 62936 6069 62945
rect 6027 62896 6028 62936
rect 6068 62896 6069 62936
rect 6027 62887 6069 62896
rect 5836 62560 5972 62600
rect 5836 62432 5876 62441
rect 5836 62189 5876 62392
rect 5835 62180 5877 62189
rect 5835 62140 5836 62180
rect 5876 62140 5877 62180
rect 5835 62131 5877 62140
rect 5739 61928 5781 61937
rect 5739 61888 5740 61928
rect 5780 61888 5781 61928
rect 5739 61879 5781 61888
rect 5644 61543 5684 61552
rect 5740 61592 5780 61879
rect 5740 61543 5780 61552
rect 5643 61088 5685 61097
rect 5643 61048 5644 61088
rect 5684 61048 5685 61088
rect 5643 61039 5685 61048
rect 5547 60416 5589 60425
rect 5547 60376 5548 60416
rect 5588 60376 5589 60416
rect 5547 60367 5589 60376
rect 5356 60080 5396 60089
rect 5260 60040 5356 60080
rect 5356 60031 5396 60040
rect 5164 59872 5396 59912
rect 4779 59863 4821 59872
rect 4588 57856 4684 57896
rect 4491 57812 4533 57821
rect 4491 57772 4492 57812
rect 4532 57772 4533 57812
rect 4491 57763 4533 57772
rect 4395 57056 4437 57065
rect 4395 57016 4396 57056
rect 4436 57016 4437 57056
rect 4395 57007 4437 57016
rect 4203 56972 4245 56981
rect 4203 56932 4204 56972
rect 4244 56932 4245 56972
rect 4203 56923 4245 56932
rect 3723 56552 3765 56561
rect 3723 56512 3724 56552
rect 3764 56512 3765 56552
rect 3723 56503 3765 56512
rect 3724 56384 3764 56393
rect 3532 56344 3724 56384
rect 3435 55628 3477 55637
rect 3435 55588 3436 55628
rect 3476 55588 3477 55628
rect 3435 55579 3477 55588
rect 3436 55544 3476 55579
rect 3436 55493 3476 55504
rect 3339 55124 3381 55133
rect 3339 55084 3340 55124
rect 3380 55084 3381 55124
rect 3339 55075 3381 55084
rect 3339 54956 3381 54965
rect 3339 54916 3340 54956
rect 3380 54916 3381 54956
rect 3339 54907 3381 54916
rect 3340 54872 3380 54907
rect 3340 54821 3380 54832
rect 3435 54788 3477 54797
rect 3435 54748 3436 54788
rect 3476 54748 3477 54788
rect 3435 54739 3477 54748
rect 3436 54654 3476 54739
rect 3340 54032 3380 54041
rect 3148 53992 3340 54032
rect 3340 53983 3380 53992
rect 3436 54032 3476 54041
rect 3148 53528 3188 53537
rect 3052 53488 3148 53528
rect 3148 53479 3188 53488
rect 2956 53444 2996 53453
rect 2996 53404 3092 53444
rect 2956 53395 2996 53404
rect 3052 53360 3092 53404
rect 3436 53369 3476 53992
rect 3435 53360 3477 53369
rect 3052 53350 3332 53360
rect 3052 53320 3292 53350
rect 2764 53285 2804 53320
rect 3435 53320 3436 53360
rect 3476 53320 3477 53360
rect 3435 53311 3477 53320
rect 3292 53301 3332 53310
rect 2763 53276 2805 53285
rect 2763 53236 2764 53276
rect 2804 53236 2805 53276
rect 2763 53227 2805 53236
rect 3532 53192 3572 56344
rect 3724 56335 3764 56344
rect 4204 56384 4244 56923
rect 4395 56468 4437 56477
rect 4395 56428 4396 56468
rect 4436 56428 4437 56468
rect 4395 56419 4437 56428
rect 4204 56335 4244 56344
rect 4299 56300 4341 56309
rect 4299 56260 4300 56300
rect 4340 56260 4341 56300
rect 4299 56251 4341 56260
rect 4300 56166 4340 56251
rect 3688 55964 4056 55973
rect 3728 55924 3770 55964
rect 3810 55924 3852 55964
rect 3892 55924 3934 55964
rect 3974 55924 4016 55964
rect 3688 55915 4056 55924
rect 4396 55460 4436 56419
rect 4300 55420 4436 55460
rect 3915 55376 3957 55385
rect 3915 55336 3916 55376
rect 3956 55336 3957 55376
rect 3915 55327 3957 55336
rect 3819 54872 3861 54881
rect 3819 54832 3820 54872
rect 3860 54832 3861 54872
rect 3819 54823 3861 54832
rect 3916 54872 3956 55327
rect 3916 54823 3956 54832
rect 3820 54738 3860 54823
rect 3688 54452 4056 54461
rect 3728 54412 3770 54452
rect 3810 54412 3852 54452
rect 3892 54412 3934 54452
rect 3974 54412 4016 54452
rect 3688 54403 4056 54412
rect 3723 54200 3765 54209
rect 3723 54160 3724 54200
rect 3764 54160 3765 54200
rect 3723 54151 3765 54160
rect 3627 53948 3669 53957
rect 3627 53908 3628 53948
rect 3668 53908 3669 53948
rect 3627 53899 3669 53908
rect 3628 53537 3668 53899
rect 3627 53528 3669 53537
rect 3627 53488 3628 53528
rect 3668 53488 3669 53528
rect 3627 53479 3669 53488
rect 3052 53152 3572 53192
rect 2763 53108 2805 53117
rect 2763 53068 2764 53108
rect 2804 53068 2805 53108
rect 2763 53059 2805 53068
rect 2667 52100 2709 52109
rect 2667 52060 2668 52100
rect 2708 52060 2709 52100
rect 2667 52051 2709 52060
rect 2572 51794 2612 51803
rect 2379 51764 2421 51773
rect 2379 51724 2380 51764
rect 2420 51724 2421 51764
rect 2379 51715 2421 51724
rect 2764 51689 2804 53059
rect 2955 52940 2997 52949
rect 2955 52900 2956 52940
rect 2996 52900 2997 52940
rect 2955 52891 2997 52900
rect 2859 52352 2901 52361
rect 2859 52312 2860 52352
rect 2900 52312 2901 52352
rect 2859 52303 2901 52312
rect 2763 51680 2805 51689
rect 2763 51640 2764 51680
rect 2804 51640 2805 51680
rect 2763 51631 2805 51640
rect 2860 51260 2900 52303
rect 2860 51211 2900 51220
rect 2763 51176 2805 51185
rect 2763 51136 2764 51176
rect 2804 51136 2805 51176
rect 2763 51127 2805 51136
rect 1996 50380 2324 50420
rect 2476 51008 2516 51017
rect 2476 50420 2516 50968
rect 2667 50840 2709 50849
rect 2667 50800 2668 50840
rect 2708 50800 2709 50840
rect 2667 50791 2709 50800
rect 2668 50706 2708 50791
rect 2476 50380 2540 50420
rect 1899 49916 1941 49925
rect 1899 49876 1900 49916
rect 1940 49876 1941 49916
rect 1899 49867 1941 49876
rect 1900 49748 1940 49757
rect 1804 49708 1900 49748
rect 1900 49699 1940 49708
rect 1708 49580 1748 49589
rect 1708 49421 1748 49540
rect 1707 49412 1749 49421
rect 1707 49372 1708 49412
rect 1748 49372 1749 49412
rect 1707 49363 1749 49372
rect 1996 48665 2036 50380
rect 2500 50336 2540 50380
rect 2667 50336 2709 50345
rect 2500 50296 2668 50336
rect 2708 50296 2709 50336
rect 2475 50084 2517 50093
rect 2475 50044 2476 50084
rect 2516 50044 2517 50084
rect 2475 50035 2517 50044
rect 2092 49580 2132 49589
rect 2132 49540 2420 49580
rect 2092 49531 2132 49540
rect 2283 49412 2325 49421
rect 2283 49372 2284 49412
rect 2324 49372 2325 49412
rect 2283 49363 2325 49372
rect 2284 49278 2324 49363
rect 2380 48917 2420 49540
rect 2476 49510 2516 50035
rect 2476 49461 2516 49470
rect 2379 48908 2421 48917
rect 2379 48868 2380 48908
rect 2420 48868 2421 48908
rect 2379 48859 2421 48868
rect 2476 48824 2516 48833
rect 2572 48824 2612 50296
rect 2667 50287 2709 50296
rect 2668 50202 2708 50287
rect 2764 48992 2804 51127
rect 2956 50765 2996 52891
rect 3052 51848 3092 53152
rect 3628 53108 3668 53479
rect 3724 53117 3764 54151
rect 3819 54032 3861 54041
rect 3819 53992 3820 54032
rect 3860 53992 3861 54032
rect 3819 53983 3861 53992
rect 3916 54032 3956 54043
rect 3820 53780 3860 53983
rect 3916 53957 3956 53992
rect 3915 53948 3957 53957
rect 3915 53908 3916 53948
rect 3956 53908 3957 53948
rect 3915 53899 3957 53908
rect 3820 53740 3956 53780
rect 3820 53360 3860 53369
rect 3532 53068 3668 53108
rect 3723 53108 3765 53117
rect 3820 53108 3860 53320
rect 3916 53117 3956 53740
rect 4300 53444 4340 55420
rect 4395 54956 4437 54965
rect 4395 54916 4396 54956
rect 4436 54916 4437 54956
rect 4395 54907 4437 54916
rect 4396 54209 4436 54907
rect 4395 54200 4437 54209
rect 4395 54160 4396 54200
rect 4436 54160 4437 54200
rect 4395 54151 4437 54160
rect 4396 54032 4436 54151
rect 4492 54041 4532 57763
rect 4396 53983 4436 53992
rect 4491 54032 4533 54041
rect 4491 53992 4492 54032
rect 4532 53992 4533 54032
rect 4491 53983 4533 53992
rect 4300 53404 4532 53444
rect 4203 53360 4245 53369
rect 4203 53320 4204 53360
rect 4244 53320 4245 53360
rect 4203 53311 4245 53320
rect 3723 53068 3724 53108
rect 3764 53068 3860 53108
rect 3915 53108 3957 53117
rect 3915 53068 3916 53108
rect 3956 53068 3957 53108
rect 3435 52940 3477 52949
rect 3435 52900 3436 52940
rect 3476 52900 3477 52940
rect 3435 52891 3477 52900
rect 3092 51808 3284 51848
rect 3052 51799 3092 51808
rect 3147 51680 3189 51689
rect 3147 51640 3148 51680
rect 3188 51640 3189 51680
rect 3147 51631 3189 51640
rect 3051 51092 3093 51101
rect 3051 51052 3052 51092
rect 3092 51052 3093 51092
rect 3051 51043 3093 51052
rect 3052 50958 3092 51043
rect 2955 50756 2997 50765
rect 2955 50716 2956 50756
rect 2996 50716 2997 50756
rect 2955 50707 2997 50716
rect 3052 50336 3092 50345
rect 2859 50084 2901 50093
rect 2859 50044 2860 50084
rect 2900 50044 2901 50084
rect 2859 50035 2901 50044
rect 2860 49950 2900 50035
rect 3052 50009 3092 50296
rect 3051 50000 3093 50009
rect 3051 49960 3052 50000
rect 3092 49960 3093 50000
rect 3051 49951 3093 49960
rect 2955 49496 2997 49505
rect 2955 49456 2956 49496
rect 2996 49456 2997 49496
rect 3148 49496 3188 51631
rect 3244 49580 3284 51808
rect 3339 51008 3381 51017
rect 3339 50968 3340 51008
rect 3380 50968 3381 51008
rect 3339 50959 3381 50968
rect 3340 50874 3380 50959
rect 3436 50504 3476 52891
rect 3532 51848 3572 53068
rect 3723 53059 3765 53068
rect 3915 53059 3957 53068
rect 3688 52940 4056 52949
rect 3728 52900 3770 52940
rect 3810 52900 3852 52940
rect 3892 52900 3934 52940
rect 3974 52900 4016 52940
rect 3688 52891 4056 52900
rect 3723 52772 3765 52781
rect 3723 52732 3724 52772
rect 3764 52732 3765 52772
rect 3723 52723 3765 52732
rect 3627 52520 3669 52529
rect 3627 52480 3628 52520
rect 3668 52480 3669 52520
rect 3627 52471 3669 52480
rect 3628 52386 3668 52471
rect 3532 51799 3572 51808
rect 3627 51764 3669 51773
rect 3724 51764 3764 52723
rect 3819 52520 3861 52529
rect 3819 52480 3820 52520
rect 3860 52480 3861 52520
rect 3819 52471 3861 52480
rect 3820 52386 3860 52471
rect 4107 52100 4149 52109
rect 4107 52060 4108 52100
rect 4148 52060 4149 52100
rect 4107 52051 4149 52060
rect 3627 51724 3628 51764
rect 3668 51724 3764 51764
rect 4012 51848 4052 51857
rect 3627 51715 3669 51724
rect 3628 51630 3668 51715
rect 4012 51596 4052 51808
rect 4108 51848 4148 52051
rect 4108 51799 4148 51808
rect 4204 51596 4244 53311
rect 4300 53276 4340 53285
rect 4300 53117 4340 53236
rect 4396 53276 4436 53285
rect 4299 53108 4341 53117
rect 4299 53068 4300 53108
rect 4340 53068 4341 53108
rect 4299 53059 4341 53068
rect 4396 52781 4436 53236
rect 4395 52772 4437 52781
rect 4395 52732 4396 52772
rect 4436 52732 4437 52772
rect 4395 52723 4437 52732
rect 4012 51556 4244 51596
rect 3688 51428 4056 51437
rect 3728 51388 3770 51428
rect 3810 51388 3852 51428
rect 3892 51388 3934 51428
rect 3974 51388 4016 51428
rect 3688 51379 4056 51388
rect 4011 51008 4053 51017
rect 4011 50968 4012 51008
rect 4052 50968 4053 51008
rect 4011 50959 4053 50968
rect 3436 50464 3572 50504
rect 3436 49580 3476 49589
rect 3244 49540 3436 49580
rect 3148 49456 3284 49496
rect 2955 49447 2997 49456
rect 2860 48992 2900 49001
rect 2764 48952 2860 48992
rect 2860 48943 2900 48952
rect 2516 48784 2612 48824
rect 1995 48656 2037 48665
rect 1995 48616 1996 48656
rect 2036 48616 2037 48656
rect 1995 48607 2037 48616
rect 2283 48572 2325 48581
rect 2283 48532 2284 48572
rect 2324 48532 2325 48572
rect 2283 48523 2325 48532
rect 1612 48187 1652 48196
rect 1707 48152 1749 48161
rect 1707 48112 1708 48152
rect 1748 48112 1749 48152
rect 1707 48103 1749 48112
rect 1708 47480 1748 48103
rect 1803 48068 1845 48077
rect 1803 48028 1804 48068
rect 1844 48028 1845 48068
rect 1803 48019 1845 48028
rect 1804 47934 1844 48019
rect 1995 47984 2037 47993
rect 1995 47944 1996 47984
rect 2036 47944 2037 47984
rect 1995 47935 2037 47944
rect 1996 47850 2036 47935
rect 1804 47480 1844 47489
rect 1708 47440 1804 47480
rect 1804 47431 1844 47440
rect 2284 47312 2324 48523
rect 2476 48161 2516 48784
rect 2667 48572 2709 48581
rect 2667 48532 2668 48572
rect 2708 48532 2709 48572
rect 2667 48523 2709 48532
rect 2668 48438 2708 48523
rect 2859 48236 2901 48245
rect 2859 48196 2860 48236
rect 2900 48196 2901 48236
rect 2859 48187 2901 48196
rect 2475 48152 2517 48161
rect 2475 48112 2476 48152
rect 2516 48112 2517 48152
rect 2475 48103 2517 48112
rect 2284 47263 2324 47272
rect 2379 47312 2421 47321
rect 2379 47272 2380 47312
rect 2420 47272 2421 47312
rect 2379 47263 2421 47272
rect 1995 47228 2037 47237
rect 1995 47188 1996 47228
rect 2036 47188 2037 47228
rect 1995 47179 2037 47188
rect 1899 47144 1941 47153
rect 1899 47104 1900 47144
rect 1940 47104 1941 47144
rect 1899 47095 1941 47104
rect 1420 46936 1556 46976
rect 1420 45632 1460 46936
rect 1515 46808 1557 46817
rect 1515 46768 1516 46808
rect 1556 46768 1557 46808
rect 1515 46759 1557 46768
rect 1516 45968 1556 46759
rect 1516 45919 1556 45928
rect 1900 45968 1940 47095
rect 1996 47094 2036 47179
rect 2380 47178 2420 47263
rect 1900 45919 1940 45928
rect 2476 46472 2516 48103
rect 2571 47984 2613 47993
rect 2571 47944 2572 47984
rect 2612 47944 2613 47984
rect 2571 47935 2613 47944
rect 2476 45809 2516 46432
rect 2283 45800 2325 45809
rect 2283 45760 2284 45800
rect 2324 45760 2325 45800
rect 2283 45751 2325 45760
rect 2475 45800 2517 45809
rect 2475 45760 2476 45800
rect 2516 45760 2517 45800
rect 2475 45751 2517 45760
rect 1707 45716 1749 45725
rect 1707 45676 1708 45716
rect 1748 45676 1749 45716
rect 1707 45667 1749 45676
rect 2092 45716 2132 45725
rect 1420 45592 1652 45632
rect 1515 45464 1557 45473
rect 1515 45424 1516 45464
rect 1556 45424 1557 45464
rect 1515 45415 1557 45424
rect 1516 45212 1556 45415
rect 1612 45296 1652 45592
rect 1708 45582 1748 45667
rect 2092 45305 2132 45676
rect 2091 45296 2133 45305
rect 1612 45256 1844 45296
rect 1516 45163 1556 45172
rect 1708 45044 1748 45053
rect 1324 45004 1708 45044
rect 1708 44995 1748 45004
rect 1228 44920 1652 44960
rect 1228 42776 1268 42785
rect 1228 42692 1268 42736
rect 1323 42692 1365 42701
rect 1228 42652 1324 42692
rect 1364 42652 1365 42692
rect 1323 42643 1365 42652
rect 1612 42188 1652 44920
rect 1804 44456 1844 45256
rect 2091 45256 2092 45296
rect 2132 45256 2133 45296
rect 2091 45247 2133 45256
rect 2091 45044 2133 45053
rect 2091 45004 2092 45044
rect 2132 45004 2133 45044
rect 2091 44995 2133 45004
rect 2092 44910 2132 44995
rect 1900 44792 1940 44801
rect 1900 44465 1940 44752
rect 1804 44407 1844 44416
rect 1899 44456 1941 44465
rect 1899 44416 1900 44456
rect 1940 44416 1941 44456
rect 1899 44407 1941 44416
rect 2284 44288 2324 45751
rect 2379 45716 2421 45725
rect 2379 45676 2380 45716
rect 2420 45676 2421 45716
rect 2379 45667 2421 45676
rect 2380 44876 2420 45667
rect 2476 45548 2516 45557
rect 2476 45078 2516 45508
rect 2572 45212 2612 47935
rect 2763 47900 2805 47909
rect 2763 47860 2764 47900
rect 2804 47860 2805 47900
rect 2763 47851 2805 47860
rect 2764 47228 2804 47851
rect 2667 46304 2709 46313
rect 2667 46264 2668 46304
rect 2708 46264 2709 46304
rect 2667 46255 2709 46264
rect 2668 46170 2708 46255
rect 2667 45800 2709 45809
rect 2667 45760 2668 45800
rect 2708 45760 2709 45800
rect 2667 45751 2709 45760
rect 2668 45666 2708 45751
rect 2572 45172 2708 45212
rect 2476 45044 2540 45078
rect 2476 45004 2564 45044
rect 2524 45002 2564 45004
rect 2524 44953 2564 44962
rect 2668 44876 2708 45172
rect 2380 44827 2420 44836
rect 2572 44836 2708 44876
rect 2380 44288 2420 44297
rect 2284 44248 2380 44288
rect 1995 44204 2037 44213
rect 1995 44164 1996 44204
rect 2036 44164 2037 44204
rect 1995 44155 2037 44164
rect 1996 44070 2036 44155
rect 2187 44036 2229 44045
rect 2187 43996 2188 44036
rect 2228 43996 2229 44036
rect 2187 43987 2229 43996
rect 2188 43902 2228 43987
rect 2284 42776 2324 44248
rect 2380 44239 2420 44248
rect 2475 44204 2517 44213
rect 2475 44164 2476 44204
rect 2516 44164 2517 44204
rect 2475 44155 2517 44164
rect 2476 43364 2516 44155
rect 2476 43315 2516 43324
rect 2476 42776 2516 42785
rect 2284 42736 2476 42776
rect 1900 42188 1940 42197
rect 1612 42148 1900 42188
rect 1900 42139 1940 42148
rect 2092 42020 2132 42029
rect 2092 41852 2132 41980
rect 2284 41852 2324 41861
rect 2092 41812 2284 41852
rect 2284 41803 2324 41812
rect 1899 41264 1941 41273
rect 1899 41224 1900 41264
rect 1940 41224 1941 41264
rect 1899 41215 1941 41224
rect 1419 41180 1461 41189
rect 1419 41140 1420 41180
rect 1460 41140 1461 41180
rect 1419 41131 1461 41140
rect 1420 40517 1460 41131
rect 1900 41130 1940 41215
rect 1419 40508 1461 40517
rect 1419 40468 1420 40508
rect 1460 40468 1461 40508
rect 1419 40459 1461 40468
rect 1707 40508 1749 40517
rect 1707 40468 1708 40508
rect 1748 40468 1749 40508
rect 1707 40459 1749 40468
rect 2380 40508 2420 42736
rect 2476 42727 2516 42736
rect 2476 41941 2516 41950
rect 2476 41525 2516 41901
rect 2475 41516 2517 41525
rect 2475 41476 2476 41516
rect 2516 41476 2517 41516
rect 2475 41467 2517 41476
rect 2380 40468 2516 40508
rect 1228 40424 1268 40433
rect 1323 40424 1365 40433
rect 1268 40384 1324 40424
rect 1364 40384 1365 40424
rect 1228 40375 1268 40384
rect 1323 40375 1365 40384
rect 1515 39920 1557 39929
rect 1515 39880 1516 39920
rect 1556 39880 1557 39920
rect 1515 39871 1557 39880
rect 1419 39752 1461 39761
rect 1419 39712 1420 39752
rect 1460 39712 1461 39752
rect 1419 39703 1461 39712
rect 939 39500 981 39509
rect 939 39460 940 39500
rect 980 39460 981 39500
rect 939 39451 981 39460
rect 75 34880 117 34889
rect 75 34840 76 34880
rect 116 34840 117 34880
rect 75 34831 117 34840
rect 76 34721 116 34831
rect 75 34712 117 34721
rect 75 34672 76 34712
rect 116 34672 117 34712
rect 75 34663 117 34672
rect 267 34124 309 34133
rect 267 34084 268 34124
rect 308 34084 309 34124
rect 267 34075 309 34084
rect 171 32864 213 32873
rect 171 32824 172 32864
rect 212 32824 213 32864
rect 171 32815 213 32824
rect 75 29168 117 29177
rect 75 29128 76 29168
rect 116 29128 117 29168
rect 75 29119 117 29128
rect 76 13217 116 29119
rect 172 18929 212 32815
rect 268 21617 308 34075
rect 747 31604 789 31613
rect 747 31564 748 31604
rect 788 31564 789 31604
rect 747 31555 789 31564
rect 748 26657 788 31555
rect 747 26648 789 26657
rect 747 26608 748 26648
rect 788 26608 789 26648
rect 747 26599 789 26608
rect 267 21608 309 21617
rect 267 21568 268 21608
rect 308 21568 309 21608
rect 267 21559 309 21568
rect 171 18920 213 18929
rect 171 18880 172 18920
rect 212 18880 213 18920
rect 171 18871 213 18880
rect 75 13208 117 13217
rect 75 13168 76 13208
rect 116 13168 117 13208
rect 75 13159 117 13168
rect 940 2885 980 39451
rect 1323 38912 1365 38921
rect 1323 38872 1324 38912
rect 1364 38872 1365 38912
rect 1323 38863 1365 38872
rect 1324 37745 1364 38863
rect 1323 37736 1365 37745
rect 1323 37696 1324 37736
rect 1364 37696 1365 37736
rect 1323 37687 1365 37696
rect 1228 36728 1268 36737
rect 1324 36728 1364 37687
rect 1420 37493 1460 39703
rect 1516 39593 1556 39871
rect 1515 39584 1557 39593
rect 1515 39544 1516 39584
rect 1556 39544 1557 39584
rect 1515 39535 1557 39544
rect 1612 38333 1652 38364
rect 1611 38324 1653 38333
rect 1611 38284 1612 38324
rect 1652 38284 1653 38324
rect 1611 38275 1653 38284
rect 1612 38240 1652 38275
rect 1612 38081 1652 38200
rect 1611 38072 1653 38081
rect 1611 38032 1612 38072
rect 1652 38032 1653 38072
rect 1611 38023 1653 38032
rect 1419 37484 1461 37493
rect 1419 37444 1420 37484
rect 1460 37444 1461 37484
rect 1419 37435 1461 37444
rect 1419 37064 1461 37073
rect 1708 37064 1748 40459
rect 2380 40349 2420 40468
rect 2476 40466 2516 40468
rect 2572 40433 2612 44836
rect 2667 44036 2709 44045
rect 2667 43996 2668 44036
rect 2708 43996 2709 44036
rect 2667 43987 2709 43996
rect 2668 43462 2708 43987
rect 2668 43413 2708 43422
rect 2667 42860 2709 42869
rect 2667 42820 2668 42860
rect 2708 42820 2709 42860
rect 2667 42811 2709 42820
rect 2668 42726 2708 42811
rect 2667 41936 2709 41945
rect 2667 41896 2668 41936
rect 2708 41896 2709 41936
rect 2667 41887 2709 41896
rect 2668 40676 2708 41887
rect 2668 40627 2708 40636
rect 2476 40417 2516 40426
rect 2571 40424 2613 40433
rect 2571 40384 2572 40424
rect 2612 40384 2613 40424
rect 2571 40375 2613 40384
rect 2379 40340 2421 40349
rect 2379 40300 2380 40340
rect 2420 40300 2421 40340
rect 2379 40291 2421 40300
rect 2572 39845 2612 40375
rect 2667 40340 2709 40349
rect 2667 40300 2668 40340
rect 2708 40300 2709 40340
rect 2667 40291 2709 40300
rect 2571 39836 2613 39845
rect 2571 39796 2572 39836
rect 2612 39796 2613 39836
rect 2571 39787 2613 39796
rect 1996 39752 2036 39761
rect 1803 39584 1845 39593
rect 1803 39544 1804 39584
rect 1844 39544 1845 39584
rect 1803 39535 1845 39544
rect 1419 37024 1420 37064
rect 1460 37024 1461 37064
rect 1419 37015 1461 37024
rect 1516 37024 1748 37064
rect 1268 36688 1364 36728
rect 1228 36679 1268 36688
rect 1228 35888 1268 35897
rect 1323 35888 1365 35897
rect 1268 35848 1324 35888
rect 1364 35848 1365 35888
rect 1228 35839 1268 35848
rect 1323 35839 1365 35848
rect 1420 35216 1460 37015
rect 1420 34805 1460 35176
rect 1227 34796 1269 34805
rect 1227 34756 1228 34796
rect 1268 34756 1269 34796
rect 1227 34747 1269 34756
rect 1419 34796 1461 34805
rect 1419 34756 1420 34796
rect 1460 34756 1461 34796
rect 1419 34747 1461 34756
rect 1131 34040 1173 34049
rect 1131 34000 1132 34040
rect 1172 34000 1173 34040
rect 1131 33991 1173 34000
rect 1132 29849 1172 33991
rect 1228 31352 1268 34747
rect 1419 33200 1461 33209
rect 1419 33160 1420 33200
rect 1460 33160 1461 33200
rect 1419 33151 1461 33160
rect 1228 31303 1268 31312
rect 1420 31100 1460 33151
rect 1324 31060 1460 31100
rect 1131 29840 1173 29849
rect 1131 29800 1132 29840
rect 1172 29800 1173 29840
rect 1131 29791 1173 29800
rect 1228 29840 1268 29849
rect 1324 29840 1364 31060
rect 1419 30680 1461 30689
rect 1419 30640 1420 30680
rect 1460 30640 1461 30680
rect 1419 30631 1461 30640
rect 1420 30269 1460 30631
rect 1419 30260 1461 30269
rect 1419 30220 1420 30260
rect 1460 30220 1461 30260
rect 1419 30211 1461 30220
rect 1268 29800 1364 29840
rect 1228 29791 1268 29800
rect 1035 29084 1077 29093
rect 1035 29044 1036 29084
rect 1076 29044 1077 29084
rect 1035 29035 1077 29044
rect 1036 26069 1076 29035
rect 1516 29000 1556 37024
rect 1611 36896 1653 36905
rect 1611 36856 1612 36896
rect 1652 36856 1653 36896
rect 1611 36847 1653 36856
rect 1324 28960 1556 29000
rect 1612 30680 1652 36847
rect 1707 33704 1749 33713
rect 1707 33664 1708 33704
rect 1748 33664 1749 33704
rect 1707 33655 1749 33664
rect 1708 33570 1748 33655
rect 1707 30932 1749 30941
rect 1707 30892 1708 30932
rect 1748 30892 1749 30932
rect 1707 30883 1749 30892
rect 1708 30848 1748 30883
rect 1708 30797 1748 30808
rect 1228 28328 1268 28337
rect 1228 28244 1268 28288
rect 1324 28253 1364 28960
rect 1612 28328 1652 30640
rect 1707 30260 1749 30269
rect 1707 30220 1708 30260
rect 1748 30220 1749 30260
rect 1707 30211 1749 30220
rect 1708 28496 1748 30211
rect 1804 28580 1844 39535
rect 1996 39089 2036 39712
rect 2092 39752 2132 39761
rect 1995 39080 2037 39089
rect 1995 39040 1996 39080
rect 2036 39040 2037 39080
rect 1995 39031 2037 39040
rect 1995 38912 2037 38921
rect 1995 38872 1996 38912
rect 2036 38872 2037 38912
rect 1995 38863 2037 38872
rect 1996 38669 2036 38863
rect 1995 38660 2037 38669
rect 1995 38620 1996 38660
rect 2036 38620 2037 38660
rect 1995 38611 2037 38620
rect 1899 37484 1941 37493
rect 1899 37444 1900 37484
rect 1940 37444 1941 37484
rect 1899 37435 1941 37444
rect 1900 35897 1940 37435
rect 2092 36401 2132 39712
rect 2476 39668 2516 39677
rect 2188 39628 2476 39668
rect 2091 36392 2133 36401
rect 2091 36352 2092 36392
rect 2132 36352 2133 36392
rect 2091 36343 2133 36352
rect 2188 36149 2228 39628
rect 2476 39619 2516 39628
rect 2572 39668 2612 39677
rect 2283 38240 2325 38249
rect 2283 38200 2284 38240
rect 2324 38200 2325 38240
rect 2283 38191 2325 38200
rect 2284 36653 2324 38191
rect 2572 37913 2612 39628
rect 2668 39416 2708 40291
rect 2764 39593 2804 47188
rect 2860 47312 2900 48187
rect 2860 43541 2900 47272
rect 2956 46640 2996 49447
rect 3051 48740 3093 48749
rect 3051 48700 3052 48740
rect 3092 48700 3093 48740
rect 3051 48691 3093 48700
rect 3052 48606 3092 48691
rect 3244 48488 3284 49456
rect 3052 48448 3284 48488
rect 3052 47321 3092 48448
rect 3147 48320 3189 48329
rect 3147 48280 3148 48320
rect 3188 48280 3189 48320
rect 3147 48271 3189 48280
rect 3051 47312 3093 47321
rect 3051 47272 3052 47312
rect 3092 47272 3093 47312
rect 3051 47263 3093 47272
rect 2956 46600 3092 46640
rect 3052 44960 3092 46600
rect 3052 44801 3092 44920
rect 3051 44792 3093 44801
rect 3051 44752 3052 44792
rect 3092 44752 3093 44792
rect 3051 44743 3093 44752
rect 3148 43625 3188 48271
rect 3243 48152 3285 48161
rect 3243 48112 3244 48152
rect 3284 48112 3285 48152
rect 3243 48103 3285 48112
rect 3244 47984 3284 48103
rect 3244 47935 3284 47944
rect 3340 47564 3380 49540
rect 3436 49531 3476 49540
rect 3532 49580 3572 50464
rect 4012 50093 4052 50959
rect 4107 50840 4149 50849
rect 4107 50800 4108 50840
rect 4148 50800 4149 50840
rect 4107 50791 4149 50800
rect 4011 50084 4053 50093
rect 4011 50044 4012 50084
rect 4052 50044 4053 50084
rect 4011 50035 4053 50044
rect 3688 49916 4056 49925
rect 3728 49876 3770 49916
rect 3810 49876 3852 49916
rect 3892 49876 3934 49916
rect 3974 49876 4016 49916
rect 3688 49867 4056 49876
rect 3435 49076 3477 49085
rect 3435 49036 3436 49076
rect 3476 49036 3477 49076
rect 3435 49027 3477 49036
rect 3436 48824 3476 49027
rect 3436 48775 3476 48784
rect 3435 47816 3477 47825
rect 3435 47776 3436 47816
rect 3476 47776 3477 47816
rect 3435 47767 3477 47776
rect 3436 47682 3476 47767
rect 3340 47524 3476 47564
rect 3339 47312 3381 47321
rect 3339 47272 3340 47312
rect 3380 47272 3381 47312
rect 3339 47263 3381 47272
rect 3340 46640 3380 47263
rect 3244 46600 3380 46640
rect 3147 43616 3189 43625
rect 3147 43576 3148 43616
rect 3188 43576 3189 43616
rect 3147 43567 3189 43576
rect 2859 43532 2901 43541
rect 2859 43492 2860 43532
rect 2900 43492 2901 43532
rect 2859 43483 2901 43492
rect 3148 43448 3188 43457
rect 3244 43448 3284 46600
rect 3436 45044 3476 47524
rect 3532 45128 3572 49540
rect 3916 49496 3956 49507
rect 3916 49421 3956 49456
rect 4012 49496 4052 49505
rect 4108 49496 4148 50791
rect 4052 49456 4148 49496
rect 4012 49447 4052 49456
rect 4204 49421 4244 51556
rect 4299 51260 4341 51269
rect 4299 51220 4300 51260
rect 4340 51220 4341 51260
rect 4299 51211 4341 51220
rect 4300 50345 4340 51211
rect 4299 50336 4341 50345
rect 4492 50336 4532 53404
rect 4588 51437 4628 57856
rect 4684 57847 4724 57856
rect 4683 56552 4725 56561
rect 4683 56512 4684 56552
rect 4724 56512 4725 56552
rect 4683 56503 4725 56512
rect 4684 56384 4724 56503
rect 4684 55721 4724 56344
rect 4780 56384 4820 59863
rect 4928 59744 5296 59753
rect 4968 59704 5010 59744
rect 5050 59704 5092 59744
rect 5132 59704 5174 59744
rect 5214 59704 5256 59744
rect 4928 59695 5296 59704
rect 5164 59408 5204 59417
rect 5356 59408 5396 59872
rect 5204 59368 5396 59408
rect 5164 59359 5204 59368
rect 5356 59249 5396 59368
rect 5451 59408 5493 59417
rect 5451 59368 5452 59408
rect 5492 59368 5493 59408
rect 5451 59359 5493 59368
rect 5355 59240 5397 59249
rect 5355 59200 5356 59240
rect 5396 59200 5397 59240
rect 5355 59191 5397 59200
rect 4971 58736 5013 58745
rect 4971 58696 4972 58736
rect 5012 58696 5013 58736
rect 4971 58687 5013 58696
rect 4972 58568 5012 58687
rect 5355 58652 5397 58661
rect 5355 58612 5356 58652
rect 5396 58612 5397 58652
rect 5355 58603 5397 58612
rect 4972 58519 5012 58528
rect 5356 58568 5396 58603
rect 5356 58517 5396 58528
rect 5164 58409 5204 58494
rect 5163 58400 5205 58409
rect 5163 58360 5164 58400
rect 5204 58360 5205 58400
rect 5163 58351 5205 58360
rect 4928 58232 5296 58241
rect 4968 58192 5010 58232
rect 5050 58192 5092 58232
rect 5132 58192 5174 58232
rect 5214 58192 5256 58232
rect 4928 58183 5296 58192
rect 5067 57980 5109 57989
rect 5067 57940 5068 57980
rect 5108 57940 5109 57980
rect 5067 57931 5109 57940
rect 5356 57980 5396 57989
rect 5452 57980 5492 59359
rect 5547 58400 5589 58409
rect 5547 58360 5548 58400
rect 5588 58360 5589 58400
rect 5547 58351 5589 58360
rect 5396 57940 5492 57980
rect 5356 57931 5396 57940
rect 5068 57056 5108 57931
rect 5212 57886 5252 57895
rect 5548 57886 5588 58351
rect 5252 57846 5588 57886
rect 5212 57837 5252 57846
rect 5452 57065 5492 57150
rect 5068 57007 5108 57016
rect 5451 57056 5493 57065
rect 5451 57016 5452 57056
rect 5492 57016 5493 57056
rect 5451 57007 5493 57016
rect 5260 56888 5300 56897
rect 5644 56888 5684 61039
rect 5835 60584 5877 60593
rect 5835 60544 5836 60584
rect 5876 60544 5877 60584
rect 5835 60535 5877 60544
rect 5739 60248 5781 60257
rect 5739 60208 5740 60248
rect 5780 60208 5781 60248
rect 5739 60199 5781 60208
rect 5740 57065 5780 60199
rect 5739 57056 5781 57065
rect 5739 57016 5740 57056
rect 5780 57016 5781 57056
rect 5739 57007 5781 57016
rect 5300 56848 5396 56888
rect 5260 56839 5300 56848
rect 4928 56720 5296 56729
rect 4968 56680 5010 56720
rect 5050 56680 5092 56720
rect 5132 56680 5174 56720
rect 5214 56680 5256 56720
rect 4928 56671 5296 56680
rect 4780 56335 4820 56344
rect 5356 56216 5396 56848
rect 5164 56176 5396 56216
rect 5452 56848 5684 56888
rect 4683 55712 4725 55721
rect 4683 55672 4684 55712
rect 4724 55672 4725 55712
rect 4683 55663 4725 55672
rect 4684 55544 4724 55555
rect 4684 55469 4724 55504
rect 5164 55544 5204 56176
rect 5259 55712 5301 55721
rect 5259 55672 5260 55712
rect 5300 55672 5301 55712
rect 5259 55663 5301 55672
rect 5164 55495 5204 55504
rect 5260 55544 5300 55663
rect 4683 55460 4725 55469
rect 4683 55420 4684 55460
rect 4724 55420 4725 55460
rect 5260 55460 5300 55504
rect 5260 55420 5396 55460
rect 4683 55411 4725 55420
rect 4587 51428 4629 51437
rect 4587 51388 4588 51428
rect 4628 51388 4629 51428
rect 4587 51379 4629 51388
rect 4587 51260 4629 51269
rect 4587 51220 4588 51260
rect 4628 51220 4629 51260
rect 4587 51211 4629 51220
rect 4588 51008 4628 51211
rect 4588 50959 4628 50968
rect 4684 50588 4724 55411
rect 4876 55376 4916 55385
rect 4780 55336 4876 55376
rect 4780 54704 4820 55336
rect 4876 55327 4916 55336
rect 4928 55208 5296 55217
rect 4968 55168 5010 55208
rect 5050 55168 5092 55208
rect 5132 55168 5174 55208
rect 5214 55168 5256 55208
rect 4928 55159 5296 55168
rect 5067 55040 5109 55049
rect 5067 55000 5068 55040
rect 5108 55000 5109 55040
rect 5067 54991 5109 55000
rect 4780 54664 4916 54704
rect 4779 54368 4821 54377
rect 4779 54328 4780 54368
rect 4820 54328 4821 54368
rect 4779 54319 4821 54328
rect 4780 53528 4820 54319
rect 4876 54046 4916 54664
rect 4876 53997 4916 54006
rect 5068 53948 5108 54991
rect 5356 54881 5396 55420
rect 5355 54872 5397 54881
rect 5355 54832 5356 54872
rect 5396 54832 5397 54872
rect 5355 54823 5397 54832
rect 5452 54872 5492 56848
rect 5739 56552 5781 56561
rect 5739 56512 5740 56552
rect 5780 56512 5781 56552
rect 5739 56503 5781 56512
rect 5740 56384 5780 56503
rect 5740 56335 5780 56344
rect 5643 56300 5685 56309
rect 5643 56260 5644 56300
rect 5684 56260 5685 56300
rect 5643 56251 5685 56260
rect 5644 55628 5684 56251
rect 5739 56132 5781 56141
rect 5739 56092 5740 56132
rect 5780 56092 5781 56132
rect 5739 56083 5781 56092
rect 5644 55579 5684 55588
rect 5740 55628 5780 56083
rect 5740 55579 5780 55588
rect 5836 55460 5876 60535
rect 5068 53899 5108 53908
rect 4928 53696 5296 53705
rect 4968 53656 5010 53696
rect 5050 53656 5092 53696
rect 5132 53656 5174 53696
rect 5214 53656 5256 53696
rect 4928 53647 5296 53656
rect 4780 53488 4916 53528
rect 4779 53360 4821 53369
rect 4779 53320 4780 53360
rect 4820 53320 4821 53360
rect 4779 53311 4821 53320
rect 4876 53360 4916 53488
rect 4876 53311 4916 53320
rect 4780 53226 4820 53311
rect 5067 53276 5109 53285
rect 5067 53236 5068 53276
rect 5108 53236 5109 53276
rect 5067 53227 5109 53236
rect 4779 53024 4821 53033
rect 4779 52984 4780 53024
rect 4820 52984 4821 53024
rect 4779 52975 4821 52984
rect 4780 51017 4820 52975
rect 5068 52520 5108 53227
rect 5452 52520 5492 54832
rect 5548 55420 5876 55460
rect 5548 53873 5588 55420
rect 5932 53957 5972 62560
rect 5931 53948 5973 53957
rect 5931 53908 5932 53948
rect 5972 53908 5973 53948
rect 5931 53899 5973 53908
rect 5547 53864 5589 53873
rect 5547 53824 5548 53864
rect 5588 53824 5589 53864
rect 5547 53815 5589 53824
rect 5548 52949 5588 53815
rect 5836 53360 5876 53369
rect 5836 53033 5876 53320
rect 5835 53024 5877 53033
rect 5835 52984 5836 53024
rect 5876 52984 5877 53024
rect 5835 52975 5877 52984
rect 5547 52940 5589 52949
rect 5547 52900 5548 52940
rect 5588 52900 5589 52940
rect 5547 52891 5589 52900
rect 5547 52520 5589 52529
rect 5452 52480 5548 52520
rect 5588 52480 5589 52520
rect 5068 52471 5108 52480
rect 5547 52471 5589 52480
rect 5260 52352 5300 52361
rect 5300 52312 5396 52352
rect 5260 52303 5300 52312
rect 4928 52184 5296 52193
rect 4968 52144 5010 52184
rect 5050 52144 5092 52184
rect 5132 52144 5174 52184
rect 5214 52144 5256 52184
rect 4928 52135 5296 52144
rect 4971 51428 5013 51437
rect 4971 51388 4972 51428
rect 5012 51388 5013 51428
rect 4971 51379 5013 51388
rect 4779 51008 4821 51017
rect 4779 50968 4780 51008
rect 4820 50968 4821 51008
rect 4779 50959 4821 50968
rect 4779 50840 4821 50849
rect 4779 50800 4780 50840
rect 4820 50800 4821 50840
rect 4972 50840 5012 51379
rect 5356 51008 5396 52312
rect 5356 50959 5396 50968
rect 5452 51008 5492 51017
rect 4972 50800 5396 50840
rect 4779 50791 4821 50800
rect 4780 50706 4820 50791
rect 4928 50672 5296 50681
rect 4968 50632 5010 50672
rect 5050 50632 5092 50672
rect 5132 50632 5174 50672
rect 5214 50632 5256 50672
rect 4928 50623 5296 50632
rect 4299 50296 4300 50336
rect 4340 50296 4341 50336
rect 4299 50287 4341 50296
rect 4396 50296 4532 50336
rect 4588 50548 4724 50588
rect 4299 50084 4341 50093
rect 4299 50044 4300 50084
rect 4340 50044 4341 50084
rect 4299 50035 4341 50044
rect 3915 49412 3957 49421
rect 3915 49372 3916 49412
rect 3956 49372 3957 49412
rect 3915 49363 3957 49372
rect 4203 49412 4245 49421
rect 4203 49372 4204 49412
rect 4244 49372 4245 49412
rect 4203 49363 4245 49372
rect 3688 48404 4056 48413
rect 3728 48364 3770 48404
rect 3810 48364 3852 48404
rect 3892 48364 3934 48404
rect 3974 48364 4016 48404
rect 3688 48355 4056 48364
rect 3627 48152 3669 48161
rect 3627 48112 3628 48152
rect 3668 48112 3669 48152
rect 3627 48103 3669 48112
rect 3628 47993 3668 48103
rect 3627 47984 3669 47993
rect 3627 47944 3628 47984
rect 3668 47944 3669 47984
rect 3627 47935 3669 47944
rect 3628 47850 3668 47935
rect 3819 47816 3861 47825
rect 3819 47776 3820 47816
rect 3860 47776 3861 47816
rect 3819 47767 3861 47776
rect 3820 47307 3860 47767
rect 3820 47258 3860 47267
rect 4012 47396 4052 47405
rect 4012 47237 4052 47356
rect 4011 47228 4053 47237
rect 4011 47188 4012 47228
rect 4052 47188 4053 47228
rect 4011 47179 4053 47188
rect 3688 46892 4056 46901
rect 3728 46852 3770 46892
rect 3810 46852 3852 46892
rect 3892 46852 3934 46892
rect 3974 46852 4016 46892
rect 3688 46843 4056 46852
rect 4011 46304 4053 46313
rect 4011 46264 4012 46304
rect 4052 46264 4053 46304
rect 4011 46255 4053 46264
rect 3916 45800 3956 45809
rect 3916 45641 3956 45760
rect 3915 45632 3957 45641
rect 3915 45592 3916 45632
rect 3956 45592 3957 45632
rect 4012 45632 4052 46255
rect 4107 45884 4149 45893
rect 4107 45844 4108 45884
rect 4148 45844 4149 45884
rect 4107 45835 4149 45844
rect 4108 45800 4148 45835
rect 4108 45749 4148 45760
rect 4012 45592 4148 45632
rect 3915 45583 3957 45592
rect 3688 45380 4056 45389
rect 3728 45340 3770 45380
rect 3810 45340 3852 45380
rect 3892 45340 3934 45380
rect 3974 45340 4016 45380
rect 3688 45331 4056 45340
rect 3532 45088 3668 45128
rect 3436 45004 3572 45044
rect 3532 44960 3572 45004
rect 3628 44969 3668 45088
rect 3532 44885 3572 44920
rect 3627 44960 3669 44969
rect 3627 44920 3628 44960
rect 3668 44920 3669 44960
rect 3627 44911 3669 44920
rect 4011 44960 4053 44969
rect 4011 44920 4012 44960
rect 4052 44920 4053 44960
rect 4011 44911 4053 44920
rect 4108 44960 4148 45592
rect 4108 44911 4148 44920
rect 3531 44876 3573 44885
rect 3531 44836 3532 44876
rect 3572 44836 3573 44876
rect 3531 44827 3573 44836
rect 3532 44796 3572 44827
rect 3628 44826 3668 44911
rect 3819 44708 3861 44717
rect 3819 44668 3820 44708
rect 3860 44668 3861 44708
rect 3819 44659 3861 44668
rect 3627 44288 3669 44297
rect 3532 44248 3628 44288
rect 3668 44248 3669 44288
rect 3435 43532 3477 43541
rect 3435 43492 3436 43532
rect 3476 43492 3477 43532
rect 3435 43483 3477 43492
rect 2956 43408 3148 43448
rect 3188 43408 3284 43448
rect 2956 42785 2996 43408
rect 3148 43399 3188 43408
rect 3243 42944 3285 42953
rect 3243 42904 3244 42944
rect 3284 42904 3285 42944
rect 3243 42895 3285 42904
rect 2955 42776 2997 42785
rect 2955 42736 2956 42776
rect 2996 42736 2997 42776
rect 2955 42727 2997 42736
rect 3244 42776 3284 42895
rect 3244 42727 3284 42736
rect 2956 41936 2996 42727
rect 3436 42020 3476 43483
rect 3532 42953 3572 44248
rect 3627 44239 3669 44248
rect 3820 44288 3860 44659
rect 3820 44239 3860 44248
rect 3628 44154 3668 44239
rect 4012 44045 4052 44911
rect 4300 44717 4340 50035
rect 4396 49085 4436 50296
rect 4491 50084 4533 50093
rect 4491 50044 4492 50084
rect 4532 50044 4533 50084
rect 4491 50035 4533 50044
rect 4492 49950 4532 50035
rect 4491 49412 4533 49421
rect 4491 49372 4492 49412
rect 4532 49372 4533 49412
rect 4491 49363 4533 49372
rect 4395 49076 4437 49085
rect 4395 49036 4396 49076
rect 4436 49036 4437 49076
rect 4395 49027 4437 49036
rect 4396 46472 4436 49027
rect 4492 46640 4532 49363
rect 4588 49337 4628 50548
rect 4683 50420 4725 50429
rect 4683 50380 4684 50420
rect 4724 50380 4725 50420
rect 4683 50371 4725 50380
rect 4684 50286 4724 50371
rect 5356 50336 5396 50800
rect 5452 50597 5492 50968
rect 5451 50588 5493 50597
rect 5451 50548 5452 50588
rect 5492 50548 5493 50588
rect 5451 50539 5493 50548
rect 4876 50322 4916 50331
rect 4876 50093 4916 50282
rect 4875 50084 4917 50093
rect 4875 50044 4876 50084
rect 4916 50044 4917 50084
rect 4875 50035 4917 50044
rect 5356 49505 5396 50296
rect 5355 49496 5397 49505
rect 5355 49456 5356 49496
rect 5396 49456 5397 49496
rect 5355 49447 5397 49456
rect 4587 49328 4629 49337
rect 4587 49288 4588 49328
rect 4628 49288 4629 49328
rect 4587 49279 4629 49288
rect 4588 48824 4628 49279
rect 4928 49160 5296 49169
rect 4968 49120 5010 49160
rect 5050 49120 5092 49160
rect 5132 49120 5174 49160
rect 5214 49120 5256 49160
rect 4928 49111 5296 49120
rect 5355 49076 5397 49085
rect 5355 49036 5356 49076
rect 5396 49036 5397 49076
rect 5355 49027 5397 49036
rect 4684 48824 4724 48833
rect 4588 48784 4684 48824
rect 4684 48775 4724 48784
rect 5067 48824 5109 48833
rect 5067 48784 5068 48824
rect 5108 48784 5109 48824
rect 5067 48775 5109 48784
rect 4876 48572 4916 48581
rect 4780 48532 4876 48572
rect 4780 47312 4820 48532
rect 4876 48523 4916 48532
rect 4875 48320 4917 48329
rect 4875 48280 4876 48320
rect 4916 48280 4917 48320
rect 4875 48271 4917 48280
rect 4876 47984 4916 48271
rect 5068 48161 5108 48775
rect 5259 48740 5301 48749
rect 5259 48700 5260 48740
rect 5300 48700 5301 48740
rect 5259 48691 5301 48700
rect 5067 48152 5109 48161
rect 5067 48112 5068 48152
rect 5108 48112 5109 48152
rect 5067 48103 5109 48112
rect 4876 47935 4916 47944
rect 5067 47900 5109 47909
rect 5067 47860 5068 47900
rect 5108 47860 5109 47900
rect 5067 47851 5109 47860
rect 5260 47900 5300 48691
rect 5356 48329 5396 49027
rect 5548 48497 5588 52471
rect 5932 51848 5972 53899
rect 5740 51808 5932 51848
rect 5740 48497 5780 51808
rect 5932 51799 5972 51808
rect 6028 51680 6068 62887
rect 6124 61592 6164 63316
rect 6220 64828 6356 64868
rect 6220 61676 6260 64828
rect 6412 64784 6452 65239
rect 6603 65204 6645 65213
rect 6603 65164 6604 65204
rect 6644 65164 6645 65204
rect 6603 65155 6645 65164
rect 6316 64744 6452 64784
rect 6316 62441 6356 64744
rect 6508 63944 6548 63953
rect 6315 62432 6357 62441
rect 6315 62392 6316 62432
rect 6356 62392 6357 62432
rect 6315 62383 6357 62392
rect 6220 61627 6260 61636
rect 6124 59912 6164 61552
rect 6124 59872 6260 59912
rect 6123 57980 6165 57989
rect 6123 57940 6124 57980
rect 6164 57940 6165 57980
rect 6123 57931 6165 57940
rect 5932 51640 6068 51680
rect 5932 51092 5972 51640
rect 6124 51269 6164 57931
rect 6220 56141 6260 59872
rect 6316 58157 6356 62383
rect 6508 61601 6548 63904
rect 6507 61592 6549 61601
rect 6507 61552 6508 61592
rect 6548 61552 6549 61592
rect 6507 61543 6549 61552
rect 6604 61097 6644 65155
rect 6795 65120 6837 65129
rect 6795 65080 6796 65120
rect 6836 65080 6837 65120
rect 6795 65071 6837 65080
rect 6699 64700 6741 64709
rect 6699 64660 6700 64700
rect 6740 64660 6741 64700
rect 6699 64651 6741 64660
rect 6700 63197 6740 64651
rect 6796 64616 6836 65071
rect 6796 64457 6836 64576
rect 6795 64448 6837 64457
rect 6795 64408 6796 64448
rect 6836 64408 6837 64448
rect 6795 64399 6837 64408
rect 6795 64112 6837 64121
rect 6795 64072 6796 64112
rect 6836 64072 6837 64112
rect 6795 64063 6837 64072
rect 6699 63188 6741 63197
rect 6699 63148 6700 63188
rect 6740 63148 6741 63188
rect 6699 63139 6741 63148
rect 6699 61592 6741 61601
rect 6699 61552 6700 61592
rect 6740 61552 6741 61592
rect 6699 61543 6741 61552
rect 6700 61458 6740 61543
rect 6699 61340 6741 61349
rect 6699 61300 6700 61340
rect 6740 61300 6741 61340
rect 6699 61291 6741 61300
rect 6603 61088 6645 61097
rect 6603 61048 6604 61088
rect 6644 61048 6645 61088
rect 6603 61039 6645 61048
rect 6604 60920 6644 60929
rect 6411 60416 6453 60425
rect 6411 60376 6412 60416
rect 6452 60376 6453 60416
rect 6411 60367 6453 60376
rect 6412 59408 6452 60367
rect 6604 60341 6644 60880
rect 6700 60761 6740 61291
rect 6796 61181 6836 64063
rect 6892 62609 6932 65668
rect 7084 65540 7124 67087
rect 7180 66893 7220 67600
rect 7371 67556 7413 67565
rect 7371 67516 7372 67556
rect 7412 67516 7413 67556
rect 7371 67507 7413 67516
rect 7179 66884 7221 66893
rect 7179 66844 7180 66884
rect 7220 66844 7221 66884
rect 7179 66835 7221 66844
rect 7180 66296 7220 66305
rect 7180 65801 7220 66256
rect 7179 65792 7221 65801
rect 7179 65752 7180 65792
rect 7220 65752 7221 65792
rect 7179 65743 7221 65752
rect 7084 65500 7220 65540
rect 6988 65456 7028 65465
rect 7028 65416 7124 65456
rect 6988 65407 7028 65416
rect 6987 65288 7029 65297
rect 6987 65248 6988 65288
rect 7028 65248 7029 65288
rect 6987 65239 7029 65248
rect 6988 65154 7028 65239
rect 6988 64448 7028 64457
rect 6988 63939 7028 64408
rect 7084 63953 7124 65416
rect 7180 65381 7220 65500
rect 7275 65456 7317 65465
rect 7275 65416 7276 65456
rect 7316 65416 7317 65456
rect 7275 65407 7317 65416
rect 7179 65372 7221 65381
rect 7179 65332 7180 65372
rect 7220 65332 7221 65372
rect 7179 65323 7221 65332
rect 7276 65322 7316 65407
rect 7372 65204 7412 67507
rect 7276 65164 7412 65204
rect 7179 64532 7221 64541
rect 7179 64492 7180 64532
rect 7220 64492 7221 64532
rect 7179 64483 7221 64492
rect 7180 64398 7220 64483
rect 7179 64112 7221 64121
rect 7179 64072 7180 64112
rect 7220 64072 7221 64112
rect 7179 64063 7221 64072
rect 7180 63978 7220 64063
rect 6988 63890 7028 63899
rect 7083 63944 7125 63953
rect 7083 63904 7084 63944
rect 7124 63904 7125 63944
rect 7083 63895 7125 63904
rect 7084 63785 7124 63895
rect 7083 63776 7125 63785
rect 7083 63736 7084 63776
rect 7124 63736 7125 63776
rect 7083 63727 7125 63736
rect 6987 63692 7029 63701
rect 6987 63652 6988 63692
rect 7028 63652 7029 63692
rect 6987 63643 7029 63652
rect 6891 62600 6933 62609
rect 6891 62560 6892 62600
rect 6932 62560 6933 62600
rect 6891 62551 6933 62560
rect 6891 62432 6933 62441
rect 6891 62392 6892 62432
rect 6932 62392 6933 62432
rect 6891 62383 6933 62392
rect 6795 61172 6837 61181
rect 6795 61132 6796 61172
rect 6836 61132 6837 61172
rect 6795 61123 6837 61132
rect 6796 61004 6836 61015
rect 6796 60929 6836 60964
rect 6795 60920 6837 60929
rect 6795 60880 6796 60920
rect 6836 60880 6837 60920
rect 6795 60871 6837 60880
rect 6699 60752 6741 60761
rect 6699 60712 6700 60752
rect 6740 60712 6741 60752
rect 6699 60703 6741 60712
rect 6603 60332 6645 60341
rect 6603 60292 6604 60332
rect 6644 60292 6645 60332
rect 6603 60283 6645 60292
rect 6604 60080 6644 60283
rect 6315 58148 6357 58157
rect 6315 58108 6316 58148
rect 6356 58108 6357 58148
rect 6315 58099 6357 58108
rect 6315 57896 6357 57905
rect 6315 57856 6316 57896
rect 6356 57856 6357 57896
rect 6315 57847 6357 57856
rect 6316 57762 6356 57847
rect 6315 57644 6357 57653
rect 6315 57604 6316 57644
rect 6356 57604 6357 57644
rect 6315 57595 6357 57604
rect 6219 56132 6261 56141
rect 6219 56092 6220 56132
rect 6260 56092 6261 56132
rect 6219 56083 6261 56092
rect 6220 55544 6260 55553
rect 6220 55133 6260 55504
rect 6316 55460 6356 57595
rect 6412 55544 6452 59368
rect 6508 60040 6604 60080
rect 6508 57056 6548 60040
rect 6604 60031 6644 60040
rect 6604 59156 6644 59165
rect 6604 58829 6644 59116
rect 6603 58820 6645 58829
rect 6603 58780 6604 58820
rect 6644 58780 6645 58820
rect 6603 58771 6645 58780
rect 6604 58568 6644 58577
rect 6604 57989 6644 58528
rect 6700 58493 6740 60703
rect 6892 60173 6932 62383
rect 6988 61685 7028 63643
rect 7179 63188 7221 63197
rect 7179 63148 7180 63188
rect 7220 63148 7221 63188
rect 7179 63139 7221 63148
rect 7180 63104 7220 63139
rect 7180 63053 7220 63064
rect 7083 62684 7125 62693
rect 7083 62644 7084 62684
rect 7124 62644 7125 62684
rect 7083 62635 7125 62644
rect 7084 62432 7124 62635
rect 7276 62441 7316 65164
rect 7372 64616 7412 64625
rect 7372 64457 7412 64576
rect 7371 64448 7413 64457
rect 7371 64408 7372 64448
rect 7412 64408 7413 64448
rect 7371 64399 7413 64408
rect 7372 63953 7412 64399
rect 7371 63944 7413 63953
rect 7371 63904 7372 63944
rect 7412 63904 7413 63944
rect 7371 63895 7413 63904
rect 7468 63701 7508 70372
rect 7852 70169 7892 73060
rect 7948 72353 7988 76504
rect 8140 76040 8180 76504
rect 8140 75991 8180 76000
rect 8235 76040 8277 76049
rect 8235 76000 8236 76040
rect 8276 76000 8277 76040
rect 8235 75991 8277 76000
rect 8043 74528 8085 74537
rect 8043 74488 8044 74528
rect 8084 74488 8085 74528
rect 8043 74479 8085 74488
rect 8044 73520 8084 74479
rect 8236 74369 8276 75991
rect 8235 74360 8277 74369
rect 8235 74320 8236 74360
rect 8276 74320 8277 74360
rect 8235 74311 8277 74320
rect 8332 74192 8372 77167
rect 8428 76712 8468 77251
rect 8428 76663 8468 76672
rect 8524 76712 8564 77503
rect 8427 76544 8469 76553
rect 8427 76504 8428 76544
rect 8468 76504 8469 76544
rect 8427 76495 8469 76504
rect 8044 73471 8084 73480
rect 8140 74152 8372 74192
rect 8043 73352 8085 73361
rect 8043 73312 8044 73352
rect 8084 73312 8085 73352
rect 8043 73303 8085 73312
rect 8044 73016 8084 73303
rect 8044 72967 8084 72976
rect 7947 72344 7989 72353
rect 7947 72304 7948 72344
rect 7988 72304 7989 72344
rect 7947 72295 7989 72304
rect 8140 72176 8180 74152
rect 8236 73688 8276 73697
rect 8428 73688 8468 76495
rect 8524 76049 8564 76672
rect 8620 76553 8660 78268
rect 8811 78224 8853 78233
rect 8811 78184 8812 78224
rect 8852 78184 8853 78224
rect 8811 78175 8853 78184
rect 8908 78224 8948 78233
rect 8812 77552 8852 78175
rect 8812 77503 8852 77512
rect 8715 77468 8757 77477
rect 8715 77428 8716 77468
rect 8756 77428 8757 77468
rect 8715 77419 8757 77428
rect 8619 76544 8661 76553
rect 8619 76504 8620 76544
rect 8660 76504 8661 76544
rect 8619 76495 8661 76504
rect 8523 76040 8565 76049
rect 8523 76000 8524 76040
rect 8564 76000 8565 76040
rect 8523 75991 8565 76000
rect 8716 76040 8756 77419
rect 8811 76880 8853 76889
rect 8811 76840 8812 76880
rect 8852 76840 8853 76880
rect 8811 76831 8853 76840
rect 8619 75956 8661 75965
rect 8619 75916 8620 75956
rect 8660 75916 8661 75956
rect 8619 75907 8661 75916
rect 8620 75822 8660 75907
rect 8716 74705 8756 76000
rect 8812 75797 8852 76831
rect 8908 76721 8948 78184
rect 9004 77477 9044 78268
rect 9003 77468 9045 77477
rect 9003 77428 9004 77468
rect 9044 77428 9045 77468
rect 9003 77419 9045 77428
rect 9004 76796 9044 77419
rect 9004 76747 9044 76756
rect 8907 76712 8949 76721
rect 8907 76672 8908 76712
rect 8948 76672 8949 76712
rect 8907 76663 8949 76672
rect 8908 75965 8948 76663
rect 8907 75956 8949 75965
rect 8907 75916 8908 75956
rect 8948 75916 8949 75956
rect 8907 75907 8949 75916
rect 8811 75788 8853 75797
rect 8811 75748 8812 75788
rect 8852 75748 8853 75788
rect 8811 75739 8853 75748
rect 8715 74696 8757 74705
rect 8715 74656 8716 74696
rect 8756 74656 8757 74696
rect 8715 74647 8757 74656
rect 8619 74612 8661 74621
rect 8619 74572 8620 74612
rect 8660 74572 8661 74612
rect 8812 74612 8852 75739
rect 9100 75713 9140 83476
rect 9196 80669 9236 83728
rect 9292 82265 9332 85936
rect 9291 82256 9333 82265
rect 9291 82216 9292 82256
rect 9332 82216 9333 82256
rect 9291 82207 9333 82216
rect 9484 82088 9524 85936
rect 9579 85784 9621 85793
rect 9579 85744 9580 85784
rect 9620 85744 9621 85784
rect 9579 85735 9621 85744
rect 9580 83768 9620 85735
rect 9676 84449 9716 85936
rect 9868 84533 9908 85936
rect 9963 85868 10005 85877
rect 9963 85828 9964 85868
rect 10004 85828 10005 85868
rect 10060 85868 10100 85936
rect 10060 85828 10196 85868
rect 9963 85819 10005 85828
rect 9867 84524 9909 84533
rect 9867 84484 9868 84524
rect 9908 84484 9909 84524
rect 9867 84475 9909 84484
rect 9675 84440 9717 84449
rect 9675 84400 9676 84440
rect 9716 84400 9717 84440
rect 9675 84391 9717 84400
rect 9964 83768 10004 85819
rect 10060 83768 10100 83777
rect 9964 83728 10060 83768
rect 9580 83719 9620 83728
rect 10060 83719 10100 83728
rect 9771 83516 9813 83525
rect 9771 83476 9772 83516
rect 9812 83476 9813 83516
rect 9771 83467 9813 83476
rect 9772 83382 9812 83467
rect 9292 82048 9524 82088
rect 9195 80660 9237 80669
rect 9195 80620 9196 80660
rect 9236 80620 9237 80660
rect 9195 80611 9237 80620
rect 9196 79736 9236 79745
rect 9196 79073 9236 79696
rect 9195 79064 9237 79073
rect 9195 79024 9196 79064
rect 9236 79024 9237 79064
rect 9195 79015 9237 79024
rect 9292 77981 9332 82048
rect 9483 81836 9525 81845
rect 9483 81796 9484 81836
rect 9524 81796 9525 81836
rect 9483 81787 9525 81796
rect 9388 79568 9428 79577
rect 9291 77972 9333 77981
rect 9291 77932 9292 77972
rect 9332 77932 9333 77972
rect 9291 77923 9333 77932
rect 9388 77552 9428 79528
rect 9484 78233 9524 81787
rect 10156 79829 10196 85828
rect 10252 84449 10292 85936
rect 10444 84449 10484 85936
rect 10636 85289 10676 85936
rect 10635 85280 10677 85289
rect 10635 85240 10636 85280
rect 10676 85240 10677 85280
rect 10635 85231 10677 85240
rect 10251 84440 10293 84449
rect 10251 84400 10252 84440
rect 10292 84400 10293 84440
rect 10251 84391 10293 84400
rect 10443 84440 10485 84449
rect 10443 84400 10444 84440
rect 10484 84400 10485 84440
rect 10443 84391 10485 84400
rect 10443 84104 10485 84113
rect 10443 84064 10444 84104
rect 10484 84064 10485 84104
rect 10443 84055 10485 84064
rect 10444 83768 10484 84055
rect 10444 83719 10484 83728
rect 10252 83516 10292 83525
rect 10252 83189 10292 83476
rect 10635 83516 10677 83525
rect 10635 83476 10636 83516
rect 10676 83476 10677 83516
rect 10635 83467 10677 83476
rect 10636 83382 10676 83467
rect 10251 83180 10293 83189
rect 10251 83140 10252 83180
rect 10292 83140 10293 83180
rect 10251 83131 10293 83140
rect 10828 80417 10868 85936
rect 10827 80408 10869 80417
rect 10827 80368 10828 80408
rect 10868 80368 10869 80408
rect 10827 80359 10869 80368
rect 10155 79820 10197 79829
rect 10155 79780 10156 79820
rect 10196 79780 10197 79820
rect 10155 79771 10197 79780
rect 9675 79400 9717 79409
rect 9675 79360 9676 79400
rect 9716 79360 9717 79400
rect 9675 79351 9717 79360
rect 9483 78224 9525 78233
rect 9483 78184 9484 78224
rect 9524 78184 9620 78224
rect 9483 78175 9525 78184
rect 9484 78090 9524 78175
rect 9340 77542 9428 77552
rect 9380 77512 9428 77542
rect 9484 77636 9524 77645
rect 9340 77493 9380 77502
rect 9484 76889 9524 77596
rect 9483 76880 9525 76889
rect 9483 76840 9484 76880
rect 9524 76840 9525 76880
rect 9483 76831 9525 76840
rect 9484 76712 9524 76721
rect 9580 76712 9620 78184
rect 9196 76672 9484 76712
rect 9524 76672 9620 76712
rect 9196 76040 9236 76672
rect 9484 76663 9524 76672
rect 9676 76544 9716 79351
rect 10155 79064 10197 79073
rect 10155 79024 10156 79064
rect 10196 79024 10197 79064
rect 10155 79015 10197 79024
rect 10539 79064 10581 79073
rect 10539 79024 10540 79064
rect 10580 79024 10581 79064
rect 10539 79015 10581 79024
rect 10156 78930 10196 79015
rect 9963 78812 10005 78821
rect 9963 78772 9964 78812
rect 10004 78772 10005 78812
rect 9963 78763 10005 78772
rect 10347 78812 10389 78821
rect 10347 78772 10348 78812
rect 10388 78772 10389 78812
rect 10347 78763 10389 78772
rect 9964 78238 10004 78763
rect 10348 78678 10388 78763
rect 9964 78189 10004 78198
rect 10156 78140 10196 78149
rect 10156 76796 10196 78100
rect 10156 76756 10484 76796
rect 10012 76721 10052 76730
rect 10052 76681 10292 76712
rect 10012 76672 10292 76681
rect 9867 76628 9909 76637
rect 9867 76588 9868 76628
rect 9908 76588 9909 76628
rect 10252 76628 10292 76672
rect 10348 76628 10388 76637
rect 10252 76588 10348 76628
rect 9867 76579 9909 76588
rect 10348 76579 10388 76588
rect 9099 75704 9141 75713
rect 9099 75664 9100 75704
rect 9140 75664 9141 75704
rect 9099 75655 9141 75664
rect 9196 75629 9236 76000
rect 9484 76504 9716 76544
rect 9195 75620 9237 75629
rect 9195 75580 9196 75620
rect 9236 75580 9237 75620
rect 9195 75571 9237 75580
rect 9099 75536 9141 75545
rect 9099 75496 9100 75536
rect 9140 75496 9141 75536
rect 9099 75487 9141 75496
rect 9100 75200 9140 75487
rect 9100 75125 9140 75160
rect 9099 75116 9141 75125
rect 9099 75076 9100 75116
rect 9140 75076 9141 75116
rect 9099 75067 9141 75076
rect 8908 74738 8948 74747
rect 8908 74696 8948 74698
rect 8908 74656 9332 74696
rect 8812 74572 8948 74612
rect 8619 74563 8661 74572
rect 8620 74528 8660 74563
rect 8620 74477 8660 74488
rect 8716 74528 8756 74537
rect 8908 74528 8948 74572
rect 9100 74528 9140 74537
rect 8756 74488 8852 74528
rect 8908 74488 9044 74528
rect 8716 74479 8756 74488
rect 8715 74360 8757 74369
rect 8715 74320 8716 74360
rect 8756 74320 8757 74360
rect 8715 74311 8757 74320
rect 8523 73772 8565 73781
rect 8523 73732 8524 73772
rect 8564 73732 8565 73772
rect 8523 73723 8565 73732
rect 8276 73648 8468 73688
rect 8236 73639 8276 73648
rect 8236 73100 8276 73109
rect 8524 73100 8564 73723
rect 8716 73109 8756 74311
rect 8812 74285 8852 74488
rect 8907 74360 8949 74369
rect 8907 74320 8908 74360
rect 8948 74320 8949 74360
rect 8907 74311 8949 74320
rect 8811 74276 8853 74285
rect 8811 74236 8812 74276
rect 8852 74236 8853 74276
rect 8811 74227 8853 74236
rect 8276 73060 8564 73100
rect 8236 73051 8276 73060
rect 8524 73016 8564 73060
rect 8715 73100 8757 73109
rect 8715 73060 8716 73100
rect 8756 73060 8757 73100
rect 8715 73051 8757 73060
rect 8524 72967 8564 72976
rect 8620 73016 8660 73025
rect 8331 72344 8373 72353
rect 8620 72344 8660 72976
rect 8716 72521 8756 73051
rect 8811 72932 8853 72941
rect 8811 72892 8812 72932
rect 8852 72892 8853 72932
rect 8811 72883 8853 72892
rect 8715 72512 8757 72521
rect 8715 72472 8716 72512
rect 8756 72472 8757 72512
rect 8715 72463 8757 72472
rect 8812 72344 8852 72883
rect 8331 72304 8332 72344
rect 8372 72304 8373 72344
rect 8331 72295 8373 72304
rect 8524 72304 8660 72344
rect 8716 72304 8852 72344
rect 8236 72176 8276 72185
rect 7948 72136 8236 72176
rect 7948 71513 7988 72136
rect 8236 72127 8276 72136
rect 8043 72008 8085 72017
rect 8043 71968 8044 72008
rect 8084 71968 8085 72008
rect 8043 71959 8085 71968
rect 7947 71504 7989 71513
rect 7947 71464 7948 71504
rect 7988 71464 7989 71504
rect 7947 71455 7989 71464
rect 7659 70160 7701 70169
rect 7659 70120 7660 70160
rect 7700 70120 7701 70160
rect 7659 70111 7701 70120
rect 7851 70160 7893 70169
rect 7851 70120 7852 70160
rect 7892 70120 7893 70160
rect 7851 70111 7893 70120
rect 7660 66137 7700 70111
rect 7755 69236 7797 69245
rect 7755 69196 7756 69236
rect 7796 69196 7797 69236
rect 7755 69187 7797 69196
rect 7659 66128 7701 66137
rect 7659 66088 7660 66128
rect 7700 66088 7701 66128
rect 7659 66079 7701 66088
rect 7660 65994 7700 66079
rect 7659 65792 7701 65801
rect 7659 65752 7660 65792
rect 7700 65752 7701 65792
rect 7659 65743 7701 65752
rect 7563 65456 7605 65465
rect 7563 65416 7564 65456
rect 7604 65416 7605 65456
rect 7563 65407 7605 65416
rect 7660 65456 7700 65743
rect 7660 65407 7700 65416
rect 7564 65322 7604 65407
rect 7756 65213 7796 69187
rect 7851 68312 7893 68321
rect 7851 68272 7852 68312
rect 7892 68272 7893 68312
rect 7851 68263 7893 68272
rect 7852 67640 7892 68263
rect 7852 67591 7892 67600
rect 7948 67472 7988 71455
rect 8044 70664 8084 71959
rect 8139 71840 8181 71849
rect 8139 71800 8140 71840
rect 8180 71800 8181 71840
rect 8139 71791 8181 71800
rect 8044 70615 8084 70624
rect 8140 70664 8180 71791
rect 8140 70615 8180 70624
rect 8235 70160 8277 70169
rect 8235 70120 8236 70160
rect 8276 70120 8277 70160
rect 8235 70111 8277 70120
rect 8236 69992 8276 70111
rect 8236 69943 8276 69952
rect 8235 69824 8277 69833
rect 8235 69784 8236 69824
rect 8276 69784 8277 69824
rect 8235 69775 8277 69784
rect 8043 69740 8085 69749
rect 8043 69700 8044 69740
rect 8084 69700 8085 69740
rect 8043 69691 8085 69700
rect 7852 67432 7988 67472
rect 7755 65204 7797 65213
rect 7755 65164 7756 65204
rect 7796 65164 7797 65204
rect 7755 65155 7797 65164
rect 7852 64280 7892 67432
rect 8044 67145 8084 69691
rect 8236 69152 8276 69775
rect 8140 69112 8236 69152
rect 8140 68741 8180 69112
rect 8236 69103 8276 69112
rect 8332 68984 8372 72295
rect 8427 72008 8469 72017
rect 8427 71968 8428 72008
rect 8468 71968 8469 72008
rect 8427 71959 8469 71968
rect 8428 71874 8468 71959
rect 8524 71849 8564 72304
rect 8620 72176 8660 72185
rect 8620 72017 8660 72136
rect 8619 72008 8661 72017
rect 8619 71968 8620 72008
rect 8660 71968 8661 72008
rect 8619 71959 8661 71968
rect 8523 71840 8565 71849
rect 8523 71800 8524 71840
rect 8564 71800 8565 71840
rect 8523 71791 8565 71800
rect 8524 70664 8564 70673
rect 8524 69581 8564 70624
rect 8619 70664 8661 70673
rect 8716 70664 8756 72304
rect 8811 72176 8853 72185
rect 8811 72136 8812 72176
rect 8852 72136 8853 72176
rect 8811 72127 8853 72136
rect 8908 72176 8948 74311
rect 9004 73100 9044 74488
rect 9100 74369 9140 74488
rect 9196 74528 9236 74537
rect 9099 74360 9141 74369
rect 9099 74320 9100 74360
rect 9140 74320 9141 74360
rect 9099 74311 9141 74320
rect 9196 74285 9236 74488
rect 9292 74528 9332 74656
rect 9292 74479 9332 74488
rect 9388 74528 9428 74537
rect 9291 74360 9333 74369
rect 9291 74320 9292 74360
rect 9332 74320 9333 74360
rect 9291 74311 9333 74320
rect 9195 74276 9237 74285
rect 9195 74236 9196 74276
rect 9236 74236 9237 74276
rect 9195 74227 9237 74236
rect 9004 73060 9140 73100
rect 9100 72941 9140 73060
rect 9292 73016 9332 74311
rect 9388 73697 9428 74488
rect 9484 73865 9524 76504
rect 9868 76208 9908 76579
rect 10156 76544 10196 76553
rect 9868 76159 9908 76168
rect 10060 76504 10156 76544
rect 9675 76124 9717 76133
rect 9675 76084 9676 76124
rect 9716 76084 9717 76124
rect 9675 76075 9717 76084
rect 9676 76035 9716 76075
rect 9676 75986 9716 75995
rect 9580 74696 9620 74705
rect 10060 74696 10100 76504
rect 10156 76495 10196 76504
rect 10444 76460 10484 76756
rect 10540 76712 10580 79015
rect 11020 78485 11060 85936
rect 11212 81920 11252 85936
rect 11307 83768 11349 83777
rect 11307 83728 11308 83768
rect 11348 83728 11349 83768
rect 11307 83719 11349 83728
rect 11308 83634 11348 83719
rect 11116 81880 11252 81920
rect 11019 78476 11061 78485
rect 11019 78436 11020 78476
rect 11060 78436 11061 78476
rect 11019 78427 11061 78436
rect 10540 76663 10580 76672
rect 10252 76420 10484 76460
rect 10155 74864 10197 74873
rect 10252 74864 10292 76420
rect 10444 76208 10484 76217
rect 10484 76168 10964 76208
rect 10444 76159 10484 76168
rect 10348 76040 10388 76049
rect 10540 76040 10580 76049
rect 10388 76000 10484 76040
rect 10348 75991 10388 76000
rect 10347 75872 10389 75881
rect 10347 75832 10348 75872
rect 10388 75832 10389 75872
rect 10347 75823 10389 75832
rect 10155 74824 10156 74864
rect 10196 74824 10292 74864
rect 10348 75200 10388 75823
rect 10155 74815 10197 74824
rect 9483 73856 9525 73865
rect 9483 73816 9484 73856
rect 9524 73816 9525 73856
rect 9483 73807 9525 73816
rect 9580 73781 9620 74656
rect 9964 74656 10100 74696
rect 9867 74612 9909 74621
rect 9867 74572 9868 74612
rect 9908 74572 9909 74612
rect 9867 74563 9909 74572
rect 9675 74528 9717 74537
rect 9675 74488 9676 74528
rect 9716 74488 9717 74528
rect 9675 74479 9717 74488
rect 9676 74394 9716 74479
rect 9868 74478 9908 74563
rect 9964 74369 10004 74656
rect 10060 74528 10100 74537
rect 9963 74360 10005 74369
rect 9963 74320 9964 74360
rect 10004 74320 10005 74360
rect 9963 74311 10005 74320
rect 10060 74285 10100 74488
rect 10156 74528 10196 74815
rect 10348 74705 10388 75160
rect 10347 74696 10389 74705
rect 10347 74656 10348 74696
rect 10388 74656 10389 74696
rect 10347 74647 10389 74656
rect 10251 74612 10293 74621
rect 10251 74572 10252 74612
rect 10292 74572 10293 74612
rect 10444 74612 10484 76000
rect 10580 76000 10772 76040
rect 10540 75991 10580 76000
rect 10539 75116 10581 75125
rect 10539 75076 10540 75116
rect 10580 75076 10581 75116
rect 10539 75067 10581 75076
rect 10540 74982 10580 75067
rect 10444 74572 10676 74612
rect 10251 74563 10293 74572
rect 10156 74479 10196 74488
rect 10252 74528 10292 74563
rect 10252 74477 10292 74488
rect 10348 74528 10388 74537
rect 10388 74488 10484 74528
rect 10348 74479 10388 74488
rect 10059 74276 10101 74285
rect 10059 74236 10060 74276
rect 10100 74236 10101 74276
rect 10059 74227 10101 74236
rect 10060 74024 10100 74227
rect 9964 73984 10100 74024
rect 9579 73772 9621 73781
rect 9579 73732 9580 73772
rect 9620 73732 9621 73772
rect 9579 73723 9621 73732
rect 9387 73688 9429 73697
rect 9387 73648 9388 73688
rect 9428 73648 9429 73688
rect 9387 73639 9429 73648
rect 9484 73688 9524 73697
rect 9484 73361 9524 73648
rect 9675 73520 9717 73529
rect 9675 73480 9676 73520
rect 9716 73480 9717 73520
rect 9964 73520 10004 73984
rect 10251 73940 10293 73949
rect 10251 73900 10252 73940
rect 10292 73900 10293 73940
rect 10251 73891 10293 73900
rect 10059 73772 10101 73781
rect 10059 73732 10060 73772
rect 10100 73732 10101 73772
rect 10059 73723 10101 73732
rect 10060 73688 10100 73723
rect 10060 73637 10100 73648
rect 10155 73688 10197 73697
rect 10155 73648 10156 73688
rect 10196 73648 10197 73688
rect 10155 73639 10197 73648
rect 10252 73688 10292 73891
rect 10252 73639 10292 73648
rect 10347 73688 10389 73697
rect 10347 73648 10348 73688
rect 10388 73648 10389 73688
rect 10347 73639 10389 73648
rect 10156 73554 10196 73639
rect 10348 73554 10388 73639
rect 10059 73520 10101 73529
rect 9964 73480 10060 73520
rect 10100 73480 10101 73520
rect 9675 73471 9717 73480
rect 10059 73471 10101 73480
rect 9676 73386 9716 73471
rect 9483 73352 9525 73361
rect 9483 73312 9484 73352
rect 9524 73312 9525 73352
rect 9483 73303 9525 73312
rect 9580 73016 9620 73025
rect 9292 72976 9580 73016
rect 9004 72932 9044 72941
rect 9004 72764 9044 72892
rect 9099 72932 9141 72941
rect 9099 72892 9100 72932
rect 9140 72892 9141 72932
rect 9099 72883 9141 72892
rect 9195 72848 9237 72857
rect 9195 72808 9196 72848
rect 9236 72808 9237 72848
rect 9195 72799 9237 72808
rect 9004 72724 9140 72764
rect 9003 72344 9045 72353
rect 9003 72304 9004 72344
rect 9044 72304 9045 72344
rect 9003 72295 9045 72304
rect 8908 72127 8948 72136
rect 8812 72042 8852 72127
rect 9004 71672 9044 72295
rect 8619 70624 8620 70664
rect 8660 70624 8756 70664
rect 8908 71632 9044 71672
rect 9100 72176 9140 72724
rect 9196 72353 9236 72799
rect 9292 72605 9332 72976
rect 9580 72967 9620 72976
rect 10060 73011 10100 73471
rect 10252 73193 10292 73195
rect 10251 73184 10293 73193
rect 10251 73144 10252 73184
rect 10292 73144 10293 73184
rect 10251 73135 10293 73144
rect 10252 73100 10292 73135
rect 10252 73051 10292 73060
rect 10060 72962 10100 72971
rect 10444 73016 10484 74488
rect 10539 73688 10581 73697
rect 10539 73648 10540 73688
rect 10580 73648 10581 73688
rect 10636 73688 10676 74572
rect 10732 74528 10772 76000
rect 10828 75872 10868 75881
rect 10828 75629 10868 75832
rect 10827 75620 10869 75629
rect 10827 75580 10828 75620
rect 10868 75580 10869 75620
rect 10827 75571 10869 75580
rect 10924 75368 10964 76168
rect 11019 76124 11061 76133
rect 11019 76084 11020 76124
rect 11060 76084 11061 76124
rect 11019 76075 11061 76084
rect 11020 75990 11060 76075
rect 10924 75328 11060 75368
rect 10828 75200 10868 75211
rect 10828 75125 10868 75160
rect 10923 75200 10965 75209
rect 10923 75160 10924 75200
rect 10964 75160 10965 75200
rect 10923 75151 10965 75160
rect 10827 75116 10869 75125
rect 10827 75076 10828 75116
rect 10868 75076 10869 75116
rect 10827 75067 10869 75076
rect 10924 75066 10964 75151
rect 10732 74488 10868 74528
rect 10731 74360 10773 74369
rect 10731 74320 10732 74360
rect 10772 74320 10773 74360
rect 10731 74311 10773 74320
rect 10732 74226 10772 74311
rect 10828 73949 10868 74488
rect 10827 73940 10869 73949
rect 10827 73900 10828 73940
rect 10868 73900 10869 73940
rect 10827 73891 10869 73900
rect 10828 73806 10868 73891
rect 11020 73856 11060 75328
rect 10924 73816 11060 73856
rect 10924 73688 10964 73816
rect 10636 73648 10772 73688
rect 10539 73639 10581 73648
rect 10540 73554 10580 73639
rect 10636 73520 10676 73529
rect 10636 73100 10676 73480
rect 10732 73193 10772 73648
rect 10828 73648 10964 73688
rect 11020 73688 11060 73697
rect 10731 73184 10773 73193
rect 10731 73144 10732 73184
rect 10772 73144 10773 73184
rect 10731 73135 10773 73144
rect 10444 72967 10484 72976
rect 10540 73060 10676 73100
rect 10540 73016 10580 73060
rect 10540 72967 10580 72976
rect 10732 73016 10772 73025
rect 10828 73016 10868 73648
rect 11020 73361 11060 73648
rect 11019 73352 11061 73361
rect 11019 73312 11020 73352
rect 11060 73312 11061 73352
rect 11019 73303 11061 73312
rect 11116 73100 11156 81880
rect 11307 78560 11349 78569
rect 11307 78520 11308 78560
rect 11348 78520 11349 78560
rect 11307 78511 11349 78520
rect 11211 76796 11253 76805
rect 11211 76756 11212 76796
rect 11252 76756 11253 76796
rect 11211 76747 11253 76756
rect 11212 76049 11252 76747
rect 11211 76040 11253 76049
rect 11211 76000 11212 76040
rect 11252 76000 11253 76040
rect 11211 75991 11253 76000
rect 11308 75872 11348 78511
rect 11404 76805 11444 85936
rect 11499 83516 11541 83525
rect 11499 83476 11500 83516
rect 11540 83476 11541 83516
rect 11499 83467 11541 83476
rect 11500 83382 11540 83467
rect 11596 82517 11636 85936
rect 11788 84449 11828 85936
rect 11787 84440 11829 84449
rect 11787 84400 11788 84440
rect 11828 84400 11829 84440
rect 11787 84391 11829 84400
rect 11595 82508 11637 82517
rect 11595 82468 11596 82508
rect 11636 82468 11637 82508
rect 11595 82459 11637 82468
rect 11980 81920 12020 85936
rect 12075 85280 12117 85289
rect 12075 85240 12076 85280
rect 12116 85240 12117 85280
rect 12075 85231 12117 85240
rect 11884 81880 12020 81920
rect 11595 80660 11637 80669
rect 11595 80620 11596 80660
rect 11636 80620 11637 80660
rect 11595 80611 11637 80620
rect 11403 76796 11445 76805
rect 11403 76756 11404 76796
rect 11444 76756 11445 76796
rect 11403 76747 11445 76756
rect 10772 72976 10868 73016
rect 10924 73058 10964 73067
rect 10732 72967 10772 72976
rect 10924 72932 10964 73018
rect 10828 72892 10964 72932
rect 11020 73060 11156 73100
rect 11212 75832 11348 75872
rect 10731 72764 10773 72773
rect 10731 72724 10732 72764
rect 10772 72724 10773 72764
rect 10731 72715 10773 72724
rect 10732 72630 10772 72715
rect 10828 72689 10868 72892
rect 10923 72764 10965 72773
rect 10923 72724 10924 72764
rect 10964 72724 10965 72764
rect 10923 72715 10965 72724
rect 10827 72680 10869 72689
rect 10827 72640 10828 72680
rect 10868 72640 10869 72680
rect 10827 72631 10869 72640
rect 9291 72596 9333 72605
rect 9291 72556 9292 72596
rect 9332 72556 9333 72596
rect 9291 72547 9333 72556
rect 9195 72344 9237 72353
rect 9195 72304 9196 72344
rect 9236 72304 9237 72344
rect 9195 72295 9237 72304
rect 9387 72344 9429 72353
rect 9387 72304 9388 72344
rect 9428 72304 9429 72344
rect 9387 72295 9429 72304
rect 9867 72344 9909 72353
rect 9867 72304 9868 72344
rect 9908 72304 9909 72344
rect 9867 72295 9909 72304
rect 8619 70615 8661 70624
rect 8620 70530 8660 70615
rect 8523 69572 8565 69581
rect 8523 69532 8524 69572
rect 8564 69532 8565 69572
rect 8523 69523 8565 69532
rect 8236 68944 8372 68984
rect 8139 68732 8181 68741
rect 8139 68692 8140 68732
rect 8180 68692 8181 68732
rect 8139 68683 8181 68692
rect 8140 68573 8180 68604
rect 8139 68564 8181 68573
rect 8139 68524 8140 68564
rect 8180 68524 8181 68564
rect 8139 68515 8181 68524
rect 8140 68480 8180 68515
rect 8043 67136 8085 67145
rect 8043 67096 8044 67136
rect 8084 67096 8085 67136
rect 8043 67087 8085 67096
rect 8044 66968 8084 66979
rect 8044 66893 8084 66928
rect 8043 66884 8085 66893
rect 8043 66844 8044 66884
rect 8084 66844 8085 66884
rect 8043 66835 8085 66844
rect 8140 66632 8180 68440
rect 8236 68396 8276 68944
rect 8332 68564 8372 68573
rect 8332 68480 8372 68524
rect 8620 68480 8660 68489
rect 8332 68440 8620 68480
rect 8620 68431 8660 68440
rect 8716 68480 8756 68489
rect 8236 68356 8372 68396
rect 8236 66800 8276 66809
rect 8236 66641 8276 66760
rect 8332 66725 8372 68356
rect 8716 68069 8756 68440
rect 8715 68060 8757 68069
rect 8715 68020 8716 68060
rect 8756 68020 8757 68060
rect 8715 68011 8757 68020
rect 8908 67481 8948 71632
rect 9003 71504 9045 71513
rect 9003 71464 9004 71504
rect 9044 71464 9045 71504
rect 9003 71455 9045 71464
rect 9004 71370 9044 71455
rect 9100 71009 9140 72136
rect 9196 72176 9236 72185
rect 9196 72017 9236 72136
rect 9292 72176 9332 72187
rect 9292 72101 9332 72136
rect 9388 72176 9428 72295
rect 9483 72260 9525 72269
rect 9483 72220 9484 72260
rect 9524 72220 9525 72260
rect 9483 72211 9525 72220
rect 9388 72127 9428 72136
rect 9291 72092 9333 72101
rect 9291 72052 9292 72092
rect 9332 72052 9333 72092
rect 9291 72043 9333 72052
rect 9195 72008 9237 72017
rect 9195 71968 9196 72008
rect 9236 71968 9237 72008
rect 9195 71959 9237 71968
rect 9195 71840 9237 71849
rect 9195 71800 9196 71840
rect 9236 71800 9237 71840
rect 9195 71791 9237 71800
rect 9196 71672 9236 71791
rect 9196 71623 9236 71632
rect 9292 71336 9332 72043
rect 9388 71336 9428 71345
rect 9292 71296 9388 71336
rect 9388 71287 9428 71296
rect 9099 71000 9141 71009
rect 9099 70960 9100 71000
rect 9140 70960 9141 71000
rect 9099 70951 9141 70960
rect 9087 70678 9127 70686
rect 9004 70677 9127 70678
rect 9004 70673 9087 70677
rect 9003 70664 9087 70673
rect 9003 70624 9004 70664
rect 9044 70638 9087 70664
rect 9044 70624 9045 70638
rect 9087 70628 9127 70637
rect 9003 70615 9045 70624
rect 8907 67472 8949 67481
rect 8907 67432 8908 67472
rect 8948 67432 8949 67472
rect 8907 67423 8949 67432
rect 8619 67136 8661 67145
rect 8619 67096 8620 67136
rect 8660 67096 8661 67136
rect 8619 67087 8661 67096
rect 8620 66968 8660 67087
rect 8908 67061 8948 67146
rect 8907 67052 8949 67061
rect 8907 67012 8908 67052
rect 8948 67012 8949 67052
rect 8907 67003 8949 67012
rect 8620 66884 8660 66928
rect 8524 66844 8660 66884
rect 8716 66968 8756 66977
rect 8331 66716 8373 66725
rect 8331 66676 8332 66716
rect 8372 66676 8373 66716
rect 8331 66667 8373 66676
rect 7948 66592 8180 66632
rect 8235 66632 8277 66641
rect 8235 66592 8236 66632
rect 8276 66592 8277 66632
rect 7948 65129 7988 66592
rect 8235 66583 8277 66592
rect 8139 66212 8181 66221
rect 8139 66172 8140 66212
rect 8180 66172 8181 66212
rect 8139 66163 8181 66172
rect 8043 65624 8085 65633
rect 8043 65584 8044 65624
rect 8084 65584 8085 65624
rect 8043 65575 8085 65584
rect 8044 65456 8084 65575
rect 8044 65407 8084 65416
rect 8140 65456 8180 66163
rect 8236 65465 8276 66583
rect 7947 65120 7989 65129
rect 7947 65080 7948 65120
rect 7988 65080 7989 65120
rect 7947 65071 7989 65080
rect 7756 64240 7892 64280
rect 7947 64280 7989 64289
rect 7947 64240 7948 64280
rect 7988 64240 7989 64280
rect 7756 64112 7796 64240
rect 7947 64231 7989 64240
rect 7660 64072 7796 64112
rect 7467 63692 7509 63701
rect 7467 63652 7468 63692
rect 7508 63652 7509 63692
rect 7467 63643 7509 63652
rect 7660 63449 7700 64072
rect 7755 63944 7797 63953
rect 7755 63904 7756 63944
rect 7796 63904 7797 63944
rect 7755 63895 7797 63904
rect 7852 63944 7892 63953
rect 7659 63440 7701 63449
rect 7659 63400 7660 63440
rect 7700 63400 7701 63440
rect 7659 63391 7701 63400
rect 7756 63272 7796 63895
rect 7852 63449 7892 63904
rect 7948 63944 7988 64231
rect 8140 64196 8180 65416
rect 8235 65456 8277 65465
rect 8235 65416 8236 65456
rect 8276 65416 8277 65456
rect 8235 65407 8277 65416
rect 7948 63895 7988 63904
rect 8044 64156 8180 64196
rect 8236 64324 8468 64364
rect 8044 63860 8084 64156
rect 8236 64112 8276 64324
rect 8332 64121 8372 64206
rect 8140 64072 8276 64112
rect 8331 64112 8373 64121
rect 8331 64072 8332 64112
rect 8372 64072 8373 64112
rect 8140 64070 8180 64072
rect 8331 64063 8373 64072
rect 8428 64070 8468 64324
rect 8140 64021 8180 64030
rect 8421 64030 8468 64070
rect 8421 63953 8461 64030
rect 8421 63944 8468 63953
rect 8421 63904 8428 63944
rect 8428 63895 8468 63904
rect 8044 63820 8276 63860
rect 7947 63608 7989 63617
rect 7947 63568 7948 63608
rect 7988 63568 7989 63608
rect 7947 63559 7989 63568
rect 7851 63440 7893 63449
rect 7851 63400 7852 63440
rect 7892 63400 7893 63440
rect 7851 63391 7893 63400
rect 7756 63232 7892 63272
rect 7371 63104 7413 63113
rect 7371 63064 7372 63104
rect 7412 63064 7413 63104
rect 7371 63055 7413 63064
rect 7659 63104 7701 63113
rect 7659 63064 7660 63104
rect 7700 63064 7701 63104
rect 7659 63055 7701 63064
rect 7756 63104 7796 63115
rect 7372 63020 7412 63055
rect 7372 62969 7412 62980
rect 7660 62970 7700 63055
rect 7756 63029 7796 63064
rect 7755 63020 7797 63029
rect 7755 62980 7756 63020
rect 7796 62980 7797 63020
rect 7755 62971 7797 62980
rect 7659 62852 7701 62861
rect 7659 62812 7660 62852
rect 7700 62812 7701 62852
rect 7659 62803 7701 62812
rect 7084 62383 7124 62392
rect 7275 62432 7317 62441
rect 7275 62392 7276 62432
rect 7316 62392 7317 62432
rect 7275 62383 7317 62392
rect 7467 62432 7509 62441
rect 7467 62392 7468 62432
rect 7508 62392 7509 62432
rect 7467 62383 7509 62392
rect 7468 62298 7508 62383
rect 7276 62180 7316 62189
rect 7276 61760 7316 62140
rect 7180 61720 7316 61760
rect 6987 61676 7029 61685
rect 6987 61636 6988 61676
rect 7028 61636 7029 61676
rect 6987 61627 7029 61636
rect 7180 61606 7220 61720
rect 7180 61557 7220 61566
rect 7563 61508 7605 61517
rect 7563 61468 7564 61508
rect 7604 61468 7605 61508
rect 7563 61459 7605 61468
rect 7372 61424 7412 61433
rect 7084 61048 7316 61088
rect 6988 60920 7028 60929
rect 6891 60164 6933 60173
rect 6891 60124 6892 60164
rect 6932 60124 6933 60164
rect 6891 60115 6933 60124
rect 6988 60080 7028 60880
rect 7084 60248 7124 61048
rect 7179 60920 7221 60929
rect 7179 60880 7180 60920
rect 7220 60880 7221 60920
rect 7179 60871 7221 60880
rect 7276 60920 7316 61048
rect 7276 60871 7316 60880
rect 7180 60786 7220 60871
rect 7276 60752 7316 60761
rect 7084 60208 7220 60248
rect 6796 59996 6836 60005
rect 6988 59996 7028 60040
rect 7083 60080 7125 60089
rect 7083 60040 7084 60080
rect 7124 60040 7125 60080
rect 7083 60031 7125 60040
rect 6836 59956 7028 59996
rect 6796 59947 6836 59956
rect 6795 59576 6837 59585
rect 6795 59536 6796 59576
rect 6836 59536 6837 59576
rect 6795 59527 6837 59536
rect 6796 59408 6836 59527
rect 6988 59417 7028 59956
rect 7084 59946 7124 60031
rect 6796 59359 6836 59368
rect 6987 59408 7029 59417
rect 6987 59368 6988 59408
rect 7028 59368 7029 59408
rect 6987 59359 7029 59368
rect 7180 59240 7220 60208
rect 7276 60089 7316 60712
rect 7275 60080 7317 60089
rect 7275 60040 7276 60080
rect 7316 60040 7317 60080
rect 7275 60031 7317 60040
rect 7275 59912 7317 59921
rect 7275 59872 7276 59912
rect 7316 59872 7317 59912
rect 7275 59863 7317 59872
rect 7276 59778 7316 59863
rect 7180 59200 7316 59240
rect 7179 58820 7221 58829
rect 7179 58780 7180 58820
rect 7220 58780 7221 58820
rect 7179 58771 7221 58780
rect 6699 58484 6741 58493
rect 6699 58444 6700 58484
rect 6740 58444 6741 58484
rect 6699 58435 6741 58444
rect 7083 58484 7125 58493
rect 7083 58444 7084 58484
rect 7124 58444 7125 58484
rect 7083 58435 7125 58444
rect 6796 58400 6836 58409
rect 6603 57980 6645 57989
rect 6603 57940 6604 57980
rect 6644 57940 6645 57980
rect 6603 57931 6645 57940
rect 6699 57056 6741 57065
rect 6508 57016 6700 57056
rect 6740 57016 6741 57056
rect 6699 57007 6741 57016
rect 6700 56922 6740 57007
rect 6796 56804 6836 58360
rect 6987 57056 7029 57065
rect 6987 57016 6988 57056
rect 7028 57016 7029 57056
rect 6987 57007 7029 57016
rect 6892 56897 6932 56982
rect 6891 56888 6933 56897
rect 6891 56848 6892 56888
rect 6932 56848 6933 56888
rect 6891 56839 6933 56848
rect 6700 56764 6836 56804
rect 6700 55558 6740 56764
rect 6988 56384 7028 57007
rect 6988 56335 7028 56344
rect 6891 55796 6933 55805
rect 6891 55756 6892 55796
rect 6932 55756 6933 55796
rect 6891 55747 6933 55756
rect 6412 55504 6644 55544
rect 6700 55509 6740 55518
rect 6604 55460 6644 55504
rect 6892 55460 6932 55747
rect 7084 55460 7124 58435
rect 7180 57056 7220 58771
rect 7276 57065 7316 59200
rect 7372 58736 7412 61384
rect 7564 61374 7604 61459
rect 7467 61172 7509 61181
rect 7467 61132 7468 61172
rect 7508 61132 7509 61172
rect 7467 61123 7509 61132
rect 7468 60920 7508 61123
rect 7468 60871 7508 60880
rect 7660 60425 7700 62803
rect 7756 61592 7796 61601
rect 7852 61592 7892 63232
rect 7948 61937 7988 63559
rect 8139 63440 8181 63449
rect 8139 63400 8140 63440
rect 8180 63400 8181 63440
rect 8139 63391 8181 63400
rect 8043 63356 8085 63365
rect 8043 63316 8044 63356
rect 8084 63316 8085 63356
rect 8043 63307 8085 63316
rect 8044 63113 8084 63307
rect 8140 63188 8180 63391
rect 8140 63139 8180 63148
rect 8236 63188 8276 63820
rect 8427 63692 8469 63701
rect 8427 63652 8428 63692
rect 8468 63652 8469 63692
rect 8427 63643 8469 63652
rect 8043 63104 8085 63113
rect 8043 63064 8044 63104
rect 8084 63064 8085 63104
rect 8043 63055 8085 63064
rect 8236 62768 8276 63148
rect 8331 63104 8373 63113
rect 8331 63064 8332 63104
rect 8372 63064 8373 63104
rect 8331 63055 8373 63064
rect 8044 62728 8276 62768
rect 7947 61928 7989 61937
rect 7947 61888 7948 61928
rect 7988 61888 7989 61928
rect 7947 61879 7989 61888
rect 7947 61760 7989 61769
rect 7947 61720 7948 61760
rect 7988 61720 7989 61760
rect 7947 61711 7989 61720
rect 7796 61552 7892 61592
rect 7756 61543 7796 61552
rect 7852 61013 7892 61552
rect 7851 61004 7893 61013
rect 7851 60964 7852 61004
rect 7892 60964 7893 61004
rect 7851 60955 7893 60964
rect 7851 60752 7893 60761
rect 7851 60712 7852 60752
rect 7892 60712 7893 60752
rect 7851 60703 7893 60712
rect 7659 60416 7701 60425
rect 7659 60376 7660 60416
rect 7700 60376 7796 60416
rect 7659 60367 7701 60376
rect 7467 60248 7509 60257
rect 7467 60208 7468 60248
rect 7508 60208 7509 60248
rect 7467 60199 7509 60208
rect 7468 60080 7508 60199
rect 7659 60164 7701 60173
rect 7659 60124 7660 60164
rect 7700 60124 7701 60164
rect 7659 60115 7701 60124
rect 7468 60031 7508 60040
rect 7372 58696 7508 58736
rect 7372 58568 7412 58579
rect 7372 58493 7412 58528
rect 7371 58484 7413 58493
rect 7371 58444 7372 58484
rect 7412 58444 7413 58484
rect 7371 58435 7413 58444
rect 7180 57007 7220 57016
rect 7275 57056 7317 57065
rect 7275 57016 7276 57056
rect 7316 57016 7317 57056
rect 7275 57007 7317 57016
rect 7468 56972 7508 58696
rect 7563 57896 7605 57905
rect 7563 57856 7564 57896
rect 7604 57856 7605 57896
rect 7563 57847 7605 57856
rect 7564 57762 7604 57847
rect 7660 57476 7700 60115
rect 7756 59249 7796 60376
rect 7755 59240 7797 59249
rect 7755 59200 7756 59240
rect 7796 59200 7797 59240
rect 7755 59191 7797 59200
rect 7852 57821 7892 60703
rect 7851 57812 7893 57821
rect 7851 57772 7852 57812
rect 7892 57772 7893 57812
rect 7851 57763 7893 57772
rect 7756 57644 7796 57653
rect 7796 57604 7892 57644
rect 7756 57595 7796 57604
rect 7660 57436 7796 57476
rect 7756 57149 7796 57436
rect 7755 57140 7797 57149
rect 7755 57100 7756 57140
rect 7796 57100 7797 57140
rect 7755 57091 7797 57100
rect 7563 57056 7605 57065
rect 7563 57016 7564 57056
rect 7604 57016 7605 57056
rect 7563 57007 7605 57016
rect 7660 57056 7700 57065
rect 7372 56932 7508 56972
rect 7179 56468 7221 56477
rect 7179 56428 7180 56468
rect 7220 56428 7221 56468
rect 7179 56419 7221 56428
rect 7180 56334 7220 56419
rect 7372 55460 7412 56932
rect 7467 56804 7509 56813
rect 7467 56764 7468 56804
rect 7508 56764 7509 56804
rect 7467 56755 7509 56764
rect 7468 56384 7508 56755
rect 7468 56335 7508 56344
rect 7564 56384 7604 57007
rect 7660 56393 7700 57016
rect 7756 57006 7796 57091
rect 6316 55420 6548 55460
rect 6604 55420 6740 55460
rect 6219 55124 6261 55133
rect 6219 55084 6220 55124
rect 6260 55084 6261 55124
rect 6219 55075 6261 55084
rect 6219 54200 6261 54209
rect 6219 54160 6220 54200
rect 6260 54160 6261 54200
rect 6219 54151 6261 54160
rect 6123 51260 6165 51269
rect 6123 51220 6124 51260
rect 6164 51220 6165 51260
rect 6123 51211 6165 51220
rect 5932 51017 5972 51052
rect 5836 51008 5876 51017
rect 5836 50420 5876 50968
rect 5931 51008 5973 51017
rect 6220 51008 6260 54151
rect 6411 53276 6453 53285
rect 6411 53236 6412 53276
rect 6452 53236 6453 53276
rect 6411 53227 6453 53236
rect 6412 52025 6452 53227
rect 6411 52016 6453 52025
rect 6411 51976 6412 52016
rect 6452 51976 6453 52016
rect 6411 51967 6453 51976
rect 6412 51008 6452 51017
rect 5931 50968 5932 51008
rect 5972 50968 5973 51008
rect 5931 50959 5973 50968
rect 6124 50968 6412 51008
rect 5932 50928 5972 50959
rect 5836 50380 5972 50420
rect 5835 50252 5877 50261
rect 5835 50212 5836 50252
rect 5876 50212 5877 50252
rect 5835 50203 5877 50212
rect 5932 50252 5972 50380
rect 5836 50118 5876 50203
rect 5835 49496 5877 49505
rect 5835 49456 5836 49496
rect 5876 49456 5877 49496
rect 5835 49447 5877 49456
rect 5836 49362 5876 49447
rect 5835 49076 5877 49085
rect 5835 49036 5836 49076
rect 5876 49036 5877 49076
rect 5835 49027 5877 49036
rect 5547 48488 5589 48497
rect 5547 48448 5548 48488
rect 5588 48448 5589 48488
rect 5547 48439 5589 48448
rect 5739 48488 5781 48497
rect 5739 48448 5740 48488
rect 5780 48448 5781 48488
rect 5739 48439 5781 48448
rect 5355 48320 5397 48329
rect 5355 48280 5356 48320
rect 5396 48280 5397 48320
rect 5355 48271 5397 48280
rect 5547 48320 5589 48329
rect 5836 48320 5876 49027
rect 5932 48581 5972 50212
rect 6027 50000 6069 50009
rect 6027 49960 6028 50000
rect 6068 49960 6069 50000
rect 6027 49951 6069 49960
rect 5931 48572 5973 48581
rect 5931 48532 5932 48572
rect 5972 48532 5973 48572
rect 5931 48523 5973 48532
rect 5547 48280 5548 48320
rect 5588 48280 5589 48320
rect 5547 48271 5589 48280
rect 5740 48280 5876 48320
rect 5355 48152 5397 48161
rect 5355 48112 5356 48152
rect 5396 48112 5397 48152
rect 5355 48103 5397 48112
rect 5260 47851 5300 47860
rect 5068 47766 5108 47851
rect 4928 47648 5296 47657
rect 4968 47608 5010 47648
rect 5050 47608 5092 47648
rect 5132 47608 5174 47648
rect 5214 47608 5256 47648
rect 4928 47599 5296 47608
rect 4972 47312 5012 47321
rect 4780 47272 4972 47312
rect 4972 47263 5012 47272
rect 5068 47312 5108 47321
rect 5356 47312 5396 48103
rect 5452 47993 5492 47998
rect 5451 47989 5493 47993
rect 5451 47944 5452 47989
rect 5492 47944 5493 47989
rect 5451 47935 5493 47944
rect 5452 47854 5492 47935
rect 5108 47272 5396 47312
rect 5068 47263 5108 47272
rect 4492 46600 4628 46640
rect 4492 46472 4532 46500
rect 4396 46432 4492 46472
rect 4299 44708 4341 44717
rect 4299 44668 4300 44708
rect 4340 44668 4341 44708
rect 4299 44659 4341 44668
rect 4011 44036 4053 44045
rect 4011 43996 4012 44036
rect 4052 43996 4053 44036
rect 4011 43987 4053 43996
rect 4396 43952 4436 46432
rect 4492 46423 4532 46432
rect 4588 44969 4628 46600
rect 4928 46136 5296 46145
rect 4968 46096 5010 46136
rect 5050 46096 5092 46136
rect 5132 46096 5174 46136
rect 5214 46096 5256 46136
rect 4928 46087 5296 46096
rect 5356 45968 5396 47272
rect 5451 47312 5493 47321
rect 5451 47272 5452 47312
rect 5492 47272 5493 47312
rect 5451 47263 5493 47272
rect 5548 47312 5588 48271
rect 5643 47648 5685 47657
rect 5643 47608 5644 47648
rect 5684 47608 5685 47648
rect 5643 47599 5685 47608
rect 5548 47263 5588 47272
rect 5452 47178 5492 47263
rect 5644 46640 5684 47599
rect 5260 45928 5396 45968
rect 5452 46600 5684 46640
rect 4587 44960 4629 44969
rect 4587 44920 4588 44960
rect 4628 44920 4629 44960
rect 4587 44911 4629 44920
rect 5260 44792 5300 45928
rect 5355 45800 5397 45809
rect 5355 45760 5356 45800
rect 5396 45760 5397 45800
rect 5355 45751 5397 45760
rect 5356 45666 5396 45751
rect 5452 45548 5492 46600
rect 5740 46472 5780 48280
rect 5931 48236 5973 48245
rect 5931 48196 5932 48236
rect 5972 48196 5973 48236
rect 5931 48187 5973 48196
rect 5932 47984 5972 48187
rect 5932 47935 5972 47944
rect 6028 47900 6068 49951
rect 6124 48245 6164 50968
rect 6412 50959 6452 50968
rect 6411 50840 6453 50849
rect 6411 50800 6412 50840
rect 6452 50800 6453 50840
rect 6411 50791 6453 50800
rect 6219 50588 6261 50597
rect 6219 50548 6220 50588
rect 6260 50548 6261 50588
rect 6219 50539 6261 50548
rect 6220 50336 6260 50539
rect 6316 50336 6356 50345
rect 6220 50296 6316 50336
rect 6123 48236 6165 48245
rect 6123 48196 6124 48236
rect 6164 48196 6165 48236
rect 6123 48187 6165 48196
rect 6028 47860 6164 47900
rect 6028 47312 6068 47321
rect 4300 43912 4436 43952
rect 4780 44752 5300 44792
rect 5356 45508 5492 45548
rect 5548 45548 5588 45557
rect 3688 43868 4056 43877
rect 3728 43828 3770 43868
rect 3810 43828 3852 43868
rect 3892 43828 3934 43868
rect 3974 43828 4016 43868
rect 3688 43819 4056 43828
rect 3723 43616 3765 43625
rect 3723 43576 3724 43616
rect 3764 43576 3765 43616
rect 3723 43567 3765 43576
rect 3627 43532 3669 43541
rect 3627 43492 3628 43532
rect 3668 43492 3669 43532
rect 3627 43483 3669 43492
rect 3628 43398 3668 43483
rect 3724 43448 3764 43567
rect 4108 43541 4148 43572
rect 4107 43532 4149 43541
rect 4107 43492 4108 43532
rect 4148 43492 4149 43532
rect 4107 43483 4149 43492
rect 3531 42944 3573 42953
rect 3531 42904 3532 42944
rect 3572 42904 3573 42944
rect 3531 42895 3573 42904
rect 3724 42524 3764 43408
rect 3436 41971 3476 41980
rect 3532 42484 3764 42524
rect 4108 43448 4148 43483
rect 2956 41887 2996 41896
rect 3532 41936 3572 42484
rect 3688 42356 4056 42365
rect 3728 42316 3770 42356
rect 3810 42316 3852 42356
rect 3892 42316 3934 42356
rect 3974 42316 4016 42356
rect 3688 42307 4056 42316
rect 3532 41861 3572 41896
rect 3916 41936 3956 41947
rect 3916 41861 3956 41896
rect 4011 41936 4053 41945
rect 4011 41896 4012 41936
rect 4052 41896 4053 41936
rect 4011 41887 4053 41896
rect 3531 41852 3573 41861
rect 3531 41812 3532 41852
rect 3572 41812 3573 41852
rect 3531 41803 3573 41812
rect 3915 41852 3957 41861
rect 3915 41812 3916 41852
rect 3956 41812 3957 41852
rect 3915 41803 3957 41812
rect 4012 41802 4052 41887
rect 4108 41861 4148 43408
rect 4204 43448 4244 43457
rect 4204 42869 4244 43408
rect 4203 42860 4245 42869
rect 4203 42820 4204 42860
rect 4244 42820 4245 42860
rect 4203 42811 4245 42820
rect 4107 41852 4149 41861
rect 4107 41812 4108 41852
rect 4148 41812 4149 41852
rect 4107 41803 4149 41812
rect 3531 41600 3573 41609
rect 3531 41560 3532 41600
rect 3572 41560 3573 41600
rect 3531 41551 3573 41560
rect 3339 41516 3381 41525
rect 3339 41476 3340 41516
rect 3380 41476 3381 41516
rect 3339 41467 3381 41476
rect 3340 41432 3380 41467
rect 3340 41381 3380 41392
rect 3148 41264 3188 41273
rect 2955 41012 2997 41021
rect 2955 40972 2956 41012
rect 2996 40972 2997 41012
rect 2955 40963 2997 40972
rect 2859 40592 2901 40601
rect 2859 40552 2860 40592
rect 2900 40552 2901 40592
rect 2859 40543 2901 40552
rect 2860 40097 2900 40543
rect 2859 40088 2901 40097
rect 2859 40048 2860 40088
rect 2900 40048 2901 40088
rect 2859 40039 2901 40048
rect 2763 39584 2805 39593
rect 2763 39544 2764 39584
rect 2804 39544 2805 39584
rect 2763 39535 2805 39544
rect 2668 39376 2804 39416
rect 2667 39080 2709 39089
rect 2667 39040 2668 39080
rect 2708 39040 2709 39080
rect 2667 39031 2709 39040
rect 2571 37904 2613 37913
rect 2571 37864 2572 37904
rect 2612 37864 2613 37904
rect 2571 37855 2613 37864
rect 2380 37400 2420 37409
rect 2283 36644 2325 36653
rect 2283 36604 2284 36644
rect 2324 36604 2325 36644
rect 2283 36595 2325 36604
rect 2380 36233 2420 37360
rect 2476 37400 2516 37409
rect 2476 36989 2516 37360
rect 2571 37400 2613 37409
rect 2571 37360 2572 37400
rect 2612 37360 2613 37400
rect 2571 37351 2613 37360
rect 2475 36980 2517 36989
rect 2475 36940 2476 36980
rect 2516 36940 2517 36980
rect 2475 36931 2517 36940
rect 2476 36728 2516 36768
rect 2476 36653 2516 36688
rect 2475 36644 2517 36653
rect 2475 36604 2476 36644
rect 2516 36604 2517 36644
rect 2475 36595 2517 36604
rect 2379 36224 2421 36233
rect 2379 36184 2380 36224
rect 2420 36184 2421 36224
rect 2379 36175 2421 36184
rect 2187 36140 2229 36149
rect 2187 36100 2188 36140
rect 2228 36100 2229 36140
rect 2187 36091 2229 36100
rect 1899 35888 1941 35897
rect 1899 35848 1900 35888
rect 1940 35848 1941 35888
rect 1899 35839 1941 35848
rect 2476 35888 2516 36595
rect 1900 30857 1940 35839
rect 1995 35048 2037 35057
rect 1995 35008 1996 35048
rect 2036 35008 2037 35048
rect 1995 34999 2037 35008
rect 1996 34469 2036 34999
rect 2379 34880 2421 34889
rect 2379 34840 2380 34880
rect 2420 34840 2421 34880
rect 2379 34831 2421 34840
rect 2092 34504 2324 34544
rect 1995 34460 2037 34469
rect 1995 34420 1996 34460
rect 2036 34420 2037 34460
rect 1995 34411 2037 34420
rect 1996 32696 2036 34411
rect 2092 32873 2132 34504
rect 2187 34376 2229 34385
rect 2187 34336 2188 34376
rect 2228 34336 2229 34376
rect 2187 34327 2229 34336
rect 2284 34376 2324 34504
rect 2284 34327 2324 34336
rect 2188 34242 2228 34327
rect 2380 34208 2420 34831
rect 2284 34168 2420 34208
rect 2187 33620 2229 33629
rect 2187 33580 2188 33620
rect 2228 33580 2229 33620
rect 2187 33571 2229 33580
rect 2188 33125 2228 33571
rect 2187 33116 2229 33125
rect 2187 33076 2188 33116
rect 2228 33076 2229 33116
rect 2187 33067 2229 33076
rect 2091 32864 2133 32873
rect 2091 32824 2092 32864
rect 2132 32824 2133 32864
rect 2091 32815 2133 32824
rect 1996 32656 2132 32696
rect 1995 31352 2037 31361
rect 1995 31312 1996 31352
rect 2036 31312 2037 31352
rect 1995 31303 2037 31312
rect 1899 30848 1941 30857
rect 1899 30808 1900 30848
rect 1940 30808 1941 30848
rect 1899 30799 1941 30808
rect 1996 30848 2036 31303
rect 2092 30857 2132 32656
rect 1996 30799 2036 30808
rect 2091 30848 2133 30857
rect 2091 30808 2092 30848
rect 2132 30808 2133 30848
rect 2188 30848 2228 33067
rect 2284 32705 2324 34168
rect 2476 33713 2516 35848
rect 2572 35813 2612 37351
rect 2668 36896 2708 39031
rect 2668 36847 2708 36856
rect 2667 36224 2709 36233
rect 2667 36184 2668 36224
rect 2708 36184 2709 36224
rect 2667 36175 2709 36184
rect 2668 36140 2708 36175
rect 2668 36089 2708 36100
rect 2667 35888 2709 35897
rect 2667 35848 2668 35888
rect 2708 35848 2709 35888
rect 2667 35839 2709 35848
rect 2571 35804 2613 35813
rect 2571 35764 2572 35804
rect 2612 35764 2613 35804
rect 2571 35755 2613 35764
rect 2572 33797 2612 35755
rect 2668 35216 2708 35839
rect 2668 35167 2708 35176
rect 2667 34544 2709 34553
rect 2667 34504 2668 34544
rect 2708 34504 2709 34544
rect 2764 34544 2804 39376
rect 2860 38408 2900 40039
rect 2956 39761 2996 40963
rect 3148 40349 3188 41224
rect 3532 40676 3572 41551
rect 4300 41273 4340 43912
rect 4780 43541 4820 44752
rect 4928 44624 5296 44633
rect 4968 44584 5010 44624
rect 5050 44584 5092 44624
rect 5132 44584 5174 44624
rect 5214 44584 5256 44624
rect 4928 44575 5296 44584
rect 5068 44288 5108 44299
rect 5068 44213 5108 44248
rect 5067 44204 5109 44213
rect 5067 44164 5068 44204
rect 5108 44164 5109 44204
rect 5067 44155 5109 44164
rect 5259 44120 5301 44129
rect 5259 44080 5260 44120
rect 5300 44080 5301 44120
rect 5259 44071 5301 44080
rect 5260 43986 5300 44071
rect 4779 43532 4821 43541
rect 4779 43492 4780 43532
rect 4820 43492 4821 43532
rect 4779 43483 4821 43492
rect 4928 43112 5296 43121
rect 4968 43072 5010 43112
rect 5050 43072 5092 43112
rect 5132 43072 5174 43112
rect 5214 43072 5256 43112
rect 4928 43063 5296 43072
rect 4684 42860 4724 42869
rect 4724 42820 5012 42860
rect 4684 42811 4724 42820
rect 4492 42776 4532 42785
rect 4492 41273 4532 42736
rect 4972 42776 5012 42820
rect 4972 42727 5012 42736
rect 5067 42776 5109 42785
rect 5067 42736 5068 42776
rect 5108 42736 5109 42776
rect 5067 42727 5109 42736
rect 4875 42692 4917 42701
rect 4875 42652 4876 42692
rect 4916 42652 4917 42692
rect 4875 42643 4917 42652
rect 4876 42104 4916 42643
rect 5068 42642 5108 42727
rect 5259 42608 5301 42617
rect 5356 42608 5396 45508
rect 5548 44960 5588 45508
rect 5643 45380 5685 45389
rect 5643 45340 5644 45380
rect 5684 45340 5685 45380
rect 5643 45331 5685 45340
rect 5644 45128 5684 45331
rect 5740 45212 5780 46432
rect 5836 47272 6028 47312
rect 5836 45464 5876 47272
rect 6028 47263 6068 47272
rect 5931 46640 5973 46649
rect 5931 46600 5932 46640
rect 5972 46600 5973 46640
rect 5931 46591 5973 46600
rect 5932 46506 5972 46591
rect 6124 46472 6164 47860
rect 6124 46423 6164 46432
rect 6220 45473 6260 50296
rect 6316 50287 6356 50296
rect 6412 50336 6452 50791
rect 6508 50345 6548 55420
rect 6603 55208 6645 55217
rect 6603 55168 6604 55208
rect 6644 55168 6645 55208
rect 6603 55159 6645 55168
rect 6412 50287 6452 50296
rect 6507 50336 6549 50345
rect 6507 50296 6508 50336
rect 6548 50296 6549 50336
rect 6507 50287 6549 50296
rect 6604 50168 6644 55159
rect 6700 54872 6740 55420
rect 6892 55411 6932 55420
rect 6988 55420 7124 55460
rect 7180 55420 7412 55460
rect 7564 55460 7604 56344
rect 7659 56384 7701 56393
rect 7659 56344 7660 56384
rect 7700 56344 7701 56384
rect 7659 56335 7701 56344
rect 7852 55544 7892 57604
rect 7948 56729 7988 61711
rect 8044 60761 8084 62728
rect 8332 62600 8372 63055
rect 8140 62560 8372 62600
rect 8043 60752 8085 60761
rect 8043 60712 8044 60752
rect 8084 60712 8085 60752
rect 8043 60703 8085 60712
rect 8044 59408 8084 59417
rect 8044 57905 8084 59368
rect 8043 57896 8085 57905
rect 8043 57856 8044 57896
rect 8084 57856 8085 57896
rect 8043 57847 8085 57856
rect 8140 57737 8180 62560
rect 8428 61853 8468 63643
rect 8524 63449 8564 66844
rect 8716 66641 8756 66928
rect 8812 66968 8852 66977
rect 8715 66632 8757 66641
rect 8715 66592 8716 66632
rect 8756 66592 8757 66632
rect 8715 66583 8757 66592
rect 8715 66296 8757 66305
rect 8715 66256 8716 66296
rect 8756 66256 8757 66296
rect 8715 66247 8757 66256
rect 8619 65540 8661 65549
rect 8619 65500 8620 65540
rect 8660 65500 8661 65540
rect 8619 65491 8661 65500
rect 8620 65456 8660 65491
rect 8620 65405 8660 65416
rect 8619 64700 8661 64709
rect 8619 64660 8620 64700
rect 8660 64660 8661 64700
rect 8619 64651 8661 64660
rect 8620 64616 8660 64651
rect 8620 64565 8660 64576
rect 8619 63692 8661 63701
rect 8619 63652 8620 63692
rect 8660 63652 8661 63692
rect 8619 63643 8661 63652
rect 8620 63558 8660 63643
rect 8523 63440 8565 63449
rect 8523 63400 8524 63440
rect 8564 63400 8565 63440
rect 8523 63391 8565 63400
rect 8716 63113 8756 66247
rect 8812 65969 8852 66928
rect 8907 66884 8949 66893
rect 8907 66844 8908 66884
rect 8948 66844 8949 66884
rect 8907 66835 8949 66844
rect 8908 66128 8948 66835
rect 8811 65960 8853 65969
rect 8811 65920 8812 65960
rect 8852 65920 8853 65960
rect 8811 65911 8853 65920
rect 8908 65885 8948 66088
rect 8907 65876 8949 65885
rect 8907 65836 8908 65876
rect 8948 65836 8949 65876
rect 8907 65827 8949 65836
rect 9004 65708 9044 70615
rect 9484 70580 9524 72211
rect 9580 72176 9620 72185
rect 9580 71849 9620 72136
rect 9771 72176 9813 72185
rect 9771 72136 9772 72176
rect 9812 72136 9813 72176
rect 9771 72127 9813 72136
rect 9868 72176 9908 72295
rect 10348 72185 10388 72270
rect 10828 72269 10868 72631
rect 10827 72260 10869 72269
rect 10827 72220 10828 72260
rect 10868 72220 10869 72260
rect 10827 72211 10869 72220
rect 9868 72127 9908 72136
rect 10060 72176 10100 72185
rect 9772 72042 9812 72127
rect 9675 72008 9717 72017
rect 9675 71968 9676 72008
rect 9716 71968 9717 72008
rect 9675 71959 9717 71968
rect 9676 71874 9716 71959
rect 9579 71840 9621 71849
rect 9579 71800 9580 71840
rect 9620 71800 9621 71840
rect 9579 71791 9621 71800
rect 9580 71672 9620 71791
rect 9771 71756 9813 71765
rect 9771 71716 9772 71756
rect 9812 71716 9813 71756
rect 9771 71707 9813 71716
rect 9580 71632 9716 71672
rect 9579 71504 9621 71513
rect 9579 71464 9580 71504
rect 9620 71464 9621 71504
rect 9579 71455 9621 71464
rect 9580 71370 9620 71455
rect 9676 70748 9716 71632
rect 9772 71513 9812 71707
rect 9771 71504 9813 71513
rect 9771 71464 9772 71504
rect 9812 71464 9813 71504
rect 9771 71455 9813 71464
rect 9628 70708 9716 70748
rect 9628 70706 9668 70708
rect 9628 70657 9668 70666
rect 9196 70540 9524 70580
rect 9772 70580 9812 70589
rect 10060 70580 10100 72136
rect 10347 72176 10389 72185
rect 10347 72136 10348 72176
rect 10388 72136 10389 72176
rect 10347 72127 10389 72136
rect 10252 72008 10292 72017
rect 10252 70664 10292 71968
rect 10347 72008 10389 72017
rect 10347 71968 10348 72008
rect 10388 71968 10389 72008
rect 10347 71959 10389 71968
rect 10348 70832 10388 71959
rect 10443 71756 10485 71765
rect 10443 71716 10444 71756
rect 10484 71716 10485 71756
rect 10443 71707 10485 71716
rect 10348 70783 10388 70792
rect 10348 70664 10388 70673
rect 10252 70624 10348 70664
rect 10348 70615 10388 70624
rect 9812 70540 10100 70580
rect 9196 68480 9236 70540
rect 9772 70531 9812 70540
rect 10444 70496 10484 71707
rect 10827 71588 10869 71597
rect 10827 71548 10828 71588
rect 10868 71548 10869 71588
rect 10827 71539 10869 71548
rect 10828 71504 10868 71539
rect 10635 71420 10677 71429
rect 10635 71380 10636 71420
rect 10676 71380 10677 71420
rect 10635 71371 10677 71380
rect 10539 70832 10581 70841
rect 10539 70792 10540 70832
rect 10580 70792 10581 70832
rect 10539 70783 10581 70792
rect 10540 70698 10580 70783
rect 10252 70456 10484 70496
rect 9867 70412 9909 70421
rect 9867 70372 9868 70412
rect 9908 70372 9909 70412
rect 9867 70363 9909 70372
rect 9483 69992 9525 70001
rect 9483 69952 9484 69992
rect 9524 69952 9525 69992
rect 9483 69943 9525 69952
rect 9868 69992 9908 70363
rect 9484 69858 9524 69943
rect 9868 69917 9908 69952
rect 9867 69908 9909 69917
rect 9867 69868 9868 69908
rect 9908 69868 9909 69908
rect 9867 69859 9909 69868
rect 9676 69740 9716 69749
rect 9716 69700 10004 69740
rect 9676 69691 9716 69700
rect 9484 69245 9524 69276
rect 9483 69236 9525 69245
rect 9483 69196 9484 69236
rect 9524 69196 9525 69236
rect 9483 69187 9525 69196
rect 9484 69152 9524 69187
rect 9484 68573 9524 69112
rect 9964 69152 10004 69700
rect 9964 69103 10004 69112
rect 10059 69152 10101 69161
rect 10059 69112 10060 69152
rect 10100 69112 10101 69152
rect 10059 69103 10101 69112
rect 9675 68984 9717 68993
rect 9675 68944 9676 68984
rect 9716 68944 9717 68984
rect 9675 68935 9717 68944
rect 9676 68850 9716 68935
rect 9483 68564 9525 68573
rect 9483 68524 9484 68564
rect 9524 68524 9525 68564
rect 9483 68515 9525 68524
rect 9100 68396 9140 68405
rect 9100 67901 9140 68356
rect 9099 67892 9141 67901
rect 9099 67852 9100 67892
rect 9140 67852 9141 67892
rect 9099 67843 9141 67852
rect 9099 67724 9141 67733
rect 9099 67684 9100 67724
rect 9140 67684 9141 67724
rect 9099 67675 9141 67684
rect 9100 67640 9140 67675
rect 9100 67589 9140 67600
rect 9196 67145 9236 68440
rect 9676 68480 9716 68491
rect 9676 68405 9716 68440
rect 9675 68396 9717 68405
rect 9675 68356 9676 68396
rect 9716 68356 9717 68396
rect 9675 68347 9717 68356
rect 9675 68060 9717 68069
rect 9675 68020 9676 68060
rect 9716 68020 9717 68060
rect 9675 68011 9717 68020
rect 9580 67640 9620 67649
rect 9292 67556 9332 67565
rect 9580 67556 9620 67600
rect 9676 67640 9716 68011
rect 10060 67901 10100 69103
rect 10155 68984 10197 68993
rect 10155 68944 10156 68984
rect 10196 68944 10197 68984
rect 10155 68935 10197 68944
rect 10156 68475 10196 68935
rect 10252 68480 10292 70456
rect 10636 70412 10676 71371
rect 10828 70673 10868 71464
rect 10348 70372 10676 70412
rect 10732 70664 10772 70673
rect 10348 68984 10388 70372
rect 10635 69908 10677 69917
rect 10635 69868 10636 69908
rect 10676 69868 10677 69908
rect 10635 69859 10677 69868
rect 10443 69320 10485 69329
rect 10443 69280 10444 69320
rect 10484 69280 10485 69320
rect 10443 69271 10485 69280
rect 10444 69236 10484 69271
rect 10444 69185 10484 69196
rect 10539 69152 10581 69161
rect 10539 69112 10540 69152
rect 10580 69112 10581 69152
rect 10636 69157 10676 69859
rect 10732 69329 10772 70624
rect 10827 70664 10869 70673
rect 10827 70624 10828 70664
rect 10868 70624 10869 70664
rect 10827 70615 10869 70624
rect 10731 69320 10773 69329
rect 10731 69280 10732 69320
rect 10772 69280 10773 69320
rect 10731 69271 10773 69280
rect 10636 69117 10772 69157
rect 10539 69103 10581 69112
rect 10540 69018 10580 69103
rect 10348 68944 10484 68984
rect 10348 68657 10388 68742
rect 10347 68648 10389 68657
rect 10347 68608 10348 68648
rect 10388 68608 10389 68648
rect 10347 68599 10389 68608
rect 10252 68440 10388 68480
rect 10156 68426 10196 68435
rect 9771 67892 9813 67901
rect 9771 67852 9772 67892
rect 9812 67852 9813 67892
rect 9771 67843 9813 67852
rect 10059 67892 10101 67901
rect 10059 67852 10060 67892
rect 10100 67852 10101 67892
rect 10059 67843 10101 67852
rect 9676 67591 9716 67600
rect 9772 67565 9812 67843
rect 10155 67724 10197 67733
rect 10155 67684 10156 67724
rect 10196 67684 10197 67724
rect 10155 67675 10197 67684
rect 10060 67640 10100 67649
rect 10060 67565 10100 67600
rect 10156 67590 10196 67675
rect 9332 67516 9620 67556
rect 9771 67556 9813 67565
rect 9771 67516 9772 67556
rect 9812 67516 9813 67556
rect 9292 67507 9332 67516
rect 9771 67507 9813 67516
rect 10059 67556 10101 67565
rect 10059 67516 10060 67556
rect 10100 67516 10101 67556
rect 10059 67507 10101 67516
rect 9675 67472 9717 67481
rect 9675 67432 9676 67472
rect 9716 67432 9717 67472
rect 9675 67423 9717 67432
rect 9195 67136 9237 67145
rect 9195 67096 9196 67136
rect 9236 67096 9237 67136
rect 9195 67087 9237 67096
rect 9676 67136 9716 67423
rect 9676 67087 9716 67096
rect 9387 67052 9429 67061
rect 9387 67012 9388 67052
rect 9428 67012 9429 67052
rect 9387 67003 9429 67012
rect 9867 67052 9909 67061
rect 9867 67012 9868 67052
rect 9908 67012 9909 67052
rect 9867 67003 9909 67012
rect 9100 66968 9140 66977
rect 9292 66968 9332 66977
rect 9100 66380 9140 66928
rect 9100 66331 9140 66340
rect 9196 66928 9292 66968
rect 8812 65668 9044 65708
rect 9100 65960 9140 65969
rect 8812 64280 8852 65668
rect 8907 65540 8949 65549
rect 8907 65500 8908 65540
rect 8948 65500 8949 65540
rect 8907 65491 8949 65500
rect 8908 64616 8948 65491
rect 9100 65451 9140 65920
rect 9100 65402 9140 65411
rect 9196 65297 9236 66928
rect 9292 66919 9332 66928
rect 9388 66968 9428 67003
rect 9388 66917 9428 66928
rect 9580 66968 9620 66977
rect 9388 66800 9428 66809
rect 9388 66305 9428 66760
rect 9387 66296 9429 66305
rect 9387 66256 9388 66296
rect 9428 66256 9429 66296
rect 9580 66296 9620 66928
rect 9772 66968 9812 66977
rect 9772 66809 9812 66928
rect 9868 66893 9908 67003
rect 9867 66884 9909 66893
rect 9867 66844 9868 66884
rect 9908 66844 9909 66884
rect 9867 66835 9909 66844
rect 9771 66800 9813 66809
rect 9771 66760 9772 66800
rect 9812 66760 9813 66800
rect 9771 66751 9813 66760
rect 9676 66380 9716 66389
rect 9716 66340 9908 66380
rect 9676 66331 9716 66340
rect 9580 66256 9621 66296
rect 9387 66247 9429 66256
rect 9581 66212 9621 66256
rect 9580 66172 9621 66212
rect 9388 66128 9428 66137
rect 9292 65624 9332 65633
rect 9388 65624 9428 66088
rect 9483 65960 9525 65969
rect 9483 65920 9484 65960
rect 9524 65920 9525 65960
rect 9483 65911 9525 65920
rect 9332 65584 9428 65624
rect 9484 65624 9524 65911
rect 9292 65575 9332 65584
rect 9484 65575 9524 65584
rect 9195 65288 9237 65297
rect 9195 65248 9196 65288
rect 9236 65248 9237 65288
rect 9195 65239 9237 65248
rect 9580 64961 9620 66172
rect 9676 66121 9716 66130
rect 9868 66128 9908 66340
rect 9964 66305 10004 66390
rect 9963 66296 10005 66305
rect 9963 66256 9964 66296
rect 10004 66256 10005 66296
rect 9963 66247 10005 66256
rect 9964 66128 10004 66137
rect 9868 66088 9964 66128
rect 9676 66053 9716 66081
rect 9964 66079 10004 66088
rect 9675 66044 9717 66053
rect 9675 66004 9676 66044
rect 9716 66004 9717 66044
rect 9675 65995 9717 66004
rect 9676 65986 9716 65995
rect 9675 65876 9717 65885
rect 9675 65836 9676 65876
rect 9716 65836 9717 65876
rect 9675 65827 9717 65836
rect 9676 65456 9716 65827
rect 9579 64952 9621 64961
rect 9579 64912 9580 64952
rect 9620 64912 9621 64952
rect 9579 64903 9621 64912
rect 8908 64567 8948 64576
rect 9004 64616 9044 64625
rect 9004 64373 9044 64576
rect 9580 64616 9620 64627
rect 9580 64541 9620 64576
rect 9579 64532 9621 64541
rect 9579 64492 9580 64532
rect 9620 64492 9621 64532
rect 9579 64483 9621 64492
rect 9196 64448 9236 64457
rect 9100 64408 9196 64448
rect 9003 64364 9045 64373
rect 9003 64324 9004 64364
rect 9044 64324 9045 64364
rect 9003 64315 9045 64324
rect 8812 64240 8948 64280
rect 8811 63944 8853 63953
rect 8811 63904 8812 63944
rect 8852 63904 8853 63944
rect 8811 63895 8853 63904
rect 8812 63810 8852 63895
rect 8811 63608 8853 63617
rect 8811 63568 8812 63608
rect 8852 63568 8853 63608
rect 8811 63559 8853 63568
rect 8812 63197 8852 63559
rect 8811 63188 8853 63197
rect 8811 63148 8812 63188
rect 8852 63148 8853 63188
rect 8811 63139 8853 63148
rect 8715 63104 8757 63113
rect 8715 63064 8716 63104
rect 8756 63064 8757 63104
rect 8715 63055 8757 63064
rect 8716 62970 8756 63055
rect 8812 62852 8852 63139
rect 8716 62812 8852 62852
rect 8716 62432 8756 62812
rect 8427 61844 8469 61853
rect 8716 61844 8756 62392
rect 8908 62348 8948 64240
rect 9100 63356 9140 64408
rect 9196 64399 9236 64408
rect 9195 64280 9237 64289
rect 9676 64280 9716 65416
rect 10060 65045 10100 67507
rect 10251 67220 10293 67229
rect 10251 67180 10252 67220
rect 10292 67180 10293 67220
rect 10251 67171 10293 67180
rect 10252 66968 10292 67171
rect 10252 66919 10292 66928
rect 10251 66380 10293 66389
rect 10251 66340 10252 66380
rect 10292 66340 10293 66380
rect 10251 66331 10293 66340
rect 10155 65960 10197 65969
rect 10155 65920 10156 65960
rect 10196 65920 10197 65960
rect 10155 65911 10197 65920
rect 10156 65826 10196 65911
rect 10059 65036 10101 65045
rect 10059 64996 10060 65036
rect 10100 64996 10101 65036
rect 10059 64987 10101 64996
rect 9195 64240 9196 64280
rect 9236 64240 9237 64280
rect 9195 64231 9237 64240
rect 9484 64240 9716 64280
rect 9004 63316 9140 63356
rect 9004 62441 9044 63316
rect 9196 63118 9236 64231
rect 9291 63692 9333 63701
rect 9291 63652 9292 63692
rect 9332 63652 9333 63692
rect 9291 63643 9333 63652
rect 9100 63078 9196 63118
rect 9003 62432 9045 62441
rect 9003 62392 9004 62432
rect 9044 62392 9045 62432
rect 9003 62383 9045 62392
rect 9100 62432 9140 63078
rect 9196 63069 9236 63078
rect 9195 62600 9237 62609
rect 9195 62560 9196 62600
rect 9236 62560 9237 62600
rect 9195 62551 9237 62560
rect 9100 62357 9140 62392
rect 9196 62432 9236 62551
rect 9099 62348 9141 62357
rect 8427 61804 8428 61844
rect 8468 61804 8469 61844
rect 8427 61795 8469 61804
rect 8524 61804 8756 61844
rect 8812 62308 8948 62348
rect 9087 62308 9100 62348
rect 9140 62308 9141 62348
rect 8331 61592 8373 61601
rect 8331 61552 8332 61592
rect 8372 61552 8373 61592
rect 8331 61543 8373 61552
rect 8332 59240 8372 61543
rect 8524 60593 8564 61804
rect 8715 61676 8757 61685
rect 8715 61636 8716 61676
rect 8756 61636 8757 61676
rect 8715 61627 8757 61636
rect 8716 61013 8756 61627
rect 8715 61004 8757 61013
rect 8715 60964 8716 61004
rect 8756 60964 8757 61004
rect 8715 60955 8757 60964
rect 8619 60920 8661 60929
rect 8619 60880 8620 60920
rect 8660 60880 8661 60920
rect 8619 60871 8661 60880
rect 8716 60920 8756 60955
rect 8523 60584 8565 60593
rect 8523 60544 8524 60584
rect 8564 60544 8565 60584
rect 8523 60535 8565 60544
rect 8427 60080 8469 60089
rect 8427 60040 8428 60080
rect 8468 60040 8469 60080
rect 8427 60031 8469 60040
rect 8428 59408 8468 60031
rect 8523 59912 8565 59921
rect 8523 59872 8524 59912
rect 8564 59872 8565 59912
rect 8523 59863 8565 59872
rect 8428 59359 8468 59368
rect 8524 59408 8564 59863
rect 8620 59408 8660 60871
rect 8716 60869 8756 60880
rect 8812 60836 8852 62308
rect 9087 62299 9141 62308
rect 9087 62264 9127 62299
rect 8908 62224 9127 62264
rect 8908 62180 8948 62224
rect 8908 62131 8948 62140
rect 9003 61760 9045 61769
rect 9003 61720 9004 61760
rect 9044 61720 9045 61760
rect 9003 61711 9045 61720
rect 9004 61592 9044 61711
rect 8908 61013 8948 61098
rect 8907 61004 8949 61013
rect 8907 60964 8908 61004
rect 8948 60964 8949 61004
rect 8907 60955 8949 60964
rect 8812 60796 8948 60836
rect 8811 60668 8853 60677
rect 8811 60628 8812 60668
rect 8852 60628 8853 60668
rect 8811 60619 8853 60628
rect 8715 60416 8757 60425
rect 8715 60376 8716 60416
rect 8756 60376 8757 60416
rect 8715 60367 8757 60376
rect 8716 60080 8756 60367
rect 8716 60031 8756 60040
rect 8716 59408 8756 59417
rect 8620 59368 8716 59408
rect 8524 59359 8564 59368
rect 8716 59359 8756 59368
rect 8812 59408 8852 60619
rect 8908 60173 8948 60796
rect 9004 60425 9044 61552
rect 9196 61088 9236 62392
rect 9292 62432 9332 63643
rect 9387 63440 9429 63449
rect 9387 63400 9388 63440
rect 9428 63400 9429 63440
rect 9387 63391 9429 63400
rect 9388 63020 9428 63391
rect 9388 62971 9428 62980
rect 9387 62600 9429 62609
rect 9387 62560 9388 62600
rect 9428 62560 9429 62600
rect 9387 62551 9429 62560
rect 9388 62466 9428 62551
rect 9292 62383 9332 62392
rect 9484 62096 9524 64240
rect 9963 64196 10005 64205
rect 9963 64156 9964 64196
rect 10004 64156 10005 64196
rect 9963 64147 10005 64156
rect 9579 63776 9621 63785
rect 9579 63736 9580 63776
rect 9620 63736 9621 63776
rect 9579 63727 9621 63736
rect 9580 62432 9620 63727
rect 9964 63281 10004 64147
rect 10059 64112 10101 64121
rect 10059 64072 10060 64112
rect 10100 64072 10101 64112
rect 10059 64063 10101 64072
rect 10060 63944 10100 64063
rect 10252 64037 10292 66331
rect 10348 64121 10388 68440
rect 10444 64625 10484 68944
rect 10732 68657 10772 69117
rect 10924 68732 10964 72715
rect 11020 69152 11060 73060
rect 11115 69992 11157 70001
rect 11115 69952 11116 69992
rect 11156 69952 11157 69992
rect 11115 69943 11157 69952
rect 11116 69749 11156 69943
rect 11115 69740 11157 69749
rect 11115 69700 11116 69740
rect 11156 69700 11157 69740
rect 11115 69691 11157 69700
rect 11020 69103 11060 69112
rect 11212 68816 11252 75832
rect 11403 75620 11445 75629
rect 11403 75580 11404 75620
rect 11444 75580 11445 75620
rect 11403 75571 11445 75580
rect 11307 75284 11349 75293
rect 11307 75244 11308 75284
rect 11348 75244 11349 75284
rect 11307 75235 11349 75244
rect 11404 75284 11444 75571
rect 11499 75536 11541 75545
rect 11499 75496 11500 75536
rect 11540 75496 11541 75536
rect 11499 75487 11541 75496
rect 11404 75235 11444 75244
rect 11308 75150 11348 75235
rect 11403 74948 11445 74957
rect 11403 74908 11404 74948
rect 11444 74908 11445 74948
rect 11403 74899 11445 74908
rect 11320 74537 11360 74556
rect 11308 74528 11360 74537
rect 11404 74528 11444 74899
rect 11348 74488 11444 74528
rect 11308 74479 11348 74488
rect 11500 74444 11540 75487
rect 11404 74404 11540 74444
rect 11307 73352 11349 73361
rect 11307 73312 11308 73352
rect 11348 73312 11349 73352
rect 11307 73303 11349 73312
rect 11308 71765 11348 73303
rect 11307 71756 11349 71765
rect 11307 71716 11308 71756
rect 11348 71716 11349 71756
rect 11307 71707 11349 71716
rect 11308 69740 11348 69749
rect 11308 69161 11348 69700
rect 11307 69152 11349 69161
rect 11307 69112 11308 69152
rect 11348 69112 11349 69152
rect 11307 69103 11349 69112
rect 11212 68776 11348 68816
rect 10924 68692 11252 68732
rect 10731 68648 10773 68657
rect 10731 68608 10732 68648
rect 10772 68608 10773 68648
rect 10731 68599 10773 68608
rect 10635 68396 10677 68405
rect 10635 68356 10636 68396
rect 10676 68356 10677 68396
rect 10635 68347 10677 68356
rect 10636 67640 10676 68347
rect 10539 64784 10581 64793
rect 10539 64744 10540 64784
rect 10580 64744 10581 64784
rect 10539 64735 10581 64744
rect 10443 64616 10485 64625
rect 10443 64576 10444 64616
rect 10484 64576 10485 64616
rect 10443 64567 10485 64576
rect 10347 64112 10389 64121
rect 10347 64072 10348 64112
rect 10388 64072 10389 64112
rect 10347 64063 10389 64072
rect 10540 64037 10580 64735
rect 10636 64121 10676 67600
rect 10635 64112 10677 64121
rect 10635 64072 10636 64112
rect 10676 64072 10677 64112
rect 10635 64063 10677 64072
rect 10251 64028 10293 64037
rect 10251 63988 10252 64028
rect 10292 63988 10293 64028
rect 10251 63979 10293 63988
rect 10539 64028 10581 64037
rect 10539 63988 10540 64028
rect 10580 63988 10581 64028
rect 10539 63979 10581 63988
rect 10060 63617 10100 63904
rect 10252 63692 10292 63701
rect 10292 63652 10484 63692
rect 10252 63643 10292 63652
rect 10059 63608 10101 63617
rect 10059 63568 10060 63608
rect 10100 63568 10101 63608
rect 10059 63559 10101 63568
rect 10251 63356 10293 63365
rect 10251 63316 10252 63356
rect 10292 63316 10293 63356
rect 10251 63307 10293 63316
rect 9963 63272 10005 63281
rect 9963 63232 9964 63272
rect 10004 63232 10005 63272
rect 9963 63223 10005 63232
rect 9867 63188 9909 63197
rect 9867 63148 9868 63188
rect 9908 63148 9909 63188
rect 9867 63139 9909 63148
rect 10252 63146 10292 63307
rect 9772 63104 9812 63113
rect 9675 62600 9717 62609
rect 9772 62600 9812 63064
rect 9868 63104 9908 63139
rect 9868 63053 9908 63064
rect 10059 63104 10101 63113
rect 10059 63064 10060 63104
rect 10100 63064 10101 63104
rect 10444 63113 10484 63652
rect 10539 63608 10581 63617
rect 10732 63608 10772 68599
rect 11116 67645 11156 67654
rect 11116 67145 11156 67605
rect 11115 67136 11157 67145
rect 11115 67096 11116 67136
rect 11156 67096 11157 67136
rect 11115 67087 11157 67096
rect 10924 65456 10964 65465
rect 10827 65372 10869 65381
rect 10827 65332 10828 65372
rect 10868 65332 10869 65372
rect 10827 65323 10869 65332
rect 10828 64616 10868 65323
rect 10924 64793 10964 65416
rect 11116 65456 11156 65465
rect 11019 64868 11061 64877
rect 11019 64828 11020 64868
rect 11060 64828 11061 64868
rect 11019 64819 11061 64828
rect 10923 64784 10965 64793
rect 10923 64744 10924 64784
rect 10964 64744 10965 64784
rect 10923 64735 10965 64744
rect 11020 64734 11060 64819
rect 10828 64567 10868 64576
rect 11019 64616 11061 64625
rect 11019 64576 11020 64616
rect 11060 64576 11061 64616
rect 11019 64567 11061 64576
rect 11020 64280 11060 64567
rect 11116 64457 11156 65416
rect 11115 64448 11157 64457
rect 11115 64408 11116 64448
rect 11156 64408 11157 64448
rect 11115 64399 11157 64408
rect 11020 64240 11156 64280
rect 10923 64028 10965 64037
rect 10923 63988 10924 64028
rect 10964 63988 10965 64028
rect 10923 63979 10965 63988
rect 10827 63944 10869 63953
rect 10827 63904 10828 63944
rect 10868 63904 10869 63944
rect 10827 63895 10869 63904
rect 10828 63810 10868 63895
rect 10539 63568 10540 63608
rect 10580 63568 10581 63608
rect 10539 63559 10581 63568
rect 10636 63568 10772 63608
rect 10252 63097 10292 63106
rect 10348 63104 10388 63113
rect 10059 63055 10101 63064
rect 9963 63020 10005 63029
rect 9963 62980 9964 63020
rect 10004 62980 10005 63020
rect 9963 62971 10005 62980
rect 9964 62886 10004 62971
rect 10060 62970 10100 63055
rect 10348 62609 10388 63064
rect 10443 63104 10485 63113
rect 10443 63064 10444 63104
rect 10484 63064 10485 63104
rect 10443 63055 10485 63064
rect 10540 63104 10580 63559
rect 10540 63055 10580 63064
rect 10444 62970 10484 63055
rect 9675 62560 9676 62600
rect 9716 62560 9812 62600
rect 9867 62600 9909 62609
rect 9867 62560 9868 62600
rect 9908 62560 9909 62600
rect 9675 62551 9717 62560
rect 9867 62551 9909 62560
rect 10347 62600 10389 62609
rect 10347 62560 10348 62600
rect 10388 62560 10389 62600
rect 10347 62551 10389 62560
rect 9868 62466 9908 62551
rect 9580 62383 9620 62392
rect 9676 62432 9716 62443
rect 9676 62357 9716 62392
rect 9771 62432 9813 62441
rect 9771 62392 9772 62432
rect 9812 62392 9813 62432
rect 9771 62383 9813 62392
rect 10155 62432 10197 62441
rect 10155 62392 10156 62432
rect 10196 62392 10197 62432
rect 10155 62383 10197 62392
rect 10252 62432 10292 62441
rect 10636 62432 10676 63568
rect 10731 63440 10773 63449
rect 10731 63400 10732 63440
rect 10772 63400 10773 63440
rect 10731 63391 10773 63400
rect 10732 63104 10772 63391
rect 10924 63281 10964 63979
rect 11019 63608 11061 63617
rect 11019 63568 11020 63608
rect 11060 63568 11061 63608
rect 11019 63559 11061 63568
rect 10923 63272 10965 63281
rect 10923 63232 10924 63272
rect 10964 63232 10965 63272
rect 10923 63223 10965 63232
rect 10732 63055 10772 63064
rect 10923 63104 10965 63113
rect 10923 63064 10924 63104
rect 10964 63064 10965 63104
rect 11020 63104 11060 63559
rect 11116 63356 11156 64240
rect 11212 63533 11252 68692
rect 11308 68573 11348 68776
rect 11307 68564 11349 68573
rect 11307 68524 11308 68564
rect 11348 68524 11349 68564
rect 11307 68515 11349 68524
rect 11404 68480 11444 74404
rect 11596 74360 11636 80611
rect 11788 76712 11828 76721
rect 11788 75461 11828 76672
rect 11787 75452 11829 75461
rect 11787 75412 11788 75452
rect 11828 75412 11829 75452
rect 11787 75403 11829 75412
rect 11884 75200 11924 81880
rect 11979 80576 12021 80585
rect 11979 80536 11980 80576
rect 12020 80536 12021 80576
rect 11979 80527 12021 80536
rect 11884 75151 11924 75160
rect 11787 74696 11829 74705
rect 11787 74656 11788 74696
rect 11828 74656 11829 74696
rect 11787 74647 11829 74656
rect 11500 74320 11636 74360
rect 11500 69320 11540 74320
rect 11595 73688 11637 73697
rect 11595 73648 11596 73688
rect 11636 73648 11637 73688
rect 11595 73639 11637 73648
rect 11596 73193 11636 73639
rect 11595 73184 11637 73193
rect 11595 73144 11596 73184
rect 11636 73144 11637 73184
rect 11595 73135 11637 73144
rect 11788 73184 11828 74647
rect 11788 73144 11924 73184
rect 11788 70664 11828 73144
rect 11884 73025 11924 73144
rect 11883 73016 11925 73025
rect 11883 72976 11884 73016
rect 11924 72976 11925 73016
rect 11883 72967 11925 72976
rect 11883 72764 11925 72773
rect 11883 72724 11884 72764
rect 11924 72724 11925 72764
rect 11883 72715 11925 72724
rect 11884 72176 11924 72715
rect 11884 72127 11924 72136
rect 11980 72176 12020 80527
rect 11980 72101 12020 72136
rect 11979 72092 12021 72101
rect 11979 72052 11980 72092
rect 12020 72052 12021 72092
rect 11979 72043 12021 72052
rect 11980 70664 12020 70673
rect 11788 70624 11980 70664
rect 11595 70496 11637 70505
rect 11595 70456 11596 70496
rect 11636 70456 11637 70496
rect 11595 70447 11637 70456
rect 11596 69992 11636 70447
rect 11883 70160 11925 70169
rect 11883 70120 11884 70160
rect 11924 70120 11925 70160
rect 11883 70111 11925 70120
rect 11596 69943 11636 69952
rect 11691 69992 11733 70001
rect 11691 69952 11692 69992
rect 11732 69952 11733 69992
rect 11691 69943 11733 69952
rect 11692 69858 11732 69943
rect 11787 69320 11829 69329
rect 11500 69280 11636 69320
rect 11500 69161 11540 69166
rect 11499 69157 11541 69161
rect 11499 69112 11500 69157
rect 11540 69112 11541 69157
rect 11499 69103 11541 69112
rect 11500 69022 11540 69103
rect 11500 68480 11540 68489
rect 11404 68440 11500 68480
rect 11307 67472 11349 67481
rect 11307 67432 11308 67472
rect 11348 67432 11349 67472
rect 11307 67423 11349 67432
rect 11308 67338 11348 67423
rect 11404 65960 11444 68440
rect 11500 68431 11540 68440
rect 11500 66977 11540 67062
rect 11499 66968 11541 66977
rect 11499 66928 11500 66968
rect 11540 66928 11541 66968
rect 11499 66919 11541 66928
rect 11404 65920 11540 65960
rect 11307 65288 11349 65297
rect 11307 65248 11308 65288
rect 11348 65248 11349 65288
rect 11307 65239 11349 65248
rect 11308 64877 11348 65239
rect 11307 64868 11349 64877
rect 11307 64828 11308 64868
rect 11348 64828 11349 64868
rect 11307 64819 11349 64828
rect 11308 64616 11348 64819
rect 11308 64567 11348 64576
rect 11404 64616 11444 64625
rect 11211 63524 11253 63533
rect 11211 63484 11212 63524
rect 11252 63484 11253 63524
rect 11211 63475 11253 63484
rect 11116 63316 11348 63356
rect 11211 63188 11253 63197
rect 11211 63148 11212 63188
rect 11252 63148 11253 63188
rect 11211 63139 11253 63148
rect 11116 63104 11156 63113
rect 11020 63064 11116 63104
rect 10923 63055 10965 63064
rect 11116 63055 11156 63064
rect 10827 63020 10869 63029
rect 10827 62980 10828 63020
rect 10868 62980 10869 63020
rect 10827 62971 10869 62980
rect 10731 62936 10773 62945
rect 10731 62896 10732 62936
rect 10772 62896 10773 62936
rect 10731 62887 10773 62896
rect 10292 62392 10676 62432
rect 10252 62383 10292 62392
rect 9675 62348 9717 62357
rect 9675 62308 9676 62348
rect 9716 62308 9717 62348
rect 9675 62299 9717 62308
rect 9772 62298 9812 62383
rect 9484 62056 10004 62096
rect 9579 61928 9621 61937
rect 9579 61888 9580 61928
rect 9620 61888 9621 61928
rect 9579 61879 9621 61888
rect 9580 61424 9620 61879
rect 9676 61601 9716 61686
rect 9675 61592 9717 61601
rect 9675 61552 9676 61592
rect 9716 61552 9717 61592
rect 9675 61543 9717 61552
rect 9580 61384 9716 61424
rect 9483 61172 9525 61181
rect 9483 61132 9484 61172
rect 9524 61132 9525 61172
rect 9483 61123 9525 61132
rect 9196 61048 9428 61088
rect 9099 61004 9141 61013
rect 9099 60964 9100 61004
rect 9140 60964 9236 61004
rect 9099 60955 9141 60964
rect 9196 60920 9236 60964
rect 9196 60871 9236 60880
rect 9292 60920 9332 60931
rect 9292 60845 9332 60880
rect 9291 60836 9333 60845
rect 9291 60796 9292 60836
rect 9332 60796 9333 60836
rect 9291 60787 9333 60796
rect 9003 60416 9045 60425
rect 9003 60376 9004 60416
rect 9044 60376 9045 60416
rect 9003 60367 9045 60376
rect 9291 60248 9333 60257
rect 9291 60208 9292 60248
rect 9332 60208 9333 60248
rect 9291 60199 9333 60208
rect 8907 60164 8949 60173
rect 8907 60124 8908 60164
rect 8948 60124 8949 60164
rect 8907 60115 8949 60124
rect 9196 60080 9236 60089
rect 9004 60040 9196 60080
rect 8908 59996 8948 60005
rect 9004 59996 9044 60040
rect 9196 60031 9236 60040
rect 9292 60080 9332 60199
rect 8948 59956 9044 59996
rect 8908 59947 8948 59956
rect 9099 59912 9141 59921
rect 9099 59872 9100 59912
rect 9140 59872 9141 59912
rect 9099 59863 9141 59872
rect 9003 59828 9045 59837
rect 9003 59788 9004 59828
rect 9044 59788 9045 59828
rect 9003 59779 9045 59788
rect 8812 59359 8852 59368
rect 8912 59408 8954 59417
rect 8912 59368 8913 59408
rect 8953 59368 8954 59408
rect 8912 59359 8954 59368
rect 8913 59274 8953 59359
rect 8619 59240 8661 59249
rect 8332 59200 8468 59240
rect 8236 59156 8276 59165
rect 8428 59156 8468 59200
rect 8619 59200 8620 59240
rect 8660 59200 8661 59240
rect 8619 59191 8661 59200
rect 8276 59116 8372 59156
rect 8236 59107 8276 59116
rect 8332 57896 8372 59116
rect 8428 59107 8468 59116
rect 8620 58568 8660 59191
rect 9004 59156 9044 59779
rect 8620 58519 8660 58528
rect 8908 59116 9044 59156
rect 8812 58400 8852 58409
rect 8716 58360 8812 58400
rect 8428 57896 8468 57905
rect 8332 57856 8428 57896
rect 8428 57847 8468 57856
rect 8523 57896 8565 57905
rect 8523 57856 8524 57896
rect 8564 57856 8565 57896
rect 8523 57847 8565 57856
rect 8524 57762 8564 57847
rect 8139 57728 8181 57737
rect 8139 57688 8140 57728
rect 8180 57688 8181 57728
rect 8139 57679 8181 57688
rect 8043 57140 8085 57149
rect 8043 57100 8044 57140
rect 8084 57100 8085 57140
rect 8043 57091 8085 57100
rect 7947 56720 7989 56729
rect 7947 56680 7948 56720
rect 7988 56680 7989 56720
rect 7947 56671 7989 56680
rect 7947 56384 7989 56393
rect 7947 56344 7948 56384
rect 7988 56344 7989 56384
rect 7947 56335 7989 56344
rect 8044 56384 8084 57091
rect 8716 57070 8756 58360
rect 8812 58351 8852 58360
rect 8908 57896 8948 59116
rect 9004 58661 9044 58692
rect 9003 58652 9045 58661
rect 9003 58612 9004 58652
rect 9044 58612 9045 58652
rect 9003 58603 9045 58612
rect 9004 58568 9044 58603
rect 9004 58493 9044 58528
rect 9003 58484 9045 58493
rect 9003 58444 9004 58484
rect 9044 58444 9045 58484
rect 9003 58435 9045 58444
rect 8908 57847 8948 57856
rect 9004 57812 9044 57821
rect 8811 57728 8853 57737
rect 9004 57728 9044 57772
rect 8811 57688 8812 57728
rect 8852 57688 9044 57728
rect 8811 57679 8853 57688
rect 8235 57056 8277 57065
rect 8523 57056 8565 57065
rect 8235 57016 8236 57056
rect 8276 57016 8372 57056
rect 8235 57007 8277 57016
rect 8236 56922 8276 57007
rect 8084 56344 8276 56384
rect 8044 56335 8084 56344
rect 7948 56048 7988 56335
rect 7948 56008 8084 56048
rect 7948 55544 7988 55553
rect 7852 55504 7948 55544
rect 7948 55495 7988 55504
rect 8044 55544 8084 56008
rect 7564 55420 7700 55460
rect 6700 54209 6740 54832
rect 6988 54788 7028 55420
rect 6796 54748 7028 54788
rect 6699 54200 6741 54209
rect 6699 54160 6700 54200
rect 6740 54160 6741 54200
rect 6699 54151 6741 54160
rect 6700 54032 6740 54043
rect 6700 53957 6740 53992
rect 6699 53948 6741 53957
rect 6699 53908 6700 53948
rect 6740 53908 6741 53948
rect 6699 53899 6741 53908
rect 6796 52772 6836 54748
rect 6412 50128 6644 50168
rect 6700 52732 6836 52772
rect 6892 54620 6932 54629
rect 6315 49328 6357 49337
rect 6315 49288 6316 49328
rect 6356 49288 6357 49328
rect 6315 49279 6357 49288
rect 6316 48824 6356 49279
rect 6316 48775 6356 48784
rect 6315 48236 6357 48245
rect 6315 48196 6316 48236
rect 6356 48196 6357 48236
rect 6315 48187 6357 48196
rect 6316 46640 6356 48187
rect 6412 48068 6452 50128
rect 6700 49505 6740 52732
rect 6795 52604 6837 52613
rect 6795 52564 6796 52604
rect 6836 52564 6837 52604
rect 6795 52555 6837 52564
rect 6796 50840 6836 52555
rect 6892 52520 6932 54580
rect 7083 54032 7125 54041
rect 7083 53992 7084 54032
rect 7124 53992 7125 54032
rect 7083 53983 7125 53992
rect 7084 53360 7124 53983
rect 7084 53311 7124 53320
rect 6892 52471 6932 52480
rect 6987 52520 7029 52529
rect 6987 52480 6988 52520
rect 7028 52480 7029 52520
rect 6987 52471 7029 52480
rect 6988 52386 7028 52471
rect 7180 52277 7220 55420
rect 7563 54872 7605 54881
rect 7563 54832 7564 54872
rect 7604 54832 7605 54872
rect 7563 54823 7605 54832
rect 7564 54125 7604 54823
rect 7563 54116 7605 54125
rect 7563 54076 7564 54116
rect 7604 54076 7605 54116
rect 7563 54067 7605 54076
rect 7564 53873 7604 54067
rect 7563 53864 7605 53873
rect 7563 53824 7564 53864
rect 7604 53824 7605 53864
rect 7563 53815 7605 53824
rect 7276 53444 7316 53453
rect 7316 53404 7604 53444
rect 7276 53395 7316 53404
rect 7564 53360 7604 53404
rect 7564 53311 7604 53320
rect 7660 53360 7700 55420
rect 7755 55124 7797 55133
rect 7755 55084 7756 55124
rect 7796 55084 7797 55124
rect 7755 55075 7797 55084
rect 7371 52940 7413 52949
rect 7371 52900 7372 52940
rect 7412 52900 7413 52940
rect 7371 52891 7413 52900
rect 7275 52772 7317 52781
rect 7275 52732 7276 52772
rect 7316 52732 7317 52772
rect 7275 52723 7317 52732
rect 7179 52268 7221 52277
rect 7179 52228 7180 52268
rect 7220 52228 7221 52268
rect 7179 52219 7221 52228
rect 7083 52100 7125 52109
rect 7083 52060 7084 52100
rect 7124 52060 7125 52100
rect 7083 52051 7125 52060
rect 6891 51596 6933 51605
rect 6891 51556 6892 51596
rect 6932 51556 6933 51596
rect 6891 51547 6933 51556
rect 6892 51022 6932 51547
rect 6892 50973 6932 50982
rect 7084 51008 7124 52051
rect 7179 52016 7221 52025
rect 7179 51976 7180 52016
rect 7220 51976 7221 52016
rect 7179 51967 7221 51976
rect 7180 51848 7220 51967
rect 7276 51941 7316 52723
rect 7372 52520 7412 52891
rect 7660 52529 7700 53320
rect 7372 52445 7412 52480
rect 7468 52520 7508 52529
rect 7371 52436 7413 52445
rect 7371 52396 7372 52436
rect 7412 52396 7413 52436
rect 7371 52387 7413 52396
rect 7468 52277 7508 52480
rect 7659 52520 7701 52529
rect 7659 52480 7660 52520
rect 7700 52480 7701 52520
rect 7659 52471 7701 52480
rect 7467 52268 7509 52277
rect 7467 52228 7468 52268
rect 7508 52228 7509 52268
rect 7467 52219 7509 52228
rect 7275 51932 7317 51941
rect 7275 51892 7276 51932
rect 7316 51892 7317 51932
rect 7275 51883 7317 51892
rect 7180 51680 7220 51808
rect 7276 51764 7316 51883
rect 7276 51724 7508 51764
rect 7180 51640 7316 51680
rect 7084 50968 7220 51008
rect 7084 50840 7124 50849
rect 6796 50800 7084 50840
rect 7084 50791 7124 50800
rect 6795 50336 6837 50345
rect 6795 50296 6796 50336
rect 6836 50296 6837 50336
rect 6795 50287 6837 50296
rect 6699 49496 6741 49505
rect 6699 49456 6700 49496
rect 6740 49456 6741 49496
rect 6699 49447 6741 49456
rect 6700 48656 6740 49447
rect 6796 49169 6836 50287
rect 7083 50000 7125 50009
rect 7083 49960 7084 50000
rect 7124 49960 7125 50000
rect 7083 49951 7125 49960
rect 7084 49496 7124 49951
rect 7084 49337 7124 49456
rect 7083 49328 7125 49337
rect 7083 49288 7084 49328
rect 7124 49288 7125 49328
rect 7083 49279 7125 49288
rect 6795 49160 6837 49169
rect 6795 49120 6796 49160
rect 6836 49120 6837 49160
rect 6795 49111 6837 49120
rect 6796 48824 6836 49111
rect 6796 48775 6836 48784
rect 6700 48616 6836 48656
rect 6508 48572 6548 48581
rect 6548 48532 6644 48572
rect 6508 48523 6548 48532
rect 6507 48236 6549 48245
rect 6507 48196 6508 48236
rect 6548 48196 6549 48236
rect 6507 48187 6549 48196
rect 6412 47321 6452 48028
rect 6508 48068 6548 48187
rect 6508 48019 6548 48028
rect 6411 47312 6453 47321
rect 6604 47312 6644 48532
rect 6699 48068 6741 48077
rect 6699 48028 6700 48068
rect 6740 48028 6741 48068
rect 6699 48019 6741 48028
rect 6700 47480 6740 48019
rect 6700 47431 6740 47440
rect 6411 47272 6412 47312
rect 6452 47272 6453 47312
rect 6411 47263 6453 47272
rect 6556 47302 6644 47312
rect 6596 47272 6644 47302
rect 6556 47253 6596 47262
rect 6796 46640 6836 48616
rect 6891 48068 6933 48077
rect 6891 48028 6892 48068
rect 6932 48028 6933 48068
rect 6891 48019 6933 48028
rect 6892 47984 6932 48019
rect 6892 47933 6932 47944
rect 6988 47984 7028 47995
rect 6988 47909 7028 47944
rect 6987 47900 7029 47909
rect 6987 47860 6988 47900
rect 7028 47860 7029 47900
rect 6987 47851 7029 47860
rect 7084 46649 7124 49279
rect 6316 46600 6452 46640
rect 6315 45968 6357 45977
rect 6315 45928 6316 45968
rect 6356 45928 6357 45968
rect 6315 45919 6357 45928
rect 6316 45800 6356 45919
rect 6316 45751 6356 45760
rect 6219 45464 6261 45473
rect 5836 45424 5972 45464
rect 5740 45172 5876 45212
rect 5644 45088 5780 45128
rect 5644 44960 5684 44969
rect 5548 44920 5644 44960
rect 5644 44911 5684 44920
rect 5740 44960 5780 45088
rect 5643 44372 5685 44381
rect 5740 44372 5780 44920
rect 5643 44332 5644 44372
rect 5684 44332 5780 44372
rect 5643 44323 5685 44332
rect 5548 44288 5588 44297
rect 5548 44129 5588 44248
rect 5644 44288 5684 44323
rect 5644 44237 5684 44248
rect 5547 44120 5589 44129
rect 5547 44080 5548 44120
rect 5588 44080 5589 44120
rect 5547 44071 5589 44080
rect 5836 43616 5876 45172
rect 5932 44885 5972 45424
rect 6219 45424 6220 45464
rect 6260 45424 6261 45464
rect 6219 45415 6261 45424
rect 6412 45296 6452 46600
rect 6700 46600 6836 46640
rect 7083 46640 7125 46649
rect 7083 46600 7084 46640
rect 7124 46600 7125 46640
rect 6700 45977 6740 46600
rect 7083 46591 7125 46600
rect 7180 46472 7220 50968
rect 7276 50840 7316 51640
rect 7371 51596 7413 51605
rect 7371 51556 7372 51596
rect 7412 51556 7413 51596
rect 7371 51547 7413 51556
rect 7372 51462 7412 51547
rect 7276 50800 7412 50840
rect 7275 50588 7317 50597
rect 7275 50548 7276 50588
rect 7316 50548 7317 50588
rect 7275 50539 7317 50548
rect 7276 49748 7316 50539
rect 7276 49699 7316 49708
rect 7275 49160 7317 49169
rect 7275 49120 7276 49160
rect 7316 49120 7317 49160
rect 7275 49111 7317 49120
rect 6796 46432 7220 46472
rect 6699 45968 6741 45977
rect 6699 45928 6700 45968
rect 6740 45928 6741 45968
rect 6699 45919 6741 45928
rect 6124 45256 6452 45296
rect 6124 45044 6164 45256
rect 6028 45004 6124 45044
rect 5931 44876 5973 44885
rect 5931 44836 5932 44876
rect 5972 44836 5973 44876
rect 5931 44827 5973 44836
rect 6028 44288 6068 45004
rect 6124 44995 6164 45004
rect 6220 44960 6260 44971
rect 6220 44885 6260 44920
rect 6700 44960 6740 44969
rect 6219 44876 6261 44885
rect 6219 44836 6220 44876
rect 6260 44836 6261 44876
rect 6219 44827 6261 44836
rect 6028 44239 6068 44248
rect 6124 44288 6164 44297
rect 6220 44288 6260 44827
rect 6700 44801 6740 44920
rect 6699 44792 6741 44801
rect 6699 44752 6700 44792
rect 6740 44752 6741 44792
rect 6699 44743 6741 44752
rect 6164 44248 6260 44288
rect 6604 44288 6644 44297
rect 6700 44288 6740 44743
rect 6644 44248 6740 44288
rect 6124 44239 6164 44248
rect 6604 44239 6644 44248
rect 6219 44036 6261 44045
rect 6219 43996 6220 44036
rect 6260 43996 6261 44036
rect 6219 43987 6261 43996
rect 5644 43576 5876 43616
rect 5259 42568 5260 42608
rect 5300 42568 5396 42608
rect 5452 42692 5492 42701
rect 5259 42559 5301 42568
rect 5163 42524 5205 42533
rect 5163 42484 5164 42524
rect 5204 42484 5205 42524
rect 5163 42475 5205 42484
rect 5164 42365 5204 42475
rect 5163 42356 5205 42365
rect 5163 42316 5164 42356
rect 5204 42316 5205 42356
rect 5163 42307 5205 42316
rect 4876 42055 4916 42064
rect 5260 41936 5300 42559
rect 5452 42533 5492 42652
rect 5548 42692 5588 42701
rect 5451 42524 5493 42533
rect 5451 42484 5452 42524
rect 5492 42484 5493 42524
rect 5451 42475 5493 42484
rect 5260 41887 5300 41896
rect 4928 41600 5296 41609
rect 4968 41560 5010 41600
rect 5050 41560 5092 41600
rect 5132 41560 5174 41600
rect 5214 41560 5256 41600
rect 4928 41551 5296 41560
rect 5068 41348 5108 41357
rect 5108 41308 5396 41348
rect 5068 41299 5108 41308
rect 3628 41264 3668 41273
rect 3628 41021 3668 41224
rect 4299 41264 4341 41273
rect 4299 41224 4300 41264
rect 4340 41224 4341 41264
rect 4299 41215 4341 41224
rect 4491 41264 4533 41273
rect 4491 41224 4492 41264
rect 4532 41224 4533 41264
rect 4491 41215 4533 41224
rect 4875 41264 4917 41273
rect 4875 41224 4876 41264
rect 4916 41224 4917 41264
rect 4875 41215 4917 41224
rect 5356 41264 5396 41308
rect 5356 41215 5396 41224
rect 5451 41264 5493 41273
rect 5451 41224 5452 41264
rect 5492 41224 5493 41264
rect 5451 41215 5493 41224
rect 3627 41012 3669 41021
rect 3627 40972 3628 41012
rect 3668 40972 3669 41012
rect 3627 40963 3669 40972
rect 3688 40844 4056 40853
rect 3728 40804 3770 40844
rect 3810 40804 3852 40844
rect 3892 40804 3934 40844
rect 3974 40804 4016 40844
rect 3688 40795 4056 40804
rect 3532 40636 3764 40676
rect 3147 40340 3189 40349
rect 3147 40300 3148 40340
rect 3188 40300 3189 40340
rect 3147 40291 3189 40300
rect 3051 39920 3093 39929
rect 3724 39920 3764 40636
rect 3915 40508 3957 40517
rect 3915 40468 3916 40508
rect 3956 40468 3957 40508
rect 3915 40459 3957 40468
rect 3916 40424 3956 40459
rect 3916 40373 3956 40384
rect 4107 40340 4149 40349
rect 4107 40300 4108 40340
rect 4148 40300 4149 40340
rect 4107 40291 4149 40300
rect 3051 39880 3052 39920
rect 3092 39880 3093 39920
rect 3051 39871 3093 39880
rect 3148 39880 3572 39920
rect 2955 39752 2997 39761
rect 2955 39712 2956 39752
rect 2996 39712 2997 39752
rect 2955 39703 2997 39712
rect 3052 39752 3092 39871
rect 3052 39703 3092 39712
rect 3052 38408 3092 38417
rect 3148 38408 3188 39880
rect 3435 39752 3477 39761
rect 3435 39712 3436 39752
rect 3476 39712 3477 39752
rect 3435 39703 3477 39712
rect 3532 39747 3572 39880
rect 3724 39871 3764 39880
rect 3339 39584 3381 39593
rect 3339 39544 3340 39584
rect 3380 39544 3381 39584
rect 3339 39535 3381 39544
rect 3243 38912 3285 38921
rect 3243 38872 3244 38912
rect 3284 38872 3285 38912
rect 3243 38863 3285 38872
rect 3244 38778 3284 38863
rect 2860 38368 2996 38408
rect 2859 38240 2901 38249
rect 2859 38200 2860 38240
rect 2900 38200 2901 38240
rect 2859 38191 2901 38200
rect 2860 38106 2900 38191
rect 2956 37820 2996 38368
rect 3092 38368 3188 38408
rect 3052 38359 3092 38368
rect 3147 38240 3189 38249
rect 3147 38200 3148 38240
rect 3188 38200 3189 38240
rect 3147 38191 3189 38200
rect 3148 37829 3188 38191
rect 3147 37820 3189 37829
rect 2956 37780 3092 37820
rect 2859 37400 2901 37409
rect 2859 37360 2860 37400
rect 2900 37360 2901 37400
rect 2859 37351 2901 37360
rect 2956 37400 2996 37409
rect 2860 37266 2900 37351
rect 2956 36905 2996 37360
rect 2955 36896 2997 36905
rect 2955 36856 2956 36896
rect 2996 36856 2997 36896
rect 2955 36847 2997 36856
rect 2860 36728 2900 36737
rect 3052 36728 3092 37780
rect 3147 37780 3148 37820
rect 3188 37780 3189 37820
rect 3147 37771 3189 37780
rect 2900 36688 3092 36728
rect 2860 36679 2900 36688
rect 2955 36560 2997 36569
rect 2955 36520 2956 36560
rect 2996 36520 2997 36560
rect 2955 36511 2997 36520
rect 2860 35888 2900 35899
rect 2860 35813 2900 35848
rect 2859 35804 2901 35813
rect 2859 35764 2860 35804
rect 2900 35764 2901 35804
rect 2859 35755 2901 35764
rect 2859 35300 2901 35309
rect 2859 35260 2860 35300
rect 2900 35260 2901 35300
rect 2859 35251 2901 35260
rect 2860 35166 2900 35251
rect 2956 34973 2996 36511
rect 3051 35216 3093 35225
rect 3051 35176 3052 35216
rect 3092 35176 3093 35216
rect 3051 35167 3093 35176
rect 3052 35082 3092 35167
rect 2955 34964 2997 34973
rect 2955 34924 2956 34964
rect 2996 34924 2997 34964
rect 2955 34915 2997 34924
rect 2764 34504 2900 34544
rect 2667 34495 2709 34504
rect 2668 34460 2708 34495
rect 2668 34217 2708 34420
rect 2764 34376 2804 34385
rect 2667 34208 2709 34217
rect 2667 34168 2668 34208
rect 2708 34168 2709 34208
rect 2667 34159 2709 34168
rect 2571 33788 2613 33797
rect 2571 33748 2572 33788
rect 2612 33748 2613 33788
rect 2571 33739 2613 33748
rect 2475 33704 2517 33713
rect 2475 33664 2476 33704
rect 2516 33664 2517 33704
rect 2475 33655 2517 33664
rect 2764 33200 2804 34336
rect 2860 33881 2900 34504
rect 3148 34460 3188 37771
rect 3340 37652 3380 39535
rect 3436 39164 3476 39703
rect 3532 39698 3572 39707
rect 4011 39752 4053 39761
rect 4011 39712 4012 39752
rect 4052 39712 4053 39752
rect 4011 39703 4053 39712
rect 4108 39752 4148 40291
rect 4012 39618 4052 39703
rect 4108 39509 4148 39712
rect 4107 39500 4149 39509
rect 4107 39460 4108 39500
rect 4148 39460 4149 39500
rect 4107 39451 4149 39460
rect 3688 39332 4056 39341
rect 3728 39292 3770 39332
rect 3810 39292 3852 39332
rect 3892 39292 3934 39332
rect 3974 39292 4016 39332
rect 3688 39283 4056 39292
rect 3436 39115 3476 39124
rect 3628 38912 3668 38921
rect 3532 38872 3628 38912
rect 3532 37736 3572 38872
rect 3628 38863 3668 38872
rect 4300 38501 4340 41215
rect 4876 40769 4916 41215
rect 5452 41130 5492 41215
rect 4875 40760 4917 40769
rect 4875 40720 4876 40760
rect 4916 40720 4917 40760
rect 4875 40711 4917 40720
rect 5163 40760 5205 40769
rect 5163 40720 5164 40760
rect 5204 40720 5205 40760
rect 5163 40711 5205 40720
rect 4395 40508 4437 40517
rect 4395 40468 4396 40508
rect 4436 40468 4437 40508
rect 4395 40459 4437 40468
rect 4299 38492 4341 38501
rect 4299 38452 4300 38492
rect 4340 38452 4341 38492
rect 4299 38443 4341 38452
rect 4396 38333 4436 40459
rect 5164 40433 5204 40711
rect 5548 40433 5588 42652
rect 5163 40424 5205 40433
rect 5163 40384 5164 40424
rect 5204 40384 5205 40424
rect 5163 40375 5205 40384
rect 5547 40424 5589 40433
rect 5547 40384 5548 40424
rect 5588 40384 5589 40424
rect 5547 40375 5589 40384
rect 5164 40290 5204 40375
rect 5356 40256 5396 40265
rect 5396 40216 5588 40256
rect 5356 40207 5396 40216
rect 4928 40088 5296 40097
rect 4968 40048 5010 40088
rect 5050 40048 5092 40088
rect 5132 40048 5174 40088
rect 5214 40048 5256 40088
rect 4928 40039 5296 40048
rect 5355 40088 5397 40097
rect 5355 40048 5356 40088
rect 5396 40048 5397 40088
rect 5355 40039 5397 40048
rect 5068 39752 5108 39761
rect 5356 39752 5396 40039
rect 5108 39712 5396 39752
rect 5548 39747 5588 40216
rect 5068 39703 5108 39712
rect 5548 39698 5588 39707
rect 4492 39668 4532 39677
rect 4492 39425 4532 39628
rect 4587 39668 4629 39677
rect 4587 39628 4588 39668
rect 4628 39628 4629 39668
rect 4587 39619 4629 39628
rect 4588 39534 4628 39619
rect 4491 39416 4533 39425
rect 4491 39376 4492 39416
rect 4532 39376 4533 39416
rect 4491 39367 4533 39376
rect 5259 38996 5301 39005
rect 5259 38956 5260 38996
rect 5300 38956 5301 38996
rect 5259 38947 5301 38956
rect 4876 38912 4916 38921
rect 4780 38872 4876 38912
rect 4395 38324 4437 38333
rect 4395 38284 4396 38324
rect 4436 38284 4437 38324
rect 4395 38275 4437 38284
rect 3723 38240 3765 38249
rect 3723 38200 3724 38240
rect 3764 38200 3765 38240
rect 3723 38191 3765 38200
rect 3724 38106 3764 38191
rect 3688 37820 4056 37829
rect 3728 37780 3770 37820
rect 3810 37780 3852 37820
rect 3892 37780 3934 37820
rect 3974 37780 4016 37820
rect 3688 37771 4056 37780
rect 3532 37696 3651 37736
rect 3244 37612 3380 37652
rect 3611 37652 3651 37696
rect 3611 37612 3668 37652
rect 3244 36065 3284 37612
rect 3531 37568 3573 37577
rect 3531 37528 3532 37568
rect 3572 37528 3573 37568
rect 3531 37519 3573 37528
rect 3436 37400 3476 37409
rect 3532 37400 3572 37519
rect 3628 37409 3668 37612
rect 3964 37409 4004 37418
rect 3476 37360 3572 37400
rect 3627 37400 3669 37409
rect 3627 37360 3628 37400
rect 3668 37360 3669 37400
rect 4300 37400 4340 37409
rect 4004 37369 4244 37400
rect 3964 37360 4244 37369
rect 3436 37351 3476 37360
rect 3627 37351 3669 37360
rect 3628 36569 3668 37351
rect 4107 37232 4149 37241
rect 4107 37192 4108 37232
rect 4148 37192 4149 37232
rect 4107 37183 4149 37192
rect 4108 37098 4148 37183
rect 4204 36896 4244 37360
rect 4300 37325 4340 37360
rect 4299 37316 4341 37325
rect 4299 37276 4300 37316
rect 4340 37276 4341 37316
rect 4299 37267 4341 37276
rect 4300 37157 4340 37267
rect 4299 37148 4341 37157
rect 4299 37108 4300 37148
rect 4340 37108 4341 37148
rect 4299 37099 4341 37108
rect 4300 36896 4340 36905
rect 4204 36856 4300 36896
rect 4300 36847 4340 36856
rect 4108 36728 4148 36739
rect 4396 36728 4436 38275
rect 4780 38165 4820 38872
rect 4876 38863 4916 38872
rect 5260 38912 5300 38947
rect 5260 38861 5300 38872
rect 5068 38744 5108 38753
rect 5108 38704 5492 38744
rect 5068 38695 5108 38704
rect 4928 38576 5296 38585
rect 4968 38536 5010 38576
rect 5050 38536 5092 38576
rect 5132 38536 5174 38576
rect 5214 38536 5256 38576
rect 4928 38527 5296 38536
rect 5163 38324 5205 38333
rect 5163 38284 5164 38324
rect 5204 38284 5205 38324
rect 5163 38275 5205 38284
rect 4972 38240 5012 38251
rect 4972 38165 5012 38200
rect 5164 38190 5204 38275
rect 5452 38240 5492 38704
rect 5452 38191 5492 38200
rect 5547 38240 5589 38249
rect 5547 38200 5548 38240
rect 5588 38200 5589 38240
rect 5547 38191 5589 38200
rect 4779 38156 4821 38165
rect 4779 38116 4780 38156
rect 4820 38116 4821 38156
rect 4779 38107 4821 38116
rect 4971 38156 5013 38165
rect 4971 38116 4972 38156
rect 5012 38116 5013 38156
rect 4971 38107 5013 38116
rect 5548 38106 5588 38191
rect 5644 37988 5684 43576
rect 6220 43448 6260 43987
rect 6220 43399 6260 43408
rect 6700 42869 6740 42954
rect 6699 42860 6741 42869
rect 6699 42820 6700 42860
rect 6740 42820 6741 42860
rect 6699 42811 6741 42820
rect 6027 42776 6069 42785
rect 6027 42736 6028 42776
rect 6068 42736 6069 42776
rect 6027 42727 6069 42736
rect 6556 42734 6596 42743
rect 6028 42642 6068 42727
rect 6556 42692 6596 42694
rect 6556 42652 6740 42692
rect 5739 42524 5781 42533
rect 5739 42484 5740 42524
rect 5780 42484 5781 42524
rect 5739 42475 5781 42484
rect 5740 40097 5780 42475
rect 6603 42440 6645 42449
rect 6603 42400 6604 42440
rect 6644 42400 6645 42440
rect 6603 42391 6645 42400
rect 6027 42356 6069 42365
rect 6027 42316 6028 42356
rect 6068 42316 6069 42356
rect 6027 42307 6069 42316
rect 5835 41180 5877 41189
rect 5835 41140 5836 41180
rect 5876 41140 5877 41180
rect 5835 41131 5877 41140
rect 5932 41180 5972 41189
rect 5836 41046 5876 41131
rect 5932 40937 5972 41140
rect 5931 40928 5973 40937
rect 5931 40888 5932 40928
rect 5972 40888 5973 40928
rect 5931 40879 5973 40888
rect 5931 40592 5973 40601
rect 5931 40552 5932 40592
rect 5972 40552 5973 40592
rect 5931 40543 5973 40552
rect 5932 40424 5972 40543
rect 5932 40375 5972 40384
rect 5739 40088 5781 40097
rect 5739 40048 5740 40088
rect 5780 40048 5781 40088
rect 5739 40039 5781 40048
rect 5739 39920 5781 39929
rect 5739 39880 5740 39920
rect 5780 39880 5781 39920
rect 5739 39871 5781 39880
rect 5548 37948 5684 37988
rect 5548 37820 5588 37948
rect 5740 37820 5780 39871
rect 5932 39752 5972 39761
rect 5932 38921 5972 39712
rect 6028 39005 6068 42307
rect 6508 41936 6548 41945
rect 6411 41264 6453 41273
rect 6411 41224 6412 41264
rect 6452 41224 6453 41264
rect 6411 41215 6453 41224
rect 6412 41130 6452 41215
rect 6508 40769 6548 41896
rect 6507 40760 6549 40769
rect 6507 40720 6508 40760
rect 6548 40720 6549 40760
rect 6507 40711 6549 40720
rect 6604 40517 6644 42391
rect 6700 42188 6740 42652
rect 6700 42139 6740 42148
rect 6603 40508 6645 40517
rect 6603 40468 6604 40508
rect 6644 40468 6645 40508
rect 6603 40459 6645 40468
rect 6796 40181 6836 46432
rect 7083 46304 7125 46313
rect 7083 46264 7084 46304
rect 7124 46264 7125 46304
rect 7083 46255 7125 46264
rect 6987 45380 7029 45389
rect 6987 45340 6988 45380
rect 7028 45340 7029 45380
rect 6987 45331 7029 45340
rect 6988 42869 7028 45331
rect 7084 44283 7124 46255
rect 7276 45893 7316 49111
rect 7372 49085 7412 50800
rect 7468 49496 7508 51724
rect 7756 51269 7796 55075
rect 7947 54872 7989 54881
rect 7947 54832 7948 54872
rect 7988 54832 7989 54872
rect 7947 54823 7989 54832
rect 7948 54738 7988 54823
rect 8044 54200 8084 55504
rect 7852 54160 8084 54200
rect 7852 53276 7892 54160
rect 7947 54032 7989 54041
rect 8236 54032 8276 56344
rect 8332 55628 8372 57016
rect 8523 57016 8524 57056
rect 8564 57016 8565 57056
rect 8716 57021 8756 57030
rect 8523 57007 8565 57016
rect 8427 56720 8469 56729
rect 8427 56680 8428 56720
rect 8468 56680 8469 56720
rect 8427 56671 8469 56680
rect 8428 56216 8468 56671
rect 8524 56384 8564 57007
rect 8524 56335 8564 56344
rect 8428 56176 8564 56216
rect 8428 55628 8468 55637
rect 8332 55588 8428 55628
rect 8331 54116 8373 54125
rect 8331 54076 8332 54116
rect 8372 54076 8373 54116
rect 8331 54067 8373 54076
rect 7947 53992 7948 54032
rect 7988 53992 7989 54032
rect 7947 53983 7989 53992
rect 8044 53992 8276 54032
rect 8332 54032 8372 54067
rect 7948 53898 7988 53983
rect 8044 53696 8084 53992
rect 8332 53981 8372 53992
rect 8428 53948 8468 55588
rect 8524 55628 8564 56176
rect 8524 55217 8564 55588
rect 8523 55208 8565 55217
rect 8523 55168 8524 55208
rect 8564 55168 8565 55208
rect 8523 55159 8565 55168
rect 8812 54452 8852 57679
rect 8907 56972 8949 56981
rect 8907 56932 8908 56972
rect 8948 56932 8949 56972
rect 8907 56923 8949 56932
rect 8908 56838 8948 56923
rect 9100 56720 9140 59863
rect 9292 59669 9332 60040
rect 9291 59660 9333 59669
rect 9291 59620 9292 59660
rect 9332 59620 9333 59660
rect 9291 59611 9333 59620
rect 9388 59492 9428 61048
rect 9484 59576 9524 61123
rect 9676 60920 9716 61384
rect 9579 60836 9621 60845
rect 9579 60796 9580 60836
rect 9620 60796 9621 60836
rect 9579 60787 9621 60796
rect 9580 60164 9620 60787
rect 9676 60584 9716 60880
rect 9771 60836 9813 60845
rect 9771 60796 9772 60836
rect 9812 60796 9813 60836
rect 9771 60787 9813 60796
rect 9772 60702 9812 60787
rect 9676 60544 9812 60584
rect 9676 60164 9716 60173
rect 9580 60124 9676 60164
rect 9676 60115 9716 60124
rect 9772 60164 9812 60544
rect 9867 60416 9909 60425
rect 9867 60376 9868 60416
rect 9908 60376 9909 60416
rect 9867 60367 9909 60376
rect 9772 60115 9812 60124
rect 9868 59585 9908 60367
rect 9867 59576 9909 59585
rect 9484 59536 9620 59576
rect 9292 59452 9428 59492
rect 9195 57896 9237 57905
rect 9195 57856 9196 57896
rect 9236 57856 9237 57896
rect 9195 57847 9237 57856
rect 8716 54412 8852 54452
rect 8908 56680 9140 56720
rect 8908 55544 8948 56680
rect 9196 56636 9236 57847
rect 9292 56981 9332 59452
rect 9483 59408 9525 59417
rect 9483 59368 9484 59408
rect 9524 59368 9525 59408
rect 9483 59359 9525 59368
rect 9484 59274 9524 59359
rect 9580 57905 9620 59536
rect 9867 59536 9868 59576
rect 9908 59536 9909 59576
rect 9867 59527 9909 59536
rect 9771 58316 9813 58325
rect 9771 58276 9772 58316
rect 9812 58276 9813 58316
rect 9771 58267 9813 58276
rect 9484 57896 9524 57905
rect 9388 57856 9484 57896
rect 9291 56972 9333 56981
rect 9291 56932 9292 56972
rect 9332 56932 9333 56972
rect 9291 56923 9333 56932
rect 9100 56596 9236 56636
rect 9003 56468 9045 56477
rect 9003 56428 9004 56468
rect 9044 56428 9045 56468
rect 9003 56419 9045 56428
rect 9004 56379 9044 56419
rect 9004 56330 9044 56339
rect 9004 55544 9044 55572
rect 8908 55504 9004 55544
rect 8428 53908 8660 53948
rect 8140 53864 8180 53873
rect 8180 53824 8468 53864
rect 8140 53815 8180 53824
rect 8044 53656 8180 53696
rect 8044 53276 8084 53285
rect 7852 53236 8044 53276
rect 8044 52949 8084 53236
rect 8140 53276 8180 53656
rect 8043 52940 8085 52949
rect 8043 52900 8044 52940
rect 8084 52900 8085 52940
rect 8043 52891 8085 52900
rect 8140 52613 8180 53236
rect 8139 52604 8181 52613
rect 8139 52564 8140 52604
rect 8180 52564 8181 52604
rect 8139 52555 8181 52564
rect 8428 52534 8468 53824
rect 8620 53360 8660 53908
rect 8716 53537 8756 54412
rect 8908 54368 8948 55504
rect 9004 55495 9044 55504
rect 8812 54328 8948 54368
rect 8715 53528 8757 53537
rect 8715 53488 8716 53528
rect 8756 53488 8757 53528
rect 8715 53479 8757 53488
rect 7851 52520 7893 52529
rect 7851 52480 7852 52520
rect 7892 52480 7893 52520
rect 7851 52471 7893 52480
rect 7948 52520 7988 52529
rect 8428 52485 8468 52494
rect 8524 53320 8620 53360
rect 7755 51260 7797 51269
rect 7755 51220 7756 51260
rect 7796 51220 7797 51260
rect 7755 51211 7797 51220
rect 7564 51008 7604 51017
rect 7564 50597 7604 50968
rect 7660 51008 7700 51017
rect 7660 50681 7700 50968
rect 7659 50672 7701 50681
rect 7659 50632 7660 50672
rect 7700 50632 7701 50672
rect 7659 50623 7701 50632
rect 7563 50588 7605 50597
rect 7563 50548 7564 50588
rect 7604 50548 7605 50588
rect 7563 50539 7605 50548
rect 7563 50336 7605 50345
rect 7563 50296 7564 50336
rect 7604 50296 7605 50336
rect 7563 50287 7605 50296
rect 7564 50202 7604 50287
rect 7468 49447 7508 49456
rect 7371 49076 7413 49085
rect 7371 49036 7372 49076
rect 7412 49036 7413 49076
rect 7371 49027 7413 49036
rect 7755 48992 7797 49001
rect 7755 48952 7756 48992
rect 7796 48952 7797 48992
rect 7755 48943 7797 48952
rect 7756 47900 7796 48943
rect 7756 47851 7796 47860
rect 7852 46640 7892 52471
rect 7948 52436 7988 52480
rect 8524 52436 8564 53320
rect 8620 53311 8660 53320
rect 8619 53108 8661 53117
rect 8619 53068 8620 53108
rect 8660 53068 8661 53108
rect 8619 53059 8661 53068
rect 7948 52396 8564 52436
rect 8620 52436 8660 53059
rect 8620 52387 8660 52396
rect 8523 52268 8565 52277
rect 8523 52228 8524 52268
rect 8564 52228 8565 52268
rect 8523 52219 8565 52228
rect 8043 51764 8085 51773
rect 8043 51724 8044 51764
rect 8084 51724 8085 51764
rect 8043 51715 8085 51724
rect 8044 51092 8084 51715
rect 8331 51680 8373 51689
rect 8331 51640 8332 51680
rect 8372 51640 8373 51680
rect 8331 51631 8373 51640
rect 7947 49076 7989 49085
rect 7947 49036 7948 49076
rect 7988 49036 7989 49076
rect 7947 49027 7989 49036
rect 7948 48824 7988 49027
rect 8044 48992 8084 51052
rect 8139 51008 8181 51017
rect 8139 50968 8140 51008
rect 8180 50968 8181 51008
rect 8139 50959 8181 50968
rect 8140 50874 8180 50959
rect 8044 48952 8180 48992
rect 8044 48824 8084 48833
rect 7948 48784 8044 48824
rect 7948 47989 7988 47998
rect 7948 47480 7988 47949
rect 8044 47816 8084 48784
rect 8140 48329 8180 48952
rect 8236 48572 8276 48581
rect 8139 48320 8181 48329
rect 8139 48280 8140 48320
rect 8180 48280 8181 48320
rect 8139 48271 8181 48280
rect 8140 48161 8180 48271
rect 8139 48152 8181 48161
rect 8139 48112 8140 48152
rect 8180 48112 8181 48152
rect 8139 48103 8181 48112
rect 8236 47993 8276 48532
rect 8235 47984 8277 47993
rect 8235 47944 8236 47984
rect 8276 47944 8277 47984
rect 8235 47935 8277 47944
rect 8044 47776 8276 47816
rect 8044 47480 8084 47489
rect 7948 47440 8044 47480
rect 8044 47431 8084 47440
rect 8236 47312 8276 47776
rect 8236 47263 8276 47272
rect 7852 46600 8084 46640
rect 7467 46556 7509 46565
rect 7467 46516 7468 46556
rect 7508 46516 7509 46556
rect 7467 46507 7509 46516
rect 7372 46472 7412 46481
rect 7372 46229 7412 46432
rect 7371 46220 7413 46229
rect 7371 46180 7372 46220
rect 7412 46180 7413 46220
rect 7371 46171 7413 46180
rect 7275 45884 7317 45893
rect 7275 45844 7276 45884
rect 7316 45844 7317 45884
rect 7275 45835 7317 45844
rect 7179 45548 7221 45557
rect 7179 45508 7180 45548
rect 7220 45508 7221 45548
rect 7179 45499 7221 45508
rect 7180 44974 7220 45499
rect 7276 45389 7316 45835
rect 7275 45380 7317 45389
rect 7275 45340 7276 45380
rect 7316 45340 7317 45380
rect 7275 45331 7317 45340
rect 7371 45212 7413 45221
rect 7371 45172 7372 45212
rect 7412 45172 7413 45212
rect 7371 45163 7413 45172
rect 7275 45044 7317 45053
rect 7275 45004 7276 45044
rect 7316 45004 7317 45044
rect 7275 44995 7317 45004
rect 7180 44925 7220 44934
rect 7276 44456 7316 44995
rect 7372 44876 7412 45163
rect 7372 44827 7412 44836
rect 7468 44708 7508 46507
rect 7563 46304 7605 46313
rect 7563 46264 7564 46304
rect 7604 46264 7605 46304
rect 7563 46255 7605 46264
rect 7564 46170 7604 46255
rect 7563 45800 7605 45809
rect 7563 45760 7564 45800
rect 7604 45760 7605 45800
rect 7563 45751 7605 45760
rect 7564 44969 7604 45751
rect 7755 45548 7797 45557
rect 7755 45508 7756 45548
rect 7796 45508 7797 45548
rect 7755 45499 7797 45508
rect 7756 45414 7796 45499
rect 7947 45044 7989 45053
rect 7947 45004 7948 45044
rect 7988 45004 7989 45044
rect 7947 44995 7989 45004
rect 7563 44960 7605 44969
rect 7563 44920 7564 44960
rect 7604 44920 7605 44960
rect 7563 44911 7605 44920
rect 7948 44960 7988 44995
rect 7948 44909 7988 44920
rect 7276 44407 7316 44416
rect 7372 44668 7508 44708
rect 7084 44234 7124 44243
rect 7372 43280 7412 44668
rect 7467 44204 7509 44213
rect 7467 44164 7468 44204
rect 7508 44164 7509 44204
rect 7467 44155 7509 44164
rect 7468 43541 7508 44155
rect 7467 43532 7509 43541
rect 7467 43492 7468 43532
rect 7508 43492 7509 43532
rect 7467 43483 7509 43492
rect 7468 43448 7508 43483
rect 7468 43397 7508 43408
rect 7948 43448 7988 43457
rect 7660 43364 7700 43373
rect 7948 43364 7988 43408
rect 7700 43324 7988 43364
rect 8044 43448 8084 46600
rect 8139 46472 8181 46481
rect 8139 46432 8140 46472
rect 8180 46432 8181 46472
rect 8139 46423 8181 46432
rect 8140 46338 8180 46423
rect 7660 43315 7700 43324
rect 7372 43240 7508 43280
rect 6987 42860 7029 42869
rect 6987 42820 6988 42860
rect 7028 42820 7029 42860
rect 6987 42811 7029 42820
rect 6988 41476 7412 41516
rect 6988 41264 7028 41476
rect 6940 41254 7028 41264
rect 6980 41224 7028 41254
rect 7084 41348 7124 41357
rect 6940 41205 6980 41214
rect 6987 40508 7029 40517
rect 6987 40468 6988 40508
rect 7028 40468 7029 40508
rect 6987 40459 7029 40468
rect 6795 40172 6837 40181
rect 6795 40132 6796 40172
rect 6836 40132 6837 40172
rect 6795 40123 6837 40132
rect 6124 39752 6164 39763
rect 6220 39761 6260 39846
rect 6124 39677 6164 39712
rect 6219 39752 6261 39761
rect 6219 39712 6220 39752
rect 6260 39712 6261 39752
rect 6219 39703 6261 39712
rect 6412 39752 6452 39761
rect 6123 39668 6165 39677
rect 6412 39668 6452 39712
rect 6123 39628 6124 39668
rect 6164 39628 6165 39668
rect 6123 39619 6165 39628
rect 6316 39628 6452 39668
rect 6508 39752 6548 39761
rect 6220 39584 6260 39593
rect 6316 39584 6356 39628
rect 6508 39593 6548 39712
rect 6699 39752 6741 39761
rect 6699 39712 6700 39752
rect 6740 39712 6741 39752
rect 6699 39703 6741 39712
rect 6796 39752 6836 39761
rect 6260 39544 6356 39584
rect 6507 39584 6549 39593
rect 6507 39544 6508 39584
rect 6548 39544 6549 39584
rect 6220 39535 6260 39544
rect 6507 39535 6549 39544
rect 6412 39500 6452 39509
rect 6027 38996 6069 39005
rect 6027 38956 6028 38996
rect 6068 38956 6260 38996
rect 6027 38947 6069 38956
rect 5931 38912 5973 38921
rect 5931 38872 5932 38912
rect 5972 38872 5973 38912
rect 5931 38863 5973 38872
rect 6123 38240 6165 38249
rect 6123 38200 6124 38240
rect 6164 38200 6165 38240
rect 6123 38191 6165 38200
rect 5356 37780 5588 37820
rect 5644 37780 5780 37820
rect 5932 38156 5972 38165
rect 4928 37064 5296 37073
rect 4968 37024 5010 37064
rect 5050 37024 5092 37064
rect 5132 37024 5174 37064
rect 5214 37024 5256 37064
rect 4928 37015 5296 37024
rect 4588 36856 5012 36896
rect 4108 36653 4148 36688
rect 4204 36688 4436 36728
rect 4492 36728 4532 36737
rect 4107 36644 4149 36653
rect 4107 36604 4108 36644
rect 4148 36604 4149 36644
rect 4107 36595 4149 36604
rect 3627 36560 3669 36569
rect 3627 36520 3628 36560
rect 3668 36520 3669 36560
rect 3627 36511 3669 36520
rect 3688 36308 4056 36317
rect 3728 36268 3770 36308
rect 3810 36268 3852 36308
rect 3892 36268 3934 36308
rect 3974 36268 4016 36308
rect 3688 36259 4056 36268
rect 3243 36056 3285 36065
rect 3243 36016 3244 36056
rect 3284 36016 3285 36056
rect 3243 36007 3285 36016
rect 4107 35888 4149 35897
rect 4107 35848 4108 35888
rect 4148 35848 4149 35888
rect 4107 35839 4149 35848
rect 4108 35754 4148 35839
rect 4107 35300 4149 35309
rect 4107 35260 4108 35300
rect 4148 35260 4149 35300
rect 4107 35251 4149 35260
rect 3244 35216 3284 35225
rect 3724 35216 3764 35225
rect 3284 35176 3380 35216
rect 3244 35167 3284 35176
rect 3340 35048 3380 35176
rect 3724 35057 3764 35176
rect 3820 35216 3860 35227
rect 3820 35141 3860 35176
rect 4108 35216 4148 35251
rect 4108 35165 4148 35176
rect 3819 35132 3861 35141
rect 3819 35092 3820 35132
rect 3860 35092 3861 35132
rect 3819 35083 3861 35092
rect 3436 35048 3476 35057
rect 3340 35008 3436 35048
rect 3436 34999 3476 35008
rect 3723 35048 3765 35057
rect 3723 35008 3724 35048
rect 3764 35008 3765 35048
rect 3723 34999 3765 35008
rect 3243 34964 3285 34973
rect 3243 34924 3244 34964
rect 3284 34924 3285 34964
rect 3243 34915 3285 34924
rect 3531 34964 3573 34973
rect 3531 34924 3532 34964
rect 3572 34924 3573 34964
rect 3531 34915 3573 34924
rect 4107 34964 4149 34973
rect 4107 34924 4108 34964
rect 4148 34924 4149 34964
rect 4107 34915 4149 34924
rect 3244 34830 3284 34915
rect 2956 34420 3188 34460
rect 2956 34301 2996 34420
rect 3244 34376 3284 34385
rect 3052 34336 3244 34376
rect 2955 34292 2997 34301
rect 2955 34252 2956 34292
rect 2996 34252 2997 34292
rect 2955 34243 2997 34252
rect 2859 33872 2901 33881
rect 2859 33832 2860 33872
rect 2900 33832 2901 33872
rect 2859 33823 2901 33832
rect 2955 33704 2997 33713
rect 2955 33664 2956 33704
rect 2996 33664 2997 33704
rect 2955 33655 2997 33664
rect 2956 33570 2996 33655
rect 2764 33160 2996 33200
rect 2763 32864 2805 32873
rect 2668 32844 2708 32853
rect 2476 32804 2668 32844
rect 2763 32824 2764 32864
rect 2804 32824 2805 32864
rect 2763 32815 2805 32824
rect 2283 32696 2325 32705
rect 2283 32656 2284 32696
rect 2324 32656 2325 32696
rect 2283 32647 2325 32656
rect 2284 31268 2324 32647
rect 2476 32360 2516 32804
rect 2668 32795 2708 32804
rect 2764 32730 2804 32815
rect 2859 32780 2901 32789
rect 2859 32740 2860 32780
rect 2900 32740 2901 32780
rect 2859 32731 2901 32740
rect 2476 32320 2612 32360
rect 2476 32192 2516 32201
rect 2476 31865 2516 32152
rect 2475 31856 2517 31865
rect 2475 31816 2476 31856
rect 2516 31816 2517 31856
rect 2475 31807 2517 31816
rect 2379 31436 2421 31445
rect 2379 31396 2380 31436
rect 2420 31396 2516 31436
rect 2379 31387 2421 31396
rect 2476 31352 2516 31396
rect 2284 31228 2420 31268
rect 2188 30808 2324 30848
rect 2091 30799 2133 30808
rect 1900 30680 1940 30689
rect 1900 29840 1940 30640
rect 2092 30680 2132 30689
rect 1995 30596 2037 30605
rect 1995 30556 1996 30596
rect 2036 30556 2037 30596
rect 1995 30547 2037 30556
rect 1996 30344 2036 30547
rect 2092 30521 2132 30640
rect 2187 30680 2229 30689
rect 2187 30640 2188 30680
rect 2228 30640 2229 30680
rect 2187 30631 2229 30640
rect 2188 30546 2228 30631
rect 2091 30512 2133 30521
rect 2091 30472 2092 30512
rect 2132 30472 2133 30512
rect 2091 30463 2133 30472
rect 1996 30304 2132 30344
rect 1900 29800 2036 29840
rect 1900 29336 1940 29345
rect 1900 29177 1940 29296
rect 1899 29168 1941 29177
rect 1899 29128 1900 29168
rect 1940 29128 1941 29168
rect 1899 29119 1941 29128
rect 1996 28673 2036 29800
rect 2092 29765 2132 30304
rect 2187 30176 2229 30185
rect 2187 30136 2188 30176
rect 2228 30136 2229 30176
rect 2187 30127 2229 30136
rect 2091 29756 2133 29765
rect 2091 29716 2092 29756
rect 2132 29716 2133 29756
rect 2091 29707 2133 29716
rect 2091 29252 2133 29261
rect 2091 29212 2092 29252
rect 2132 29212 2133 29252
rect 2091 29203 2133 29212
rect 2092 29084 2132 29203
rect 2092 29035 2132 29044
rect 1995 28664 2037 28673
rect 1995 28624 1996 28664
rect 2036 28624 2037 28664
rect 1995 28615 2037 28624
rect 1804 28540 1940 28580
rect 1900 28496 1940 28540
rect 1708 28456 1844 28496
rect 1900 28456 2132 28496
rect 1707 28328 1749 28337
rect 1612 28288 1708 28328
rect 1748 28288 1749 28328
rect 1804 28328 1844 28456
rect 1804 28288 2036 28328
rect 1707 28279 1749 28288
rect 1323 28244 1365 28253
rect 1228 28204 1324 28244
rect 1364 28204 1365 28244
rect 1323 28195 1365 28204
rect 1323 27740 1365 27749
rect 1228 27700 1324 27740
rect 1364 27700 1365 27740
rect 1228 27656 1268 27700
rect 1323 27691 1365 27700
rect 1228 27607 1268 27616
rect 1420 26816 1460 26825
rect 1131 26648 1173 26657
rect 1131 26608 1132 26648
rect 1172 26608 1173 26648
rect 1131 26599 1173 26608
rect 1035 26060 1077 26069
rect 1035 26020 1036 26060
rect 1076 26020 1077 26060
rect 1035 26011 1077 26020
rect 1035 23456 1077 23465
rect 1035 23416 1036 23456
rect 1076 23416 1077 23456
rect 1035 23407 1077 23416
rect 939 2876 981 2885
rect 939 2836 940 2876
rect 980 2836 981 2876
rect 939 2827 981 2836
rect 1036 1289 1076 23407
rect 1035 1280 1077 1289
rect 1035 1240 1036 1280
rect 1076 1240 1077 1280
rect 1035 1231 1077 1240
rect 1132 1205 1172 26599
rect 1420 25976 1460 26776
rect 1516 26816 1556 26825
rect 1556 26776 1652 26816
rect 1516 26767 1556 26776
rect 1515 26144 1557 26153
rect 1515 26104 1516 26144
rect 1556 26104 1557 26144
rect 1515 26095 1557 26104
rect 1516 26010 1556 26095
rect 1228 25936 1460 25976
rect 1228 25724 1268 25936
rect 1515 25724 1557 25733
rect 1228 25684 1364 25724
rect 1324 25136 1364 25684
rect 1515 25684 1516 25724
rect 1556 25684 1557 25724
rect 1515 25675 1557 25684
rect 1324 25096 1460 25136
rect 1323 24968 1365 24977
rect 1323 24928 1324 24968
rect 1364 24928 1365 24968
rect 1323 24919 1365 24928
rect 1324 24632 1364 24919
rect 1324 24557 1364 24592
rect 1323 24548 1365 24557
rect 1323 24508 1324 24548
rect 1364 24508 1365 24548
rect 1323 24499 1365 24508
rect 1420 24128 1460 25096
rect 1324 24088 1460 24128
rect 1228 24044 1268 24053
rect 1324 24044 1364 24088
rect 1268 24004 1364 24044
rect 1228 23995 1268 24004
rect 1419 23792 1461 23801
rect 1419 23752 1420 23792
rect 1460 23752 1461 23792
rect 1419 23743 1461 23752
rect 1323 23708 1365 23717
rect 1323 23668 1324 23708
rect 1364 23668 1365 23708
rect 1323 23659 1365 23668
rect 1228 22280 1268 22289
rect 1324 22280 1364 23659
rect 1420 23658 1460 23743
rect 1420 23120 1460 23129
rect 1420 22877 1460 23080
rect 1419 22868 1461 22877
rect 1419 22828 1420 22868
rect 1460 22828 1461 22868
rect 1419 22819 1461 22828
rect 1268 22240 1364 22280
rect 1228 22231 1268 22240
rect 1324 20525 1364 22240
rect 1516 21272 1556 25675
rect 1420 21232 1556 21272
rect 1323 20516 1365 20525
rect 1323 20476 1324 20516
rect 1364 20476 1365 20516
rect 1323 20467 1365 20476
rect 1323 19760 1365 19769
rect 1323 19720 1324 19760
rect 1364 19720 1365 19760
rect 1323 19711 1365 19720
rect 1324 19256 1364 19711
rect 1324 19207 1364 19216
rect 1228 18584 1268 18593
rect 1420 18584 1460 21232
rect 1515 20768 1557 20777
rect 1515 20728 1516 20768
rect 1556 20728 1557 20768
rect 1515 20719 1557 20728
rect 1612 20768 1652 26776
rect 1708 24137 1748 28279
rect 1803 27488 1845 27497
rect 1803 27448 1804 27488
rect 1844 27448 1845 27488
rect 1803 27439 1845 27448
rect 1804 24977 1844 27439
rect 1996 26900 2036 28288
rect 1996 26851 2036 26860
rect 1900 26816 1940 26825
rect 1803 24968 1845 24977
rect 1803 24928 1804 24968
rect 1844 24928 1845 24968
rect 1803 24919 1845 24928
rect 1803 24800 1845 24809
rect 1803 24760 1804 24800
rect 1844 24760 1845 24800
rect 1803 24751 1845 24760
rect 1707 24128 1749 24137
rect 1707 24088 1708 24128
rect 1748 24088 1749 24128
rect 1707 24079 1749 24088
rect 1707 23540 1749 23549
rect 1707 23500 1708 23540
rect 1748 23500 1749 23540
rect 1707 23491 1749 23500
rect 1708 23120 1748 23491
rect 1708 23071 1748 23080
rect 1708 22868 1748 22877
rect 1708 22205 1748 22828
rect 1707 22196 1749 22205
rect 1707 22156 1708 22196
rect 1748 22156 1749 22196
rect 1707 22147 1749 22156
rect 1707 21608 1749 21617
rect 1707 21568 1708 21608
rect 1748 21568 1749 21608
rect 1707 21559 1749 21568
rect 1516 20634 1556 20719
rect 1612 19937 1652 20728
rect 1611 19928 1653 19937
rect 1611 19888 1612 19928
rect 1652 19888 1653 19928
rect 1611 19879 1653 19888
rect 1708 19853 1748 21559
rect 1707 19844 1749 19853
rect 1707 19804 1708 19844
rect 1748 19804 1749 19844
rect 1707 19795 1749 19804
rect 1804 19769 1844 24751
rect 1900 22625 1940 26776
rect 1995 25640 2037 25649
rect 1995 25600 1996 25640
rect 2036 25600 2037 25640
rect 1995 25591 2037 25600
rect 1996 23381 2036 25591
rect 2092 23960 2132 28456
rect 2188 26153 2228 30127
rect 2284 29168 2324 30808
rect 2380 30680 2420 31228
rect 2476 31109 2516 31312
rect 2475 31100 2517 31109
rect 2475 31060 2476 31100
rect 2516 31060 2517 31100
rect 2475 31051 2517 31060
rect 2380 30631 2420 30640
rect 2475 30512 2517 30521
rect 2475 30472 2476 30512
rect 2516 30472 2517 30512
rect 2475 30463 2517 30472
rect 2476 30008 2516 30463
rect 2572 30092 2612 32320
rect 2860 31529 2900 32731
rect 2667 31520 2709 31529
rect 2667 31480 2668 31520
rect 2708 31480 2709 31520
rect 2667 31471 2709 31480
rect 2859 31520 2901 31529
rect 2859 31480 2860 31520
rect 2900 31480 2901 31520
rect 2956 31520 2996 33160
rect 3052 32789 3092 34336
rect 3244 34327 3284 34336
rect 3243 34208 3285 34217
rect 3243 34168 3244 34208
rect 3284 34168 3285 34208
rect 3243 34159 3285 34168
rect 3147 33956 3189 33965
rect 3147 33916 3148 33956
rect 3188 33916 3189 33956
rect 3147 33907 3189 33916
rect 3148 33872 3188 33907
rect 3148 33821 3188 33832
rect 3244 33704 3284 34159
rect 3435 33788 3477 33797
rect 3435 33748 3436 33788
rect 3476 33748 3477 33788
rect 3435 33739 3477 33748
rect 3148 33664 3284 33704
rect 3339 33704 3381 33713
rect 3339 33664 3340 33704
rect 3380 33664 3381 33704
rect 3148 32948 3188 33664
rect 3339 33655 3381 33664
rect 3148 32899 3188 32908
rect 3340 32873 3380 33655
rect 3244 32864 3284 32873
rect 3051 32780 3093 32789
rect 3051 32740 3052 32780
rect 3092 32740 3093 32780
rect 3051 32731 3093 32740
rect 3244 32705 3284 32824
rect 3339 32864 3381 32873
rect 3339 32824 3340 32864
rect 3380 32824 3381 32864
rect 3339 32815 3381 32824
rect 3243 32696 3285 32705
rect 3243 32656 3244 32696
rect 3284 32656 3285 32696
rect 3243 32647 3285 32656
rect 3244 32033 3284 32647
rect 3436 32612 3476 33739
rect 3532 33704 3572 34915
rect 3688 34796 4056 34805
rect 3728 34756 3770 34796
rect 3810 34756 3852 34796
rect 3892 34756 3934 34796
rect 3974 34756 4016 34796
rect 3688 34747 4056 34756
rect 3724 34381 3764 34390
rect 3724 33965 3764 34341
rect 3819 34376 3861 34385
rect 3819 34336 3820 34376
rect 3860 34336 3861 34376
rect 3819 34327 3861 34336
rect 4108 34376 4148 34915
rect 4204 34544 4244 36688
rect 4492 36644 4532 36688
rect 4300 36604 4532 36644
rect 4300 36140 4340 36604
rect 4492 36476 4532 36485
rect 4492 36140 4532 36436
rect 4300 36091 4340 36100
rect 4396 36100 4532 36140
rect 4300 35720 4340 35729
rect 4300 35225 4340 35680
rect 4299 35216 4341 35225
rect 4299 35176 4300 35216
rect 4340 35176 4341 35216
rect 4299 35167 4341 35176
rect 4204 34504 4340 34544
rect 4108 34327 4148 34336
rect 4203 34376 4245 34385
rect 4203 34336 4204 34376
rect 4244 34336 4245 34376
rect 4203 34327 4245 34336
rect 3723 33956 3765 33965
rect 3723 33916 3724 33956
rect 3764 33916 3765 33956
rect 3723 33907 3765 33916
rect 3532 33655 3572 33664
rect 3820 33704 3860 34327
rect 3915 34292 3957 34301
rect 3915 34252 3916 34292
rect 3956 34252 3957 34292
rect 3915 34243 3957 34252
rect 3916 34158 3956 34243
rect 4204 34242 4244 34327
rect 3820 33655 3860 33664
rect 4204 33704 4244 33713
rect 4204 33545 4244 33664
rect 4203 33536 4245 33545
rect 4203 33496 4204 33536
rect 4244 33496 4245 33536
rect 4203 33487 4245 33496
rect 3532 33452 3572 33461
rect 3532 32789 3572 33412
rect 3688 33284 4056 33293
rect 3728 33244 3770 33284
rect 3810 33244 3852 33284
rect 3892 33244 3934 33284
rect 3974 33244 4016 33284
rect 3688 33235 4056 33244
rect 4204 33041 4244 33487
rect 4203 33032 4245 33041
rect 4203 32992 4204 33032
rect 4244 32992 4245 33032
rect 4203 32983 4245 32992
rect 3724 32864 3764 32875
rect 3724 32789 3764 32824
rect 4204 32869 4244 32878
rect 3531 32780 3573 32789
rect 3531 32740 3532 32780
rect 3572 32740 3573 32780
rect 3531 32731 3573 32740
rect 3723 32780 3765 32789
rect 3723 32740 3724 32780
rect 3764 32740 3765 32780
rect 3723 32731 3765 32740
rect 3436 32572 3572 32612
rect 3243 32024 3285 32033
rect 3243 31984 3244 32024
rect 3284 31984 3285 32024
rect 3243 31975 3285 31984
rect 3051 31520 3093 31529
rect 2956 31480 3052 31520
rect 3092 31480 3093 31520
rect 2859 31471 2901 31480
rect 3051 31471 3093 31480
rect 3435 31520 3477 31529
rect 3435 31480 3436 31520
rect 3476 31480 3477 31520
rect 3435 31471 3477 31480
rect 2668 31386 2708 31471
rect 2859 31352 2901 31361
rect 2859 31312 2860 31352
rect 2900 31312 2901 31352
rect 2859 31303 2901 31312
rect 2956 31352 2996 31361
rect 2860 31218 2900 31303
rect 2956 31193 2996 31312
rect 3051 31352 3093 31361
rect 3051 31312 3052 31352
rect 3092 31312 3093 31352
rect 3051 31303 3093 31312
rect 3148 31352 3188 31361
rect 2955 31184 2997 31193
rect 2955 31144 2956 31184
rect 2996 31144 2997 31184
rect 2955 31135 2997 31144
rect 3052 31184 3092 31303
rect 3052 31135 3092 31144
rect 3148 30773 3188 31312
rect 3244 31352 3284 31361
rect 3345 31352 3385 31361
rect 3244 30941 3284 31312
rect 3340 31312 3345 31352
rect 3340 31303 3385 31312
rect 3340 31025 3380 31303
rect 3339 31016 3381 31025
rect 3339 30976 3340 31016
rect 3380 30976 3381 31016
rect 3339 30967 3381 30976
rect 3243 30932 3285 30941
rect 3243 30892 3244 30932
rect 3284 30892 3285 30932
rect 3243 30883 3285 30892
rect 2763 30764 2805 30773
rect 2763 30724 2764 30764
rect 2804 30724 2805 30764
rect 2763 30715 2805 30724
rect 3147 30764 3189 30773
rect 3147 30724 3148 30764
rect 3188 30724 3189 30764
rect 3147 30715 3189 30724
rect 2668 30092 2708 30101
rect 2572 30052 2668 30092
rect 2668 30043 2708 30052
rect 2476 29968 2612 30008
rect 2476 29840 2516 29849
rect 2380 29168 2420 29177
rect 2284 29128 2380 29168
rect 2380 29119 2420 29128
rect 2476 29009 2516 29800
rect 2283 29000 2325 29009
rect 2475 29000 2517 29009
rect 2283 28960 2284 29000
rect 2324 28960 2420 29000
rect 2283 28951 2325 28960
rect 2283 27740 2325 27749
rect 2283 27700 2284 27740
rect 2324 27700 2325 27740
rect 2283 27691 2325 27700
rect 2187 26144 2229 26153
rect 2187 26104 2188 26144
rect 2228 26104 2229 26144
rect 2187 26095 2229 26104
rect 2188 25901 2228 26095
rect 2187 25892 2229 25901
rect 2187 25852 2188 25892
rect 2228 25852 2229 25892
rect 2187 25843 2229 25852
rect 2187 25472 2229 25481
rect 2187 25432 2188 25472
rect 2228 25432 2229 25472
rect 2187 25423 2229 25432
rect 2188 25136 2228 25423
rect 2188 25087 2228 25096
rect 2284 23960 2324 27691
rect 2380 25817 2420 28960
rect 2475 28960 2476 29000
rect 2516 28960 2517 29000
rect 2475 28951 2517 28960
rect 2572 28580 2612 29968
rect 2667 29168 2709 29177
rect 2667 29128 2668 29168
rect 2708 29128 2709 29168
rect 2667 29119 2709 29128
rect 2668 29009 2708 29119
rect 2667 29000 2709 29009
rect 2667 28960 2668 29000
rect 2708 28960 2709 29000
rect 2667 28951 2709 28960
rect 2668 28580 2708 28589
rect 2572 28540 2668 28580
rect 2668 28531 2708 28540
rect 2476 28328 2516 28337
rect 2476 27656 2516 28288
rect 2571 27824 2613 27833
rect 2571 27784 2572 27824
rect 2612 27784 2613 27824
rect 2571 27775 2613 27784
rect 2476 27413 2516 27616
rect 2475 27404 2517 27413
rect 2475 27364 2476 27404
rect 2516 27364 2517 27404
rect 2475 27355 2517 27364
rect 2475 26816 2517 26825
rect 2475 26776 2476 26816
rect 2516 26776 2517 26816
rect 2475 26767 2517 26776
rect 2476 26682 2516 26767
rect 2379 25808 2421 25817
rect 2379 25768 2380 25808
rect 2420 25768 2421 25808
rect 2379 25759 2421 25768
rect 2475 25556 2517 25565
rect 2475 25516 2476 25556
rect 2516 25516 2517 25556
rect 2475 25507 2517 25516
rect 2379 25304 2421 25313
rect 2379 25264 2380 25304
rect 2420 25264 2421 25304
rect 2379 25255 2421 25264
rect 2476 25304 2516 25507
rect 2380 25170 2420 25255
rect 2476 25061 2516 25264
rect 2475 25052 2517 25061
rect 2475 25012 2476 25052
rect 2516 25012 2517 25052
rect 2475 25003 2517 25012
rect 2572 24800 2612 27775
rect 2668 27740 2708 27749
rect 2764 27740 2804 30715
rect 3051 30680 3093 30689
rect 3051 30640 3052 30680
rect 3092 30640 3093 30680
rect 3051 30631 3093 30640
rect 2955 30596 2997 30605
rect 2955 30556 2956 30596
rect 2996 30556 2997 30596
rect 2955 30547 2997 30556
rect 2859 30428 2901 30437
rect 2859 30388 2860 30428
rect 2900 30388 2901 30428
rect 2859 30379 2901 30388
rect 2860 27833 2900 30379
rect 2956 29849 2996 30547
rect 2955 29840 2997 29849
rect 2955 29800 2956 29840
rect 2996 29800 2997 29840
rect 2955 29791 2997 29800
rect 2955 29588 2997 29597
rect 2955 29548 2956 29588
rect 2996 29548 2997 29588
rect 2955 29539 2997 29548
rect 2956 29093 2996 29539
rect 2955 29084 2997 29093
rect 2955 29044 2956 29084
rect 2996 29044 2997 29084
rect 2955 29035 2997 29044
rect 2859 27824 2901 27833
rect 2859 27784 2860 27824
rect 2900 27784 2901 27824
rect 2859 27775 2901 27784
rect 2708 27700 2804 27740
rect 2668 27691 2708 27700
rect 2860 27656 2900 27665
rect 2956 27656 2996 29035
rect 2900 27616 2996 27656
rect 2860 27497 2900 27616
rect 2859 27488 2901 27497
rect 2859 27448 2860 27488
rect 2900 27448 2901 27488
rect 2859 27439 2901 27448
rect 2763 27404 2805 27413
rect 2763 27364 2764 27404
rect 2804 27364 2805 27404
rect 2763 27355 2805 27364
rect 2764 26144 2804 27355
rect 3052 26984 3092 30631
rect 3340 30521 3380 30967
rect 3339 30512 3381 30521
rect 3339 30472 3340 30512
rect 3380 30472 3381 30512
rect 3339 30463 3381 30472
rect 3436 29681 3476 31471
rect 3435 29672 3477 29681
rect 3435 29632 3436 29672
rect 3476 29632 3477 29672
rect 3435 29623 3477 29632
rect 3436 29093 3476 29623
rect 3435 29084 3477 29093
rect 3435 29044 3436 29084
rect 3476 29044 3477 29084
rect 3435 29035 3477 29044
rect 3147 28916 3189 28925
rect 3147 28876 3148 28916
rect 3188 28876 3189 28916
rect 3147 28867 3189 28876
rect 3148 28328 3188 28867
rect 3243 28412 3285 28421
rect 3243 28372 3244 28412
rect 3284 28372 3285 28412
rect 3243 28363 3285 28372
rect 3148 27488 3188 28288
rect 3244 28328 3284 28363
rect 3244 28277 3284 28288
rect 3435 28160 3477 28169
rect 3435 28120 3436 28160
rect 3476 28120 3477 28160
rect 3435 28111 3477 28120
rect 3436 28026 3476 28111
rect 3148 27448 3476 27488
rect 3052 26944 3284 26984
rect 3004 26825 3044 26834
rect 3044 26785 3092 26816
rect 3004 26776 3092 26785
rect 2955 26480 2997 26489
rect 2955 26440 2956 26480
rect 2996 26440 2997 26480
rect 2955 26431 2997 26440
rect 2956 26312 2996 26431
rect 2956 26263 2996 26272
rect 2764 26095 2804 26104
rect 2859 26144 2901 26153
rect 2859 26104 2860 26144
rect 2900 26104 2901 26144
rect 2859 26095 2901 26104
rect 2763 25556 2805 25565
rect 2763 25516 2764 25556
rect 2804 25516 2805 25556
rect 2763 25507 2805 25516
rect 2764 25304 2804 25507
rect 2860 25397 2900 26095
rect 2859 25388 2901 25397
rect 2859 25348 2860 25388
rect 2900 25348 2901 25388
rect 2859 25339 2901 25348
rect 2764 25255 2804 25264
rect 2860 25304 2900 25339
rect 2860 25254 2900 25264
rect 3052 25136 3092 26776
rect 3147 26732 3189 26741
rect 3147 26692 3148 26732
rect 3188 26692 3189 26732
rect 3147 26683 3189 26692
rect 3148 26598 3188 26683
rect 3147 26228 3189 26237
rect 3147 26188 3148 26228
rect 3188 26188 3189 26228
rect 3147 26179 3189 26188
rect 3148 25976 3188 26179
rect 3244 26153 3284 26944
rect 3436 26816 3476 27448
rect 3436 26489 3476 26776
rect 3435 26480 3477 26489
rect 3435 26440 3436 26480
rect 3476 26440 3477 26480
rect 3435 26431 3477 26440
rect 3532 26312 3572 32572
rect 3916 32360 3956 32369
rect 4204 32360 4244 32829
rect 3956 32320 4244 32360
rect 3916 32311 3956 32320
rect 3724 32192 3764 32201
rect 3724 31949 3764 32152
rect 4108 32192 4148 32201
rect 4300 32192 4340 34504
rect 4396 34385 4436 36100
rect 4588 36056 4628 36856
rect 4684 36728 4724 36737
rect 4684 36224 4724 36688
rect 4780 36728 4820 36737
rect 4780 36560 4820 36688
rect 4972 36728 5012 36856
rect 5163 36812 5205 36821
rect 5163 36772 5164 36812
rect 5204 36772 5205 36812
rect 5163 36763 5205 36772
rect 4972 36679 5012 36688
rect 5164 36728 5204 36763
rect 5164 36677 5204 36688
rect 5068 36560 5108 36569
rect 4780 36520 5068 36560
rect 5068 36511 5108 36520
rect 4684 36184 4820 36224
rect 4492 36016 4628 36056
rect 4492 35888 4532 36016
rect 4492 35393 4532 35848
rect 4588 35888 4628 35897
rect 4588 35645 4628 35848
rect 4683 35888 4725 35897
rect 4683 35848 4684 35888
rect 4724 35848 4725 35888
rect 4683 35839 4725 35848
rect 4587 35636 4629 35645
rect 4587 35596 4588 35636
rect 4628 35596 4629 35636
rect 4587 35587 4629 35596
rect 4491 35384 4533 35393
rect 4491 35344 4492 35384
rect 4532 35344 4533 35384
rect 4491 35335 4533 35344
rect 4492 35216 4532 35225
rect 4532 35176 4628 35216
rect 4492 35167 4532 35176
rect 4491 35048 4533 35057
rect 4491 35008 4492 35048
rect 4532 35008 4533 35048
rect 4491 34999 4533 35008
rect 4395 34376 4437 34385
rect 4395 34336 4396 34376
rect 4436 34336 4437 34376
rect 4395 34327 4437 34336
rect 4395 34208 4437 34217
rect 4395 34168 4396 34208
rect 4436 34168 4437 34208
rect 4395 34159 4437 34168
rect 4396 34074 4436 34159
rect 4395 32780 4437 32789
rect 4395 32740 4396 32780
rect 4436 32740 4437 32780
rect 4395 32731 4437 32740
rect 4396 32646 4436 32731
rect 4395 32360 4437 32369
rect 4395 32320 4396 32360
rect 4436 32320 4437 32360
rect 4395 32311 4437 32320
rect 4148 32152 4340 32192
rect 4108 32143 4148 32152
rect 4203 32024 4245 32033
rect 4203 31984 4204 32024
rect 4244 31984 4245 32024
rect 4203 31975 4245 31984
rect 3723 31940 3765 31949
rect 3723 31900 3724 31940
rect 3764 31900 3765 31940
rect 3723 31891 3765 31900
rect 3688 31772 4056 31781
rect 3728 31732 3770 31772
rect 3810 31732 3852 31772
rect 3892 31732 3934 31772
rect 3974 31732 4016 31772
rect 3688 31723 4056 31732
rect 3724 31445 3764 31452
rect 3723 31436 3765 31445
rect 3723 31396 3724 31436
rect 3764 31396 3769 31436
rect 3723 31387 3769 31396
rect 3729 31362 3769 31387
rect 3628 31352 3668 31361
rect 3729 31313 3769 31322
rect 3628 31268 3668 31312
rect 4204 31268 4244 31975
rect 4300 31781 4340 32152
rect 4299 31772 4341 31781
rect 4299 31732 4300 31772
rect 4340 31732 4341 31772
rect 4299 31723 4341 31732
rect 3628 31228 3764 31268
rect 4204 31228 4340 31268
rect 3627 31100 3669 31109
rect 3627 31060 3628 31100
rect 3668 31060 3669 31100
rect 3627 31051 3669 31060
rect 3628 30680 3668 31051
rect 3724 31025 3764 31228
rect 3915 31184 3957 31193
rect 3915 31144 3916 31184
rect 3956 31144 3957 31184
rect 3915 31135 3957 31144
rect 3916 31050 3956 31135
rect 3723 31016 3765 31025
rect 3723 30976 3724 31016
rect 3764 30976 3765 31016
rect 3723 30967 3765 30976
rect 3819 30848 3861 30857
rect 3819 30808 3820 30848
rect 3860 30808 3861 30848
rect 3819 30799 3861 30808
rect 3820 30714 3860 30799
rect 3628 30521 3668 30640
rect 4108 30680 4148 30689
rect 3627 30512 3669 30521
rect 3627 30472 3628 30512
rect 3668 30472 3669 30512
rect 3627 30463 3669 30472
rect 3688 30260 4056 30269
rect 3728 30220 3770 30260
rect 3810 30220 3852 30260
rect 3892 30220 3934 30260
rect 3974 30220 4016 30260
rect 3688 30211 4056 30220
rect 3627 29840 3669 29849
rect 4108 29840 4148 30640
rect 4203 30680 4245 30689
rect 4203 30640 4204 30680
rect 4244 30640 4245 30680
rect 4203 30631 4245 30640
rect 4204 30546 4244 30631
rect 3627 29800 3628 29840
rect 3668 29800 3669 29840
rect 3627 29791 3669 29800
rect 3820 29800 4148 29840
rect 4203 29840 4245 29849
rect 4203 29800 4204 29840
rect 4244 29800 4245 29840
rect 3628 29177 3668 29791
rect 3820 29336 3860 29800
rect 4203 29791 4245 29800
rect 4204 29706 4244 29791
rect 3820 29287 3860 29296
rect 3627 29168 3669 29177
rect 3627 29128 3628 29168
rect 3668 29128 3669 29168
rect 3627 29119 3669 29128
rect 4012 29168 4052 29177
rect 3628 29034 3668 29119
rect 4012 28925 4052 29128
rect 4203 29168 4245 29177
rect 4203 29128 4204 29168
rect 4244 29128 4245 29168
rect 4203 29119 4245 29128
rect 4204 29034 4244 29119
rect 4011 28916 4053 28925
rect 4011 28876 4012 28916
rect 4052 28876 4053 28916
rect 4011 28867 4053 28876
rect 4108 28916 4148 28925
rect 3688 28748 4056 28757
rect 3728 28708 3770 28748
rect 3810 28708 3852 28748
rect 3892 28708 3934 28748
rect 3974 28708 4016 28748
rect 3688 28699 4056 28708
rect 4108 28505 4148 28876
rect 3627 28496 3669 28505
rect 3627 28456 3628 28496
rect 3668 28456 3669 28496
rect 3627 28447 3669 28456
rect 4107 28496 4149 28505
rect 4107 28456 4108 28496
rect 4148 28456 4149 28496
rect 4107 28447 4149 28456
rect 3628 28328 3668 28447
rect 3628 28279 3668 28288
rect 3724 28328 3764 28337
rect 3916 28328 3956 28337
rect 3724 28169 3764 28288
rect 3820 28288 3916 28328
rect 3723 28160 3765 28169
rect 3723 28120 3724 28160
rect 3764 28120 3765 28160
rect 3723 28111 3765 28120
rect 3820 27749 3860 28288
rect 3916 28279 3956 28288
rect 4107 28328 4149 28337
rect 4107 28288 4108 28328
rect 4148 28288 4149 28328
rect 4107 28279 4149 28288
rect 4108 28194 4148 28279
rect 4300 28169 4340 31228
rect 4396 30260 4436 32311
rect 4492 32033 4532 34999
rect 4588 34889 4628 35176
rect 4587 34880 4629 34889
rect 4587 34840 4588 34880
rect 4628 34840 4629 34880
rect 4587 34831 4629 34840
rect 4684 33377 4724 35839
rect 4780 35720 4820 36184
rect 4971 35888 5013 35897
rect 4971 35848 4972 35888
rect 5012 35848 5013 35888
rect 4971 35839 5013 35848
rect 4972 35754 5012 35839
rect 4780 35671 4820 35680
rect 4928 35552 5296 35561
rect 4968 35512 5010 35552
rect 5050 35512 5092 35552
rect 5132 35512 5174 35552
rect 5214 35512 5256 35552
rect 4928 35503 5296 35512
rect 5163 35384 5205 35393
rect 5163 35344 5164 35384
rect 5204 35344 5205 35384
rect 5163 35335 5205 35344
rect 4779 35048 4821 35057
rect 4779 35008 4780 35048
rect 4820 35008 4821 35048
rect 4779 34999 4821 35008
rect 4683 33368 4725 33377
rect 4683 33328 4684 33368
rect 4724 33328 4725 33368
rect 4683 33319 4725 33328
rect 4491 32024 4533 32033
rect 4491 31984 4492 32024
rect 4532 31984 4533 32024
rect 4491 31975 4533 31984
rect 4780 31445 4820 34999
rect 5068 34385 5108 34470
rect 5067 34376 5109 34385
rect 5067 34336 5068 34376
rect 5108 34336 5109 34376
rect 5067 34327 5109 34336
rect 5164 34376 5204 35335
rect 5259 34712 5301 34721
rect 5259 34672 5260 34712
rect 5300 34672 5301 34712
rect 5259 34663 5301 34672
rect 5164 34327 5204 34336
rect 5260 34376 5300 34663
rect 5260 34327 5300 34336
rect 4972 34208 5012 34217
rect 5067 34208 5109 34217
rect 5012 34168 5068 34208
rect 5108 34168 5109 34208
rect 4972 34159 5012 34168
rect 5067 34159 5109 34168
rect 4928 34040 5296 34049
rect 4968 34000 5010 34040
rect 5050 34000 5092 34040
rect 5132 34000 5174 34040
rect 5214 34000 5256 34040
rect 4928 33991 5296 34000
rect 4928 32528 5296 32537
rect 4968 32488 5010 32528
rect 5050 32488 5092 32528
rect 5132 32488 5174 32528
rect 5214 32488 5256 32528
rect 4928 32479 5296 32488
rect 5356 32360 5396 37780
rect 5451 37484 5493 37493
rect 5451 37444 5452 37484
rect 5492 37444 5493 37484
rect 5451 37435 5493 37444
rect 5452 35393 5492 37435
rect 5548 37400 5588 37409
rect 5548 36653 5588 37360
rect 5547 36644 5589 36653
rect 5547 36604 5548 36644
rect 5588 36604 5589 36644
rect 5547 36595 5589 36604
rect 5451 35384 5493 35393
rect 5451 35344 5452 35384
rect 5492 35344 5493 35384
rect 5451 35335 5493 35344
rect 5451 35216 5493 35225
rect 5548 35216 5588 36595
rect 5451 35176 5452 35216
rect 5492 35176 5588 35216
rect 5451 35167 5493 35176
rect 5452 33704 5492 35167
rect 5644 34544 5684 37780
rect 5835 37484 5877 37493
rect 5932 37484 5972 38116
rect 6027 38156 6069 38165
rect 6027 38116 6028 38156
rect 6068 38116 6069 38156
rect 6027 38107 6069 38116
rect 6028 38022 6068 38107
rect 5835 37444 5836 37484
rect 5876 37444 5972 37484
rect 5835 37435 5877 37444
rect 6028 37400 6068 37409
rect 5932 37360 6028 37399
rect 5932 37359 6068 37360
rect 5740 37316 5780 37325
rect 5932 37316 5972 37359
rect 6028 37351 6068 37359
rect 6124 37400 6164 38191
rect 5780 37276 5972 37316
rect 5740 37267 5780 37276
rect 5836 36728 5876 36737
rect 5836 35981 5876 36688
rect 5835 35972 5877 35981
rect 5835 35932 5836 35972
rect 5876 35932 5877 35972
rect 5835 35923 5877 35932
rect 5835 35300 5877 35309
rect 5835 35260 5836 35300
rect 5876 35260 5877 35300
rect 5835 35251 5877 35260
rect 6027 35300 6069 35309
rect 6027 35260 6028 35300
rect 6068 35260 6069 35300
rect 6027 35251 6069 35260
rect 5739 35216 5781 35225
rect 5739 35176 5740 35216
rect 5780 35176 5781 35216
rect 5739 35167 5781 35176
rect 5740 35082 5780 35167
rect 5644 34504 5780 34544
rect 5547 34376 5589 34385
rect 5547 34336 5548 34376
rect 5588 34336 5589 34376
rect 5547 34327 5589 34336
rect 5644 34376 5684 34385
rect 5548 33788 5588 34327
rect 5644 33965 5684 34336
rect 5643 33956 5685 33965
rect 5643 33916 5644 33956
rect 5684 33916 5685 33956
rect 5643 33907 5685 33916
rect 5643 33788 5685 33797
rect 5548 33748 5644 33788
rect 5684 33748 5685 33788
rect 5643 33739 5685 33748
rect 5452 32780 5492 33664
rect 5644 33654 5684 33739
rect 5452 32740 5684 32780
rect 5547 32444 5589 32453
rect 5547 32404 5548 32444
rect 5588 32404 5589 32444
rect 5547 32395 5589 32404
rect 5548 32360 5588 32395
rect 5356 32320 5492 32360
rect 5356 32192 5396 32201
rect 5356 31529 5396 32152
rect 5067 31520 5109 31529
rect 5067 31480 5068 31520
rect 5108 31480 5109 31520
rect 5067 31471 5109 31480
rect 5355 31520 5397 31529
rect 5355 31480 5356 31520
rect 5396 31480 5397 31520
rect 5355 31471 5397 31480
rect 4779 31436 4821 31445
rect 4779 31396 4780 31436
rect 4820 31396 4821 31436
rect 4779 31387 4821 31396
rect 5068 31436 5108 31471
rect 4492 31352 4532 31361
rect 4492 30857 4532 31312
rect 4588 31352 4628 31361
rect 4491 30848 4533 30857
rect 4491 30808 4492 30848
rect 4532 30808 4533 30848
rect 4491 30799 4533 30808
rect 4588 30773 4628 31312
rect 4780 31268 4820 31387
rect 5068 31385 5108 31396
rect 4777 31228 4820 31268
rect 4972 31352 5012 31361
rect 4683 31184 4725 31193
rect 4683 31144 4684 31184
rect 4724 31144 4725 31184
rect 4777 31184 4817 31228
rect 4972 31193 5012 31312
rect 5355 31352 5397 31361
rect 5355 31312 5356 31352
rect 5396 31312 5397 31352
rect 5355 31303 5397 31312
rect 4971 31184 5013 31193
rect 4777 31144 4820 31184
rect 4683 31135 4725 31144
rect 4587 30764 4629 30773
rect 4587 30724 4588 30764
rect 4628 30724 4629 30764
rect 4587 30715 4629 30724
rect 4684 30680 4724 31135
rect 4588 30596 4628 30605
rect 4588 30437 4628 30556
rect 4587 30428 4629 30437
rect 4587 30388 4588 30428
rect 4628 30388 4629 30428
rect 4587 30379 4629 30388
rect 4396 30220 4628 30260
rect 4395 30092 4437 30101
rect 4395 30052 4396 30092
rect 4436 30052 4437 30092
rect 4395 30043 4437 30052
rect 4396 29958 4436 30043
rect 4588 29840 4628 30220
rect 3916 28160 3956 28169
rect 4299 28160 4341 28169
rect 3956 28120 4052 28160
rect 3916 28111 3956 28120
rect 4012 28076 4052 28120
rect 4299 28120 4300 28160
rect 4340 28120 4341 28160
rect 4299 28111 4341 28120
rect 4107 28076 4149 28085
rect 4012 28036 4108 28076
rect 4148 28036 4149 28076
rect 4107 28027 4149 28036
rect 4012 27868 4244 27908
rect 4012 27749 4052 27868
rect 3819 27740 3861 27749
rect 3819 27700 3820 27740
rect 3860 27700 3861 27740
rect 3819 27691 3861 27700
rect 4011 27740 4053 27749
rect 4011 27700 4012 27740
rect 4052 27700 4053 27740
rect 4204 27740 4244 27868
rect 4492 27824 4532 27833
rect 4300 27740 4340 27749
rect 4204 27700 4300 27740
rect 4011 27691 4053 27700
rect 4300 27691 4340 27700
rect 4108 27656 4148 27665
rect 4148 27616 4244 27656
rect 4108 27607 4148 27616
rect 4107 27488 4149 27497
rect 4107 27448 4108 27488
rect 4148 27448 4149 27488
rect 4107 27439 4149 27448
rect 3688 27236 4056 27245
rect 3728 27196 3770 27236
rect 3810 27196 3852 27236
rect 3892 27196 3934 27236
rect 3974 27196 4016 27236
rect 3688 27187 4056 27196
rect 4108 27068 4148 27439
rect 4204 27329 4244 27616
rect 4299 27488 4341 27497
rect 4299 27448 4300 27488
rect 4340 27448 4341 27488
rect 4299 27439 4341 27448
rect 4203 27320 4245 27329
rect 4203 27280 4204 27320
rect 4244 27280 4245 27320
rect 4203 27271 4245 27280
rect 4108 27019 4148 27028
rect 4204 26993 4244 27271
rect 4203 26984 4245 26993
rect 4203 26944 4204 26984
rect 4244 26944 4245 26984
rect 4203 26935 4245 26944
rect 3724 26825 3764 26910
rect 3723 26816 3765 26825
rect 3723 26776 3724 26816
rect 3764 26776 3765 26816
rect 3723 26767 3765 26776
rect 3820 26732 3860 26741
rect 3723 26648 3765 26657
rect 3820 26648 3860 26692
rect 3723 26608 3724 26648
rect 3764 26608 3860 26648
rect 3723 26599 3765 26608
rect 3436 26272 3572 26312
rect 3243 26144 3285 26153
rect 3243 26104 3244 26144
rect 3284 26104 3285 26144
rect 3243 26095 3285 26104
rect 3148 25936 3284 25976
rect 3147 25556 3189 25565
rect 3147 25516 3148 25556
rect 3188 25516 3189 25556
rect 3147 25507 3189 25516
rect 3148 25313 3188 25507
rect 3147 25304 3189 25313
rect 3147 25264 3148 25304
rect 3188 25264 3189 25304
rect 3147 25255 3189 25264
rect 3244 25304 3284 25936
rect 2764 25096 3092 25136
rect 2667 25052 2709 25061
rect 2667 25012 2668 25052
rect 2708 25012 2709 25052
rect 2667 25003 2709 25012
rect 2476 24760 2612 24800
rect 2476 24473 2516 24760
rect 2572 24632 2612 24641
rect 2668 24632 2708 25003
rect 2764 24800 2804 25096
rect 2764 24751 2804 24760
rect 2956 24800 2996 24809
rect 3148 24800 3188 25255
rect 2996 24760 3188 24800
rect 2956 24751 2996 24760
rect 3148 24632 3188 24643
rect 2668 24592 2804 24632
rect 2475 24464 2517 24473
rect 2475 24424 2476 24464
rect 2516 24424 2517 24464
rect 2475 24415 2517 24424
rect 2572 24044 2612 24592
rect 2476 24004 2612 24044
rect 2092 23920 2228 23960
rect 2284 23920 2420 23960
rect 2188 23717 2228 23920
rect 2283 23792 2325 23801
rect 2283 23752 2284 23792
rect 2324 23752 2325 23792
rect 2283 23743 2325 23752
rect 2187 23708 2229 23717
rect 2187 23668 2188 23708
rect 2228 23668 2229 23708
rect 2187 23659 2229 23668
rect 1995 23372 2037 23381
rect 1995 23332 1996 23372
rect 2036 23332 2037 23372
rect 1995 23323 2037 23332
rect 1996 23120 2036 23129
rect 1996 22877 2036 23080
rect 2092 23120 2132 23129
rect 2092 22961 2132 23080
rect 2284 22961 2324 23743
rect 2091 22952 2133 22961
rect 2091 22912 2092 22952
rect 2132 22912 2133 22952
rect 2091 22903 2133 22912
rect 2283 22952 2325 22961
rect 2283 22912 2284 22952
rect 2324 22912 2325 22952
rect 2283 22903 2325 22912
rect 1995 22868 2037 22877
rect 1995 22828 1996 22868
rect 2036 22828 2037 22868
rect 1995 22819 2037 22828
rect 1899 22616 1941 22625
rect 1899 22576 1900 22616
rect 1940 22576 1941 22616
rect 1899 22567 1941 22576
rect 1900 20852 1940 22567
rect 2092 21617 2132 22903
rect 2091 21608 2133 21617
rect 2091 21568 2092 21608
rect 2132 21568 2133 21608
rect 2091 21559 2133 21568
rect 2091 21440 2133 21449
rect 2091 21400 2092 21440
rect 2132 21400 2133 21440
rect 2091 21391 2133 21400
rect 1996 20852 2036 20861
rect 1900 20812 1996 20852
rect 1996 20803 2036 20812
rect 2092 20852 2132 21391
rect 2092 20803 2132 20812
rect 2380 20180 2420 23920
rect 2476 23801 2516 24004
rect 2667 23960 2709 23969
rect 2667 23920 2668 23960
rect 2708 23920 2709 23960
rect 2667 23911 2709 23920
rect 2571 23876 2613 23885
rect 2571 23836 2572 23876
rect 2612 23836 2613 23876
rect 2571 23827 2613 23836
rect 2475 23792 2517 23801
rect 2475 23752 2476 23792
rect 2516 23752 2517 23792
rect 2475 23743 2517 23752
rect 2475 23372 2517 23381
rect 2475 23332 2476 23372
rect 2516 23332 2517 23372
rect 2475 23323 2517 23332
rect 2476 23120 2516 23323
rect 2476 23071 2516 23080
rect 2572 23120 2612 23827
rect 2572 23071 2612 23080
rect 2668 23792 2708 23911
rect 2668 23045 2708 23752
rect 2667 23036 2709 23045
rect 2667 22996 2668 23036
rect 2708 22996 2709 23036
rect 2667 22987 2709 22996
rect 2571 22784 2613 22793
rect 2571 22744 2572 22784
rect 2612 22744 2613 22784
rect 2571 22735 2613 22744
rect 2475 22280 2517 22289
rect 2475 22240 2476 22280
rect 2516 22240 2517 22280
rect 2475 22231 2517 22240
rect 2476 22146 2516 22231
rect 2572 20768 2612 22735
rect 2668 22532 2708 22541
rect 2764 22532 2804 24592
rect 3148 24557 3188 24592
rect 3147 24548 3189 24557
rect 3147 24508 3148 24548
rect 3188 24508 3189 24548
rect 3147 24499 3189 24508
rect 3051 24464 3093 24473
rect 3051 24424 3052 24464
rect 3092 24424 3093 24464
rect 3051 24415 3093 24424
rect 2859 23792 2901 23801
rect 2859 23752 2860 23792
rect 2900 23752 2901 23792
rect 2859 23743 2901 23752
rect 2708 22492 2804 22532
rect 2860 22532 2900 23743
rect 3052 23120 3092 24415
rect 3244 24389 3284 25264
rect 3340 25304 3380 25313
rect 3243 24380 3285 24389
rect 3243 24340 3244 24380
rect 3284 24340 3285 24380
rect 3243 24331 3285 24340
rect 3340 24305 3380 25264
rect 3339 24296 3381 24305
rect 3339 24256 3340 24296
rect 3380 24256 3381 24296
rect 3339 24247 3381 24256
rect 3436 23960 3476 26272
rect 3531 26144 3573 26153
rect 3531 26104 3532 26144
rect 3572 26104 3573 26144
rect 3531 26095 3573 26104
rect 3532 26010 3572 26095
rect 3531 25892 3573 25901
rect 4300 25892 4340 27439
rect 4492 26984 4532 27784
rect 4588 27068 4628 29800
rect 4684 29345 4724 30640
rect 4683 29336 4725 29345
rect 4683 29296 4684 29336
rect 4724 29296 4725 29336
rect 4683 29287 4725 29296
rect 4780 28757 4820 31144
rect 4971 31144 4972 31184
rect 5012 31144 5013 31184
rect 4971 31135 5013 31144
rect 4928 31016 5296 31025
rect 4968 30976 5010 31016
rect 5050 30976 5092 31016
rect 5132 30976 5174 31016
rect 5214 30976 5256 31016
rect 4928 30967 5296 30976
rect 5067 30848 5109 30857
rect 5067 30808 5068 30848
rect 5108 30808 5109 30848
rect 5067 30799 5109 30808
rect 5068 30353 5108 30799
rect 5164 30680 5204 30689
rect 5356 30680 5396 31303
rect 5204 30640 5396 30680
rect 5164 30631 5204 30640
rect 5067 30344 5109 30353
rect 5067 30304 5068 30344
rect 5108 30304 5109 30344
rect 5067 30295 5109 30304
rect 5452 30269 5492 32320
rect 5548 32309 5588 32320
rect 5547 31352 5589 31361
rect 5547 31312 5548 31352
rect 5588 31312 5589 31352
rect 5547 31303 5589 31312
rect 5548 31218 5588 31303
rect 5644 31100 5684 32740
rect 5548 31060 5684 31100
rect 5451 30260 5493 30269
rect 5451 30220 5452 30260
rect 5492 30220 5493 30260
rect 5451 30211 5493 30220
rect 5548 29849 5588 31060
rect 5644 30666 5684 30675
rect 5644 30101 5684 30626
rect 5643 30092 5685 30101
rect 5643 30052 5644 30092
rect 5684 30052 5685 30092
rect 5643 30043 5685 30052
rect 5547 29840 5589 29849
rect 5547 29800 5548 29840
rect 5588 29800 5589 29840
rect 5547 29791 5589 29800
rect 5355 29756 5397 29765
rect 5355 29716 5356 29756
rect 5396 29716 5397 29756
rect 5355 29707 5397 29716
rect 4928 29504 5296 29513
rect 4968 29464 5010 29504
rect 5050 29464 5092 29504
rect 5132 29464 5174 29504
rect 5214 29464 5256 29504
rect 4928 29455 5296 29464
rect 5356 29177 5396 29707
rect 5164 29168 5204 29177
rect 5355 29168 5397 29177
rect 5204 29128 5356 29168
rect 5396 29128 5397 29168
rect 5164 29119 5204 29128
rect 5355 29119 5397 29128
rect 5356 29034 5396 29119
rect 4779 28748 4821 28757
rect 4779 28708 4780 28748
rect 4820 28708 4821 28748
rect 4779 28699 4821 28708
rect 5451 28580 5493 28589
rect 5451 28540 5452 28580
rect 5492 28540 5493 28580
rect 5451 28531 5493 28540
rect 5356 28328 5396 28339
rect 5356 28253 5396 28288
rect 5355 28244 5397 28253
rect 5355 28204 5356 28244
rect 5396 28204 5397 28244
rect 5452 28244 5492 28531
rect 5547 28496 5589 28505
rect 5547 28456 5548 28496
rect 5588 28456 5589 28496
rect 5547 28447 5589 28456
rect 5548 28362 5588 28447
rect 5452 28204 5588 28244
rect 5355 28195 5397 28204
rect 4683 28076 4725 28085
rect 4683 28036 4684 28076
rect 4724 28036 4725 28076
rect 4683 28027 4725 28036
rect 4684 27824 4724 28027
rect 4928 27992 5296 28001
rect 4968 27952 5010 27992
rect 5050 27952 5092 27992
rect 5132 27952 5174 27992
rect 5214 27952 5256 27992
rect 4928 27943 5296 27952
rect 4684 27784 5012 27824
rect 4684 27656 4724 27784
rect 4684 27607 4724 27616
rect 4779 27656 4821 27665
rect 4779 27616 4780 27656
rect 4820 27616 4821 27656
rect 4779 27607 4821 27616
rect 4972 27656 5012 27784
rect 5260 27665 5300 27750
rect 5452 27665 5492 27750
rect 4972 27607 5012 27616
rect 5259 27656 5301 27665
rect 5451 27656 5493 27665
rect 5259 27616 5260 27656
rect 5300 27616 5396 27656
rect 5259 27607 5301 27616
rect 4780 27522 4820 27607
rect 5356 27488 5396 27616
rect 5451 27616 5452 27656
rect 5492 27616 5493 27656
rect 5451 27607 5493 27616
rect 5452 27488 5492 27497
rect 5356 27448 5452 27488
rect 5452 27439 5492 27448
rect 5260 27404 5300 27413
rect 4779 27320 4821 27329
rect 4779 27280 4780 27320
rect 4820 27280 4821 27320
rect 4779 27271 4821 27280
rect 4588 27028 4724 27068
rect 4492 26944 4628 26984
rect 4491 26816 4533 26825
rect 4491 26776 4492 26816
rect 4532 26776 4533 26816
rect 4491 26767 4533 26776
rect 4492 26682 4532 26767
rect 4395 26480 4437 26489
rect 4395 26440 4396 26480
rect 4436 26440 4437 26480
rect 4395 26431 4437 26440
rect 3531 25852 3532 25892
rect 3572 25852 3573 25892
rect 3531 25843 3573 25852
rect 4108 25852 4340 25892
rect 3532 23969 3572 25843
rect 3688 25724 4056 25733
rect 3728 25684 3770 25724
rect 3810 25684 3852 25724
rect 3892 25684 3934 25724
rect 3974 25684 4016 25724
rect 3688 25675 4056 25684
rect 3819 25304 3861 25313
rect 3819 25264 3820 25304
rect 3860 25264 3861 25304
rect 3819 25255 3861 25264
rect 3820 25170 3860 25255
rect 3688 24212 4056 24221
rect 3728 24172 3770 24212
rect 3810 24172 3852 24212
rect 3892 24172 3934 24212
rect 3974 24172 4016 24212
rect 3688 24163 4056 24172
rect 3819 24044 3861 24053
rect 3819 24004 3820 24044
rect 3860 24004 3861 24044
rect 3819 23995 3861 24004
rect 3244 23920 3476 23960
rect 3531 23960 3573 23969
rect 3531 23920 3532 23960
rect 3572 23920 3573 23960
rect 3148 23801 3188 23886
rect 3147 23792 3189 23801
rect 3147 23752 3148 23792
rect 3188 23752 3189 23792
rect 3147 23743 3189 23752
rect 2668 22483 2708 22492
rect 2860 22483 2900 22492
rect 2956 23080 3052 23120
rect 2956 21953 2996 23080
rect 3052 23071 3092 23080
rect 3051 22280 3093 22289
rect 3051 22240 3052 22280
rect 3092 22240 3093 22280
rect 3051 22231 3093 22240
rect 2955 21944 2997 21953
rect 2955 21904 2956 21944
rect 2996 21904 2997 21944
rect 2955 21895 2997 21904
rect 2956 21776 2996 21895
rect 2860 21736 2996 21776
rect 2763 21692 2805 21701
rect 2763 21652 2764 21692
rect 2804 21652 2805 21692
rect 2763 21643 2805 21652
rect 2764 21113 2804 21643
rect 2860 21449 2900 21736
rect 2956 21608 2996 21617
rect 3052 21608 3092 22231
rect 3147 21776 3189 21785
rect 3147 21736 3148 21776
rect 3188 21736 3189 21776
rect 3147 21727 3189 21736
rect 3148 21642 3188 21727
rect 2996 21568 3092 21608
rect 2956 21559 2996 21568
rect 3244 21524 3284 23920
rect 3531 23911 3573 23920
rect 3820 23910 3860 23995
rect 3436 23792 3476 23801
rect 3436 23456 3476 23752
rect 4012 23792 4052 23801
rect 3531 23708 3573 23717
rect 3531 23668 3532 23708
rect 3572 23668 3573 23708
rect 3531 23659 3573 23668
rect 3532 23574 3572 23659
rect 3436 23416 3764 23456
rect 3724 23288 3764 23416
rect 3724 23239 3764 23248
rect 3916 23120 3956 23131
rect 4012 23129 4052 23752
rect 4108 23465 4148 25852
rect 4203 25724 4245 25733
rect 4203 25684 4204 25724
rect 4244 25684 4245 25724
rect 4203 25675 4245 25684
rect 4204 25313 4244 25675
rect 4203 25304 4245 25313
rect 4203 25264 4204 25304
rect 4244 25264 4245 25304
rect 4203 25255 4245 25264
rect 4300 25309 4340 25318
rect 4300 25229 4340 25269
rect 4299 25220 4341 25229
rect 4299 25180 4300 25220
rect 4340 25180 4341 25220
rect 4299 25171 4341 25180
rect 4203 24884 4245 24893
rect 4203 24844 4204 24884
rect 4244 24844 4245 24884
rect 4203 24835 4245 24844
rect 4204 24725 4244 24835
rect 4396 24800 4436 26431
rect 4491 26144 4533 26153
rect 4491 26104 4492 26144
rect 4532 26104 4533 26144
rect 4491 26095 4533 26104
rect 4492 25220 4532 26095
rect 4492 25171 4532 25180
rect 4396 24760 4532 24800
rect 4203 24716 4245 24725
rect 4203 24676 4204 24716
rect 4244 24676 4245 24716
rect 4203 24667 4245 24676
rect 4396 24632 4436 24643
rect 4396 24557 4436 24592
rect 4395 24548 4437 24557
rect 4395 24508 4396 24548
rect 4436 24508 4437 24548
rect 4395 24499 4437 24508
rect 4395 24128 4437 24137
rect 4395 24088 4396 24128
rect 4436 24088 4437 24128
rect 4395 24079 4437 24088
rect 4299 23960 4341 23969
rect 4299 23920 4300 23960
rect 4340 23920 4341 23960
rect 4299 23911 4341 23920
rect 4107 23456 4149 23465
rect 4107 23416 4108 23456
rect 4148 23416 4149 23456
rect 4107 23407 4149 23416
rect 3532 23106 3572 23115
rect 3435 22952 3477 22961
rect 3435 22912 3436 22952
rect 3476 22912 3477 22952
rect 3435 22903 3477 22912
rect 3148 21484 3284 21524
rect 2859 21440 2901 21449
rect 2859 21400 2860 21440
rect 2900 21400 2901 21440
rect 2859 21391 2901 21400
rect 2763 21104 2805 21113
rect 2763 21064 2764 21104
rect 2804 21064 2805 21104
rect 2763 21055 2805 21064
rect 2284 20140 2516 20180
rect 1803 19760 1845 19769
rect 1803 19720 1804 19760
rect 1844 19720 1845 19760
rect 1803 19711 1845 19720
rect 1268 18544 1460 18584
rect 1803 18584 1845 18593
rect 1803 18544 1804 18584
rect 1844 18544 1845 18584
rect 1228 18535 1268 18544
rect 1803 18535 1845 18544
rect 1323 17996 1365 18005
rect 1323 17956 1324 17996
rect 1364 17956 1365 17996
rect 1323 17947 1365 17956
rect 1324 17744 1364 17947
rect 1324 17695 1364 17704
rect 1515 17744 1557 17753
rect 1515 17704 1516 17744
rect 1556 17704 1557 17744
rect 1515 17695 1557 17704
rect 1612 17744 1652 17753
rect 1516 17610 1556 17695
rect 1420 17576 1460 17585
rect 1420 17081 1460 17536
rect 1612 17165 1652 17704
rect 1804 17744 1844 18535
rect 1804 17660 1844 17704
rect 1708 17620 1844 17660
rect 1611 17156 1653 17165
rect 1611 17116 1612 17156
rect 1652 17116 1653 17156
rect 1611 17107 1653 17116
rect 1228 17072 1268 17081
rect 1419 17072 1461 17081
rect 1268 17032 1364 17072
rect 1228 17023 1268 17032
rect 1324 16904 1364 17032
rect 1419 17032 1420 17072
rect 1460 17032 1461 17072
rect 1419 17023 1461 17032
rect 1708 16904 1748 17620
rect 1803 17492 1845 17501
rect 1803 17452 1804 17492
rect 1844 17452 1845 17492
rect 1803 17443 1845 17452
rect 1324 16864 1748 16904
rect 1227 16820 1269 16829
rect 1227 16780 1228 16820
rect 1268 16780 1269 16820
rect 1227 16771 1269 16780
rect 1228 16232 1268 16771
rect 1228 16183 1268 16192
rect 1515 15896 1557 15905
rect 1515 15856 1516 15896
rect 1556 15856 1557 15896
rect 1515 15847 1557 15856
rect 1420 15392 1460 15401
rect 1228 15352 1420 15392
rect 1228 13553 1268 15352
rect 1420 15343 1460 15352
rect 1323 15224 1365 15233
rect 1323 15184 1324 15224
rect 1364 15184 1365 15224
rect 1323 15175 1365 15184
rect 1324 14216 1364 15175
rect 1420 14972 1460 14981
rect 1516 14972 1556 15847
rect 1611 15644 1653 15653
rect 1611 15604 1612 15644
rect 1652 15604 1653 15644
rect 1611 15595 1653 15604
rect 1804 15602 1844 17443
rect 2284 16493 2324 20140
rect 2476 20096 2516 20140
rect 2476 20047 2516 20056
rect 2475 19844 2517 19853
rect 2475 19804 2476 19844
rect 2516 19804 2517 19844
rect 2475 19795 2517 19804
rect 2476 19270 2516 19795
rect 2572 19433 2612 20728
rect 2667 20768 2709 20777
rect 2667 20728 2668 20768
rect 2708 20728 2709 20768
rect 2667 20719 2709 20728
rect 2571 19424 2613 19433
rect 2571 19384 2572 19424
rect 2612 19384 2613 19424
rect 2571 19375 2613 19384
rect 2476 19265 2611 19270
rect 2476 19256 2612 19265
rect 2476 19230 2572 19256
rect 2476 18584 2516 19230
rect 2571 19216 2572 19230
rect 2572 19207 2612 19216
rect 2571 18752 2613 18761
rect 2571 18712 2572 18752
rect 2612 18712 2613 18752
rect 2571 18703 2613 18712
rect 2668 18752 2708 20719
rect 2764 20180 2804 21055
rect 2955 20936 2997 20945
rect 2955 20896 2956 20936
rect 2996 20896 2997 20936
rect 2955 20887 2997 20896
rect 2956 20357 2996 20887
rect 3052 20773 3092 20782
rect 2955 20348 2997 20357
rect 2955 20308 2956 20348
rect 2996 20308 2997 20348
rect 2955 20299 2997 20308
rect 2764 20140 2900 20180
rect 2763 19508 2805 19517
rect 2763 19468 2764 19508
rect 2804 19468 2805 19508
rect 2763 19459 2805 19468
rect 2764 19374 2804 19459
rect 2860 18752 2900 20140
rect 3052 19517 3092 20733
rect 3051 19508 3093 19517
rect 3051 19468 3052 19508
rect 3092 19468 3093 19508
rect 3051 19459 3093 19468
rect 2955 19424 2997 19433
rect 2955 19384 2956 19424
rect 2996 19384 2997 19424
rect 2955 19375 2997 19384
rect 2668 18703 2708 18712
rect 2764 18712 2900 18752
rect 2956 18752 2996 19375
rect 3148 18929 3188 21484
rect 3339 21020 3381 21029
rect 3339 20980 3340 21020
rect 3380 20980 3381 21020
rect 3339 20971 3381 20980
rect 3244 20600 3284 20609
rect 3147 18920 3189 18929
rect 3147 18880 3148 18920
rect 3188 18880 3189 18920
rect 3147 18871 3189 18880
rect 3148 18752 3188 18761
rect 2956 18712 3092 18752
rect 2476 18535 2516 18544
rect 2572 17324 2612 18703
rect 2667 17660 2709 17669
rect 2667 17620 2668 17660
rect 2708 17620 2709 17660
rect 2667 17611 2709 17620
rect 2380 17284 2612 17324
rect 1899 16484 1941 16493
rect 1899 16444 1900 16484
rect 1940 16444 1941 16484
rect 1899 16435 1941 16444
rect 2283 16484 2325 16493
rect 2283 16444 2284 16484
rect 2324 16444 2325 16484
rect 2283 16435 2325 16444
rect 1612 15476 1652 15595
rect 1707 15560 1749 15569
rect 1707 15520 1708 15560
rect 1748 15520 1749 15560
rect 1804 15553 1844 15562
rect 1707 15511 1749 15520
rect 1612 15427 1652 15436
rect 1611 15224 1653 15233
rect 1611 15184 1612 15224
rect 1652 15184 1653 15224
rect 1611 15175 1653 15184
rect 1460 14932 1556 14972
rect 1420 14923 1460 14932
rect 1612 14804 1652 15175
rect 1612 14755 1652 14764
rect 1708 14636 1748 15511
rect 1900 15476 1940 16435
rect 2380 15560 2420 17284
rect 2668 17240 2708 17611
rect 2668 17191 2708 17200
rect 2571 17156 2613 17165
rect 2571 17116 2572 17156
rect 2612 17116 2613 17156
rect 2571 17107 2613 17116
rect 2476 17072 2516 17081
rect 2476 16232 2516 17032
rect 2572 16484 2612 17107
rect 2668 16484 2708 16493
rect 2572 16444 2668 16484
rect 2668 16435 2708 16444
rect 2764 16241 2804 18712
rect 2860 18584 2900 18593
rect 2860 17669 2900 18544
rect 2956 18584 2996 18593
rect 2956 18089 2996 18544
rect 2955 18080 2997 18089
rect 2955 18040 2956 18080
rect 2996 18040 2997 18080
rect 2955 18031 2997 18040
rect 3052 17912 3092 18712
rect 2956 17872 3092 17912
rect 2859 17660 2901 17669
rect 2859 17620 2860 17660
rect 2900 17620 2901 17660
rect 2859 17611 2901 17620
rect 2860 17333 2900 17611
rect 2956 17501 2996 17872
rect 3052 17744 3092 17755
rect 3052 17669 3092 17704
rect 3051 17660 3093 17669
rect 3051 17620 3052 17660
rect 3092 17620 3093 17660
rect 3051 17611 3093 17620
rect 3052 17580 3092 17611
rect 2955 17492 2997 17501
rect 2955 17452 2956 17492
rect 2996 17452 2997 17492
rect 2955 17443 2997 17452
rect 2859 17324 2901 17333
rect 2859 17284 2860 17324
rect 2900 17284 2901 17324
rect 2859 17275 2901 17284
rect 2860 17081 2900 17166
rect 2955 17156 2997 17165
rect 2955 17116 2956 17156
rect 2996 17116 2997 17156
rect 2955 17107 2997 17116
rect 2859 17072 2901 17081
rect 2859 17032 2860 17072
rect 2900 17032 2901 17072
rect 2859 17023 2901 17032
rect 2956 17072 2996 17107
rect 2956 17021 2996 17032
rect 3148 17072 3188 18712
rect 3244 17837 3284 20560
rect 3340 18761 3380 20971
rect 3436 20945 3476 22903
rect 3532 22373 3572 23066
rect 3916 23045 3956 23080
rect 4011 23120 4053 23129
rect 4011 23080 4012 23120
rect 4052 23080 4053 23120
rect 4011 23071 4053 23080
rect 3915 23036 3957 23045
rect 3915 22996 3916 23036
rect 3956 22996 3957 23036
rect 3915 22987 3957 22996
rect 3688 22700 4056 22709
rect 3728 22660 3770 22700
rect 3810 22660 3852 22700
rect 3892 22660 3934 22700
rect 3974 22660 4016 22700
rect 3688 22651 4056 22660
rect 3531 22364 3573 22373
rect 3531 22324 3532 22364
rect 3572 22324 3573 22364
rect 3531 22315 3573 22324
rect 3532 21785 3572 22315
rect 4300 22280 4340 23911
rect 4300 22231 4340 22240
rect 4107 21944 4149 21953
rect 4107 21904 4108 21944
rect 4148 21904 4149 21944
rect 4107 21895 4149 21904
rect 3531 21776 3573 21785
rect 3531 21736 3532 21776
rect 3572 21736 3573 21776
rect 3531 21727 3573 21736
rect 3723 21692 3765 21701
rect 3723 21652 3724 21692
rect 3764 21652 3765 21692
rect 3723 21643 3765 21652
rect 3628 21608 3668 21617
rect 3532 21568 3628 21608
rect 3435 20936 3477 20945
rect 3435 20896 3436 20936
rect 3476 20896 3477 20936
rect 3435 20887 3477 20896
rect 3532 20861 3572 21568
rect 3628 21559 3668 21568
rect 3724 21608 3764 21643
rect 3724 21557 3764 21568
rect 4108 21608 4148 21895
rect 4108 21559 4148 21568
rect 4203 21608 4245 21617
rect 4203 21568 4204 21608
rect 4244 21568 4245 21608
rect 4203 21559 4245 21568
rect 4204 21474 4244 21559
rect 3688 21188 4056 21197
rect 3728 21148 3770 21188
rect 3810 21148 3852 21188
rect 3892 21148 3934 21188
rect 3974 21148 4016 21188
rect 3688 21139 4056 21148
rect 3723 20936 3765 20945
rect 3723 20896 3724 20936
rect 3764 20896 3765 20936
rect 3723 20887 3765 20896
rect 3531 20852 3573 20861
rect 3531 20812 3532 20852
rect 3572 20812 3573 20852
rect 3531 20803 3573 20812
rect 3435 20768 3477 20777
rect 3435 20728 3436 20768
rect 3476 20728 3477 20768
rect 3435 20719 3477 20728
rect 3436 20634 3476 20719
rect 3724 20096 3764 20887
rect 3915 20852 3957 20861
rect 3915 20812 3916 20852
rect 3956 20812 3957 20852
rect 3915 20803 3957 20812
rect 3916 20180 3956 20803
rect 3916 20131 3956 20140
rect 3724 20047 3764 20056
rect 4396 20096 4436 24079
rect 4492 22448 4532 24760
rect 4588 24137 4628 26944
rect 4684 26825 4724 27028
rect 4683 26816 4725 26825
rect 4683 26776 4684 26816
rect 4724 26776 4725 26816
rect 4683 26767 4725 26776
rect 4780 26144 4820 27271
rect 5260 26741 5300 27364
rect 5259 26732 5301 26741
rect 5259 26692 5260 26732
rect 5300 26692 5301 26732
rect 5259 26683 5301 26692
rect 5548 26648 5588 28204
rect 5643 27740 5685 27749
rect 5643 27700 5644 27740
rect 5684 27700 5685 27740
rect 5643 27691 5685 27700
rect 5644 27656 5684 27691
rect 5644 27605 5684 27616
rect 5740 27152 5780 34504
rect 5836 32612 5876 35251
rect 5932 34964 5972 34973
rect 5932 34721 5972 34924
rect 5931 34712 5973 34721
rect 5931 34672 5932 34712
rect 5972 34672 5973 34712
rect 5931 34663 5973 34672
rect 5932 34124 5972 34663
rect 6028 34460 6068 35251
rect 6124 34544 6164 37360
rect 6220 36569 6260 38956
rect 6412 38240 6452 39460
rect 6700 39164 6740 39703
rect 6700 39115 6740 39124
rect 6796 39089 6836 39712
rect 6896 39752 6938 39761
rect 6896 39712 6897 39752
rect 6937 39712 6938 39752
rect 6896 39703 6938 39712
rect 6897 39618 6937 39703
rect 6795 39080 6837 39089
rect 6795 39040 6796 39080
rect 6836 39040 6837 39080
rect 6795 39031 6837 39040
rect 6891 38996 6933 39005
rect 6891 38956 6892 38996
rect 6932 38956 6933 38996
rect 6891 38947 6933 38956
rect 6508 38912 6548 38923
rect 6508 38837 6548 38872
rect 6892 38912 6932 38947
rect 6892 38861 6932 38872
rect 6507 38828 6549 38837
rect 6507 38788 6508 38828
rect 6548 38788 6549 38828
rect 6507 38779 6549 38788
rect 6988 38744 7028 40459
rect 6892 38704 7028 38744
rect 6508 38240 6548 38249
rect 6412 38200 6508 38240
rect 6508 37652 6548 38200
rect 6699 37904 6741 37913
rect 6699 37864 6700 37904
rect 6740 37864 6741 37904
rect 6699 37855 6741 37864
rect 6700 37736 6740 37855
rect 6700 37696 6836 37736
rect 6508 37612 6740 37652
rect 6700 37493 6740 37612
rect 6699 37484 6741 37493
rect 6699 37444 6700 37484
rect 6740 37444 6741 37484
rect 6699 37435 6741 37444
rect 6508 37400 6548 37409
rect 6219 36560 6261 36569
rect 6219 36520 6220 36560
rect 6260 36520 6261 36560
rect 6219 36511 6261 36520
rect 6220 35888 6260 35897
rect 6220 35225 6260 35848
rect 6412 35720 6452 35729
rect 6316 35680 6412 35720
rect 6219 35216 6261 35225
rect 6219 35176 6220 35216
rect 6260 35176 6261 35216
rect 6219 35167 6261 35176
rect 6124 34504 6260 34544
rect 6028 34301 6068 34420
rect 6123 34376 6165 34385
rect 6123 34336 6124 34376
rect 6164 34336 6165 34376
rect 6123 34327 6165 34336
rect 6027 34292 6069 34301
rect 6027 34252 6028 34292
rect 6068 34252 6069 34292
rect 6027 34243 6069 34252
rect 6124 34242 6164 34327
rect 5932 34084 6164 34124
rect 5931 33956 5973 33965
rect 5931 33916 5932 33956
rect 5972 33916 5973 33956
rect 5931 33907 5973 33916
rect 5932 32696 5972 33907
rect 6028 33704 6068 33715
rect 6124 33713 6164 34084
rect 6220 34049 6260 34504
rect 6316 34385 6356 35680
rect 6412 35671 6452 35680
rect 6508 35393 6548 37360
rect 6603 37400 6645 37409
rect 6603 37360 6604 37400
rect 6644 37360 6645 37400
rect 6603 37351 6645 37360
rect 6604 37266 6644 37351
rect 6603 35888 6645 35897
rect 6603 35848 6604 35888
rect 6644 35848 6645 35888
rect 6603 35839 6645 35848
rect 6604 35754 6644 35839
rect 6507 35384 6549 35393
rect 6507 35344 6508 35384
rect 6548 35344 6549 35384
rect 6507 35335 6549 35344
rect 6603 35300 6645 35309
rect 6603 35260 6604 35300
rect 6644 35260 6645 35300
rect 6603 35251 6645 35260
rect 6412 35216 6452 35225
rect 6412 34637 6452 35176
rect 6508 35216 6548 35225
rect 6411 34628 6453 34637
rect 6411 34588 6412 34628
rect 6452 34588 6453 34628
rect 6411 34579 6453 34588
rect 6315 34376 6357 34385
rect 6315 34336 6316 34376
rect 6356 34336 6357 34376
rect 6315 34327 6357 34336
rect 6315 34208 6357 34217
rect 6315 34168 6316 34208
rect 6356 34168 6357 34208
rect 6315 34159 6357 34168
rect 6219 34040 6261 34049
rect 6219 34000 6220 34040
rect 6260 34000 6261 34040
rect 6219 33991 6261 34000
rect 6219 33872 6261 33881
rect 6219 33832 6220 33872
rect 6260 33832 6261 33872
rect 6219 33823 6261 33832
rect 6220 33738 6260 33823
rect 6028 33629 6068 33664
rect 6123 33704 6165 33713
rect 6123 33664 6124 33704
rect 6164 33664 6165 33704
rect 6123 33655 6165 33664
rect 6316 33704 6356 34159
rect 6508 34049 6548 35176
rect 6604 35166 6644 35251
rect 6700 35216 6740 35225
rect 6700 34721 6740 35176
rect 6796 35141 6836 37696
rect 6892 35897 6932 38704
rect 6987 38324 7029 38333
rect 6987 38284 6988 38324
rect 7028 38284 7029 38324
rect 6987 38275 7029 38284
rect 6988 38235 7028 38275
rect 6988 38186 7028 38195
rect 6987 38072 7029 38081
rect 6987 38032 6988 38072
rect 7028 38032 7029 38072
rect 6987 38023 7029 38032
rect 6891 35888 6933 35897
rect 6891 35848 6892 35888
rect 6932 35848 6933 35888
rect 6891 35839 6933 35848
rect 6892 35393 6932 35839
rect 6891 35384 6933 35393
rect 6891 35344 6892 35384
rect 6932 35344 6933 35384
rect 6891 35335 6933 35344
rect 6892 35258 6932 35267
rect 6988 35225 7028 38023
rect 7084 37820 7124 41308
rect 7275 41096 7317 41105
rect 7275 41056 7276 41096
rect 7316 41056 7317 41096
rect 7275 41047 7317 41056
rect 7179 40760 7221 40769
rect 7179 40720 7180 40760
rect 7220 40720 7221 40760
rect 7179 40711 7221 40720
rect 7180 40433 7220 40711
rect 7179 40424 7221 40433
rect 7179 40384 7180 40424
rect 7220 40384 7221 40424
rect 7179 40375 7221 40384
rect 7179 40172 7221 40181
rect 7179 40132 7180 40172
rect 7220 40132 7221 40172
rect 7179 40123 7221 40132
rect 7180 38744 7220 40123
rect 7276 39005 7316 41047
rect 7372 40676 7412 41476
rect 7372 40627 7412 40636
rect 7468 40508 7508 43240
rect 8044 42692 8084 43408
rect 8140 42785 8180 42870
rect 8139 42776 8181 42785
rect 8139 42736 8140 42776
rect 8180 42736 8181 42776
rect 8139 42727 8181 42736
rect 7948 42652 8084 42692
rect 7948 42524 7988 42652
rect 7948 42484 8276 42524
rect 7564 41936 7604 41945
rect 7564 41693 7604 41896
rect 7563 41684 7605 41693
rect 7563 41644 7564 41684
rect 7604 41644 7605 41684
rect 7563 41635 7605 41644
rect 7660 41264 7700 41273
rect 7700 41224 7988 41264
rect 7660 41215 7700 41224
rect 7659 40592 7701 40601
rect 7659 40552 7660 40592
rect 7700 40552 7701 40592
rect 7659 40543 7701 40552
rect 7372 40468 7508 40508
rect 7275 38996 7317 39005
rect 7275 38956 7276 38996
rect 7316 38956 7317 38996
rect 7275 38947 7317 38956
rect 7180 38704 7316 38744
rect 7179 38576 7221 38585
rect 7179 38536 7180 38576
rect 7220 38536 7221 38576
rect 7179 38527 7221 38536
rect 7180 38408 7220 38527
rect 7180 38359 7220 38368
rect 7276 38081 7316 38704
rect 7275 38072 7317 38081
rect 7275 38032 7276 38072
rect 7316 38032 7317 38072
rect 7275 38023 7317 38032
rect 7372 37820 7412 40468
rect 7564 40340 7604 40349
rect 7564 39761 7604 40300
rect 7563 39752 7605 39761
rect 7563 39712 7564 39752
rect 7604 39712 7605 39752
rect 7563 39703 7605 39712
rect 7660 39752 7700 40543
rect 7755 40424 7797 40433
rect 7755 40384 7756 40424
rect 7796 40384 7797 40424
rect 7755 40375 7797 40384
rect 7756 40290 7796 40375
rect 7700 39712 7892 39752
rect 7660 39703 7700 39712
rect 7467 39584 7509 39593
rect 7467 39544 7468 39584
rect 7508 39544 7509 39584
rect 7467 39535 7509 39544
rect 7468 38408 7508 39535
rect 7564 39500 7604 39703
rect 7564 39460 7796 39500
rect 7659 38996 7701 39005
rect 7659 38956 7660 38996
rect 7700 38956 7701 38996
rect 7659 38947 7701 38956
rect 7468 38359 7508 38368
rect 7660 38240 7700 38947
rect 7660 38191 7700 38200
rect 7756 38240 7796 39460
rect 7756 38191 7796 38200
rect 7852 37820 7892 39712
rect 7948 39425 7988 41224
rect 8139 39752 8181 39761
rect 8139 39712 8140 39752
rect 8180 39712 8181 39752
rect 8139 39703 8181 39712
rect 7947 39416 7989 39425
rect 7947 39376 7948 39416
rect 7988 39376 7989 39416
rect 7947 39367 7989 39376
rect 8043 39080 8085 39089
rect 8043 39040 8044 39080
rect 8084 39040 8085 39080
rect 8043 39031 8085 39040
rect 8044 38408 8084 39031
rect 8044 38359 8084 38368
rect 8140 38912 8180 39703
rect 7948 38240 7988 38249
rect 7948 37913 7988 38200
rect 7947 37904 7989 37913
rect 7947 37864 7948 37904
rect 7988 37864 7989 37904
rect 7947 37855 7989 37864
rect 7084 37780 7316 37820
rect 7372 37780 7508 37820
rect 7276 37577 7316 37780
rect 7275 37568 7317 37577
rect 7275 37528 7276 37568
rect 7316 37528 7412 37568
rect 7275 37519 7317 37528
rect 7082 37484 7124 37493
rect 7082 37444 7083 37484
rect 7123 37444 7124 37484
rect 7082 37435 7124 37444
rect 7084 37400 7124 37435
rect 7084 37351 7124 37360
rect 7179 37064 7221 37073
rect 7179 37024 7180 37064
rect 7220 37024 7221 37064
rect 7179 37015 7221 37024
rect 7084 36728 7124 36739
rect 7084 36653 7124 36688
rect 7083 36644 7125 36653
rect 7083 36604 7084 36644
rect 7124 36604 7125 36644
rect 7083 36595 7125 36604
rect 6892 35216 6932 35218
rect 6887 35176 6932 35216
rect 6987 35216 7029 35225
rect 6987 35176 6988 35216
rect 7028 35176 7029 35216
rect 6795 35132 6837 35141
rect 6795 35092 6796 35132
rect 6836 35092 6837 35132
rect 6887 35132 6927 35176
rect 6987 35167 7029 35176
rect 6887 35092 6932 35132
rect 6795 35083 6837 35092
rect 6892 35048 6932 35092
rect 6892 35008 6935 35048
rect 6895 34964 6935 35008
rect 6892 34924 6935 34964
rect 6892 34805 6932 34924
rect 6891 34796 6933 34805
rect 6891 34756 6892 34796
rect 6932 34756 6933 34796
rect 6891 34747 6933 34756
rect 6699 34712 6741 34721
rect 6699 34672 6700 34712
rect 6740 34672 6741 34712
rect 6699 34663 6741 34672
rect 6604 34376 6644 34385
rect 6604 34217 6644 34336
rect 7084 34381 7124 34390
rect 6795 34292 6837 34301
rect 6795 34252 6796 34292
rect 6836 34252 6837 34292
rect 6795 34243 6837 34252
rect 6603 34208 6645 34217
rect 6603 34168 6604 34208
rect 6644 34168 6740 34208
rect 6603 34159 6645 34168
rect 6507 34040 6549 34049
rect 6507 34000 6508 34040
rect 6548 34000 6549 34040
rect 6507 33991 6549 34000
rect 6316 33655 6356 33664
rect 6603 33704 6645 33713
rect 6603 33664 6604 33704
rect 6644 33664 6645 33704
rect 6603 33655 6645 33664
rect 6027 33620 6069 33629
rect 6027 33580 6028 33620
rect 6068 33580 6069 33620
rect 6027 33571 6069 33580
rect 6124 33570 6164 33655
rect 6604 33570 6644 33655
rect 6123 33200 6165 33209
rect 6123 33160 6124 33200
rect 6164 33160 6165 33200
rect 6123 33151 6165 33160
rect 6124 32864 6164 33151
rect 6700 33032 6740 34168
rect 6124 32815 6164 32824
rect 6604 32992 6740 33032
rect 5932 32656 6164 32696
rect 5836 32572 6068 32612
rect 5835 32444 5877 32453
rect 5835 32404 5836 32444
rect 5876 32404 5877 32444
rect 5835 32395 5877 32404
rect 5836 32192 5876 32395
rect 5932 32285 5972 32307
rect 5931 32276 5973 32285
rect 5931 32236 5932 32276
rect 5972 32236 5973 32276
rect 5931 32227 5973 32236
rect 5932 32212 5972 32227
rect 5932 32163 5972 32172
rect 5836 32143 5876 32152
rect 6028 32024 6068 32572
rect 5836 31984 6068 32024
rect 5836 30941 5876 31984
rect 5931 31772 5973 31781
rect 5931 31732 5932 31772
rect 5972 31732 5973 31772
rect 5931 31723 5973 31732
rect 5835 30932 5877 30941
rect 5835 30892 5836 30932
rect 5876 30892 5877 30932
rect 5835 30883 5877 30892
rect 5835 30764 5877 30773
rect 5835 30724 5836 30764
rect 5876 30724 5877 30764
rect 5835 30715 5877 30724
rect 5836 30630 5876 30715
rect 5835 30512 5877 30521
rect 5835 30472 5836 30512
rect 5876 30472 5877 30512
rect 5835 30463 5877 30472
rect 5836 29840 5876 30463
rect 5836 29513 5876 29800
rect 5835 29504 5877 29513
rect 5835 29464 5836 29504
rect 5876 29464 5877 29504
rect 5835 29455 5877 29464
rect 5932 29000 5972 31723
rect 6028 31357 6068 31366
rect 6028 30092 6068 31317
rect 6124 30689 6164 32656
rect 6219 32612 6261 32621
rect 6219 32572 6220 32612
rect 6260 32572 6261 32612
rect 6219 32563 6261 32572
rect 6220 31268 6260 32563
rect 6507 32444 6549 32453
rect 6507 32404 6508 32444
rect 6548 32404 6549 32444
rect 6507 32395 6549 32404
rect 6316 32108 6356 32117
rect 6316 31613 6356 32068
rect 6411 32108 6453 32117
rect 6411 32068 6412 32108
rect 6452 32068 6453 32108
rect 6411 32059 6453 32068
rect 6315 31604 6357 31613
rect 6315 31564 6316 31604
rect 6356 31564 6357 31604
rect 6315 31555 6357 31564
rect 6412 31436 6452 32059
rect 6220 31219 6260 31228
rect 6316 31396 6452 31436
rect 6123 30680 6165 30689
rect 6123 30640 6124 30680
rect 6164 30640 6165 30680
rect 6123 30631 6165 30640
rect 6028 30043 6068 30052
rect 6123 29840 6165 29849
rect 6123 29800 6124 29840
rect 6164 29800 6165 29840
rect 6123 29791 6165 29800
rect 5932 28960 6068 29000
rect 5931 28664 5973 28673
rect 5931 28624 5932 28664
rect 5972 28624 5973 28664
rect 5931 28615 5973 28624
rect 5835 28496 5877 28505
rect 5835 28456 5836 28496
rect 5876 28456 5877 28496
rect 5835 28447 5877 28456
rect 5836 28328 5876 28447
rect 5836 28279 5876 28288
rect 5932 28328 5972 28615
rect 5932 28085 5972 28288
rect 5931 28076 5973 28085
rect 5931 28036 5932 28076
rect 5972 28036 5973 28076
rect 5931 28027 5973 28036
rect 5931 27908 5973 27917
rect 5931 27868 5932 27908
rect 5972 27868 5973 27908
rect 5931 27859 5973 27868
rect 5932 27656 5972 27859
rect 5932 27607 5972 27616
rect 5740 27112 5876 27152
rect 5739 26984 5781 26993
rect 5739 26944 5740 26984
rect 5780 26944 5781 26984
rect 5739 26935 5781 26944
rect 5740 26816 5780 26935
rect 5740 26767 5780 26776
rect 5548 26608 5780 26648
rect 4928 26480 5296 26489
rect 4968 26440 5010 26480
rect 5050 26440 5092 26480
rect 5132 26440 5174 26480
rect 5214 26440 5256 26480
rect 4928 26431 5296 26440
rect 5547 26480 5589 26489
rect 5547 26440 5548 26480
rect 5588 26440 5589 26480
rect 5547 26431 5589 26440
rect 5067 26312 5109 26321
rect 5067 26272 5068 26312
rect 5108 26272 5109 26312
rect 5067 26263 5109 26272
rect 5451 26312 5493 26321
rect 5451 26272 5452 26312
rect 5492 26272 5493 26312
rect 5451 26263 5493 26272
rect 4780 25985 4820 26104
rect 4779 25976 4821 25985
rect 4779 25936 4780 25976
rect 4820 25936 4821 25976
rect 4779 25927 4821 25936
rect 4972 25892 5012 25901
rect 4972 25649 5012 25852
rect 4971 25640 5013 25649
rect 4971 25600 4972 25640
rect 5012 25600 5013 25640
rect 4971 25591 5013 25600
rect 4683 25472 4725 25481
rect 4683 25432 4684 25472
rect 4724 25432 4725 25472
rect 4683 25423 4725 25432
rect 4684 25304 4724 25423
rect 4780 25313 4820 25398
rect 4684 25255 4724 25264
rect 4779 25304 4821 25313
rect 4779 25264 4780 25304
rect 4820 25264 4821 25304
rect 4779 25255 4821 25264
rect 4876 25304 4916 25313
rect 5068 25304 5108 26263
rect 5452 26178 5492 26263
rect 5164 26144 5204 26153
rect 5164 25565 5204 26104
rect 5259 26144 5301 26153
rect 5259 26104 5260 26144
rect 5300 26104 5301 26144
rect 5259 26095 5301 26104
rect 5260 26010 5300 26095
rect 5163 25556 5205 25565
rect 5163 25516 5164 25556
rect 5204 25516 5205 25556
rect 5163 25507 5205 25516
rect 5259 25472 5301 25481
rect 5259 25432 5260 25472
rect 5300 25432 5301 25472
rect 5259 25423 5301 25432
rect 5163 25388 5205 25397
rect 5163 25348 5164 25388
rect 5204 25348 5205 25388
rect 5163 25339 5205 25348
rect 4916 25264 5108 25304
rect 5164 25304 5204 25339
rect 4876 25255 4916 25264
rect 5164 25253 5204 25264
rect 5260 25304 5300 25423
rect 5260 25255 5300 25264
rect 5356 25304 5396 25313
rect 4972 25136 5012 25145
rect 5067 25136 5109 25145
rect 5012 25096 5068 25136
rect 5108 25096 5109 25136
rect 4972 25087 5012 25096
rect 5067 25087 5109 25096
rect 4928 24968 5296 24977
rect 4968 24928 5010 24968
rect 5050 24928 5092 24968
rect 5132 24928 5174 24968
rect 5214 24928 5256 24968
rect 4928 24919 5296 24928
rect 5356 24809 5396 25264
rect 5452 25283 5492 25292
rect 5452 25229 5492 25243
rect 5451 25220 5493 25229
rect 5451 25180 5452 25220
rect 5492 25180 5493 25220
rect 5451 25171 5493 25180
rect 5452 25148 5492 25171
rect 4875 24800 4917 24809
rect 4875 24760 4876 24800
rect 4916 24760 4917 24800
rect 4875 24751 4917 24760
rect 5355 24800 5397 24809
rect 5355 24760 5356 24800
rect 5396 24760 5397 24800
rect 5355 24751 5397 24760
rect 4876 24632 4916 24751
rect 4876 24583 4916 24592
rect 5355 24464 5397 24473
rect 5355 24424 5356 24464
rect 5396 24424 5397 24464
rect 5355 24415 5397 24424
rect 4587 24128 4629 24137
rect 4587 24088 4588 24128
rect 4628 24088 4629 24128
rect 4587 24079 4629 24088
rect 5259 24128 5301 24137
rect 5259 24088 5260 24128
rect 5300 24088 5301 24128
rect 5259 24079 5301 24088
rect 5260 23792 5300 24079
rect 5260 23743 5300 23752
rect 4928 23456 5296 23465
rect 4968 23416 5010 23456
rect 5050 23416 5092 23456
rect 5132 23416 5174 23456
rect 5214 23416 5256 23456
rect 4928 23407 5296 23416
rect 5164 23120 5204 23129
rect 5356 23120 5396 24415
rect 5451 23792 5493 23801
rect 5451 23752 5452 23792
rect 5492 23752 5493 23792
rect 5451 23743 5493 23752
rect 5452 23708 5492 23743
rect 5452 23657 5492 23668
rect 5204 23080 5396 23120
rect 5164 23071 5204 23080
rect 5355 22868 5397 22877
rect 5355 22828 5356 22868
rect 5396 22828 5397 22868
rect 5355 22819 5397 22828
rect 5356 22734 5396 22819
rect 4492 22408 4628 22448
rect 4491 22280 4533 22289
rect 4491 22240 4492 22280
rect 4532 22240 4533 22280
rect 4491 22231 4533 22240
rect 4492 22146 4532 22231
rect 4396 20021 4436 20056
rect 4491 20096 4533 20105
rect 4491 20056 4492 20096
rect 4532 20056 4533 20096
rect 4491 20047 4533 20056
rect 3435 20012 3477 20021
rect 3435 19972 3436 20012
rect 3476 19972 3477 20012
rect 3435 19963 3477 19972
rect 4395 20012 4437 20021
rect 4395 19972 4396 20012
rect 4436 19972 4437 20012
rect 4395 19963 4437 19972
rect 3339 18752 3381 18761
rect 3339 18712 3340 18752
rect 3380 18712 3381 18752
rect 3339 18703 3381 18712
rect 3339 18164 3381 18173
rect 3339 18124 3340 18164
rect 3380 18124 3381 18164
rect 3339 18115 3381 18124
rect 3243 17828 3285 17837
rect 3243 17788 3244 17828
rect 3284 17788 3285 17828
rect 3243 17779 3285 17788
rect 3244 17660 3284 17669
rect 3340 17660 3380 18115
rect 3284 17620 3380 17660
rect 3244 17611 3284 17620
rect 3243 17324 3285 17333
rect 3243 17284 3244 17324
rect 3284 17284 3285 17324
rect 3243 17275 3285 17284
rect 3148 17023 3188 17032
rect 3244 17072 3284 17275
rect 3345 17072 3385 17081
rect 3436 17072 3476 19963
rect 4396 19932 4436 19963
rect 4492 19962 4532 20047
rect 4588 19844 4628 22408
rect 5451 22280 5493 22289
rect 5451 22240 5452 22280
rect 5492 22240 5493 22280
rect 5451 22231 5493 22240
rect 4683 22112 4725 22121
rect 4683 22072 4684 22112
rect 4724 22072 4725 22112
rect 4683 22063 4725 22072
rect 4684 21608 4724 22063
rect 4779 22028 4821 22037
rect 4779 21988 4780 22028
rect 4820 21988 4821 22028
rect 4779 21979 4821 21988
rect 4684 21559 4724 21568
rect 4683 20936 4725 20945
rect 4683 20896 4684 20936
rect 4724 20896 4725 20936
rect 4683 20887 4725 20896
rect 4684 20768 4724 20887
rect 4684 20719 4724 20728
rect 4780 20180 4820 21979
rect 4928 21944 5296 21953
rect 4968 21904 5010 21944
rect 5050 21904 5092 21944
rect 5132 21904 5174 21944
rect 5214 21904 5256 21944
rect 4928 21895 5296 21904
rect 5163 21776 5205 21785
rect 5163 21736 5164 21776
rect 5204 21736 5205 21776
rect 5163 21727 5205 21736
rect 5164 21617 5204 21727
rect 5355 21692 5397 21701
rect 5355 21652 5356 21692
rect 5396 21652 5397 21692
rect 5355 21643 5397 21652
rect 5163 21608 5205 21617
rect 5163 21563 5164 21608
rect 5204 21563 5205 21608
rect 5163 21559 5205 21563
rect 5164 21104 5204 21559
rect 5356 21558 5396 21643
rect 5452 21440 5492 22231
rect 5548 21869 5588 26431
rect 5643 25472 5685 25481
rect 5643 25432 5644 25472
rect 5684 25432 5685 25472
rect 5643 25423 5685 25432
rect 5644 25136 5684 25423
rect 5644 25087 5684 25096
rect 5740 24977 5780 26608
rect 5836 25565 5876 27112
rect 5931 26732 5973 26741
rect 5931 26692 5932 26732
rect 5972 26692 5973 26732
rect 5931 26683 5973 26692
rect 5932 26598 5972 26683
rect 6028 26144 6068 28960
rect 6124 26480 6164 29791
rect 6316 29429 6356 31396
rect 6508 31352 6548 32395
rect 6604 31352 6644 32992
rect 6699 32864 6741 32873
rect 6699 32824 6700 32864
rect 6740 32824 6741 32864
rect 6699 32815 6741 32824
rect 6700 31520 6740 32815
rect 6796 32705 6836 34243
rect 7084 33965 7124 34341
rect 7083 33956 7125 33965
rect 7083 33916 7084 33956
rect 7124 33916 7125 33956
rect 7083 33907 7125 33916
rect 6988 33788 7028 33797
rect 7028 33748 7124 33788
rect 6988 33739 7028 33748
rect 6892 33704 6932 33715
rect 6892 33629 6932 33664
rect 6891 33620 6933 33629
rect 6891 33580 6892 33620
rect 6932 33580 6933 33620
rect 6891 33571 6933 33580
rect 7084 33125 7124 33748
rect 7083 33116 7125 33125
rect 7083 33076 7084 33116
rect 7124 33076 7125 33116
rect 7180 33116 7220 37015
rect 7275 36644 7317 36653
rect 7275 36604 7276 36644
rect 7316 36604 7317 36644
rect 7275 36595 7317 36604
rect 7276 36560 7316 36595
rect 7276 36509 7316 36520
rect 7275 34292 7317 34301
rect 7275 34252 7276 34292
rect 7316 34252 7317 34292
rect 7275 34243 7317 34252
rect 7276 34158 7316 34243
rect 7275 33956 7317 33965
rect 7275 33916 7276 33956
rect 7316 33916 7317 33956
rect 7275 33907 7317 33916
rect 7276 33713 7316 33907
rect 7275 33704 7317 33713
rect 7275 33664 7276 33704
rect 7316 33664 7317 33704
rect 7275 33655 7317 33664
rect 7275 33452 7317 33461
rect 7275 33412 7276 33452
rect 7316 33412 7317 33452
rect 7275 33403 7317 33412
rect 7276 33318 7316 33403
rect 7372 33293 7412 37528
rect 7468 37073 7508 37780
rect 7660 37780 7892 37820
rect 7564 37405 7604 37414
rect 7467 37064 7509 37073
rect 7467 37024 7468 37064
rect 7508 37024 7509 37064
rect 7467 37015 7509 37024
rect 7467 36728 7509 36737
rect 7467 36688 7468 36728
rect 7508 36688 7509 36728
rect 7467 36679 7509 36688
rect 7468 36594 7508 36679
rect 7564 36653 7604 37365
rect 7563 36644 7605 36653
rect 7563 36604 7564 36644
rect 7604 36604 7605 36644
rect 7563 36595 7605 36604
rect 7563 36476 7605 36485
rect 7563 36436 7564 36476
rect 7604 36436 7605 36476
rect 7563 36427 7605 36436
rect 7564 35813 7604 36427
rect 7563 35804 7605 35813
rect 7563 35764 7564 35804
rect 7604 35764 7605 35804
rect 7563 35755 7605 35764
rect 7468 34637 7508 34722
rect 7467 34628 7509 34637
rect 7467 34588 7468 34628
rect 7508 34588 7509 34628
rect 7467 34579 7509 34588
rect 7468 34376 7508 34385
rect 7468 33881 7508 34336
rect 7564 33965 7604 35755
rect 7563 33956 7605 33965
rect 7563 33916 7564 33956
rect 7604 33916 7605 33956
rect 7563 33907 7605 33916
rect 7467 33872 7509 33881
rect 7467 33832 7468 33872
rect 7508 33832 7509 33872
rect 7467 33823 7509 33832
rect 7467 33704 7509 33713
rect 7467 33664 7468 33704
rect 7508 33664 7509 33704
rect 7467 33655 7509 33664
rect 7564 33704 7604 33713
rect 7468 33570 7508 33655
rect 7564 33461 7604 33664
rect 7563 33452 7605 33461
rect 7563 33412 7564 33452
rect 7604 33412 7605 33452
rect 7563 33403 7605 33412
rect 7371 33284 7413 33293
rect 7371 33244 7372 33284
rect 7412 33244 7413 33284
rect 7371 33235 7413 33244
rect 7180 33076 7316 33116
rect 7083 33067 7125 33076
rect 6795 32696 6837 32705
rect 6795 32656 6796 32696
rect 6836 32656 6837 32696
rect 6795 32647 6837 32656
rect 6796 32192 6836 32647
rect 6892 32192 6932 32201
rect 6796 32152 6892 32192
rect 6892 32143 6932 32152
rect 6891 31856 6933 31865
rect 6891 31816 6892 31856
rect 6932 31816 6933 31856
rect 6891 31807 6933 31816
rect 6892 31613 6932 31807
rect 6891 31604 6933 31613
rect 6891 31564 6892 31604
rect 6932 31564 6933 31604
rect 6891 31555 6933 31564
rect 6700 31471 6740 31480
rect 6699 31352 6741 31361
rect 6604 31312 6700 31352
rect 6740 31312 6741 31352
rect 6508 31303 6548 31312
rect 6699 31303 6741 31312
rect 6892 31352 6932 31555
rect 6892 31303 6932 31312
rect 6700 31218 6740 31303
rect 7084 31193 7124 33067
rect 7179 32948 7221 32957
rect 7179 32908 7180 32948
rect 7220 32908 7221 32948
rect 7179 32899 7221 32908
rect 7083 31184 7125 31193
rect 7083 31144 7084 31184
rect 7124 31144 7125 31184
rect 7083 31135 7125 31144
rect 7084 30680 7124 30691
rect 7084 30605 7124 30640
rect 7083 30596 7125 30605
rect 7083 30556 7084 30596
rect 7124 30556 7125 30596
rect 7083 30547 7125 30556
rect 6411 30260 6453 30269
rect 6411 30220 6412 30260
rect 6452 30220 6453 30260
rect 6411 30211 6453 30220
rect 6987 30260 7029 30269
rect 6987 30220 6988 30260
rect 7028 30220 7029 30260
rect 6987 30211 7029 30220
rect 6412 29849 6452 30211
rect 6411 29840 6453 29849
rect 6411 29800 6412 29840
rect 6452 29800 6453 29840
rect 6411 29791 6453 29800
rect 6315 29420 6357 29429
rect 6315 29380 6316 29420
rect 6356 29380 6357 29420
rect 6315 29371 6357 29380
rect 6412 29168 6452 29791
rect 6604 29252 6644 29261
rect 6644 29212 6932 29252
rect 6604 29203 6644 29212
rect 6412 29009 6452 29128
rect 6892 29168 6932 29212
rect 6988 29177 7028 30211
rect 7084 29840 7124 29849
rect 7180 29840 7220 32899
rect 7276 32864 7316 33076
rect 7660 32957 7700 37780
rect 7851 37568 7893 37577
rect 7851 37528 7852 37568
rect 7892 37528 7893 37568
rect 7851 37519 7893 37528
rect 7755 37232 7797 37241
rect 7755 37192 7756 37232
rect 7796 37192 7797 37232
rect 7755 37183 7797 37192
rect 7756 37098 7796 37183
rect 7852 37157 7892 37519
rect 7851 37148 7893 37157
rect 7851 37108 7852 37148
rect 7892 37108 7893 37148
rect 7851 37099 7893 37108
rect 8140 36056 8180 38872
rect 7852 36016 8180 36056
rect 7852 35888 7892 36016
rect 8236 35972 8276 42484
rect 8332 39005 8372 51631
rect 8427 49412 8469 49421
rect 8427 49372 8428 49412
rect 8468 49372 8469 49412
rect 8427 49363 8469 49372
rect 8428 47984 8468 49363
rect 8428 47935 8468 47944
rect 8524 43532 8564 52219
rect 8620 51848 8660 51857
rect 8620 51689 8660 51808
rect 8619 51680 8661 51689
rect 8619 51640 8620 51680
rect 8660 51640 8661 51680
rect 8619 51631 8661 51640
rect 8619 51260 8661 51269
rect 8619 51220 8620 51260
rect 8660 51220 8661 51260
rect 8619 51211 8661 51220
rect 8620 51008 8660 51211
rect 8620 50959 8660 50968
rect 8812 50504 8852 54328
rect 9100 54284 9140 56596
rect 9196 56468 9236 56477
rect 9388 56468 9428 57856
rect 9484 57847 9524 57856
rect 9579 57896 9621 57905
rect 9579 57856 9580 57896
rect 9620 57856 9621 57896
rect 9579 57847 9621 57856
rect 9580 57569 9620 57847
rect 9579 57560 9621 57569
rect 9579 57520 9580 57560
rect 9620 57520 9621 57560
rect 9579 57511 9621 57520
rect 9675 57140 9717 57149
rect 9675 57100 9676 57140
rect 9716 57100 9717 57140
rect 9675 57091 9717 57100
rect 9676 57006 9716 57091
rect 9772 57056 9812 58267
rect 9868 57485 9908 59527
rect 9964 58745 10004 62056
rect 10059 59828 10101 59837
rect 10059 59788 10060 59828
rect 10100 59788 10101 59828
rect 10059 59779 10101 59788
rect 9963 58736 10005 58745
rect 9963 58696 9964 58736
rect 10004 58696 10005 58736
rect 9963 58687 10005 58696
rect 9963 58400 10005 58409
rect 9963 58360 9964 58400
rect 10004 58360 10005 58400
rect 9963 58351 10005 58360
rect 9964 57891 10004 58351
rect 9964 57842 10004 57851
rect 9867 57476 9909 57485
rect 9867 57436 9868 57476
rect 9908 57436 9909 57476
rect 9867 57427 9909 57436
rect 9868 57056 9908 57065
rect 9772 57016 9868 57056
rect 9236 56428 9428 56468
rect 9484 56888 9524 56897
rect 9196 56141 9236 56428
rect 9291 56300 9333 56309
rect 9291 56260 9292 56300
rect 9332 56260 9333 56300
rect 9291 56251 9333 56260
rect 9195 56132 9237 56141
rect 9195 56092 9196 56132
rect 9236 56092 9237 56132
rect 9195 56083 9237 56092
rect 9195 54872 9237 54881
rect 9195 54832 9196 54872
rect 9236 54832 9237 54872
rect 9292 54872 9332 56251
rect 9484 56225 9524 56848
rect 9483 56216 9525 56225
rect 9483 56176 9484 56216
rect 9524 56176 9525 56216
rect 9483 56167 9525 56176
rect 9579 56048 9621 56057
rect 9579 56008 9580 56048
rect 9620 56008 9621 56048
rect 9579 55999 9621 56008
rect 9484 55549 9524 55558
rect 9388 55040 9428 55049
rect 9484 55040 9524 55509
rect 9428 55000 9524 55040
rect 9580 55040 9620 55999
rect 9675 55712 9717 55721
rect 9675 55672 9676 55712
rect 9716 55672 9717 55712
rect 9675 55663 9717 55672
rect 9676 55460 9716 55663
rect 9868 55553 9908 57016
rect 10060 55796 10100 59779
rect 10156 59249 10196 62383
rect 10251 62264 10293 62273
rect 10251 62224 10252 62264
rect 10292 62224 10293 62264
rect 10251 62215 10293 62224
rect 10252 60920 10292 62215
rect 10252 60080 10292 60880
rect 10443 60500 10485 60509
rect 10443 60460 10444 60500
rect 10484 60460 10485 60500
rect 10443 60451 10485 60460
rect 10155 59240 10197 59249
rect 10155 59200 10156 59240
rect 10196 59200 10197 59240
rect 10155 59191 10197 59200
rect 10252 59072 10292 60040
rect 10347 59912 10389 59921
rect 10347 59872 10348 59912
rect 10388 59872 10389 59912
rect 10347 59863 10389 59872
rect 10156 59032 10292 59072
rect 10156 58157 10196 59032
rect 10252 58568 10292 58577
rect 10155 58148 10197 58157
rect 10155 58108 10156 58148
rect 10196 58108 10197 58148
rect 10155 58099 10197 58108
rect 10156 57980 10196 57989
rect 10156 57149 10196 57940
rect 10252 57821 10292 58528
rect 10251 57812 10293 57821
rect 10251 57772 10252 57812
rect 10292 57772 10293 57812
rect 10251 57763 10293 57772
rect 10348 57644 10388 59863
rect 10444 59417 10484 60451
rect 10443 59408 10485 59417
rect 10443 59368 10444 59408
rect 10484 59368 10485 59408
rect 10443 59359 10485 59368
rect 10443 58400 10485 58409
rect 10443 58360 10444 58400
rect 10484 58360 10485 58400
rect 10443 58351 10485 58360
rect 10444 58266 10484 58351
rect 10540 58148 10580 62392
rect 10732 61004 10772 62887
rect 10828 62886 10868 62971
rect 10924 62970 10964 63055
rect 11212 63054 11252 63139
rect 11211 62936 11253 62945
rect 11211 62896 11212 62936
rect 11252 62896 11253 62936
rect 11211 62887 11253 62896
rect 10923 61676 10965 61685
rect 10923 61636 10924 61676
rect 10964 61636 10965 61676
rect 10923 61627 10965 61636
rect 10924 61592 10964 61627
rect 11212 61601 11252 62887
rect 10924 61541 10964 61552
rect 11211 61592 11253 61601
rect 11211 61552 11212 61592
rect 11252 61552 11253 61592
rect 11211 61543 11253 61552
rect 11116 61424 11156 61433
rect 11116 61256 11156 61384
rect 10636 60964 10772 61004
rect 10828 61216 11156 61256
rect 10636 58241 10676 60964
rect 10828 60920 10868 61216
rect 10923 61088 10965 61097
rect 10923 61048 10924 61088
rect 10964 61048 10965 61088
rect 10923 61039 10965 61048
rect 11115 61088 11157 61097
rect 11115 61048 11116 61088
rect 11156 61048 11157 61088
rect 11115 61039 11157 61048
rect 10924 60954 10964 61039
rect 11116 60920 11156 61039
rect 10780 60910 10868 60920
rect 10820 60880 10868 60910
rect 11020 60880 11116 60920
rect 10780 60861 10820 60870
rect 10923 60752 10965 60761
rect 10923 60712 10924 60752
rect 10964 60712 10965 60752
rect 10923 60703 10965 60712
rect 10732 60089 10772 60175
rect 10924 60173 10964 60703
rect 10923 60164 10965 60173
rect 10923 60124 10924 60164
rect 10964 60124 10965 60164
rect 10923 60115 10965 60124
rect 10731 60040 10732 60089
rect 10772 60040 10773 60089
rect 10731 60031 10773 60040
rect 10827 59996 10869 60005
rect 10827 59956 10828 59996
rect 10868 59956 10869 59996
rect 10827 59947 10869 59956
rect 10828 59576 10868 59947
rect 10923 59912 10965 59921
rect 10923 59872 10924 59912
rect 10964 59872 10965 59912
rect 10923 59863 10965 59872
rect 10924 59778 10964 59863
rect 10924 59576 10964 59585
rect 10828 59536 10924 59576
rect 10924 59527 10964 59536
rect 10731 59408 10773 59417
rect 10731 59368 10732 59408
rect 10772 59368 10964 59408
rect 10731 59359 10773 59368
rect 10732 59274 10772 59359
rect 10635 58232 10677 58241
rect 10635 58192 10636 58232
rect 10676 58192 10677 58232
rect 10635 58183 10677 58192
rect 10252 57604 10388 57644
rect 10444 58108 10580 58148
rect 10155 57140 10197 57149
rect 10155 57100 10156 57140
rect 10196 57100 10197 57140
rect 10155 57091 10197 57100
rect 10060 55756 10196 55796
rect 9963 55712 10005 55721
rect 9963 55672 9964 55712
rect 10004 55672 10100 55712
rect 9963 55663 10005 55672
rect 10060 55639 10100 55672
rect 10060 55590 10100 55599
rect 9867 55544 9909 55553
rect 9867 55504 9868 55544
rect 9908 55504 9909 55544
rect 9867 55495 9909 55504
rect 9676 55411 9716 55420
rect 9868 55376 9908 55387
rect 9868 55301 9908 55336
rect 9867 55292 9909 55301
rect 9867 55252 9868 55292
rect 9908 55252 9909 55292
rect 9867 55243 9909 55252
rect 10156 55133 10196 55756
rect 9867 55124 9909 55133
rect 9867 55084 9868 55124
rect 9908 55084 9909 55124
rect 9867 55075 9909 55084
rect 10155 55124 10197 55133
rect 10155 55084 10156 55124
rect 10196 55084 10197 55124
rect 10155 55075 10197 55084
rect 9580 55000 9716 55040
rect 9388 54991 9428 55000
rect 9580 54872 9620 54881
rect 9292 54832 9580 54872
rect 9195 54823 9237 54832
rect 8716 50464 8852 50504
rect 8908 54244 9140 54284
rect 8716 50261 8756 50464
rect 8812 50336 8852 50345
rect 8715 50252 8757 50261
rect 8715 50212 8716 50252
rect 8756 50212 8757 50252
rect 8715 50203 8757 50212
rect 8812 50009 8852 50296
rect 8811 50000 8853 50009
rect 8811 49960 8812 50000
rect 8852 49960 8853 50000
rect 8811 49951 8853 49960
rect 8715 49580 8757 49589
rect 8715 49540 8716 49580
rect 8756 49540 8757 49580
rect 8715 49531 8757 49540
rect 8619 49496 8661 49505
rect 8619 49456 8620 49496
rect 8660 49456 8661 49496
rect 8619 49447 8661 49456
rect 8716 49496 8756 49531
rect 8908 49505 8948 54244
rect 9099 53360 9141 53369
rect 9099 53315 9100 53360
rect 9140 53315 9141 53360
rect 9099 53311 9141 53315
rect 9100 53225 9140 53311
rect 9196 53285 9236 54823
rect 9291 53528 9333 53537
rect 9291 53488 9292 53528
rect 9332 53488 9333 53528
rect 9291 53479 9333 53488
rect 9292 53394 9332 53479
rect 9195 53276 9237 53285
rect 9388 53276 9428 54832
rect 9580 54823 9620 54832
rect 9580 54032 9620 54043
rect 9580 53957 9620 53992
rect 9579 53948 9621 53957
rect 9579 53908 9580 53948
rect 9620 53908 9621 53948
rect 9579 53899 9621 53908
rect 9195 53236 9196 53276
rect 9236 53236 9237 53276
rect 9195 53227 9237 53236
rect 9292 53236 9428 53276
rect 9484 53360 9524 53369
rect 9676 53360 9716 55000
rect 9772 53864 9812 53873
rect 9772 53369 9812 53824
rect 9524 53320 9716 53360
rect 9771 53360 9813 53369
rect 9771 53320 9772 53360
rect 9812 53320 9813 53360
rect 9292 51689 9332 53236
rect 9387 51764 9429 51773
rect 9387 51724 9388 51764
rect 9428 51724 9429 51764
rect 9387 51715 9429 51724
rect 9291 51680 9333 51689
rect 9291 51640 9292 51680
rect 9332 51640 9333 51680
rect 9291 51631 9333 51640
rect 9195 51344 9237 51353
rect 9195 51304 9196 51344
rect 9236 51304 9237 51344
rect 9195 51295 9237 51304
rect 9100 51013 9140 51022
rect 9004 50504 9044 50513
rect 9100 50504 9140 50973
rect 9044 50464 9140 50504
rect 9004 50455 9044 50464
rect 9196 50336 9236 51295
rect 9291 51092 9333 51101
rect 9291 51052 9292 51092
rect 9332 51052 9333 51092
rect 9291 51043 9333 51052
rect 9292 50924 9332 51043
rect 9292 50875 9332 50884
rect 9196 50287 9236 50296
rect 9388 50252 9428 51715
rect 9292 50212 9428 50252
rect 8620 46481 8660 49447
rect 8716 46640 8756 49456
rect 8907 49496 8949 49505
rect 8907 49456 8908 49496
rect 8948 49456 8949 49496
rect 8907 49447 8949 49456
rect 8908 49328 8948 49337
rect 8812 49288 8908 49328
rect 8812 48824 8852 49288
rect 8908 49279 8948 49288
rect 8812 48775 8852 48784
rect 8907 48824 8949 48833
rect 8907 48784 8908 48824
rect 8948 48784 8949 48824
rect 8907 48775 8949 48784
rect 9099 48824 9141 48833
rect 9099 48784 9100 48824
rect 9140 48784 9141 48824
rect 9099 48775 9141 48784
rect 9292 48824 9332 50212
rect 9292 48775 9332 48784
rect 9387 48824 9429 48833
rect 9387 48784 9388 48824
rect 9428 48784 9429 48824
rect 9387 48775 9429 48784
rect 8908 48690 8948 48775
rect 9003 48236 9045 48245
rect 9003 48196 9004 48236
rect 9044 48196 9045 48236
rect 9003 48187 9045 48196
rect 8907 48152 8949 48161
rect 8907 48112 8908 48152
rect 8948 48112 8949 48152
rect 8907 48103 8949 48112
rect 8908 48068 8948 48103
rect 8908 48017 8948 48028
rect 9004 48068 9044 48187
rect 9004 48019 9044 48028
rect 9003 47816 9045 47825
rect 9003 47776 9004 47816
rect 9044 47776 9045 47816
rect 9003 47767 9045 47776
rect 8716 46600 8948 46640
rect 8619 46472 8661 46481
rect 8619 46432 8620 46472
rect 8660 46432 8661 46472
rect 8619 46423 8661 46432
rect 8908 46229 8948 46600
rect 8907 46220 8949 46229
rect 8907 46180 8908 46220
rect 8948 46180 8949 46220
rect 8907 46171 8949 46180
rect 8811 46052 8853 46061
rect 8811 46012 8812 46052
rect 8852 46012 8853 46052
rect 8811 46003 8853 46012
rect 8812 45221 8852 46003
rect 8811 45212 8853 45221
rect 8811 45172 8812 45212
rect 8852 45172 8853 45212
rect 8811 45163 8853 45172
rect 8908 44120 8948 46171
rect 9004 45053 9044 47767
rect 9003 45044 9045 45053
rect 9003 45004 9004 45044
rect 9044 45004 9045 45044
rect 9003 44995 9045 45004
rect 8812 44080 8948 44120
rect 8812 43541 8852 44080
rect 9004 44036 9044 44045
rect 8908 43996 9004 44036
rect 8524 43483 8564 43492
rect 8811 43532 8853 43541
rect 8811 43492 8812 43532
rect 8852 43492 8853 43532
rect 8811 43483 8853 43492
rect 8428 43448 8468 43459
rect 8428 43373 8468 43408
rect 8427 43364 8469 43373
rect 8427 43324 8428 43364
rect 8468 43324 8469 43364
rect 8427 43315 8469 43324
rect 8908 43205 8948 43996
rect 9004 43987 9044 43996
rect 9004 43448 9044 43457
rect 9004 43289 9044 43408
rect 9003 43280 9045 43289
rect 9003 43240 9004 43280
rect 9044 43240 9045 43280
rect 9003 43231 9045 43240
rect 8907 43196 8949 43205
rect 8907 43156 8908 43196
rect 8948 43156 8949 43196
rect 8907 43147 8949 43156
rect 8811 42104 8853 42113
rect 8811 42064 8812 42104
rect 8852 42064 8853 42104
rect 8811 42055 8853 42064
rect 8812 41936 8852 42055
rect 9100 42020 9140 48775
rect 9388 48690 9428 48775
rect 9484 48572 9524 53320
rect 9771 53311 9813 53320
rect 9868 52016 9908 55075
rect 9963 54200 10005 54209
rect 9963 54160 9964 54200
rect 10004 54160 10005 54200
rect 9963 54151 10005 54160
rect 9964 54116 10004 54151
rect 9964 54065 10004 54076
rect 10059 54032 10101 54041
rect 10059 53992 10060 54032
rect 10100 53992 10101 54032
rect 10059 53983 10101 53992
rect 9963 53276 10005 53285
rect 9963 53236 9964 53276
rect 10004 53236 10005 53276
rect 9963 53227 10005 53236
rect 9772 51976 9908 52016
rect 9579 51680 9621 51689
rect 9579 51640 9580 51680
rect 9620 51640 9621 51680
rect 9579 51631 9621 51640
rect 9292 48532 9524 48572
rect 9292 47825 9332 48532
rect 9387 48068 9429 48077
rect 9387 48028 9388 48068
rect 9428 48028 9429 48068
rect 9387 48019 9429 48028
rect 9388 47984 9428 48019
rect 9388 47933 9428 47944
rect 9483 47984 9525 47993
rect 9483 47944 9484 47984
rect 9524 47944 9525 47984
rect 9483 47935 9525 47944
rect 9484 47850 9524 47935
rect 9291 47816 9333 47825
rect 9291 47776 9292 47816
rect 9332 47776 9333 47816
rect 9291 47767 9333 47776
rect 9484 47312 9524 47321
rect 9196 47272 9484 47312
rect 9196 45977 9236 47272
rect 9484 47263 9524 47272
rect 9580 46640 9620 51631
rect 9292 46600 9620 46640
rect 9195 45968 9237 45977
rect 9195 45928 9196 45968
rect 9236 45928 9237 45968
rect 9195 45919 9237 45928
rect 9195 44960 9237 44969
rect 9195 44920 9196 44960
rect 9236 44920 9237 44960
rect 9195 44911 9237 44920
rect 9196 44826 9236 44911
rect 9196 44204 9236 44213
rect 9196 43784 9236 44164
rect 9292 43961 9332 46600
rect 9388 46472 9428 46481
rect 9388 46229 9428 46432
rect 9483 46472 9525 46481
rect 9483 46432 9484 46472
rect 9524 46432 9525 46472
rect 9483 46423 9525 46432
rect 9387 46220 9429 46229
rect 9387 46180 9388 46220
rect 9428 46180 9429 46220
rect 9387 46171 9429 46180
rect 9484 46136 9524 46423
rect 9580 46313 9620 46398
rect 9579 46304 9621 46313
rect 9579 46264 9580 46304
rect 9620 46264 9621 46304
rect 9579 46255 9621 46264
rect 9675 46220 9717 46229
rect 9675 46180 9676 46220
rect 9716 46180 9717 46220
rect 9675 46171 9717 46180
rect 9484 46096 9620 46136
rect 9484 45800 9524 45809
rect 9388 45212 9428 45221
rect 9484 45212 9524 45760
rect 9428 45172 9524 45212
rect 9580 45800 9620 46096
rect 9676 45893 9716 46171
rect 9675 45884 9717 45893
rect 9675 45844 9676 45884
rect 9716 45844 9717 45884
rect 9675 45835 9717 45844
rect 9388 45163 9428 45172
rect 9580 45128 9620 45760
rect 9484 45088 9620 45128
rect 9484 44045 9524 45088
rect 9580 44960 9620 44969
rect 9676 44960 9716 45835
rect 9620 44920 9716 44960
rect 9580 44911 9620 44920
rect 9675 44456 9717 44465
rect 9675 44416 9676 44456
rect 9716 44416 9717 44456
rect 9675 44407 9717 44416
rect 9676 44322 9716 44407
rect 9483 44036 9525 44045
rect 9483 43996 9484 44036
rect 9524 43996 9525 44036
rect 9483 43987 9525 43996
rect 9291 43952 9333 43961
rect 9291 43912 9292 43952
rect 9332 43912 9333 43952
rect 9291 43903 9333 43912
rect 9772 43877 9812 51976
rect 9868 51848 9908 51857
rect 9964 51848 10004 53227
rect 9908 51808 10004 51848
rect 9868 51605 9908 51808
rect 10060 51764 10100 53983
rect 10155 53864 10197 53873
rect 10155 53824 10156 53864
rect 10196 53824 10197 53864
rect 10155 53815 10197 53824
rect 10156 53730 10196 53815
rect 10252 52016 10292 57604
rect 10347 57476 10389 57485
rect 10347 57436 10348 57476
rect 10388 57436 10389 57476
rect 10347 57427 10389 57436
rect 10348 56300 10388 57427
rect 10348 56251 10388 56260
rect 10347 55964 10389 55973
rect 10347 55924 10348 55964
rect 10388 55924 10389 55964
rect 10347 55915 10389 55924
rect 10348 54209 10388 55915
rect 10444 54881 10484 58108
rect 10636 56384 10676 58183
rect 10732 56384 10772 56393
rect 10636 56344 10732 56384
rect 10539 56132 10581 56141
rect 10539 56092 10540 56132
rect 10580 56092 10581 56132
rect 10539 56083 10581 56092
rect 10540 55998 10580 56083
rect 10636 55973 10676 56344
rect 10732 56335 10772 56344
rect 10635 55964 10677 55973
rect 10635 55924 10636 55964
rect 10676 55924 10677 55964
rect 10635 55915 10677 55924
rect 10540 55756 10868 55796
rect 10443 54872 10485 54881
rect 10443 54832 10444 54872
rect 10484 54832 10485 54872
rect 10443 54823 10485 54832
rect 10347 54200 10389 54209
rect 10347 54160 10348 54200
rect 10388 54160 10389 54200
rect 10347 54151 10389 54160
rect 10347 54032 10389 54041
rect 10347 53992 10348 54032
rect 10388 53992 10389 54032
rect 10347 53983 10389 53992
rect 10348 53898 10388 53983
rect 10347 53108 10389 53117
rect 10347 53068 10348 53108
rect 10388 53068 10389 53108
rect 10347 53059 10389 53068
rect 10348 52520 10388 53059
rect 10348 52471 10388 52480
rect 10444 52520 10484 52529
rect 10540 52520 10580 55756
rect 10732 55553 10772 55638
rect 10731 55544 10773 55553
rect 10731 55504 10732 55544
rect 10772 55504 10773 55544
rect 10731 55495 10773 55504
rect 10828 55544 10868 55756
rect 10828 55495 10868 55504
rect 10924 55376 10964 59368
rect 11020 58913 11060 60880
rect 11116 60871 11156 60880
rect 11212 60761 11252 61543
rect 11211 60752 11253 60761
rect 11211 60712 11212 60752
rect 11252 60712 11253 60752
rect 11211 60703 11253 60712
rect 11308 60332 11348 63316
rect 11404 63281 11444 64576
rect 11403 63272 11445 63281
rect 11403 63232 11404 63272
rect 11444 63232 11445 63272
rect 11403 63223 11445 63232
rect 11500 62600 11540 65920
rect 11596 62861 11636 69280
rect 11787 69280 11788 69320
rect 11828 69280 11829 69320
rect 11787 69271 11829 69280
rect 11692 68984 11732 68995
rect 11692 68909 11732 68944
rect 11691 68900 11733 68909
rect 11691 68860 11692 68900
rect 11732 68860 11733 68900
rect 11691 68851 11733 68860
rect 11788 68741 11828 69271
rect 11787 68732 11829 68741
rect 11787 68692 11788 68732
rect 11828 68692 11829 68732
rect 11787 68683 11829 68692
rect 11787 67808 11829 67817
rect 11787 67768 11788 67808
rect 11828 67768 11829 67808
rect 11787 67759 11829 67768
rect 11691 67220 11733 67229
rect 11691 67180 11692 67220
rect 11732 67180 11733 67220
rect 11691 67171 11733 67180
rect 11692 67136 11732 67171
rect 11692 67085 11732 67096
rect 11788 66977 11828 67759
rect 11787 66968 11829 66977
rect 11692 66928 11788 66968
rect 11828 66928 11829 66968
rect 11692 66221 11732 66928
rect 11787 66919 11829 66928
rect 11787 66800 11829 66809
rect 11787 66760 11788 66800
rect 11828 66760 11829 66800
rect 11787 66751 11829 66760
rect 11788 66641 11828 66751
rect 11787 66632 11829 66641
rect 11787 66592 11788 66632
rect 11828 66592 11829 66632
rect 11787 66583 11829 66592
rect 11691 66212 11733 66221
rect 11691 66172 11692 66212
rect 11732 66172 11733 66212
rect 11691 66163 11733 66172
rect 11691 66044 11733 66053
rect 11691 66004 11692 66044
rect 11732 66004 11733 66044
rect 11691 65995 11733 66004
rect 11595 62852 11637 62861
rect 11595 62812 11596 62852
rect 11636 62812 11637 62852
rect 11595 62803 11637 62812
rect 11692 62684 11732 65995
rect 11788 64700 11828 66583
rect 11884 66557 11924 70111
rect 11980 69749 12020 70624
rect 12076 69908 12116 85231
rect 12172 77636 12212 85936
rect 12364 83105 12404 85936
rect 12363 83096 12405 83105
rect 12363 83056 12364 83096
rect 12404 83056 12405 83096
rect 12363 83047 12405 83056
rect 12172 77596 12404 77636
rect 12364 76889 12404 77596
rect 12363 76880 12405 76889
rect 12363 76840 12364 76880
rect 12404 76840 12405 76880
rect 12363 76831 12405 76840
rect 12556 76208 12596 85936
rect 12748 77552 12788 85936
rect 12940 84449 12980 85936
rect 12939 84440 12981 84449
rect 12939 84400 12940 84440
rect 12980 84400 12981 84440
rect 12939 84391 12981 84400
rect 13132 83516 13172 85936
rect 13324 84449 13364 85936
rect 13516 85625 13556 85936
rect 13515 85616 13557 85625
rect 13515 85576 13516 85616
rect 13556 85576 13557 85616
rect 13515 85567 13557 85576
rect 13708 84533 13748 85936
rect 13707 84524 13749 84533
rect 13707 84484 13708 84524
rect 13748 84484 13749 84524
rect 13707 84475 13749 84484
rect 13900 84449 13940 85936
rect 14092 85912 14142 85936
rect 14102 85868 14142 85912
rect 14092 85828 14142 85868
rect 14092 84944 14132 85828
rect 13996 84904 14132 84944
rect 13323 84440 13365 84449
rect 13323 84400 13324 84440
rect 13364 84400 13365 84440
rect 13323 84391 13365 84400
rect 13899 84440 13941 84449
rect 13899 84400 13900 84440
rect 13940 84400 13941 84440
rect 13899 84391 13941 84400
rect 13996 84281 14036 84904
rect 14091 84776 14133 84785
rect 14091 84736 14092 84776
rect 14132 84736 14133 84776
rect 14091 84727 14133 84736
rect 13323 84272 13365 84281
rect 13323 84232 13324 84272
rect 13364 84232 13365 84272
rect 13323 84223 13365 84232
rect 13995 84272 14037 84281
rect 13995 84232 13996 84272
rect 14036 84232 14037 84272
rect 13995 84223 14037 84232
rect 13036 83476 13172 83516
rect 13324 83516 13364 84223
rect 13995 83600 14037 83609
rect 13995 83560 13996 83600
rect 14036 83560 14037 83600
rect 13995 83551 14037 83560
rect 13036 81929 13076 83476
rect 13324 83467 13364 83476
rect 13707 83516 13749 83525
rect 13707 83476 13708 83516
rect 13748 83476 13749 83516
rect 13707 83467 13749 83476
rect 13708 83382 13748 83467
rect 13131 83348 13173 83357
rect 13131 83308 13132 83348
rect 13172 83308 13173 83348
rect 13131 83299 13173 83308
rect 13516 83348 13556 83357
rect 13132 83214 13172 83299
rect 13516 83189 13556 83308
rect 13899 83348 13941 83357
rect 13899 83308 13900 83348
rect 13940 83308 13941 83348
rect 13899 83299 13941 83308
rect 13900 83214 13940 83299
rect 13515 83180 13557 83189
rect 13515 83140 13516 83180
rect 13556 83140 13557 83180
rect 13515 83131 13557 83140
rect 13035 81920 13077 81929
rect 13035 81880 13036 81920
rect 13076 81880 13077 81920
rect 13035 81871 13077 81880
rect 12748 77512 13076 77552
rect 12843 76880 12885 76889
rect 12843 76840 12844 76880
rect 12884 76840 12885 76880
rect 12843 76831 12885 76840
rect 12172 76168 12596 76208
rect 12172 73940 12212 76168
rect 12460 76040 12500 76049
rect 12268 76000 12460 76040
rect 12268 74024 12308 76000
rect 12460 75991 12500 76000
rect 12412 75209 12452 75218
rect 12452 75169 12788 75200
rect 12412 75160 12788 75169
rect 12556 75032 12596 75041
rect 12596 74992 12692 75032
rect 12556 74983 12596 74992
rect 12555 74696 12597 74705
rect 12555 74656 12556 74696
rect 12596 74656 12597 74696
rect 12555 74647 12597 74656
rect 12556 74528 12596 74647
rect 12556 74479 12596 74488
rect 12268 73984 12596 74024
rect 12172 73900 12500 73940
rect 12267 73688 12309 73697
rect 12267 73648 12268 73688
rect 12308 73648 12309 73688
rect 12267 73639 12309 73648
rect 12268 73554 12308 73639
rect 12171 73016 12213 73025
rect 12171 72976 12172 73016
rect 12212 72976 12213 73016
rect 12171 72967 12213 72976
rect 12172 72882 12212 72967
rect 12363 72764 12405 72773
rect 12363 72724 12364 72764
rect 12404 72724 12405 72764
rect 12363 72715 12405 72724
rect 12364 72630 12404 72715
rect 12460 72344 12500 73900
rect 12268 72304 12500 72344
rect 12171 71504 12213 71513
rect 12171 71464 12172 71504
rect 12212 71464 12213 71504
rect 12171 71455 12213 71464
rect 12172 71370 12212 71455
rect 12171 70496 12213 70505
rect 12171 70456 12172 70496
rect 12212 70456 12213 70496
rect 12171 70447 12213 70456
rect 12172 70362 12212 70447
rect 12076 69833 12116 69868
rect 12171 69908 12213 69917
rect 12171 69868 12172 69908
rect 12212 69868 12213 69908
rect 12171 69859 12213 69868
rect 12075 69824 12117 69833
rect 12075 69784 12076 69824
rect 12116 69784 12117 69824
rect 12075 69775 12117 69784
rect 12172 69774 12212 69859
rect 11979 69740 12021 69749
rect 11979 69700 11980 69740
rect 12020 69700 12021 69740
rect 11979 69691 12021 69700
rect 11980 69152 12020 69161
rect 12020 69112 12116 69152
rect 11980 69103 12020 69112
rect 11979 68732 12021 68741
rect 11979 68692 11980 68732
rect 12020 68692 12021 68732
rect 11979 68683 12021 68692
rect 11980 67640 12020 68683
rect 12076 68489 12116 69112
rect 12075 68480 12117 68489
rect 12075 68440 12076 68480
rect 12116 68440 12117 68480
rect 12075 68431 12117 68440
rect 12076 68153 12116 68431
rect 12075 68144 12117 68153
rect 12075 68104 12076 68144
rect 12116 68104 12117 68144
rect 12075 68095 12117 68104
rect 12076 67640 12116 67649
rect 11980 67600 12076 67640
rect 11883 66548 11925 66557
rect 11883 66508 11884 66548
rect 11924 66508 11925 66548
rect 11883 66499 11925 66508
rect 11883 66212 11925 66221
rect 11883 66172 11884 66212
rect 11924 66172 11925 66212
rect 11883 66163 11925 66172
rect 11884 65381 11924 66163
rect 11883 65372 11925 65381
rect 11883 65332 11884 65372
rect 11924 65332 11925 65372
rect 11883 65323 11925 65332
rect 11788 64651 11828 64660
rect 11883 64700 11925 64709
rect 11883 64660 11884 64700
rect 11924 64660 11925 64700
rect 11883 64651 11925 64660
rect 11884 64566 11924 64651
rect 11980 64280 12020 67600
rect 12076 67591 12116 67600
rect 12075 66968 12117 66977
rect 12075 66928 12076 66968
rect 12116 66928 12117 66968
rect 12075 66919 12117 66928
rect 12172 66968 12212 66977
rect 12076 66834 12116 66919
rect 12172 66809 12212 66928
rect 12171 66800 12213 66809
rect 12171 66760 12172 66800
rect 12212 66760 12213 66800
rect 12171 66751 12213 66760
rect 12171 66548 12213 66557
rect 12171 66508 12172 66548
rect 12212 66508 12213 66548
rect 12171 66499 12213 66508
rect 11884 64240 12020 64280
rect 11787 62852 11829 62861
rect 11787 62812 11788 62852
rect 11828 62812 11829 62852
rect 11787 62803 11829 62812
rect 11116 60292 11348 60332
rect 11404 62560 11540 62600
rect 11596 62644 11732 62684
rect 11019 58904 11061 58913
rect 11019 58864 11020 58904
rect 11060 58864 11061 58904
rect 11019 58855 11061 58864
rect 11019 58736 11061 58745
rect 11019 58696 11020 58736
rect 11060 58696 11061 58736
rect 11019 58687 11061 58696
rect 11020 57989 11060 58687
rect 11116 58568 11156 60292
rect 11211 60164 11253 60173
rect 11211 60124 11212 60164
rect 11252 60124 11253 60164
rect 11211 60115 11253 60124
rect 11212 58913 11252 60115
rect 11308 59408 11348 59419
rect 11308 59333 11348 59368
rect 11307 59324 11349 59333
rect 11307 59284 11308 59324
rect 11348 59284 11349 59324
rect 11307 59275 11349 59284
rect 11211 58904 11253 58913
rect 11211 58864 11212 58904
rect 11252 58864 11253 58904
rect 11211 58855 11253 58864
rect 11116 58409 11156 58528
rect 11115 58400 11157 58409
rect 11115 58360 11116 58400
rect 11156 58360 11157 58400
rect 11115 58351 11157 58360
rect 11019 57980 11061 57989
rect 11019 57940 11020 57980
rect 11060 57940 11061 57980
rect 11019 57931 11061 57940
rect 11020 57056 11060 57931
rect 11116 57056 11156 57065
rect 11020 57016 11116 57056
rect 11020 56309 11060 57016
rect 11116 57007 11156 57016
rect 11212 56813 11252 58855
rect 11307 58568 11349 58577
rect 11307 58528 11308 58568
rect 11348 58528 11349 58568
rect 11307 58519 11349 58528
rect 11308 57728 11348 58519
rect 11308 57679 11348 57688
rect 11307 56972 11349 56981
rect 11307 56932 11308 56972
rect 11348 56932 11349 56972
rect 11307 56923 11349 56932
rect 11308 56838 11348 56923
rect 11211 56804 11253 56813
rect 11211 56764 11212 56804
rect 11252 56764 11253 56804
rect 11211 56755 11253 56764
rect 11115 56636 11157 56645
rect 11115 56596 11116 56636
rect 11156 56596 11157 56636
rect 11115 56587 11157 56596
rect 11019 56300 11061 56309
rect 11019 56260 11020 56300
rect 11060 56260 11061 56300
rect 11019 56251 11061 56260
rect 11116 55628 11156 56587
rect 11307 55712 11349 55721
rect 11307 55672 11308 55712
rect 11348 55672 11349 55712
rect 11307 55663 11349 55672
rect 11212 55628 11252 55656
rect 11116 55588 11212 55628
rect 11019 55544 11061 55553
rect 11019 55504 11020 55544
rect 11060 55504 11061 55544
rect 11019 55495 11061 55504
rect 10484 52480 10580 52520
rect 10444 52471 10484 52480
rect 9964 51724 10100 51764
rect 10156 51976 10292 52016
rect 9867 51596 9909 51605
rect 9867 51556 9868 51596
rect 9908 51556 9909 51596
rect 9867 51547 9909 51556
rect 9964 50840 10004 51724
rect 10060 51596 10100 51605
rect 10060 51017 10100 51556
rect 10059 51008 10101 51017
rect 10059 50968 10060 51008
rect 10100 50968 10101 51008
rect 10059 50959 10101 50968
rect 9964 50800 10100 50840
rect 9867 49496 9909 49505
rect 9867 49456 9868 49496
rect 9908 49456 9909 49496
rect 9867 49447 9909 49456
rect 9868 49362 9908 49447
rect 9868 48824 9908 48833
rect 9868 48077 9908 48784
rect 9867 48068 9909 48077
rect 9867 48028 9868 48068
rect 9908 48028 9909 48068
rect 9867 48019 9909 48028
rect 9964 46481 10004 46566
rect 9868 46472 9908 46481
rect 9868 46313 9908 46432
rect 9963 46472 10005 46481
rect 9963 46432 9964 46472
rect 10004 46432 10005 46472
rect 9963 46423 10005 46432
rect 10060 46313 10100 50800
rect 10156 46640 10196 51976
rect 10252 51848 10292 51857
rect 10252 51689 10292 51808
rect 10251 51680 10293 51689
rect 10251 51640 10252 51680
rect 10292 51640 10293 51680
rect 10251 51631 10293 51640
rect 10443 51008 10485 51017
rect 10443 50968 10444 51008
rect 10484 50968 10485 51008
rect 10443 50959 10485 50968
rect 10540 51008 10580 52480
rect 10444 50874 10484 50959
rect 10540 50597 10580 50968
rect 10636 55336 10964 55376
rect 10539 50588 10581 50597
rect 10539 50548 10540 50588
rect 10580 50548 10581 50588
rect 10539 50539 10581 50548
rect 10251 50336 10293 50345
rect 10251 50296 10252 50336
rect 10292 50296 10293 50336
rect 10251 50287 10293 50296
rect 10444 50336 10484 50347
rect 10252 47984 10292 50287
rect 10444 50261 10484 50296
rect 10636 50261 10676 55336
rect 11020 55040 11060 55495
rect 11020 54991 11060 55000
rect 10827 54956 10869 54965
rect 10827 54916 10828 54956
rect 10868 54916 10869 54956
rect 10827 54907 10869 54916
rect 10828 54872 10868 54907
rect 10828 54545 10868 54832
rect 10827 54536 10869 54545
rect 10827 54496 10828 54536
rect 10868 54496 10869 54536
rect 10827 54487 10869 54496
rect 11116 53528 11156 55588
rect 11212 55579 11252 55588
rect 11308 55628 11348 55663
rect 11308 55577 11348 55588
rect 11307 54872 11349 54881
rect 11307 54832 11308 54872
rect 11348 54832 11349 54872
rect 11307 54823 11349 54832
rect 11308 54461 11348 54823
rect 11404 54713 11444 62560
rect 11500 62432 11540 62441
rect 11500 61601 11540 62392
rect 11499 61592 11541 61601
rect 11499 61552 11500 61592
rect 11540 61552 11541 61592
rect 11499 61543 11541 61552
rect 11596 60845 11636 62644
rect 11691 62264 11733 62273
rect 11691 62224 11692 62264
rect 11732 62224 11733 62264
rect 11691 62215 11733 62224
rect 11692 62130 11732 62215
rect 11595 60836 11637 60845
rect 11595 60796 11596 60836
rect 11636 60796 11637 60836
rect 11595 60787 11637 60796
rect 11691 60416 11733 60425
rect 11691 60376 11692 60416
rect 11732 60376 11733 60416
rect 11691 60367 11733 60376
rect 11692 59921 11732 60367
rect 11691 59912 11733 59921
rect 11691 59872 11692 59912
rect 11732 59872 11733 59912
rect 11691 59863 11733 59872
rect 11595 59072 11637 59081
rect 11595 59032 11596 59072
rect 11636 59032 11637 59072
rect 11595 59023 11637 59032
rect 11500 57812 11540 57821
rect 11500 57485 11540 57772
rect 11499 57476 11541 57485
rect 11499 57436 11500 57476
rect 11540 57436 11541 57476
rect 11499 57427 11541 57436
rect 11596 57308 11636 59023
rect 11692 57905 11732 59863
rect 11788 59408 11828 62803
rect 11884 61004 11924 64240
rect 12075 63944 12117 63953
rect 12075 63904 12076 63944
rect 12116 63904 12117 63944
rect 12075 63895 12117 63904
rect 12076 63810 12116 63895
rect 12075 63272 12117 63281
rect 12075 63232 12076 63272
rect 12116 63232 12117 63272
rect 12075 63223 12117 63232
rect 11980 62432 12020 62441
rect 11980 62273 12020 62392
rect 12076 62432 12116 63223
rect 11979 62264 12021 62273
rect 11979 62224 11980 62264
rect 12020 62224 12021 62264
rect 11979 62215 12021 62224
rect 12076 61013 12116 62392
rect 12172 61592 12212 66499
rect 12268 64448 12308 72304
rect 12364 72176 12404 72185
rect 12364 71849 12404 72136
rect 12459 72176 12501 72185
rect 12459 72136 12460 72176
rect 12500 72136 12501 72176
rect 12459 72127 12501 72136
rect 12460 72042 12500 72127
rect 12363 71840 12405 71849
rect 12363 71800 12364 71840
rect 12404 71800 12405 71840
rect 12363 71791 12405 71800
rect 12459 71672 12501 71681
rect 12459 71632 12460 71672
rect 12500 71632 12501 71672
rect 12459 71623 12501 71632
rect 12363 66716 12405 66725
rect 12363 66676 12364 66716
rect 12404 66676 12405 66716
rect 12363 66667 12405 66676
rect 12364 66380 12404 66667
rect 12364 66331 12404 66340
rect 12364 66128 12404 66137
rect 12364 65633 12404 66088
rect 12460 66053 12500 71623
rect 12556 71513 12596 73984
rect 12555 71504 12597 71513
rect 12555 71464 12556 71504
rect 12596 71464 12597 71504
rect 12555 71455 12597 71464
rect 12652 71093 12692 74992
rect 12748 74696 12788 75160
rect 12748 74647 12788 74656
rect 12651 71084 12693 71093
rect 12651 71044 12652 71084
rect 12692 71044 12693 71084
rect 12651 71035 12693 71044
rect 12652 69992 12692 70001
rect 12844 69992 12884 76831
rect 12939 76796 12981 76805
rect 12939 76756 12940 76796
rect 12980 76756 12981 76796
rect 12939 76747 12981 76756
rect 12940 72176 12980 76747
rect 13036 73100 13076 77512
rect 13996 73100 14036 83551
rect 14092 83516 14132 84727
rect 14284 83525 14324 85936
rect 14476 84785 14516 85936
rect 14475 84776 14517 84785
rect 14475 84736 14476 84776
rect 14516 84736 14517 84776
rect 14475 84727 14517 84736
rect 14379 84356 14421 84365
rect 14379 84316 14380 84356
rect 14420 84316 14421 84356
rect 14379 84307 14421 84316
rect 14092 83467 14132 83476
rect 14283 83516 14325 83525
rect 14283 83476 14284 83516
rect 14324 83476 14325 83516
rect 14283 83467 14325 83476
rect 14283 83348 14325 83357
rect 14283 83308 14284 83348
rect 14324 83308 14325 83348
rect 14283 83299 14325 83308
rect 14284 83214 14324 83299
rect 14380 82844 14420 84307
rect 14476 83516 14516 83525
rect 14668 83516 14708 85936
rect 14763 84440 14805 84449
rect 14763 84400 14764 84440
rect 14804 84400 14805 84440
rect 14763 84391 14805 84400
rect 14516 83476 14708 83516
rect 14476 83467 14516 83476
rect 14667 83348 14709 83357
rect 14667 83308 14668 83348
rect 14708 83308 14709 83348
rect 14667 83299 14709 83308
rect 14571 83264 14613 83273
rect 14571 83224 14572 83264
rect 14612 83224 14613 83264
rect 14571 83215 14613 83224
rect 14380 82795 14420 82804
rect 14572 82760 14612 83215
rect 14668 83214 14708 83299
rect 14764 82844 14804 84391
rect 14860 83516 14900 85936
rect 15052 84365 15092 85936
rect 15051 84356 15093 84365
rect 15051 84316 15052 84356
rect 15092 84316 15093 84356
rect 15051 84307 15093 84316
rect 14860 83467 14900 83476
rect 15244 83516 15284 85936
rect 15436 84449 15476 85936
rect 15435 84440 15477 84449
rect 15435 84400 15436 84440
rect 15476 84400 15477 84440
rect 15435 84391 15477 84400
rect 15628 83768 15668 85936
rect 15724 83768 15764 83777
rect 15628 83728 15724 83768
rect 15724 83719 15764 83728
rect 15244 83467 15284 83476
rect 15051 83348 15093 83357
rect 15051 83308 15052 83348
rect 15092 83308 15093 83348
rect 15051 83299 15093 83308
rect 15052 83214 15092 83299
rect 14764 82795 14804 82804
rect 14572 82720 14708 82760
rect 14187 82592 14229 82601
rect 14187 82552 14188 82592
rect 14228 82552 14229 82592
rect 14187 82543 14229 82552
rect 14572 82592 14612 82601
rect 14188 82458 14228 82543
rect 14572 81929 14612 82552
rect 14571 81920 14613 81929
rect 14571 81880 14572 81920
rect 14612 81880 14613 81920
rect 14571 81871 14613 81880
rect 13036 73060 13748 73100
rect 13468 72185 13508 72194
rect 13508 72145 13556 72176
rect 13468 72136 13556 72145
rect 12940 72127 12980 72136
rect 13131 72008 13173 72017
rect 13131 71968 13132 72008
rect 13172 71968 13173 72008
rect 13131 71959 13173 71968
rect 13035 70664 13077 70673
rect 13035 70624 13036 70664
rect 13076 70624 13077 70664
rect 13035 70615 13077 70624
rect 13036 70530 13076 70615
rect 13132 70076 13172 71959
rect 13516 71672 13556 72136
rect 13611 72008 13653 72017
rect 13611 71968 13612 72008
rect 13652 71968 13653 72008
rect 13611 71959 13653 71968
rect 13612 71874 13652 71959
rect 13612 71672 13652 71681
rect 13516 71632 13612 71672
rect 13612 71623 13652 71632
rect 13420 71504 13460 71513
rect 13460 71464 13556 71504
rect 13420 71455 13460 71464
rect 12692 69952 12884 69992
rect 13036 70036 13172 70076
rect 13228 70204 13460 70244
rect 12652 69943 12692 69952
rect 13036 68993 13076 70036
rect 13228 69992 13268 70204
rect 13180 69982 13268 69992
rect 13220 69952 13268 69982
rect 13324 70076 13364 70085
rect 13180 69933 13220 69942
rect 13131 69740 13173 69749
rect 13131 69700 13132 69740
rect 13172 69700 13173 69740
rect 13131 69691 13173 69700
rect 13132 69152 13172 69691
rect 13228 69152 13268 69161
rect 13132 69112 13228 69152
rect 13035 68984 13077 68993
rect 13035 68944 13036 68984
rect 13076 68944 13077 68984
rect 13035 68935 13077 68944
rect 12843 68900 12885 68909
rect 12843 68860 12844 68900
rect 12884 68860 12885 68900
rect 12843 68851 12885 68860
rect 12748 68480 12788 68489
rect 12748 68069 12788 68440
rect 12747 68060 12789 68069
rect 12747 68020 12748 68060
rect 12788 68020 12789 68060
rect 12747 68011 12789 68020
rect 12747 67388 12789 67397
rect 12747 67348 12748 67388
rect 12788 67348 12789 67388
rect 12747 67339 12789 67348
rect 12555 66884 12597 66893
rect 12555 66844 12556 66884
rect 12596 66844 12597 66884
rect 12555 66835 12597 66844
rect 12652 66884 12692 66893
rect 12556 66750 12596 66835
rect 12556 66128 12596 66137
rect 12459 66044 12501 66053
rect 12459 66004 12460 66044
rect 12500 66004 12501 66044
rect 12459 65995 12501 66004
rect 12363 65624 12405 65633
rect 12363 65584 12364 65624
rect 12404 65584 12405 65624
rect 12363 65575 12405 65584
rect 12556 65549 12596 66088
rect 12555 65540 12597 65549
rect 12555 65500 12556 65540
rect 12596 65500 12597 65540
rect 12555 65491 12597 65500
rect 12364 65456 12404 65465
rect 12364 65381 12404 65416
rect 12363 65372 12405 65381
rect 12363 65332 12364 65372
rect 12404 65332 12405 65372
rect 12363 65323 12405 65332
rect 12555 65372 12597 65381
rect 12555 65332 12556 65372
rect 12596 65332 12597 65372
rect 12555 65323 12597 65332
rect 12364 65213 12404 65323
rect 12556 65288 12596 65323
rect 12556 65237 12596 65248
rect 12363 65204 12405 65213
rect 12363 65164 12364 65204
rect 12404 65164 12500 65204
rect 12363 65155 12405 65164
rect 12363 64868 12405 64877
rect 12363 64828 12364 64868
rect 12404 64828 12405 64868
rect 12363 64819 12405 64828
rect 12364 64616 12404 64819
rect 12364 64567 12404 64576
rect 12268 64408 12404 64448
rect 12267 64280 12309 64289
rect 12267 64240 12268 64280
rect 12308 64240 12309 64280
rect 12267 64231 12309 64240
rect 12268 64112 12308 64231
rect 12268 64063 12308 64072
rect 12267 63944 12309 63953
rect 12267 63904 12268 63944
rect 12308 63904 12309 63944
rect 12267 63895 12309 63904
rect 12075 61004 12117 61013
rect 11884 60964 12020 61004
rect 11883 60836 11925 60845
rect 11883 60796 11884 60836
rect 11924 60796 11925 60836
rect 11883 60787 11925 60796
rect 11884 60080 11924 60787
rect 11980 60761 12020 60964
rect 12075 60964 12076 61004
rect 12116 60964 12117 61004
rect 12075 60955 12117 60964
rect 11979 60752 12021 60761
rect 11979 60712 11980 60752
rect 12020 60712 12021 60752
rect 11979 60703 12021 60712
rect 11884 60031 11924 60040
rect 11980 59912 12020 59921
rect 11788 59368 11924 59408
rect 11787 59240 11829 59249
rect 11787 59200 11788 59240
rect 11828 59200 11829 59240
rect 11787 59191 11829 59200
rect 11691 57896 11733 57905
rect 11691 57856 11692 57896
rect 11732 57856 11733 57896
rect 11691 57847 11733 57856
rect 11692 57762 11732 57847
rect 11500 57268 11636 57308
rect 11403 54704 11445 54713
rect 11403 54664 11404 54704
rect 11444 54664 11445 54704
rect 11403 54655 11445 54664
rect 11307 54452 11349 54461
rect 11307 54412 11308 54452
rect 11348 54412 11349 54452
rect 11307 54403 11349 54412
rect 11500 54284 11540 57268
rect 11595 57056 11637 57065
rect 11595 57016 11596 57056
rect 11636 57016 11637 57056
rect 11595 57007 11637 57016
rect 11692 57056 11732 57065
rect 11596 56922 11636 57007
rect 11595 56804 11637 56813
rect 11595 56764 11596 56804
rect 11636 56764 11637 56804
rect 11595 56755 11637 56764
rect 11404 54244 11540 54284
rect 11211 54200 11253 54209
rect 11211 54160 11212 54200
rect 11252 54160 11253 54200
rect 11211 54151 11253 54160
rect 11020 53488 11156 53528
rect 10732 53360 10772 53371
rect 10732 53285 10772 53320
rect 10731 53276 10773 53285
rect 10731 53236 10732 53276
rect 10772 53236 10773 53276
rect 10731 53227 10773 53236
rect 10923 53108 10965 53117
rect 10923 53068 10924 53108
rect 10964 53068 10965 53108
rect 10923 53059 10965 53068
rect 10924 52974 10964 53059
rect 10924 52604 10964 52613
rect 11020 52604 11060 53488
rect 11115 53360 11157 53369
rect 11115 53320 11116 53360
rect 11156 53320 11157 53360
rect 11115 53311 11157 53320
rect 11116 53226 11156 53311
rect 10964 52564 11060 52604
rect 10924 52555 10964 52564
rect 10828 52520 10868 52529
rect 10828 51008 10868 52480
rect 11212 51689 11252 54151
rect 11404 54125 11444 54244
rect 11596 54200 11636 56755
rect 11692 55301 11732 57016
rect 11788 55544 11828 59191
rect 11884 58745 11924 59368
rect 11883 58736 11925 58745
rect 11883 58696 11884 58736
rect 11924 58696 11925 58736
rect 11883 58687 11925 58696
rect 11980 58577 12020 59872
rect 12076 59501 12116 60955
rect 12075 59492 12117 59501
rect 12075 59452 12076 59492
rect 12116 59452 12117 59492
rect 12075 59443 12117 59452
rect 11979 58568 12021 58577
rect 11979 58528 11980 58568
rect 12020 58528 12021 58568
rect 11979 58519 12021 58528
rect 11883 57896 11925 57905
rect 11883 57856 11884 57896
rect 11924 57856 11925 57896
rect 11883 57847 11925 57856
rect 11884 56057 11924 57847
rect 12172 57812 12212 61552
rect 12268 60910 12308 63895
rect 12364 61097 12404 64408
rect 12460 63953 12500 65164
rect 12555 64448 12597 64457
rect 12555 64408 12556 64448
rect 12596 64408 12597 64448
rect 12555 64399 12597 64408
rect 12459 63944 12501 63953
rect 12459 63904 12460 63944
rect 12500 63904 12501 63944
rect 12459 63895 12501 63904
rect 12556 63944 12596 64399
rect 12652 64280 12692 66844
rect 12748 66128 12788 67339
rect 12844 66473 12884 68851
rect 13036 68405 13076 68935
rect 13035 68396 13077 68405
rect 13035 68356 13036 68396
rect 13076 68356 13077 68396
rect 13035 68347 13077 68356
rect 12940 68228 12980 68237
rect 13132 68228 13172 69112
rect 13228 69103 13268 69112
rect 13324 69077 13364 70036
rect 13420 69404 13460 70204
rect 13516 69749 13556 71464
rect 13515 69740 13557 69749
rect 13515 69700 13516 69740
rect 13556 69700 13557 69740
rect 13515 69691 13557 69700
rect 13420 69355 13460 69364
rect 13708 69329 13748 73060
rect 13900 73060 14036 73100
rect 13803 71504 13845 71513
rect 13803 71464 13804 71504
rect 13844 71464 13845 71504
rect 13803 71455 13845 71464
rect 13804 71370 13844 71455
rect 13803 71084 13845 71093
rect 13803 71044 13804 71084
rect 13844 71044 13845 71084
rect 13803 71035 13845 71044
rect 13707 69320 13749 69329
rect 13707 69280 13708 69320
rect 13748 69280 13749 69320
rect 13707 69271 13749 69280
rect 13708 69152 13748 69161
rect 13323 69068 13365 69077
rect 13323 69028 13324 69068
rect 13364 69028 13365 69068
rect 13323 69019 13365 69028
rect 13324 68732 13364 69019
rect 13708 68825 13748 69112
rect 13707 68816 13749 68825
rect 13707 68776 13708 68816
rect 13748 68776 13749 68816
rect 13707 68767 13749 68776
rect 12940 66977 12980 68188
rect 13036 68188 13172 68228
rect 13228 68692 13364 68732
rect 12939 66968 12981 66977
rect 12939 66928 12940 66968
rect 12980 66928 12981 66968
rect 12939 66919 12981 66928
rect 12843 66464 12885 66473
rect 12843 66424 12844 66464
rect 12884 66424 12885 66464
rect 12843 66415 12885 66424
rect 12940 66380 12980 66919
rect 13036 66641 13076 68188
rect 13132 66968 13172 66977
rect 13035 66632 13077 66641
rect 13035 66592 13036 66632
rect 13076 66592 13077 66632
rect 13035 66583 13077 66592
rect 13132 66557 13172 66928
rect 13131 66548 13173 66557
rect 13131 66508 13132 66548
rect 13172 66508 13173 66548
rect 13131 66499 13173 66508
rect 13228 66473 13268 68692
rect 13708 68480 13748 68489
rect 13708 68237 13748 68440
rect 13707 68228 13749 68237
rect 13707 68188 13708 68228
rect 13748 68188 13749 68228
rect 13707 68179 13749 68188
rect 13804 68069 13844 71035
rect 13323 68060 13365 68069
rect 13323 68020 13324 68060
rect 13364 68020 13365 68060
rect 13323 68011 13365 68020
rect 13803 68060 13845 68069
rect 13803 68020 13804 68060
rect 13844 68020 13845 68060
rect 13803 68011 13845 68020
rect 13324 67640 13364 68011
rect 13324 66977 13364 67600
rect 13516 67472 13556 67481
rect 13556 67432 13652 67472
rect 13516 67423 13556 67432
rect 13323 66968 13365 66977
rect 13323 66928 13324 66968
rect 13364 66928 13365 66968
rect 13323 66919 13365 66928
rect 13612 66963 13652 67432
rect 13803 67388 13845 67397
rect 13803 67348 13804 67388
rect 13844 67348 13845 67388
rect 13803 67339 13845 67348
rect 13804 67136 13844 67339
rect 13900 67229 13940 73060
rect 14283 72344 14325 72353
rect 14283 72304 14284 72344
rect 14324 72304 14325 72344
rect 14283 72295 14325 72304
rect 13996 72176 14036 72185
rect 13996 71429 14036 72136
rect 13995 71420 14037 71429
rect 13995 71380 13996 71420
rect 14036 71380 14037 71420
rect 13995 71371 14037 71380
rect 14284 70664 14324 72295
rect 14284 69161 14324 70624
rect 14475 70664 14517 70673
rect 14475 70624 14476 70664
rect 14516 70624 14517 70664
rect 14475 70615 14517 70624
rect 14476 70496 14516 70615
rect 14379 70244 14421 70253
rect 14379 70204 14380 70244
rect 14420 70204 14421 70244
rect 14379 70195 14421 70204
rect 14380 69572 14420 70195
rect 14476 69992 14516 70456
rect 14476 69943 14516 69952
rect 14572 69992 14612 70001
rect 14572 69749 14612 69952
rect 14571 69740 14613 69749
rect 14571 69700 14572 69740
rect 14612 69700 14613 69740
rect 14571 69691 14613 69700
rect 14380 69532 14612 69572
rect 14283 69152 14325 69161
rect 14283 69112 14284 69152
rect 14324 69112 14325 69152
rect 14283 69103 14325 69112
rect 14188 67768 14516 67808
rect 14188 67724 14228 67768
rect 14188 67675 14228 67684
rect 14092 67640 14132 67649
rect 14092 67397 14132 67600
rect 14284 67640 14324 67649
rect 14091 67388 14133 67397
rect 14091 67348 14092 67388
rect 14132 67348 14133 67388
rect 14091 67339 14133 67348
rect 13899 67220 13941 67229
rect 13899 67180 13900 67220
rect 13940 67180 13941 67220
rect 13899 67171 13941 67180
rect 13804 67087 13844 67096
rect 14188 66977 14228 67062
rect 13612 66884 13652 66923
rect 14187 66968 14229 66977
rect 14187 66928 14188 66968
rect 14228 66928 14229 66968
rect 14187 66919 14229 66928
rect 13612 66844 13844 66884
rect 13227 66464 13269 66473
rect 13227 66424 13228 66464
rect 13268 66424 13269 66464
rect 13227 66415 13269 66424
rect 12940 66340 13172 66380
rect 13132 66296 13172 66340
rect 13132 66256 13556 66296
rect 12748 65801 12788 66088
rect 12843 66128 12885 66137
rect 12843 66088 12844 66128
rect 12884 66088 12885 66128
rect 12843 66079 12885 66088
rect 13036 66128 13076 66139
rect 12844 65994 12884 66079
rect 13036 66053 13076 66088
rect 13132 66128 13172 66256
rect 13516 66147 13556 66256
rect 13132 66079 13172 66088
rect 13228 66128 13268 66139
rect 13612 66137 13652 66222
rect 13516 66098 13556 66107
rect 13611 66128 13653 66137
rect 13228 66053 13268 66088
rect 13611 66088 13612 66128
rect 13652 66088 13653 66128
rect 13611 66079 13653 66088
rect 13708 66053 13748 66138
rect 13804 66128 13844 66844
rect 13996 66800 14036 66809
rect 14284 66800 14324 67600
rect 14036 66760 14324 66800
rect 13996 66751 14036 66760
rect 13804 66079 13844 66088
rect 14188 66128 14228 66137
rect 13035 66044 13077 66053
rect 13035 66004 13036 66044
rect 13076 66004 13077 66044
rect 13035 65995 13077 66004
rect 13227 66044 13269 66053
rect 13227 66004 13228 66044
rect 13268 66004 13269 66044
rect 13227 65995 13269 66004
rect 13707 66044 13749 66053
rect 13707 66004 13708 66044
rect 13748 66004 13749 66044
rect 13707 65995 13749 66004
rect 14188 65969 14228 66088
rect 14284 66128 14324 66760
rect 14284 66079 14324 66088
rect 14476 66128 14516 67768
rect 14476 66079 14516 66088
rect 13323 65960 13365 65969
rect 13323 65920 13324 65960
rect 13364 65920 13365 65960
rect 13323 65911 13365 65920
rect 14187 65960 14229 65969
rect 14187 65920 14188 65960
rect 14228 65920 14229 65960
rect 14187 65911 14229 65920
rect 14379 65960 14421 65969
rect 14379 65920 14380 65960
rect 14420 65920 14421 65960
rect 14379 65911 14421 65920
rect 13324 65826 13364 65911
rect 13611 65876 13653 65885
rect 13611 65836 13612 65876
rect 13652 65836 13653 65876
rect 13611 65827 13653 65836
rect 12747 65792 12789 65801
rect 12747 65752 12748 65792
rect 12788 65752 12789 65792
rect 12747 65743 12789 65752
rect 13036 65624 13076 65633
rect 13076 65584 13175 65624
rect 13036 65575 13076 65584
rect 12940 65477 12980 65486
rect 12748 65456 12788 65465
rect 12748 65297 12788 65416
rect 12844 65456 12884 65465
rect 13135 65465 13175 65584
rect 13228 65465 13268 65550
rect 13323 65540 13365 65549
rect 13323 65500 13324 65540
rect 13364 65500 13365 65540
rect 13323 65491 13365 65500
rect 13131 65456 13175 65465
rect 12980 65437 13075 65456
rect 12940 65416 13075 65437
rect 12747 65288 12789 65297
rect 12747 65248 12748 65288
rect 12788 65248 12789 65288
rect 12747 65239 12789 65248
rect 12747 64952 12789 64961
rect 12747 64912 12748 64952
rect 12788 64912 12789 64952
rect 12844 64952 12884 65416
rect 13035 65381 13075 65416
rect 13131 65416 13132 65456
rect 13172 65416 13175 65456
rect 13131 65411 13175 65416
rect 13227 65456 13269 65465
rect 13227 65416 13228 65456
rect 13268 65416 13269 65456
rect 13131 65407 13173 65411
rect 13227 65407 13269 65416
rect 13324 65406 13364 65491
rect 13420 65456 13460 65465
rect 13035 65372 13077 65381
rect 13035 65332 13036 65372
rect 13076 65332 13077 65372
rect 13035 65323 13077 65332
rect 13420 65297 13460 65416
rect 13516 65456 13556 65465
rect 13419 65288 13461 65297
rect 13419 65248 13420 65288
rect 13460 65248 13461 65288
rect 13419 65239 13461 65248
rect 13516 65045 13556 65416
rect 13035 65036 13077 65045
rect 13035 64996 13036 65036
rect 13076 64996 13077 65036
rect 13035 64987 13077 64996
rect 13515 65036 13557 65045
rect 13515 64996 13516 65036
rect 13556 64996 13557 65036
rect 13515 64987 13557 64996
rect 12844 64912 12980 64952
rect 12747 64903 12789 64912
rect 12748 64541 12788 64903
rect 12844 64621 12884 64630
rect 12940 64625 12980 64912
rect 13036 64868 13076 64987
rect 13036 64828 13172 64868
rect 12747 64532 12789 64541
rect 12747 64492 12748 64532
rect 12788 64492 12789 64532
rect 12747 64483 12789 64492
rect 12844 64457 12884 64581
rect 12939 64616 12981 64625
rect 12939 64576 12940 64616
rect 12980 64576 12981 64616
rect 12939 64567 12981 64576
rect 13035 64532 13077 64541
rect 13035 64492 13036 64532
rect 13076 64492 13077 64532
rect 13035 64483 13077 64492
rect 12843 64448 12885 64457
rect 12843 64408 12844 64448
rect 12884 64408 12885 64448
rect 12843 64399 12885 64408
rect 13036 64398 13076 64483
rect 12652 64240 12788 64280
rect 12748 63944 12788 64240
rect 12939 64028 12981 64037
rect 12939 63988 12940 64028
rect 12980 63988 12981 64028
rect 12939 63979 12981 63988
rect 12844 63944 12884 63953
rect 12596 63904 12692 63944
rect 12556 63895 12596 63904
rect 12555 63776 12597 63785
rect 12555 63736 12556 63776
rect 12596 63736 12597 63776
rect 12555 63727 12597 63736
rect 12556 63104 12596 63727
rect 12459 62768 12501 62777
rect 12459 62728 12460 62768
rect 12500 62728 12501 62768
rect 12459 62719 12501 62728
rect 12460 62441 12500 62719
rect 12459 62432 12501 62441
rect 12459 62392 12460 62432
rect 12500 62392 12501 62432
rect 12459 62383 12501 62392
rect 12460 62298 12500 62383
rect 12556 62348 12596 63064
rect 12652 63104 12692 63904
rect 12652 63055 12692 63064
rect 12748 63904 12844 63944
rect 12556 62273 12596 62308
rect 12555 62264 12597 62273
rect 12555 62224 12556 62264
rect 12596 62224 12597 62264
rect 12555 62215 12597 62224
rect 12748 61097 12788 63904
rect 12844 63895 12884 63904
rect 12940 63894 12980 63979
rect 13132 63776 13172 64828
rect 13228 64616 13268 64625
rect 13228 64289 13268 64576
rect 13324 64616 13364 64625
rect 13324 64457 13364 64576
rect 13420 64616 13460 64625
rect 13323 64448 13365 64457
rect 13323 64408 13324 64448
rect 13364 64408 13365 64448
rect 13323 64399 13365 64408
rect 13227 64280 13269 64289
rect 13227 64240 13228 64280
rect 13268 64240 13269 64280
rect 13227 64231 13269 64240
rect 13228 63776 13268 63785
rect 13132 63736 13228 63776
rect 13228 63727 13268 63736
rect 13420 63608 13460 64576
rect 13515 64616 13557 64625
rect 13515 64576 13516 64616
rect 13556 64576 13557 64616
rect 13515 64567 13557 64576
rect 13516 64482 13556 64567
rect 13515 64364 13557 64373
rect 13515 64324 13516 64364
rect 13556 64324 13557 64364
rect 13515 64315 13557 64324
rect 12844 63568 13460 63608
rect 12844 62936 12884 63568
rect 13131 63440 13173 63449
rect 13131 63400 13132 63440
rect 13172 63400 13173 63440
rect 13131 63391 13173 63400
rect 12844 62887 12884 62896
rect 13132 62516 13172 63391
rect 13227 63104 13269 63113
rect 13227 63064 13228 63104
rect 13268 63064 13269 63104
rect 13227 63055 13269 63064
rect 13228 62970 13268 63055
rect 13516 62516 13556 64315
rect 13132 62476 13268 62516
rect 13036 62432 13076 62441
rect 13076 62392 13172 62432
rect 13036 62383 13076 62392
rect 12363 61088 12405 61097
rect 12363 61048 12364 61088
rect 12404 61048 12405 61088
rect 12363 61039 12405 61048
rect 12747 61088 12789 61097
rect 12747 61048 12748 61088
rect 12788 61048 12789 61088
rect 12747 61039 12789 61048
rect 12364 60929 12404 60994
rect 13036 60929 13076 61014
rect 12363 60920 12405 60929
rect 12363 60910 12364 60920
rect 12268 60870 12364 60910
rect 12404 60871 12405 60920
rect 12651 60920 12693 60929
rect 12651 60880 12652 60920
rect 12692 60880 12693 60920
rect 12651 60871 12693 60880
rect 12748 60920 12788 60929
rect 12364 60850 12404 60859
rect 12556 60668 12596 60677
rect 12556 60500 12596 60628
rect 12268 60460 12596 60500
rect 12268 60080 12308 60460
rect 12555 60332 12597 60341
rect 12555 60292 12556 60332
rect 12596 60292 12597 60332
rect 12555 60283 12597 60292
rect 12459 60164 12501 60173
rect 12459 60124 12460 60164
rect 12500 60124 12501 60164
rect 12459 60115 12501 60124
rect 12268 60031 12308 60040
rect 12364 60080 12404 60089
rect 12364 59501 12404 60040
rect 12363 59492 12405 59501
rect 12363 59452 12364 59492
rect 12404 59452 12405 59492
rect 12363 59443 12405 59452
rect 12363 59072 12405 59081
rect 12363 59032 12364 59072
rect 12404 59032 12405 59072
rect 12363 59023 12405 59032
rect 12364 58568 12404 59023
rect 12364 58519 12404 58528
rect 12172 57772 12308 57812
rect 12171 57644 12213 57653
rect 12171 57604 12172 57644
rect 12212 57604 12213 57644
rect 12171 57595 12213 57604
rect 12172 57140 12212 57595
rect 12172 57091 12212 57100
rect 12076 57056 12116 57065
rect 12076 56645 12116 57016
rect 12268 56729 12308 57772
rect 12363 57224 12405 57233
rect 12363 57184 12364 57224
rect 12404 57184 12405 57224
rect 12363 57175 12405 57184
rect 12267 56720 12309 56729
rect 12267 56680 12268 56720
rect 12308 56680 12309 56720
rect 12267 56671 12309 56680
rect 12075 56636 12117 56645
rect 12075 56596 12076 56636
rect 12116 56596 12117 56636
rect 12075 56587 12117 56596
rect 12364 56552 12404 57175
rect 12460 57149 12500 60115
rect 12556 59408 12596 60283
rect 12652 59576 12692 60871
rect 12748 60248 12788 60880
rect 12843 60920 12885 60929
rect 12843 60880 12844 60920
rect 12884 60880 12885 60920
rect 12843 60871 12885 60880
rect 13035 60920 13077 60929
rect 13035 60880 13036 60920
rect 13076 60880 13077 60920
rect 13035 60871 13077 60880
rect 12844 60786 12884 60871
rect 12940 60752 12980 60761
rect 12980 60712 13076 60752
rect 12940 60703 12980 60712
rect 12748 60208 12980 60248
rect 12747 60080 12789 60089
rect 12747 60040 12748 60080
rect 12788 60040 12789 60080
rect 12747 60031 12789 60040
rect 12844 60080 12884 60091
rect 12748 59946 12788 60031
rect 12844 60005 12884 60040
rect 12843 59996 12885 60005
rect 12843 59956 12844 59996
rect 12884 59956 12885 59996
rect 12843 59947 12885 59956
rect 12748 59576 12788 59585
rect 12940 59576 12980 60208
rect 12652 59536 12748 59576
rect 12748 59527 12788 59536
rect 12844 59536 12980 59576
rect 12556 59081 12596 59368
rect 12844 59324 12884 59536
rect 13036 59501 13076 60712
rect 13132 60080 13172 62392
rect 13228 60425 13268 62476
rect 13324 62476 13556 62516
rect 13227 60416 13269 60425
rect 13227 60376 13228 60416
rect 13268 60376 13269 60416
rect 13227 60367 13269 60376
rect 13324 60248 13364 62476
rect 13516 62418 13556 62427
rect 13612 62418 13652 65827
rect 14380 65826 14420 65911
rect 13707 65624 13749 65633
rect 13707 65584 13708 65624
rect 13748 65584 13749 65624
rect 13707 65575 13749 65584
rect 13708 64868 13748 65575
rect 14476 65456 14516 65465
rect 13899 65372 13941 65381
rect 13899 65332 13900 65372
rect 13940 65332 13941 65372
rect 13899 65323 13941 65332
rect 13803 64952 13845 64961
rect 13803 64912 13804 64952
rect 13844 64912 13845 64952
rect 13803 64903 13845 64912
rect 13708 64819 13748 64828
rect 13708 64616 13748 64627
rect 13708 64541 13748 64576
rect 13707 64532 13749 64541
rect 13707 64492 13708 64532
rect 13748 64492 13749 64532
rect 13707 64483 13749 64492
rect 13804 64373 13844 64903
rect 13900 64616 13940 65323
rect 14476 65129 14516 65416
rect 14475 65120 14517 65129
rect 14475 65080 14476 65120
rect 14516 65080 14517 65120
rect 14475 65071 14517 65080
rect 14283 64868 14325 64877
rect 14283 64828 14284 64868
rect 14324 64828 14325 64868
rect 14283 64819 14325 64828
rect 14475 64868 14517 64877
rect 14475 64828 14476 64868
rect 14516 64828 14517 64868
rect 14475 64819 14517 64828
rect 14091 64784 14133 64793
rect 14091 64744 14092 64784
rect 14132 64744 14133 64784
rect 14091 64735 14133 64744
rect 13900 64567 13940 64576
rect 14092 64616 14132 64735
rect 14187 64700 14229 64709
rect 14187 64660 14188 64700
rect 14228 64660 14229 64700
rect 14187 64651 14229 64660
rect 14092 64567 14132 64576
rect 13803 64364 13845 64373
rect 14188 64364 14228 64651
rect 13803 64324 13804 64364
rect 13844 64324 13845 64364
rect 13803 64315 13845 64324
rect 14092 64324 14228 64364
rect 13803 63944 13845 63953
rect 13803 63904 13804 63944
rect 13844 63904 13845 63944
rect 13803 63895 13845 63904
rect 13900 63944 13940 63953
rect 13804 63810 13844 63895
rect 13900 63272 13940 63904
rect 13900 63232 14036 63272
rect 13707 62600 13749 62609
rect 13707 62560 13708 62600
rect 13748 62560 13749 62600
rect 13707 62551 13749 62560
rect 13708 62466 13748 62551
rect 13612 62378 13748 62418
rect 13516 61844 13556 62378
rect 13612 61844 13652 61853
rect 13516 61804 13612 61844
rect 13612 61795 13652 61804
rect 13419 61592 13461 61601
rect 13419 61552 13420 61592
rect 13460 61552 13652 61592
rect 13419 61543 13461 61552
rect 13420 61458 13460 61543
rect 13515 60920 13557 60929
rect 13515 60880 13516 60920
rect 13556 60880 13557 60920
rect 13515 60871 13557 60880
rect 13324 60208 13460 60248
rect 13324 60080 13364 60089
rect 13132 60040 13324 60080
rect 13035 59492 13077 59501
rect 13035 59452 13036 59492
rect 13076 59452 13077 59492
rect 13035 59443 13077 59452
rect 12939 59408 12981 59417
rect 12939 59368 12940 59408
rect 12980 59368 12981 59408
rect 12939 59359 12981 59368
rect 12652 59284 12884 59324
rect 12555 59072 12597 59081
rect 12555 59032 12556 59072
rect 12596 59032 12597 59072
rect 12555 59023 12597 59032
rect 12556 58736 12596 58747
rect 12556 58661 12596 58696
rect 12555 58652 12597 58661
rect 12555 58612 12556 58652
rect 12596 58612 12597 58652
rect 12555 58603 12597 58612
rect 12555 58148 12597 58157
rect 12555 58108 12556 58148
rect 12596 58108 12597 58148
rect 12652 58148 12692 59284
rect 12940 59274 12980 59359
rect 12748 59156 12788 59165
rect 12788 59116 13076 59156
rect 12748 59107 12788 59116
rect 12838 58652 12880 58661
rect 12838 58612 12839 58652
rect 12879 58612 12880 58652
rect 12838 58603 12880 58612
rect 12839 58568 12879 58603
rect 12839 58517 12879 58528
rect 12939 58568 12981 58577
rect 12939 58528 12940 58568
rect 12980 58528 12981 58568
rect 12939 58519 12981 58528
rect 13036 58568 13076 59116
rect 13036 58519 13076 58528
rect 12940 58434 12980 58519
rect 13035 58400 13077 58409
rect 13035 58360 13036 58400
rect 13076 58360 13077 58400
rect 13035 58351 13077 58360
rect 13132 58400 13172 60040
rect 13324 60031 13364 60040
rect 13323 59492 13365 59501
rect 13323 59452 13324 59492
rect 13364 59452 13365 59492
rect 13323 59443 13365 59452
rect 13228 58568 13268 58577
rect 13228 58409 13268 58528
rect 13324 58568 13364 59443
rect 13324 58519 13364 58528
rect 13132 58351 13172 58360
rect 13227 58400 13269 58409
rect 13227 58360 13228 58400
rect 13268 58360 13269 58400
rect 13227 58351 13269 58360
rect 13036 58232 13076 58351
rect 13036 58192 13268 58232
rect 12652 58108 13076 58148
rect 12555 58099 12597 58108
rect 12556 57980 12596 58099
rect 12939 57980 12981 57989
rect 12556 57940 12692 57980
rect 12459 57140 12501 57149
rect 12459 57100 12460 57140
rect 12500 57100 12501 57140
rect 12459 57091 12501 57100
rect 12364 56503 12404 56512
rect 12652 57056 12692 57940
rect 12939 57940 12940 57980
rect 12980 57940 12981 57980
rect 12939 57931 12981 57940
rect 12940 57896 12980 57931
rect 12940 57845 12980 57856
rect 11980 56342 12020 56351
rect 11979 56302 11980 56309
rect 12020 56302 12021 56309
rect 11979 56300 12021 56302
rect 11979 56260 11980 56300
rect 12020 56260 12021 56300
rect 11979 56251 12021 56260
rect 12556 56300 12596 56309
rect 11980 56207 12020 56251
rect 12172 56132 12212 56141
rect 12212 56092 12308 56132
rect 12172 56083 12212 56092
rect 11883 56048 11925 56057
rect 11883 56008 11884 56048
rect 11924 56008 11925 56048
rect 11883 55999 11925 56008
rect 12268 55558 12308 56092
rect 12268 55509 12308 55518
rect 11691 55292 11733 55301
rect 11691 55252 11692 55292
rect 11732 55252 11733 55292
rect 11691 55243 11733 55252
rect 11788 54377 11828 55504
rect 12460 55460 12500 55469
rect 12556 55460 12596 56260
rect 12500 55420 12596 55460
rect 12460 55411 12500 55420
rect 12363 55292 12405 55301
rect 12363 55252 12364 55292
rect 12404 55252 12405 55292
rect 12363 55243 12405 55252
rect 12075 54704 12117 54713
rect 12075 54664 12076 54704
rect 12116 54664 12117 54704
rect 12075 54655 12117 54664
rect 11787 54368 11829 54377
rect 11787 54328 11788 54368
rect 11828 54328 11829 54368
rect 11787 54319 11829 54328
rect 12076 54200 12116 54655
rect 12267 54368 12309 54377
rect 12267 54328 12268 54368
rect 12308 54328 12309 54368
rect 12267 54319 12309 54328
rect 11500 54160 11636 54200
rect 11980 54160 12116 54200
rect 11403 54116 11445 54125
rect 11403 54076 11404 54116
rect 11444 54076 11445 54116
rect 11403 54067 11445 54076
rect 11403 52604 11445 52613
rect 11403 52564 11404 52604
rect 11444 52564 11445 52604
rect 11403 52555 11445 52564
rect 11404 52520 11444 52555
rect 11404 52469 11444 52480
rect 11500 52016 11540 54160
rect 11980 54041 12020 54160
rect 12172 54116 12212 54125
rect 12076 54076 12172 54116
rect 11596 54032 11636 54041
rect 11596 53285 11636 53992
rect 11979 54032 12021 54041
rect 11979 53992 11980 54032
rect 12020 53992 12021 54032
rect 11979 53983 12021 53992
rect 11788 53864 11828 53873
rect 11980 53864 12020 53873
rect 11828 53824 11924 53864
rect 11788 53815 11828 53824
rect 11787 53696 11829 53705
rect 11787 53656 11788 53696
rect 11828 53656 11829 53696
rect 11787 53647 11829 53656
rect 11595 53276 11637 53285
rect 11595 53236 11596 53276
rect 11636 53236 11637 53276
rect 11595 53227 11637 53236
rect 11500 51976 11636 52016
rect 11500 51848 11540 51857
rect 11500 51689 11540 51808
rect 11211 51680 11253 51689
rect 11211 51640 11212 51680
rect 11252 51640 11253 51680
rect 11211 51631 11253 51640
rect 11499 51680 11541 51689
rect 11499 51640 11500 51680
rect 11540 51640 11541 51680
rect 11499 51631 11541 51640
rect 10924 51008 10964 51017
rect 10732 50968 10924 51008
rect 10443 50252 10485 50261
rect 10348 50212 10444 50252
rect 10484 50212 10485 50252
rect 10348 49589 10388 50212
rect 10443 50203 10485 50212
rect 10635 50252 10677 50261
rect 10635 50212 10636 50252
rect 10676 50212 10677 50252
rect 10635 50203 10677 50212
rect 10636 50084 10676 50093
rect 10444 50044 10636 50084
rect 10347 49580 10389 49589
rect 10347 49540 10348 49580
rect 10388 49540 10389 49580
rect 10347 49531 10389 49540
rect 10444 48824 10484 50044
rect 10636 50035 10676 50044
rect 10396 48814 10484 48824
rect 10436 48784 10484 48814
rect 10540 48908 10580 48917
rect 10396 48765 10436 48774
rect 10252 47935 10292 47944
rect 10540 46640 10580 48868
rect 10635 47732 10677 47741
rect 10635 47692 10636 47732
rect 10676 47692 10677 47732
rect 10635 47683 10677 47692
rect 10636 47480 10676 47683
rect 10636 47431 10676 47440
rect 10156 46600 10292 46640
rect 10540 46600 10676 46640
rect 9867 46304 9909 46313
rect 9867 46264 9868 46304
rect 9908 46264 9909 46304
rect 9867 46255 9909 46264
rect 10059 46304 10101 46313
rect 10059 46264 10060 46304
rect 10100 46264 10101 46304
rect 10059 46255 10101 46264
rect 10059 46136 10101 46145
rect 10059 46096 10060 46136
rect 10100 46096 10101 46136
rect 10059 46087 10101 46096
rect 10060 45800 10100 46087
rect 10060 45751 10100 45760
rect 9963 45716 10005 45725
rect 9963 45676 9964 45716
rect 10004 45676 10005 45716
rect 9963 45667 10005 45676
rect 9964 45582 10004 45667
rect 10059 44288 10101 44297
rect 10059 44248 10060 44288
rect 10100 44248 10101 44288
rect 10059 44239 10101 44248
rect 9867 44204 9909 44213
rect 9867 44164 9868 44204
rect 9908 44164 9909 44204
rect 9867 44155 9909 44164
rect 9868 44070 9908 44155
rect 10060 44154 10100 44239
rect 9867 43952 9909 43961
rect 9867 43912 9868 43952
rect 9908 43912 9909 43952
rect 9867 43903 9909 43912
rect 9771 43868 9813 43877
rect 9771 43828 9772 43868
rect 9812 43828 9813 43868
rect 9771 43819 9813 43828
rect 9196 43744 9716 43784
rect 9387 43532 9429 43541
rect 9387 43492 9388 43532
rect 9428 43492 9429 43532
rect 9387 43483 9429 43492
rect 9388 42776 9428 43483
rect 9532 43457 9572 43466
rect 9572 43417 9620 43448
rect 9532 43408 9620 43417
rect 9580 42944 9620 43408
rect 9676 43364 9716 43744
rect 9868 43448 9908 43903
rect 9964 43448 10004 43457
rect 9676 43315 9716 43324
rect 9772 43408 9964 43448
rect 9580 42895 9620 42904
rect 9428 42736 9620 42776
rect 9388 42727 9428 42736
rect 9195 42440 9237 42449
rect 9195 42400 9196 42440
rect 9236 42400 9237 42440
rect 9195 42391 9237 42400
rect 8812 41609 8852 41896
rect 8908 41980 9140 42020
rect 8811 41600 8853 41609
rect 8811 41560 8812 41600
rect 8852 41560 8853 41600
rect 8811 41551 8853 41560
rect 8908 41432 8948 41980
rect 9196 41936 9236 42391
rect 9004 41777 9044 41862
rect 9003 41768 9045 41777
rect 9003 41728 9004 41768
rect 9044 41728 9045 41768
rect 9003 41719 9045 41728
rect 9003 41600 9045 41609
rect 9003 41560 9004 41600
rect 9044 41560 9045 41600
rect 9003 41551 9045 41560
rect 8812 41392 8948 41432
rect 8331 38996 8373 39005
rect 8331 38956 8332 38996
rect 8372 38956 8373 38996
rect 8331 38947 8373 38956
rect 8620 38912 8660 38921
rect 8332 38828 8372 38837
rect 8620 38828 8660 38872
rect 8715 38912 8757 38921
rect 8715 38872 8716 38912
rect 8756 38872 8757 38912
rect 8715 38863 8757 38872
rect 8372 38788 8660 38828
rect 8332 38779 8372 38788
rect 8523 38240 8565 38249
rect 8523 38200 8524 38240
rect 8564 38200 8565 38240
rect 8523 38191 8565 38200
rect 8620 38240 8660 38249
rect 8716 38240 8756 38863
rect 8812 38585 8852 41392
rect 8908 41264 8948 41273
rect 9004 41264 9044 41551
rect 9099 41348 9141 41357
rect 9099 41308 9100 41348
rect 9140 41308 9141 41348
rect 9099 41299 9141 41308
rect 8948 41224 9044 41264
rect 8908 40433 8948 41224
rect 9100 41214 9140 41299
rect 9003 40760 9045 40769
rect 9003 40720 9004 40760
rect 9044 40720 9045 40760
rect 9003 40711 9045 40720
rect 9004 40517 9044 40711
rect 9003 40508 9045 40517
rect 9003 40468 9004 40508
rect 9044 40468 9045 40508
rect 9003 40459 9045 40468
rect 8907 40424 8949 40433
rect 8907 40384 8908 40424
rect 8948 40384 8949 40424
rect 8907 40375 8949 40384
rect 9004 40424 9044 40459
rect 9004 40373 9044 40384
rect 8907 39752 8949 39761
rect 8907 39712 8908 39752
rect 8948 39712 8949 39752
rect 8907 39703 8949 39712
rect 8908 39618 8948 39703
rect 9100 39500 9140 39509
rect 9100 39089 9140 39460
rect 9196 39332 9236 41896
rect 9387 41768 9429 41777
rect 9387 41728 9388 41768
rect 9428 41728 9429 41768
rect 9387 41719 9429 41728
rect 9291 41600 9333 41609
rect 9291 41560 9292 41600
rect 9332 41560 9333 41600
rect 9291 41551 9333 41560
rect 9292 41432 9332 41551
rect 9292 41383 9332 41392
rect 9388 40424 9428 41719
rect 9483 41600 9525 41609
rect 9483 41560 9484 41600
rect 9524 41560 9525 41600
rect 9483 41551 9525 41560
rect 9388 40375 9428 40384
rect 9484 40424 9524 41551
rect 9388 39920 9428 39929
rect 9484 39920 9524 40384
rect 9428 39880 9524 39920
rect 9388 39871 9428 39880
rect 9580 39836 9620 42736
rect 9772 40181 9812 43408
rect 9964 43399 10004 43408
rect 10252 42692 10292 46600
rect 10348 46565 10388 46596
rect 10347 46556 10389 46565
rect 10347 46516 10348 46556
rect 10388 46516 10389 46556
rect 10347 46507 10389 46516
rect 10348 46472 10388 46507
rect 10348 45725 10388 46432
rect 10444 46472 10484 46481
rect 10444 46145 10484 46432
rect 10539 46472 10581 46481
rect 10539 46432 10540 46472
rect 10580 46432 10581 46472
rect 10539 46423 10581 46432
rect 10443 46136 10485 46145
rect 10443 46096 10444 46136
rect 10484 46096 10485 46136
rect 10443 46087 10485 46096
rect 10540 45800 10580 46423
rect 10540 45751 10580 45760
rect 10347 45716 10389 45725
rect 10347 45676 10348 45716
rect 10388 45676 10389 45716
rect 10347 45667 10389 45676
rect 10636 44213 10676 46600
rect 10732 46565 10772 50968
rect 10924 50959 10964 50968
rect 11020 51008 11060 51017
rect 11020 50849 11060 50968
rect 11019 50840 11061 50849
rect 11019 50800 11020 50840
rect 11060 50800 11061 50840
rect 11019 50791 11061 50800
rect 11115 49496 11157 49505
rect 11115 49456 11116 49496
rect 11156 49456 11157 49496
rect 11115 49447 11157 49456
rect 11116 49362 11156 49447
rect 11116 47312 11156 47321
rect 10828 47228 10868 47237
rect 10828 46640 10868 47188
rect 11116 46817 11156 47272
rect 11115 46808 11157 46817
rect 11115 46768 11116 46808
rect 11156 46768 11157 46808
rect 11115 46759 11157 46768
rect 11212 46640 11252 51631
rect 11499 51008 11541 51017
rect 11499 50968 11500 51008
rect 11540 50968 11541 51008
rect 11499 50959 11541 50968
rect 11500 50874 11540 50959
rect 11596 50345 11636 51976
rect 11788 51680 11828 53647
rect 11884 52534 11924 53824
rect 11980 53201 12020 53824
rect 11979 53192 12021 53201
rect 11979 53152 11980 53192
rect 12020 53152 12021 53192
rect 11979 53143 12021 53152
rect 11979 52940 12021 52949
rect 11979 52900 11980 52940
rect 12020 52900 12021 52940
rect 11979 52891 12021 52900
rect 11884 52485 11924 52494
rect 11884 51848 11924 51857
rect 11980 51848 12020 52891
rect 12076 52436 12116 54076
rect 12172 54067 12212 54076
rect 12171 53528 12213 53537
rect 12171 53488 12172 53528
rect 12212 53488 12213 53528
rect 12171 53479 12213 53488
rect 12076 52387 12116 52396
rect 11924 51808 12020 51848
rect 11884 51799 11924 51808
rect 11788 51640 12116 51680
rect 11692 51596 11732 51605
rect 11732 51556 12020 51596
rect 11692 51547 11732 51556
rect 11691 51092 11733 51101
rect 11691 51052 11692 51092
rect 11732 51052 11733 51092
rect 11691 51043 11733 51052
rect 11595 50336 11637 50345
rect 11595 50296 11596 50336
rect 11636 50296 11637 50336
rect 11595 50287 11637 50296
rect 11403 50252 11445 50261
rect 11403 50212 11404 50252
rect 11444 50212 11445 50252
rect 11403 50203 11445 50212
rect 11307 49664 11349 49673
rect 11307 49624 11308 49664
rect 11348 49624 11349 49664
rect 11307 49615 11349 49624
rect 11308 49530 11348 49615
rect 11404 47984 11444 50203
rect 11596 50202 11636 50287
rect 11595 49664 11637 49673
rect 11595 49624 11596 49664
rect 11636 49624 11637 49664
rect 11595 49615 11637 49624
rect 11596 49496 11636 49615
rect 11596 49447 11636 49456
rect 11692 49496 11732 51043
rect 11980 51022 12020 51556
rect 11787 51008 11829 51017
rect 11787 50968 11788 51008
rect 11828 50968 11829 51008
rect 11980 50973 12020 50982
rect 11787 50959 11829 50968
rect 11499 48824 11541 48833
rect 11499 48784 11500 48824
rect 11540 48784 11541 48824
rect 11499 48775 11541 48784
rect 11500 48690 11540 48775
rect 11500 47984 11540 47993
rect 11692 47984 11732 49456
rect 11404 47944 11500 47984
rect 11500 47237 11540 47944
rect 11596 47944 11732 47984
rect 11499 47228 11541 47237
rect 11499 47188 11500 47228
rect 11540 47188 11541 47228
rect 11499 47179 11541 47188
rect 11403 46724 11445 46733
rect 11596 46724 11636 47944
rect 11403 46684 11404 46724
rect 11444 46684 11636 46724
rect 11692 47816 11732 47825
rect 11403 46675 11445 46684
rect 10828 46600 11156 46640
rect 11212 46600 11348 46640
rect 10731 46556 10773 46565
rect 10731 46516 10732 46556
rect 10772 46516 10773 46556
rect 10731 46507 10773 46516
rect 10923 46472 10965 46481
rect 10923 46432 10924 46472
rect 10964 46432 10965 46472
rect 10923 46423 10965 46432
rect 10924 46229 10964 46423
rect 10923 46220 10965 46229
rect 10923 46180 10924 46220
rect 10964 46180 10965 46220
rect 10923 46171 10965 46180
rect 11116 45968 11156 46600
rect 11212 45968 11252 45977
rect 11116 45928 11212 45968
rect 11212 45919 11252 45928
rect 11020 45786 11060 45795
rect 11020 45212 11060 45746
rect 11020 45163 11060 45172
rect 10827 44960 10869 44969
rect 10827 44920 10828 44960
rect 10868 44920 10869 44960
rect 10827 44911 10869 44920
rect 11211 44960 11253 44969
rect 11211 44920 11212 44960
rect 11252 44920 11253 44960
rect 11211 44911 11253 44920
rect 10828 44826 10868 44911
rect 11212 44288 11252 44911
rect 11308 44465 11348 46600
rect 11452 46481 11492 46490
rect 11692 46472 11732 47776
rect 11788 47069 11828 50959
rect 12076 50756 12116 51640
rect 12172 51101 12212 53479
rect 12268 52109 12308 54319
rect 12364 53537 12404 55243
rect 12555 54872 12597 54881
rect 12555 54823 12556 54872
rect 12596 54823 12597 54872
rect 12556 53957 12596 54811
rect 12555 53948 12597 53957
rect 12555 53908 12556 53948
rect 12596 53908 12597 53948
rect 12555 53899 12597 53908
rect 12363 53528 12405 53537
rect 12363 53488 12364 53528
rect 12404 53488 12405 53528
rect 12363 53479 12405 53488
rect 12556 53444 12596 53899
rect 12460 53404 12596 53444
rect 12364 53360 12404 53369
rect 12460 53360 12500 53404
rect 12404 53320 12500 53360
rect 12364 53311 12404 53320
rect 12363 52604 12405 52613
rect 12363 52564 12364 52604
rect 12404 52564 12405 52604
rect 12363 52555 12405 52564
rect 12267 52100 12309 52109
rect 12267 52060 12268 52100
rect 12308 52060 12309 52100
rect 12364 52100 12404 52555
rect 12460 52352 12500 53320
rect 12556 53108 12596 53117
rect 12556 52520 12596 53068
rect 12652 52697 12692 57016
rect 13036 55040 13076 58108
rect 13132 57644 13172 57653
rect 13132 57070 13172 57604
rect 13132 57021 13172 57030
rect 13131 56720 13173 56729
rect 13131 56680 13132 56720
rect 13172 56680 13173 56720
rect 13131 56671 13173 56680
rect 13132 55544 13172 56671
rect 13132 55495 13172 55504
rect 13228 56384 13268 58192
rect 13324 57737 13364 57822
rect 13323 57728 13365 57737
rect 13323 57688 13324 57728
rect 13364 57688 13365 57728
rect 13323 57679 13365 57688
rect 13323 57476 13365 57485
rect 13323 57436 13324 57476
rect 13364 57436 13365 57476
rect 13323 57427 13365 57436
rect 13324 56972 13364 57427
rect 13324 56923 13364 56932
rect 13323 56804 13365 56813
rect 13323 56764 13324 56804
rect 13364 56764 13365 56804
rect 13323 56755 13365 56764
rect 13036 55000 13172 55040
rect 12748 54956 12788 54965
rect 12788 54916 13076 54956
rect 12748 54907 12788 54916
rect 13036 54872 13076 54916
rect 13036 54823 13076 54832
rect 13132 54872 13172 55000
rect 13132 54536 13172 54832
rect 12844 54496 13172 54536
rect 12747 54032 12789 54041
rect 12747 53992 12748 54032
rect 12788 53992 12789 54032
rect 12747 53983 12789 53992
rect 12748 53360 12788 53983
rect 12748 53033 12788 53320
rect 12747 53024 12789 53033
rect 12747 52984 12748 53024
rect 12788 52984 12789 53024
rect 12747 52975 12789 52984
rect 12651 52688 12693 52697
rect 12651 52648 12652 52688
rect 12692 52648 12693 52688
rect 12651 52639 12693 52648
rect 12652 52520 12692 52529
rect 12556 52480 12652 52520
rect 12652 52471 12692 52480
rect 12748 52520 12788 52529
rect 12844 52520 12884 54496
rect 12939 54368 12981 54377
rect 12939 54328 12940 54368
rect 12980 54328 12981 54368
rect 12939 54319 12981 54328
rect 12788 52480 12884 52520
rect 12460 52312 12692 52352
rect 12364 52060 12500 52100
rect 12267 52051 12309 52060
rect 12363 51932 12405 51941
rect 12363 51892 12364 51932
rect 12404 51892 12405 51932
rect 12363 51883 12405 51892
rect 12364 51260 12404 51883
rect 12460 51680 12500 52060
rect 12652 51857 12692 52312
rect 12651 51848 12693 51857
rect 12651 51808 12652 51848
rect 12692 51808 12693 51848
rect 12651 51799 12693 51808
rect 12460 51640 12692 51680
rect 12364 51211 12404 51220
rect 12171 51092 12213 51101
rect 12171 51052 12172 51092
rect 12212 51052 12213 51092
rect 12171 51043 12213 51052
rect 12556 51092 12596 51101
rect 12556 51008 12596 51052
rect 12268 50968 12596 51008
rect 12172 50924 12212 50933
rect 12268 50924 12308 50968
rect 12212 50884 12308 50924
rect 12172 50875 12212 50884
rect 12076 50716 12500 50756
rect 12267 50588 12309 50597
rect 12267 50548 12268 50588
rect 12308 50548 12309 50588
rect 12267 50539 12309 50548
rect 12075 49832 12117 49841
rect 12075 49792 12076 49832
rect 12116 49792 12117 49832
rect 12075 49783 12117 49792
rect 12076 49580 12116 49783
rect 11883 48656 11925 48665
rect 11883 48616 11884 48656
rect 11924 48616 11925 48656
rect 11883 48607 11925 48616
rect 11787 47060 11829 47069
rect 11787 47020 11788 47060
rect 11828 47020 11829 47060
rect 11787 47011 11829 47020
rect 11884 46556 11924 48607
rect 12076 46640 12116 49540
rect 12171 49580 12213 49589
rect 12171 49540 12172 49580
rect 12212 49540 12213 49580
rect 12171 49531 12213 49540
rect 12172 49446 12212 49531
rect 12076 46600 12212 46640
rect 11884 46507 11924 46516
rect 11492 46441 11732 46472
rect 11452 46432 11732 46441
rect 11596 46304 11636 46313
rect 11596 45716 11636 46264
rect 12076 46304 12116 46313
rect 12076 46061 12116 46264
rect 12075 46052 12117 46061
rect 12075 46012 12076 46052
rect 12116 46012 12117 46052
rect 12075 46003 12117 46012
rect 11596 45667 11636 45676
rect 11404 45548 11444 45557
rect 11404 45137 11444 45508
rect 11883 45380 11925 45389
rect 11883 45340 11884 45380
rect 11924 45340 11925 45380
rect 11883 45331 11925 45340
rect 11403 45128 11445 45137
rect 11403 45088 11404 45128
rect 11444 45088 11445 45128
rect 11403 45079 11445 45088
rect 11307 44456 11349 44465
rect 11307 44416 11308 44456
rect 11348 44416 11349 44456
rect 11307 44407 11349 44416
rect 11308 44288 11348 44297
rect 11788 44288 11828 44297
rect 11212 44248 11308 44288
rect 10635 44204 10677 44213
rect 10635 44164 10636 44204
rect 10676 44164 10677 44204
rect 10635 44155 10677 44164
rect 11212 43448 11252 44248
rect 11308 44239 11348 44248
rect 11404 44248 11788 44288
rect 11404 43700 11444 44248
rect 11788 44239 11828 44248
rect 11884 44288 11924 45331
rect 12075 45128 12117 45137
rect 12075 45088 12076 45128
rect 12116 45088 12117 45128
rect 12075 45079 12117 45088
rect 12076 44960 12116 45079
rect 12076 44911 12116 44920
rect 11500 44036 11540 44045
rect 11540 43996 11732 44036
rect 11500 43987 11540 43996
rect 11404 43651 11444 43660
rect 11212 43399 11252 43408
rect 11692 43448 11732 43996
rect 11692 43399 11732 43408
rect 11788 43448 11828 43457
rect 11884 43448 11924 44248
rect 11828 43408 11924 43448
rect 12172 44204 12212 46600
rect 12268 46565 12308 50539
rect 12364 47312 12404 47323
rect 12364 47237 12404 47272
rect 12363 47228 12405 47237
rect 12363 47188 12364 47228
rect 12404 47188 12405 47228
rect 12363 47179 12405 47188
rect 12363 47060 12405 47069
rect 12363 47020 12364 47060
rect 12404 47020 12405 47060
rect 12363 47011 12405 47020
rect 12364 46733 12404 47011
rect 12363 46724 12405 46733
rect 12363 46684 12364 46724
rect 12404 46684 12405 46724
rect 12363 46675 12405 46684
rect 12267 46556 12309 46565
rect 12267 46516 12268 46556
rect 12308 46516 12309 46556
rect 12267 46507 12309 46516
rect 12268 45389 12308 46507
rect 12267 45380 12309 45389
rect 12267 45340 12268 45380
rect 12308 45340 12309 45380
rect 12267 45331 12309 45340
rect 12364 44288 12404 46675
rect 12460 44624 12500 50716
rect 12652 49496 12692 51640
rect 12748 51017 12788 52480
rect 12747 51008 12789 51017
rect 12747 50968 12748 51008
rect 12788 50968 12789 51008
rect 12747 50959 12789 50968
rect 12843 50336 12885 50345
rect 12843 50296 12844 50336
rect 12884 50296 12885 50336
rect 12843 50287 12885 50296
rect 12747 49748 12789 49757
rect 12747 49708 12748 49748
rect 12788 49708 12789 49748
rect 12747 49699 12789 49708
rect 12652 49447 12692 49456
rect 12748 48824 12788 49699
rect 12844 49421 12884 50287
rect 12940 49505 12980 54319
rect 13131 53948 13173 53957
rect 13131 53908 13132 53948
rect 13172 53908 13173 53948
rect 13131 53899 13173 53908
rect 13132 52772 13172 53899
rect 13228 52949 13268 56344
rect 13227 52940 13269 52949
rect 13227 52900 13228 52940
rect 13268 52900 13269 52940
rect 13227 52891 13269 52900
rect 13132 52732 13268 52772
rect 13035 52688 13077 52697
rect 13035 52648 13036 52688
rect 13076 52648 13077 52688
rect 13035 52639 13077 52648
rect 13036 52193 13076 52639
rect 13132 52520 13172 52529
rect 13132 52277 13172 52480
rect 13228 52520 13268 52732
rect 13228 52361 13268 52480
rect 13227 52352 13269 52361
rect 13227 52312 13228 52352
rect 13268 52312 13269 52352
rect 13227 52303 13269 52312
rect 13131 52268 13173 52277
rect 13131 52228 13132 52268
rect 13172 52228 13173 52268
rect 13131 52219 13173 52228
rect 13035 52184 13077 52193
rect 13035 52144 13036 52184
rect 13076 52144 13077 52184
rect 13035 52135 13077 52144
rect 13324 51941 13364 56755
rect 13420 54377 13460 60208
rect 13516 58661 13556 60871
rect 13612 58829 13652 61552
rect 13611 58820 13653 58829
rect 13611 58780 13612 58820
rect 13652 58780 13653 58820
rect 13611 58771 13653 58780
rect 13515 58652 13557 58661
rect 13515 58612 13516 58652
rect 13556 58612 13557 58652
rect 13515 58603 13557 58612
rect 13516 58568 13556 58603
rect 13516 58518 13556 58528
rect 13611 58568 13653 58577
rect 13611 58528 13612 58568
rect 13652 58528 13653 58568
rect 13611 58519 13653 58528
rect 13516 57896 13556 57907
rect 13516 57821 13556 57856
rect 13515 57812 13557 57821
rect 13515 57772 13516 57812
rect 13556 57772 13557 57812
rect 13515 57763 13557 57772
rect 13612 55544 13652 58519
rect 13516 55504 13652 55544
rect 13516 55040 13556 55504
rect 13708 55385 13748 62378
rect 13899 61676 13941 61685
rect 13899 61636 13900 61676
rect 13940 61636 13941 61676
rect 13899 61627 13941 61636
rect 13900 60920 13940 61627
rect 13996 61013 14036 63232
rect 13995 61004 14037 61013
rect 13995 60964 13996 61004
rect 14036 60964 14037 61004
rect 13995 60955 14037 60964
rect 13900 60332 13940 60880
rect 13996 60920 14036 60955
rect 13996 60869 14036 60880
rect 14092 60836 14132 64324
rect 14284 64280 14324 64819
rect 14379 64700 14421 64709
rect 14379 64660 14380 64700
rect 14420 64660 14421 64700
rect 14379 64651 14421 64660
rect 14188 64240 14324 64280
rect 14188 61181 14228 64240
rect 14380 63944 14420 64651
rect 14380 63895 14420 63904
rect 14283 63860 14325 63869
rect 14283 63820 14284 63860
rect 14324 63820 14325 63860
rect 14283 63811 14325 63820
rect 14284 63726 14324 63811
rect 14476 63104 14516 64819
rect 14476 63055 14516 63064
rect 14572 62432 14612 69532
rect 14668 64373 14708 82720
rect 15820 81500 15860 85936
rect 15820 81451 15860 81460
rect 15916 83516 15956 83525
rect 15627 81332 15669 81341
rect 15627 81292 15628 81332
rect 15668 81292 15669 81332
rect 15627 81283 15669 81292
rect 15628 81198 15668 81283
rect 15820 79820 15860 79829
rect 15820 79073 15860 79780
rect 15819 79064 15861 79073
rect 15819 79024 15820 79064
rect 15860 79024 15861 79064
rect 15819 79015 15861 79024
rect 15339 75704 15381 75713
rect 15339 75664 15340 75704
rect 15380 75664 15381 75704
rect 15339 75655 15381 75664
rect 15051 72344 15093 72353
rect 15051 72304 15052 72344
rect 15092 72304 15093 72344
rect 15051 72295 15093 72304
rect 15052 71504 15092 72295
rect 15244 72176 15284 72185
rect 15148 72136 15244 72176
rect 15148 71849 15188 72136
rect 15244 72127 15284 72136
rect 15147 71840 15189 71849
rect 15147 71800 15148 71840
rect 15188 71800 15189 71840
rect 15147 71791 15189 71800
rect 15052 71455 15092 71464
rect 15052 70841 15092 70926
rect 15051 70832 15093 70841
rect 15051 70792 15052 70832
rect 15092 70792 15093 70832
rect 15051 70783 15093 70792
rect 14764 70664 14804 70673
rect 14764 69329 14804 70624
rect 14859 70664 14901 70673
rect 14859 70624 14860 70664
rect 14900 70624 14901 70664
rect 14859 70615 14901 70624
rect 15051 70664 15093 70673
rect 15051 70624 15052 70664
rect 15092 70624 15093 70664
rect 15051 70615 15093 70624
rect 14860 70530 14900 70615
rect 15052 70530 15092 70615
rect 14956 69908 14996 69917
rect 14860 69868 14956 69908
rect 14763 69320 14805 69329
rect 14763 69280 14764 69320
rect 14804 69280 14805 69320
rect 14763 69271 14805 69280
rect 14763 69152 14805 69161
rect 14763 69112 14764 69152
rect 14804 69112 14805 69152
rect 14763 69103 14805 69112
rect 14764 67136 14804 69103
rect 14860 68312 14900 69868
rect 14956 69859 14996 69868
rect 15052 69908 15092 69919
rect 15052 69833 15092 69868
rect 15051 69824 15093 69833
rect 15051 69784 15052 69824
rect 15092 69784 15093 69824
rect 15051 69775 15093 69784
rect 15148 69572 15188 71791
rect 15340 71672 15380 75655
rect 15916 73100 15956 83476
rect 16012 79988 16052 85936
rect 16012 79939 16052 79948
rect 15916 73060 16148 73100
rect 16012 72932 16052 72941
rect 15915 72260 15957 72269
rect 15915 72220 15916 72260
rect 15956 72220 15957 72260
rect 15915 72211 15957 72220
rect 15724 72176 15764 72185
rect 15436 72092 15476 72101
rect 15724 72092 15764 72136
rect 15476 72052 15764 72092
rect 15820 72176 15860 72185
rect 15436 72043 15476 72052
rect 15820 71765 15860 72136
rect 15819 71756 15861 71765
rect 15819 71716 15820 71756
rect 15860 71716 15861 71756
rect 15819 71707 15861 71716
rect 15340 71632 15668 71672
rect 15244 71588 15284 71597
rect 15284 71548 15572 71588
rect 15244 71539 15284 71548
rect 15244 70664 15284 70675
rect 15244 70589 15284 70624
rect 15340 70664 15380 70673
rect 15243 70580 15285 70589
rect 15243 70540 15244 70580
rect 15284 70540 15285 70580
rect 15243 70531 15285 70540
rect 15340 70169 15380 70624
rect 15436 70664 15476 71548
rect 15532 71504 15572 71548
rect 15532 71455 15572 71464
rect 15436 70615 15476 70624
rect 15531 70664 15573 70673
rect 15531 70624 15532 70664
rect 15572 70624 15573 70664
rect 15531 70615 15573 70624
rect 15532 70530 15572 70615
rect 15628 70496 15668 71632
rect 15724 71504 15764 71513
rect 15916 71504 15956 72211
rect 15764 71464 15860 71504
rect 15724 71455 15764 71464
rect 15724 71252 15764 71261
rect 15724 70664 15764 71212
rect 15820 71093 15860 71464
rect 15916 71455 15956 71464
rect 15819 71084 15861 71093
rect 15819 71044 15820 71084
rect 15860 71044 15861 71084
rect 15819 71035 15861 71044
rect 16012 71009 16052 72892
rect 16108 71597 16148 73060
rect 16204 72848 16244 85936
rect 16396 84449 16436 85936
rect 16588 84449 16628 85936
rect 16395 84440 16437 84449
rect 16395 84400 16396 84440
rect 16436 84400 16437 84440
rect 16395 84391 16437 84400
rect 16587 84440 16629 84449
rect 16587 84400 16588 84440
rect 16628 84400 16629 84440
rect 16587 84391 16629 84400
rect 16780 83768 16820 85936
rect 16875 85868 16917 85877
rect 16875 85828 16876 85868
rect 16916 85828 16917 85868
rect 16875 85819 16917 85828
rect 16780 83719 16820 83728
rect 16204 72799 16244 72808
rect 16588 83516 16628 83525
rect 16204 72176 16244 72185
rect 16204 71933 16244 72136
rect 16300 72176 16340 72185
rect 16203 71924 16245 71933
rect 16203 71884 16204 71924
rect 16244 71884 16245 71924
rect 16203 71875 16245 71884
rect 16203 71756 16245 71765
rect 16203 71716 16204 71756
rect 16244 71716 16245 71756
rect 16203 71707 16245 71716
rect 16107 71588 16149 71597
rect 16107 71548 16108 71588
rect 16148 71548 16149 71588
rect 16107 71539 16149 71548
rect 16204 71420 16244 71707
rect 16108 71380 16244 71420
rect 16011 71000 16053 71009
rect 16011 70960 16012 71000
rect 16052 70960 16053 71000
rect 16011 70951 16053 70960
rect 15724 70615 15764 70624
rect 15915 70664 15957 70673
rect 15915 70624 15916 70664
rect 15956 70624 15957 70664
rect 15915 70615 15957 70624
rect 15820 70580 15860 70589
rect 15820 70496 15860 70540
rect 15916 70530 15956 70615
rect 15628 70456 15860 70496
rect 15915 70412 15957 70421
rect 15915 70372 15916 70412
rect 15956 70372 15957 70412
rect 15915 70363 15957 70372
rect 15723 70328 15765 70337
rect 15723 70288 15724 70328
rect 15764 70288 15765 70328
rect 15723 70279 15765 70288
rect 15339 70160 15381 70169
rect 15339 70120 15340 70160
rect 15380 70120 15381 70160
rect 15339 70111 15381 70120
rect 15532 69992 15572 70001
rect 15532 69917 15572 69952
rect 15531 69908 15573 69917
rect 15531 69868 15532 69908
rect 15572 69868 15573 69908
rect 15531 69859 15573 69868
rect 15052 69532 15188 69572
rect 15052 69245 15092 69532
rect 15243 69488 15285 69497
rect 15243 69448 15244 69488
rect 15284 69448 15285 69488
rect 15243 69439 15285 69448
rect 15147 69404 15189 69413
rect 15147 69364 15148 69404
rect 15188 69364 15189 69404
rect 15147 69355 15189 69364
rect 15148 69270 15188 69355
rect 15051 69236 15093 69245
rect 15051 69196 15052 69236
rect 15092 69196 15093 69236
rect 15051 69187 15093 69196
rect 14955 69152 14997 69161
rect 14955 69112 14956 69152
rect 14996 69112 14997 69152
rect 14955 69103 14997 69112
rect 14956 69018 14996 69103
rect 14956 68489 14996 68574
rect 14955 68480 14997 68489
rect 14955 68440 14956 68480
rect 14996 68440 14997 68480
rect 14955 68431 14997 68440
rect 14860 68272 14996 68312
rect 14859 67724 14901 67733
rect 14859 67684 14860 67724
rect 14900 67684 14901 67724
rect 14859 67675 14901 67684
rect 14860 67640 14900 67675
rect 14860 67589 14900 67600
rect 14956 67640 14996 68272
rect 15148 68228 15188 68237
rect 15051 68060 15093 68069
rect 15051 68020 15052 68060
rect 15092 68020 15093 68060
rect 15051 68011 15093 68020
rect 14764 67096 14900 67136
rect 14763 66968 14805 66977
rect 14763 66928 14764 66968
rect 14804 66928 14805 66968
rect 14763 66919 14805 66928
rect 14764 64877 14804 66919
rect 14860 65465 14900 67096
rect 14956 66389 14996 67600
rect 15052 67556 15092 68011
rect 15148 67733 15188 68188
rect 15244 67808 15284 69439
rect 15339 69320 15381 69329
rect 15339 69280 15340 69320
rect 15380 69280 15381 69320
rect 15339 69271 15381 69280
rect 15340 69186 15380 69271
rect 15340 68480 15380 68489
rect 15340 68321 15380 68440
rect 15339 68312 15381 68321
rect 15339 68272 15340 68312
rect 15380 68272 15381 68312
rect 15339 68263 15381 68272
rect 15244 67768 15380 67808
rect 15147 67724 15189 67733
rect 15147 67684 15148 67724
rect 15188 67684 15189 67724
rect 15147 67675 15189 67684
rect 15340 67724 15380 67768
rect 15340 67675 15380 67684
rect 15435 67724 15477 67733
rect 15435 67684 15436 67724
rect 15476 67684 15477 67724
rect 15435 67675 15477 67684
rect 15436 67590 15476 67675
rect 15532 67565 15572 69859
rect 15724 69152 15764 70279
rect 15628 69068 15668 69079
rect 15628 68993 15668 69028
rect 15627 68984 15669 68993
rect 15627 68944 15628 68984
rect 15668 68944 15669 68984
rect 15627 68935 15669 68944
rect 15627 68144 15669 68153
rect 15627 68104 15628 68144
rect 15668 68104 15669 68144
rect 15627 68095 15669 68104
rect 15531 67556 15573 67565
rect 15052 67516 15284 67556
rect 14955 66380 14997 66389
rect 14955 66340 14956 66380
rect 14996 66340 14997 66380
rect 14955 66331 14997 66340
rect 14859 65456 14901 65465
rect 14859 65416 14860 65456
rect 14900 65416 14901 65456
rect 14859 65407 14901 65416
rect 14860 65213 14900 65407
rect 14859 65204 14901 65213
rect 14859 65164 14860 65204
rect 14900 65164 14901 65204
rect 14859 65155 14901 65164
rect 14763 64868 14805 64877
rect 14763 64828 14764 64868
rect 14804 64828 14805 64868
rect 14763 64819 14805 64828
rect 14859 64700 14901 64709
rect 14859 64660 14860 64700
rect 14900 64660 14901 64700
rect 14859 64651 14901 64660
rect 14667 64364 14709 64373
rect 14667 64324 14668 64364
rect 14708 64324 14709 64364
rect 14667 64315 14709 64324
rect 14763 64196 14805 64205
rect 14763 64156 14764 64196
rect 14804 64156 14805 64196
rect 14763 64147 14805 64156
rect 14667 63944 14709 63953
rect 14667 63904 14668 63944
rect 14708 63904 14709 63944
rect 14667 63895 14709 63904
rect 14668 63356 14708 63895
rect 14764 63356 14804 64147
rect 14860 64112 14900 64651
rect 15244 64280 15284 67516
rect 15531 67516 15532 67556
rect 15572 67516 15573 67556
rect 15531 67507 15573 67516
rect 15628 67481 15668 68095
rect 15724 67733 15764 69112
rect 15819 68480 15861 68489
rect 15819 68440 15820 68480
rect 15860 68440 15861 68480
rect 15819 68431 15861 68440
rect 15723 67724 15765 67733
rect 15723 67684 15724 67724
rect 15764 67684 15765 67724
rect 15723 67675 15765 67684
rect 15435 67472 15477 67481
rect 15435 67432 15436 67472
rect 15476 67432 15477 67472
rect 15435 67423 15477 67432
rect 15627 67472 15669 67481
rect 15627 67432 15628 67472
rect 15668 67432 15669 67472
rect 15627 67423 15669 67432
rect 15436 66968 15476 67423
rect 15627 67304 15669 67313
rect 15627 67264 15628 67304
rect 15668 67264 15669 67304
rect 15627 67255 15669 67264
rect 15339 64700 15381 64709
rect 15339 64660 15340 64700
rect 15380 64660 15381 64700
rect 15339 64651 15381 64660
rect 15340 64616 15380 64651
rect 15340 64565 15380 64576
rect 15436 64280 15476 66928
rect 15628 66968 15668 67255
rect 15628 66919 15668 66928
rect 15724 66884 15764 67675
rect 15820 66977 15860 68431
rect 15916 67808 15956 70363
rect 16012 70001 16052 70102
rect 16011 69992 16053 70001
rect 16011 69943 16012 69992
rect 16052 69943 16053 69992
rect 16012 69413 16052 69938
rect 16108 69749 16148 71380
rect 16203 71084 16245 71093
rect 16203 71044 16204 71084
rect 16244 71044 16245 71084
rect 16203 71035 16245 71044
rect 16204 70160 16244 71035
rect 16204 70111 16244 70120
rect 16300 70085 16340 72136
rect 16588 71681 16628 83476
rect 16876 83348 16916 85819
rect 16972 83516 17012 85936
rect 17164 83684 17204 85936
rect 17356 83768 17396 85936
rect 17548 84440 17588 85936
rect 17740 84524 17780 85936
rect 17740 84484 17876 84524
rect 17548 84400 17780 84440
rect 17356 83719 17396 83728
rect 17740 83768 17780 84400
rect 17740 83719 17780 83728
rect 17836 83684 17876 84484
rect 17932 83861 17972 85936
rect 18124 84272 18164 85936
rect 18124 84232 18260 84272
rect 18124 84104 18164 84113
rect 17931 83852 17973 83861
rect 17931 83812 17932 83852
rect 17972 83812 17973 83852
rect 17931 83803 17973 83812
rect 17164 83644 17300 83684
rect 17836 83644 18068 83684
rect 17164 83516 17204 83525
rect 16972 83476 17108 83516
rect 16972 83348 17012 83357
rect 16876 83308 16972 83348
rect 16972 83299 17012 83308
rect 16972 79232 17012 79241
rect 17068 79232 17108 83476
rect 17012 79192 17108 79232
rect 16972 79183 17012 79192
rect 16780 78980 16820 78989
rect 16780 72353 16820 78940
rect 17164 77552 17204 83476
rect 17068 77512 17204 77552
rect 16972 76796 17012 76805
rect 16972 73100 17012 76756
rect 17068 76712 17108 77512
rect 17164 76880 17204 76889
rect 17260 76880 17300 83644
rect 17548 83516 17588 83525
rect 17452 82928 17492 82937
rect 17548 82928 17588 83476
rect 17932 83516 17972 83525
rect 17492 82888 17588 82928
rect 17836 82928 17876 82937
rect 17932 82928 17972 83476
rect 18028 83348 18068 83644
rect 18124 83525 18164 84064
rect 18123 83516 18165 83525
rect 18123 83476 18124 83516
rect 18164 83476 18165 83516
rect 18123 83467 18165 83476
rect 18124 83348 18164 83357
rect 18028 83308 18124 83348
rect 18124 83299 18164 83308
rect 18220 83012 18260 84232
rect 18316 83777 18356 85936
rect 18508 84272 18548 85936
rect 18508 84232 18644 84272
rect 18508 84104 18548 84113
rect 18411 83852 18453 83861
rect 18411 83812 18412 83852
rect 18452 83812 18453 83852
rect 18411 83803 18453 83812
rect 18315 83768 18357 83777
rect 18315 83728 18316 83768
rect 18356 83728 18357 83768
rect 18315 83719 18357 83728
rect 18315 83516 18357 83525
rect 18315 83476 18316 83516
rect 18356 83476 18357 83516
rect 18315 83467 18357 83476
rect 18316 83382 18356 83467
rect 18412 83348 18452 83803
rect 18508 83525 18548 84064
rect 18507 83516 18549 83525
rect 18507 83476 18508 83516
rect 18548 83476 18549 83516
rect 18507 83467 18549 83476
rect 18508 83348 18548 83357
rect 18412 83308 18508 83348
rect 18508 83299 18548 83308
rect 18220 82963 18260 82972
rect 18604 83012 18644 84232
rect 18700 83684 18740 85936
rect 18892 84860 18932 85936
rect 19084 85037 19124 85936
rect 19083 85028 19125 85037
rect 19083 84988 19084 85028
rect 19124 84988 19125 85028
rect 19083 84979 19125 84988
rect 19276 84944 19316 85936
rect 19468 85196 19508 85936
rect 19468 85156 19988 85196
rect 19659 85028 19701 85037
rect 19659 84988 19660 85028
rect 19700 84988 19701 85028
rect 19659 84979 19701 84988
rect 19276 84904 19604 84944
rect 18892 84820 19412 84860
rect 18808 84692 19176 84701
rect 18848 84652 18890 84692
rect 18930 84652 18972 84692
rect 19012 84652 19054 84692
rect 19094 84652 19136 84692
rect 18808 84643 19176 84652
rect 18988 84104 19028 84113
rect 19276 84104 19316 84113
rect 19028 84064 19124 84104
rect 18988 84055 19028 84064
rect 18891 83768 18933 83777
rect 18891 83728 18892 83768
rect 18932 83728 18933 83768
rect 18891 83719 18933 83728
rect 18700 83644 18836 83684
rect 18699 83516 18741 83525
rect 18699 83476 18700 83516
rect 18740 83476 18741 83516
rect 18699 83467 18741 83476
rect 18700 83382 18740 83467
rect 18796 83357 18836 83644
rect 18892 83634 18932 83719
rect 19084 83525 19124 84064
rect 19276 83525 19316 84064
rect 19083 83516 19125 83525
rect 19083 83476 19084 83516
rect 19124 83476 19125 83516
rect 19083 83467 19125 83476
rect 19275 83516 19317 83525
rect 19275 83476 19276 83516
rect 19316 83476 19317 83516
rect 19275 83467 19317 83476
rect 19084 83382 19124 83467
rect 18795 83348 18837 83357
rect 18795 83308 18796 83348
rect 18836 83308 18837 83348
rect 18795 83299 18837 83308
rect 19275 83348 19317 83357
rect 19275 83308 19276 83348
rect 19316 83308 19317 83348
rect 19275 83299 19317 83308
rect 19276 83214 19316 83299
rect 18808 83180 19176 83189
rect 18848 83140 18890 83180
rect 18930 83140 18972 83180
rect 19012 83140 19054 83180
rect 19094 83140 19136 83180
rect 18808 83131 19176 83140
rect 19372 83096 19412 84820
rect 19467 83516 19509 83525
rect 19467 83476 19468 83516
rect 19508 83476 19509 83516
rect 19467 83467 19509 83476
rect 19468 83382 19508 83467
rect 19276 83056 19412 83096
rect 18604 82963 18644 82972
rect 18988 83012 19028 83021
rect 19276 83012 19316 83056
rect 19028 82972 19316 83012
rect 18988 82963 19028 82972
rect 17876 82888 17972 82928
rect 19372 82928 19412 82937
rect 19564 82928 19604 84904
rect 19660 83768 19700 84979
rect 19948 83768 19988 85156
rect 20048 83936 20416 83945
rect 20088 83896 20130 83936
rect 20170 83896 20212 83936
rect 20252 83896 20294 83936
rect 20334 83896 20376 83936
rect 20048 83887 20416 83896
rect 20044 83768 20084 83777
rect 19948 83728 20044 83768
rect 19660 83719 19700 83728
rect 20044 83719 20084 83728
rect 19852 83516 19892 83525
rect 19412 82888 19604 82928
rect 19756 82928 19796 82937
rect 19852 82928 19892 83476
rect 20236 83516 20276 83525
rect 19796 82888 19892 82928
rect 20140 82928 20180 82937
rect 20236 82928 20276 83476
rect 20180 82888 20276 82928
rect 17452 82879 17492 82888
rect 17836 82879 17876 82888
rect 19372 82879 19412 82888
rect 19756 82879 19796 82888
rect 20140 82879 20180 82888
rect 18028 82844 18068 82853
rect 17355 82592 17397 82601
rect 17355 82552 17356 82592
rect 17396 82552 17397 82592
rect 17355 82543 17397 82552
rect 17739 82592 17781 82601
rect 17739 82552 17740 82592
rect 17780 82552 17781 82592
rect 17739 82543 17781 82552
rect 17356 82458 17396 82543
rect 17740 82458 17780 82543
rect 18028 82256 18068 82804
rect 18028 82207 18068 82216
rect 18412 82844 18452 82853
rect 18412 82256 18452 82804
rect 18412 82207 18452 82216
rect 18796 82844 18836 82853
rect 18699 82088 18741 82097
rect 18699 82048 18700 82088
rect 18740 82048 18741 82088
rect 18699 82039 18741 82048
rect 18123 81920 18165 81929
rect 18123 81880 18124 81920
rect 18164 81880 18165 81920
rect 18123 81871 18165 81880
rect 18507 81920 18549 81929
rect 18507 81880 18508 81920
rect 18548 81880 18549 81920
rect 18507 81871 18549 81880
rect 18124 81786 18164 81871
rect 18508 81786 18548 81871
rect 17204 76840 17300 76880
rect 17164 76831 17204 76840
rect 17068 76672 17300 76712
rect 17260 73100 17300 76672
rect 16972 73060 17204 73100
rect 17260 73060 17492 73100
rect 16779 72344 16821 72353
rect 16779 72304 16780 72344
rect 16820 72304 16821 72344
rect 16779 72295 16821 72304
rect 16780 72176 16820 72185
rect 16820 72136 17108 72176
rect 16780 72127 16820 72136
rect 16587 71672 16629 71681
rect 16587 71632 16588 71672
rect 16628 71632 16629 71672
rect 16587 71623 16629 71632
rect 16395 71588 16437 71597
rect 16395 71548 16396 71588
rect 16436 71548 16437 71588
rect 16395 71539 16437 71548
rect 16396 70916 16436 71539
rect 16396 70867 16436 70876
rect 16972 70664 17012 70673
rect 16395 70160 16437 70169
rect 16876 70160 16916 70169
rect 16395 70120 16396 70160
rect 16436 70120 16437 70160
rect 16395 70111 16437 70120
rect 16492 70120 16876 70160
rect 16299 70076 16341 70085
rect 16299 70036 16300 70076
rect 16340 70036 16341 70076
rect 16299 70027 16341 70036
rect 16396 70026 16436 70111
rect 16492 69992 16532 70120
rect 16876 70111 16916 70120
rect 16492 69943 16532 69952
rect 16587 69992 16629 70001
rect 16587 69952 16588 69992
rect 16628 69952 16629 69992
rect 16587 69943 16629 69952
rect 16684 69992 16724 70001
rect 16588 69858 16628 69943
rect 16107 69740 16149 69749
rect 16107 69700 16108 69740
rect 16148 69700 16149 69740
rect 16107 69691 16149 69700
rect 16299 69656 16341 69665
rect 16299 69616 16300 69656
rect 16340 69616 16341 69656
rect 16299 69607 16341 69616
rect 16011 69404 16053 69413
rect 16011 69364 16012 69404
rect 16052 69364 16053 69404
rect 16011 69355 16053 69364
rect 16012 69152 16052 69355
rect 16012 69103 16052 69112
rect 16300 68489 16340 69607
rect 16684 69581 16724 69952
rect 16972 69824 17012 70624
rect 17068 70244 17108 72136
rect 17164 71849 17204 73060
rect 17308 72185 17348 72194
rect 17348 72145 17396 72176
rect 17308 72136 17396 72145
rect 17163 71840 17205 71849
rect 17163 71800 17164 71840
rect 17204 71800 17205 71840
rect 17163 71791 17205 71800
rect 17164 71504 17204 71791
rect 17356 71672 17396 72136
rect 17452 72092 17492 73060
rect 17452 72043 17492 72052
rect 18315 71924 18357 71933
rect 18315 71884 18316 71924
rect 18356 71884 18357 71924
rect 18315 71875 18357 71884
rect 17356 71623 17396 71632
rect 17164 71455 17204 71464
rect 17548 71504 17588 71515
rect 17548 71429 17588 71464
rect 17547 71420 17589 71429
rect 17547 71380 17548 71420
rect 17588 71380 17589 71420
rect 17547 71371 17589 71380
rect 18123 70916 18165 70925
rect 18123 70876 18124 70916
rect 18164 70876 18165 70916
rect 18123 70867 18165 70876
rect 17644 70664 17684 70673
rect 17644 70505 17684 70624
rect 17643 70496 17685 70505
rect 17643 70456 17644 70496
rect 17684 70456 17685 70496
rect 17643 70447 17685 70456
rect 18124 70244 18164 70867
rect 17068 70204 17492 70244
rect 17068 70001 17108 70086
rect 17163 70076 17205 70085
rect 17163 70036 17164 70076
rect 17204 70036 17205 70076
rect 17163 70027 17205 70036
rect 17067 69992 17109 70001
rect 17067 69952 17068 69992
rect 17108 69952 17109 69992
rect 17067 69943 17109 69952
rect 17164 69992 17204 70027
rect 17164 69941 17204 69952
rect 16972 69784 17204 69824
rect 16683 69572 16725 69581
rect 16683 69532 16684 69572
rect 16724 69532 16725 69572
rect 16683 69523 16725 69532
rect 16396 69152 16436 69161
rect 16396 68657 16436 69112
rect 16395 68648 16437 68657
rect 16395 68608 16396 68648
rect 16436 68608 16437 68648
rect 16395 68599 16437 68608
rect 16299 68480 16341 68489
rect 16588 68480 16628 68489
rect 16972 68480 17012 68489
rect 16299 68440 16300 68480
rect 16340 68440 16588 68480
rect 16299 68431 16341 68440
rect 16588 68431 16628 68440
rect 16876 68440 16972 68480
rect 16300 68346 16340 68431
rect 16780 68228 16820 68237
rect 16299 67808 16341 67817
rect 15916 67768 16052 67808
rect 15916 67640 15956 67651
rect 15916 67565 15956 67600
rect 15915 67556 15957 67565
rect 15915 67516 15916 67556
rect 15956 67516 15957 67556
rect 15915 67507 15957 67516
rect 15819 66968 15861 66977
rect 15819 66928 15820 66968
rect 15860 66928 15861 66968
rect 15819 66919 15861 66928
rect 15703 66844 15764 66884
rect 15703 66800 15743 66844
rect 15628 66760 15743 66800
rect 15628 65204 15668 66760
rect 16012 66557 16052 67768
rect 16299 67768 16300 67808
rect 16340 67768 16341 67808
rect 16299 67759 16341 67768
rect 16107 67640 16149 67649
rect 16107 67600 16108 67640
rect 16148 67600 16149 67640
rect 16107 67591 16149 67600
rect 16011 66548 16053 66557
rect 16011 66508 16012 66548
rect 16052 66508 16053 66548
rect 16011 66499 16053 66508
rect 16108 66380 16148 67591
rect 16203 67556 16245 67565
rect 16203 67516 16204 67556
rect 16244 67516 16245 67556
rect 16203 67507 16245 67516
rect 16108 66331 16148 66340
rect 16011 66128 16053 66137
rect 16011 66088 16012 66128
rect 16052 66088 16053 66128
rect 16011 66079 16053 66088
rect 16012 65994 16052 66079
rect 16204 65876 16244 67507
rect 16300 67388 16340 67759
rect 16396 67645 16436 67654
rect 16780 67640 16820 68188
rect 16876 67733 16916 68440
rect 16972 68431 17012 68440
rect 17067 67808 17109 67817
rect 17067 67768 17068 67808
rect 17108 67768 17109 67808
rect 17067 67759 17109 67768
rect 16875 67724 16917 67733
rect 16875 67684 16876 67724
rect 16916 67684 16917 67724
rect 16875 67675 16917 67684
rect 16436 67605 16780 67640
rect 16396 67600 16780 67605
rect 16396 67596 16436 67600
rect 16780 67591 16820 67600
rect 16971 67640 17013 67649
rect 16971 67600 16972 67640
rect 17012 67600 17013 67640
rect 16971 67591 17013 67600
rect 17068 67640 17108 67759
rect 17068 67591 17108 67600
rect 16972 67506 17012 67591
rect 16491 67472 16533 67481
rect 16491 67432 16492 67472
rect 16532 67432 16533 67472
rect 16491 67423 16533 67432
rect 16588 67472 16628 67481
rect 16300 67348 16436 67388
rect 16299 66548 16341 66557
rect 16299 66508 16300 66548
rect 16340 66508 16341 66548
rect 16299 66499 16341 66508
rect 16300 66128 16340 66499
rect 16300 65960 16340 66088
rect 16396 66128 16436 67348
rect 16396 66079 16436 66088
rect 16492 66128 16532 67423
rect 16588 66389 16628 67432
rect 16875 67472 16917 67481
rect 16875 67432 16876 67472
rect 16916 67432 16917 67472
rect 16875 67423 16917 67432
rect 16876 67338 16916 67423
rect 16875 66968 16917 66977
rect 16875 66928 16876 66968
rect 16916 66928 16917 66968
rect 16875 66919 16917 66928
rect 16876 66834 16916 66919
rect 17067 66716 17109 66725
rect 16972 66676 17068 66716
rect 17108 66676 17109 66716
rect 16587 66380 16629 66389
rect 16587 66340 16588 66380
rect 16628 66340 16629 66380
rect 16587 66331 16629 66340
rect 16779 66380 16821 66389
rect 16779 66340 16780 66380
rect 16820 66340 16821 66380
rect 16779 66331 16821 66340
rect 16492 66079 16532 66088
rect 16587 66128 16629 66137
rect 16587 66088 16588 66128
rect 16628 66088 16629 66128
rect 16587 66079 16629 66088
rect 16780 66128 16820 66331
rect 16875 66212 16917 66221
rect 16875 66172 16876 66212
rect 16916 66172 16917 66212
rect 16875 66163 16917 66172
rect 16780 66079 16820 66088
rect 16588 65994 16628 66079
rect 16876 66078 16916 66163
rect 16972 66128 17012 66676
rect 17067 66667 17109 66676
rect 17068 66582 17108 66667
rect 16972 66079 17012 66088
rect 16683 66044 16725 66053
rect 16683 66004 16684 66044
rect 16724 66004 16725 66044
rect 16683 65995 16725 66004
rect 16300 65920 16436 65960
rect 16204 65836 16340 65876
rect 15819 65708 15861 65717
rect 15819 65668 15820 65708
rect 15860 65668 15861 65708
rect 15819 65659 15861 65668
rect 15723 65456 15765 65465
rect 15723 65416 15724 65456
rect 15764 65416 15765 65456
rect 15723 65407 15765 65416
rect 15724 65322 15764 65407
rect 15820 65288 15860 65659
rect 15916 65540 15956 65549
rect 15956 65500 16244 65540
rect 15916 65491 15956 65500
rect 16204 65456 16244 65500
rect 16204 65407 16244 65416
rect 16300 65456 16340 65836
rect 15820 65248 16148 65288
rect 15628 65164 15860 65204
rect 15724 64616 15764 64625
rect 15628 64576 15724 64616
rect 15531 64448 15573 64457
rect 15531 64408 15532 64448
rect 15572 64408 15573 64448
rect 15531 64399 15573 64408
rect 15532 64314 15572 64399
rect 15148 64240 15284 64280
rect 15340 64240 15476 64280
rect 14860 64072 15092 64112
rect 14860 63944 14900 63953
rect 14860 63785 14900 63904
rect 14859 63776 14901 63785
rect 14859 63736 14860 63776
rect 14900 63736 14901 63776
rect 14859 63727 14901 63736
rect 14860 63356 14900 63365
rect 14764 63316 14860 63356
rect 14668 63307 14708 63316
rect 14860 63307 14900 63316
rect 15052 63104 15092 64072
rect 15052 63055 15092 63064
rect 14668 62936 14708 62945
rect 14860 62936 14900 62945
rect 14708 62896 14804 62936
rect 14668 62887 14708 62896
rect 14764 62768 14804 62896
rect 14900 62896 14996 62936
rect 14860 62887 14900 62896
rect 14764 62728 14900 62768
rect 14764 62432 14804 62441
rect 14284 62392 14764 62432
rect 14187 61172 14229 61181
rect 14187 61132 14188 61172
rect 14228 61132 14229 61172
rect 14187 61123 14229 61132
rect 14284 60920 14324 62392
rect 14764 62383 14804 62392
rect 14860 62432 14900 62728
rect 14860 62383 14900 62392
rect 14956 62432 14996 62896
rect 15051 62600 15093 62609
rect 15051 62560 15052 62600
rect 15092 62560 15093 62600
rect 15051 62551 15093 62560
rect 15052 62466 15092 62551
rect 14956 62383 14996 62392
rect 14667 62264 14709 62273
rect 14667 62224 14668 62264
rect 14708 62224 14709 62264
rect 14667 62215 14709 62224
rect 15051 62264 15093 62273
rect 15051 62224 15052 62264
rect 15092 62224 15093 62264
rect 15051 62215 15093 62224
rect 14380 61592 14420 61601
rect 14380 61517 14420 61552
rect 14572 61592 14612 61601
rect 14379 61508 14421 61517
rect 14379 61468 14380 61508
rect 14420 61468 14421 61508
rect 14379 61459 14421 61468
rect 14380 61097 14420 61459
rect 14476 61424 14516 61433
rect 14379 61088 14421 61097
rect 14379 61048 14380 61088
rect 14420 61048 14421 61088
rect 14379 61039 14421 61048
rect 14476 61013 14516 61384
rect 14572 61097 14612 61552
rect 14668 61592 14708 62215
rect 14955 61676 14997 61685
rect 14955 61636 14956 61676
rect 14996 61636 14997 61676
rect 14955 61627 14997 61636
rect 14764 61592 14804 61601
rect 14668 61552 14764 61592
rect 14571 61088 14613 61097
rect 14571 61048 14572 61088
rect 14612 61048 14613 61088
rect 14571 61039 14613 61048
rect 14475 61004 14517 61013
rect 14475 60964 14476 61004
rect 14516 60964 14517 61004
rect 14475 60955 14517 60964
rect 14380 60920 14420 60929
rect 14284 60880 14380 60920
rect 14380 60871 14420 60880
rect 14571 60920 14613 60929
rect 14571 60880 14572 60920
rect 14612 60880 14613 60920
rect 14571 60871 14613 60880
rect 14476 60836 14516 60845
rect 14092 60796 14324 60836
rect 14284 60752 14324 60796
rect 14476 60752 14516 60796
rect 14284 60712 14516 60752
rect 14379 60500 14421 60509
rect 14379 60460 14380 60500
rect 14420 60460 14421 60500
rect 14379 60451 14421 60460
rect 14188 60332 14228 60341
rect 13900 60292 14188 60332
rect 14188 60283 14228 60292
rect 13804 60085 13844 60094
rect 14380 60089 14420 60451
rect 13804 59585 13844 60045
rect 14379 60080 14421 60089
rect 14379 60040 14380 60080
rect 14420 60040 14421 60080
rect 14379 60031 14421 60040
rect 13899 59996 13941 60005
rect 13899 59956 13900 59996
rect 13940 59956 13941 59996
rect 13899 59947 13941 59956
rect 13803 59576 13845 59585
rect 13803 59536 13804 59576
rect 13844 59536 13845 59576
rect 13803 59527 13845 59536
rect 13803 58400 13845 58409
rect 13803 58360 13804 58400
rect 13844 58360 13845 58400
rect 13803 58351 13845 58360
rect 13804 58266 13844 58351
rect 13803 57728 13845 57737
rect 13803 57688 13804 57728
rect 13844 57688 13845 57728
rect 13803 57679 13845 57688
rect 13804 57056 13844 57679
rect 13900 57233 13940 59947
rect 14380 59946 14420 60031
rect 13996 59912 14036 59921
rect 13899 57224 13941 57233
rect 13899 57184 13900 57224
rect 13940 57184 13941 57224
rect 13899 57175 13941 57184
rect 13804 57007 13844 57016
rect 13900 57056 13940 57065
rect 13900 56981 13940 57016
rect 13899 56972 13941 56981
rect 13899 56932 13900 56972
rect 13940 56932 13941 56972
rect 13899 56923 13941 56932
rect 13803 56720 13845 56729
rect 13803 56680 13804 56720
rect 13844 56680 13845 56720
rect 13803 56671 13845 56680
rect 13707 55376 13749 55385
rect 13707 55336 13708 55376
rect 13748 55336 13749 55376
rect 13707 55327 13749 55336
rect 13707 55124 13749 55133
rect 13707 55084 13708 55124
rect 13748 55084 13749 55124
rect 13707 55075 13749 55084
rect 13516 55000 13652 55040
rect 13612 54872 13652 55000
rect 13515 54788 13557 54797
rect 13515 54748 13516 54788
rect 13556 54748 13557 54788
rect 13515 54739 13557 54748
rect 13419 54368 13461 54377
rect 13419 54328 13420 54368
rect 13460 54328 13461 54368
rect 13419 54319 13461 54328
rect 13419 54032 13461 54041
rect 13419 53992 13420 54032
rect 13460 53992 13461 54032
rect 13419 53983 13461 53992
rect 13323 51932 13365 51941
rect 13323 51892 13324 51932
rect 13364 51892 13365 51932
rect 13323 51883 13365 51892
rect 13131 51848 13173 51857
rect 13131 51808 13132 51848
rect 13172 51808 13173 51848
rect 13131 51799 13173 51808
rect 13132 51714 13172 51799
rect 13324 51596 13364 51605
rect 13228 51556 13324 51596
rect 13228 51008 13268 51556
rect 13324 51547 13364 51556
rect 13228 50959 13268 50968
rect 13323 51008 13365 51017
rect 13323 50968 13324 51008
rect 13364 50968 13365 51008
rect 13323 50959 13365 50968
rect 13227 50504 13269 50513
rect 13227 50464 13228 50504
rect 13268 50464 13269 50504
rect 13227 50455 13269 50464
rect 13228 50168 13268 50455
rect 13228 50119 13268 50128
rect 13036 50084 13076 50093
rect 13076 50044 13172 50084
rect 13036 50035 13076 50044
rect 13132 49510 13172 50044
rect 13324 50000 13364 50959
rect 13420 50420 13460 53983
rect 13516 52277 13556 54739
rect 13612 53957 13652 54832
rect 13611 53948 13653 53957
rect 13611 53908 13612 53948
rect 13652 53908 13653 53948
rect 13611 53899 13653 53908
rect 13708 52772 13748 55075
rect 13804 54041 13844 56671
rect 13803 54032 13845 54041
rect 13803 53992 13804 54032
rect 13844 53992 13845 54032
rect 13803 53983 13845 53992
rect 13804 53898 13844 53983
rect 13612 52732 13748 52772
rect 13515 52268 13557 52277
rect 13515 52228 13516 52268
rect 13556 52228 13557 52268
rect 13515 52219 13557 52228
rect 13612 52100 13652 52732
rect 13803 52688 13845 52697
rect 13803 52648 13804 52688
rect 13844 52648 13845 52688
rect 13803 52639 13845 52648
rect 13719 52520 13759 52528
rect 13804 52520 13844 52639
rect 13719 52519 13844 52520
rect 13759 52480 13844 52519
rect 13719 52470 13759 52479
rect 13803 52352 13845 52361
rect 13803 52312 13804 52352
rect 13844 52312 13845 52352
rect 13803 52303 13845 52312
rect 13707 52268 13749 52277
rect 13707 52228 13708 52268
rect 13748 52228 13749 52268
rect 13707 52219 13749 52228
rect 13516 52060 13652 52100
rect 13516 51848 13556 52060
rect 13611 51932 13653 51941
rect 13611 51892 13612 51932
rect 13652 51892 13653 51932
rect 13611 51883 13653 51892
rect 13516 51799 13556 51808
rect 13420 50380 13556 50420
rect 12939 49496 12981 49505
rect 12939 49456 12940 49496
rect 12980 49456 12981 49496
rect 13132 49461 13172 49470
rect 13228 49960 13364 50000
rect 13420 50252 13460 50261
rect 12939 49447 12981 49456
rect 12843 49412 12885 49421
rect 12843 49372 12844 49412
rect 12884 49372 12885 49412
rect 12843 49363 12885 49372
rect 12843 49244 12885 49253
rect 12843 49204 12844 49244
rect 12884 49204 12885 49244
rect 13228 49244 13268 49960
rect 13420 49832 13460 50212
rect 13324 49792 13460 49832
rect 13324 49412 13364 49792
rect 13516 49673 13556 50380
rect 13515 49664 13557 49673
rect 13515 49624 13516 49664
rect 13556 49624 13557 49664
rect 13515 49615 13557 49624
rect 13515 49496 13557 49505
rect 13515 49456 13516 49496
rect 13556 49456 13557 49496
rect 13515 49447 13557 49456
rect 13324 49363 13364 49372
rect 13516 49362 13556 49447
rect 13228 49204 13364 49244
rect 12843 49195 12885 49204
rect 12748 48656 12788 48784
rect 12844 48740 12884 49195
rect 12940 48908 12980 48917
rect 12980 48868 13268 48908
rect 12940 48859 12980 48868
rect 13228 48824 13268 48868
rect 13228 48775 13268 48784
rect 13324 48824 13364 49204
rect 13515 49160 13557 49169
rect 13515 49120 13516 49160
rect 13556 49120 13557 49160
rect 13515 49111 13557 49120
rect 13131 48740 13173 48749
rect 12844 48700 12980 48740
rect 12748 48616 12884 48656
rect 12747 47312 12789 47321
rect 12747 47272 12748 47312
rect 12788 47272 12789 47312
rect 12747 47263 12789 47272
rect 12748 47178 12788 47263
rect 12556 47060 12596 47069
rect 12556 46472 12596 47020
rect 12556 46423 12596 46432
rect 12652 46472 12692 46481
rect 12652 46313 12692 46432
rect 12651 46304 12693 46313
rect 12651 46264 12652 46304
rect 12692 46264 12693 46304
rect 12651 46255 12693 46264
rect 12460 44584 12596 44624
rect 12459 44456 12501 44465
rect 12459 44416 12460 44456
rect 12500 44416 12501 44456
rect 12459 44407 12501 44416
rect 12268 44204 12308 44213
rect 12172 44164 12268 44204
rect 12172 43448 12212 44164
rect 12268 44155 12308 44164
rect 12268 43532 12308 43541
rect 12364 43532 12404 44248
rect 12308 43492 12404 43532
rect 12268 43483 12308 43492
rect 10252 42652 11060 42692
rect 10443 42104 10485 42113
rect 10443 42064 10444 42104
rect 10484 42064 10485 42104
rect 10443 42055 10485 42064
rect 10444 41936 10484 42055
rect 10828 41945 10868 42030
rect 10444 41887 10484 41896
rect 10827 41936 10869 41945
rect 10827 41896 10828 41936
rect 10868 41896 10869 41936
rect 10827 41887 10869 41896
rect 10059 41852 10101 41861
rect 10059 41812 10060 41852
rect 10100 41812 10101 41852
rect 10059 41803 10101 41812
rect 9963 40508 10005 40517
rect 9963 40468 9964 40508
rect 10004 40468 10005 40508
rect 9963 40459 10005 40468
rect 9867 40424 9909 40433
rect 9867 40384 9868 40424
rect 9908 40384 9909 40424
rect 9867 40375 9909 40384
rect 9868 40290 9908 40375
rect 9771 40172 9813 40181
rect 9771 40132 9772 40172
rect 9812 40132 9813 40172
rect 9771 40123 9813 40132
rect 9964 40097 10004 40459
rect 9963 40088 10005 40097
rect 9963 40048 9964 40088
rect 10004 40048 10005 40088
rect 9963 40039 10005 40048
rect 10060 40013 10100 41803
rect 10636 41768 10676 41777
rect 10676 41728 10868 41768
rect 10636 41719 10676 41728
rect 10539 41516 10581 41525
rect 10539 41476 10540 41516
rect 10580 41476 10581 41516
rect 10539 41467 10581 41476
rect 10443 41348 10485 41357
rect 10443 41308 10444 41348
rect 10484 41308 10485 41348
rect 10443 41299 10485 41308
rect 10444 41264 10484 41299
rect 10444 41213 10484 41224
rect 10540 41264 10580 41467
rect 10540 41215 10580 41224
rect 10828 40928 10868 41728
rect 11020 41264 11060 42652
rect 11115 42104 11157 42113
rect 11115 42064 11116 42104
rect 11156 42064 11157 42104
rect 11115 42055 11157 42064
rect 11116 41945 11156 42055
rect 11115 41936 11157 41945
rect 11115 41896 11116 41936
rect 11156 41896 11157 41936
rect 11115 41887 11157 41896
rect 11595 41516 11637 41525
rect 11595 41476 11596 41516
rect 11636 41476 11637 41516
rect 11595 41467 11637 41476
rect 10923 41180 10965 41189
rect 10923 41140 10924 41180
rect 10964 41140 10965 41180
rect 10923 41131 10965 41140
rect 10924 41046 10964 41131
rect 10828 40888 10964 40928
rect 10635 40760 10677 40769
rect 10635 40720 10636 40760
rect 10676 40720 10677 40760
rect 10635 40711 10677 40720
rect 10636 40433 10676 40711
rect 10924 40438 10964 40888
rect 10443 40424 10485 40433
rect 10443 40384 10444 40424
rect 10484 40384 10485 40424
rect 10443 40375 10485 40384
rect 10635 40424 10677 40433
rect 10635 40384 10636 40424
rect 10676 40384 10677 40424
rect 10924 40389 10964 40398
rect 10635 40375 10677 40384
rect 10444 40290 10484 40375
rect 11020 40265 11060 41224
rect 11499 41264 11541 41273
rect 11499 41224 11500 41264
rect 11540 41224 11541 41264
rect 11499 41215 11541 41224
rect 11500 41130 11540 41215
rect 11499 40508 11541 40517
rect 11499 40468 11500 40508
rect 11540 40468 11541 40508
rect 11499 40459 11541 40468
rect 11019 40256 11061 40265
rect 11019 40216 11020 40256
rect 11060 40216 11061 40256
rect 11019 40207 11061 40216
rect 11116 40256 11156 40265
rect 10059 40004 10101 40013
rect 10059 39964 10060 40004
rect 10100 39964 10101 40004
rect 10059 39955 10101 39964
rect 9484 39796 9620 39836
rect 9291 39584 9333 39593
rect 9291 39544 9292 39584
rect 9332 39544 9333 39584
rect 9291 39535 9333 39544
rect 9292 39450 9332 39535
rect 9196 39292 9332 39332
rect 9099 39080 9141 39089
rect 9099 39040 9100 39080
rect 9140 39040 9141 39080
rect 9099 39031 9141 39040
rect 9195 38996 9237 39005
rect 9195 38956 9196 38996
rect 9236 38956 9237 38996
rect 9195 38947 9237 38956
rect 9100 38912 9140 38921
rect 9004 38872 9100 38912
rect 8811 38576 8853 38585
rect 8811 38536 8812 38576
rect 8852 38536 8853 38576
rect 8811 38527 8853 38536
rect 9004 38408 9044 38872
rect 9100 38863 9140 38872
rect 8660 38200 8756 38240
rect 8812 38368 9044 38408
rect 8524 38106 8564 38191
rect 7756 35848 7852 35888
rect 7756 35561 7796 35848
rect 7852 35839 7892 35848
rect 7948 35932 8276 35972
rect 7948 35720 7988 35932
rect 8332 35888 8372 35897
rect 8044 35804 8084 35813
rect 8332 35804 8372 35848
rect 8084 35764 8372 35804
rect 8428 35888 8468 35897
rect 8620 35888 8660 38200
rect 8715 36896 8757 36905
rect 8715 36856 8716 36896
rect 8756 36856 8757 36896
rect 8715 36847 8757 36856
rect 8716 36728 8756 36847
rect 8716 36679 8756 36688
rect 8715 36560 8757 36569
rect 8715 36520 8716 36560
rect 8756 36520 8757 36560
rect 8715 36511 8757 36520
rect 8468 35848 8660 35888
rect 8044 35755 8084 35764
rect 7852 35680 7988 35720
rect 7755 35552 7797 35561
rect 7755 35512 7756 35552
rect 7796 35512 7797 35552
rect 7755 35503 7797 35512
rect 7755 34376 7797 34385
rect 7755 34336 7756 34376
rect 7796 34336 7797 34376
rect 7755 34327 7797 34336
rect 7756 34242 7796 34327
rect 7755 34040 7797 34049
rect 7755 34000 7756 34040
rect 7796 34000 7797 34040
rect 7755 33991 7797 34000
rect 7756 33872 7796 33991
rect 7756 33823 7796 33832
rect 7659 32948 7701 32957
rect 7659 32908 7660 32948
rect 7700 32908 7701 32948
rect 7659 32899 7701 32908
rect 7372 32864 7412 32873
rect 7276 32824 7372 32864
rect 7276 31445 7316 32824
rect 7372 32815 7412 32824
rect 7756 32864 7796 32873
rect 7756 32705 7796 32824
rect 7563 32696 7605 32705
rect 7563 32656 7564 32696
rect 7604 32656 7605 32696
rect 7563 32647 7605 32656
rect 7755 32696 7797 32705
rect 7755 32656 7756 32696
rect 7796 32656 7797 32696
rect 7755 32647 7797 32656
rect 7564 32562 7604 32647
rect 7852 32621 7892 35680
rect 8139 35552 8181 35561
rect 8139 35512 8140 35552
rect 8180 35512 8181 35552
rect 8139 35503 8181 35512
rect 8043 35384 8085 35393
rect 8043 35344 8044 35384
rect 8084 35344 8085 35384
rect 8043 35335 8085 35344
rect 7947 34712 7989 34721
rect 7947 34672 7948 34712
rect 7988 34672 7989 34712
rect 7947 34663 7989 34672
rect 7948 34628 7988 34663
rect 7948 34577 7988 34588
rect 7948 34376 7988 34387
rect 7948 34301 7988 34336
rect 7947 34292 7989 34301
rect 7947 34252 7948 34292
rect 7988 34252 7989 34292
rect 7947 34243 7989 34252
rect 7947 33200 7989 33209
rect 7947 33160 7948 33200
rect 7988 33160 7989 33200
rect 7947 33151 7989 33160
rect 7948 33032 7988 33151
rect 8044 33116 8084 35335
rect 8140 35216 8180 35503
rect 8180 35176 8276 35216
rect 8140 35167 8180 35176
rect 8139 34376 8181 34385
rect 8139 34336 8140 34376
rect 8180 34336 8181 34376
rect 8139 34327 8181 34336
rect 8140 34242 8180 34327
rect 8236 33713 8276 35176
rect 8332 34964 8372 34973
rect 8332 34376 8372 34924
rect 8428 34544 8468 35848
rect 8524 35216 8564 35225
rect 8716 35216 8756 36511
rect 8564 35176 8756 35216
rect 8812 35888 8852 38368
rect 8907 38240 8949 38249
rect 8907 38200 8908 38240
rect 8948 38200 8949 38240
rect 8907 38191 8949 38200
rect 9004 38240 9044 38368
rect 9004 38191 9044 38200
rect 9100 38240 9140 38249
rect 9196 38240 9236 38947
rect 9140 38200 9236 38240
rect 8908 36896 8948 38191
rect 9004 37400 9044 37409
rect 9004 37241 9044 37360
rect 9003 37232 9045 37241
rect 9003 37192 9004 37232
rect 9044 37192 9045 37232
rect 9003 37183 9045 37192
rect 8908 36847 8948 36856
rect 8524 35167 8564 35176
rect 8428 34504 8564 34544
rect 8524 34385 8564 34504
rect 8428 34376 8468 34385
rect 8332 34336 8428 34376
rect 8428 34327 8468 34336
rect 8523 34376 8565 34385
rect 8523 34336 8524 34376
rect 8564 34336 8565 34376
rect 8523 34327 8565 34336
rect 8524 34242 8564 34327
rect 8331 33956 8373 33965
rect 8331 33916 8332 33956
rect 8372 33916 8373 33956
rect 8331 33907 8373 33916
rect 8235 33704 8277 33713
rect 8235 33664 8236 33704
rect 8276 33664 8277 33704
rect 8235 33655 8277 33664
rect 8332 33704 8372 33907
rect 8332 33655 8372 33664
rect 8331 33200 8373 33209
rect 8331 33160 8332 33200
rect 8372 33160 8373 33200
rect 8331 33151 8373 33160
rect 8044 33076 8180 33116
rect 7948 32983 7988 32992
rect 8043 32948 8085 32957
rect 8043 32908 8044 32948
rect 8084 32908 8085 32948
rect 8043 32899 8085 32908
rect 7948 32860 7988 32869
rect 7948 32789 7988 32820
rect 8044 32864 8084 32899
rect 8044 32813 8084 32824
rect 7948 32780 7990 32789
rect 7948 32740 7949 32780
rect 7989 32740 7990 32780
rect 7948 32731 7990 32740
rect 7949 32726 7989 32731
rect 7851 32612 7893 32621
rect 7851 32572 7852 32612
rect 7892 32572 7893 32612
rect 7851 32563 7893 32572
rect 7755 32528 7797 32537
rect 7755 32488 7756 32528
rect 7796 32488 7797 32528
rect 7755 32479 7797 32488
rect 7563 32276 7605 32285
rect 7563 32236 7564 32276
rect 7604 32236 7605 32276
rect 7563 32227 7605 32236
rect 7372 32178 7412 32187
rect 7564 32142 7604 32227
rect 7659 32192 7701 32201
rect 7659 32152 7660 32192
rect 7700 32152 7701 32192
rect 7659 32143 7701 32152
rect 7372 32033 7412 32138
rect 7371 32024 7413 32033
rect 7371 31984 7372 32024
rect 7412 31984 7413 32024
rect 7371 31975 7413 31984
rect 7275 31436 7317 31445
rect 7275 31396 7276 31436
rect 7316 31396 7317 31436
rect 7275 31387 7317 31396
rect 7275 31184 7317 31193
rect 7275 31144 7276 31184
rect 7316 31144 7317 31184
rect 7275 31135 7317 31144
rect 7124 29800 7220 29840
rect 6892 29119 6932 29128
rect 6987 29168 7029 29177
rect 6987 29128 6988 29168
rect 7028 29128 7029 29168
rect 6987 29119 7029 29128
rect 6988 29034 7028 29119
rect 6411 29000 6453 29009
rect 6411 28960 6412 29000
rect 6452 28960 6453 29000
rect 6411 28951 6453 28960
rect 6603 29000 6645 29009
rect 6603 28960 6604 29000
rect 6644 28960 6645 29000
rect 6603 28951 6645 28960
rect 6411 28748 6453 28757
rect 6411 28708 6412 28748
rect 6452 28708 6453 28748
rect 6411 28699 6453 28708
rect 6412 28412 6452 28699
rect 6315 28328 6357 28337
rect 6315 28288 6316 28328
rect 6356 28288 6357 28328
rect 6315 28279 6357 28288
rect 6316 28194 6356 28279
rect 6315 28076 6357 28085
rect 6315 28036 6316 28076
rect 6356 28036 6357 28076
rect 6315 28027 6357 28036
rect 6220 26816 6260 26827
rect 6220 26741 6260 26776
rect 6316 26816 6356 28027
rect 6412 26909 6452 28372
rect 6604 28328 6644 28951
rect 6891 28496 6933 28505
rect 6891 28456 6892 28496
rect 6932 28456 6933 28496
rect 6891 28447 6933 28456
rect 6508 28288 6644 28328
rect 6699 28328 6741 28337
rect 6699 28288 6700 28328
rect 6740 28288 6741 28328
rect 6411 26900 6453 26909
rect 6411 26860 6412 26900
rect 6452 26860 6453 26900
rect 6411 26851 6453 26860
rect 6219 26732 6261 26741
rect 6219 26692 6220 26732
rect 6260 26692 6261 26732
rect 6219 26683 6261 26692
rect 6124 26440 6260 26480
rect 6124 26144 6164 26153
rect 6028 26104 6124 26144
rect 6028 25901 6068 26104
rect 6124 26095 6164 26104
rect 6027 25892 6069 25901
rect 6027 25852 6028 25892
rect 6068 25852 6069 25892
rect 6027 25843 6069 25852
rect 5835 25556 5877 25565
rect 5835 25516 5836 25556
rect 5876 25516 5877 25556
rect 5835 25507 5877 25516
rect 6220 25472 6260 26440
rect 6028 25432 6260 25472
rect 5835 25388 5877 25397
rect 5835 25348 5836 25388
rect 5876 25348 5877 25388
rect 5835 25339 5877 25348
rect 5836 25304 5876 25339
rect 5836 25253 5876 25264
rect 5932 25304 5972 25313
rect 5739 24968 5781 24977
rect 5739 24928 5740 24968
rect 5780 24928 5781 24968
rect 5739 24919 5781 24928
rect 5932 24557 5972 25264
rect 5931 24548 5973 24557
rect 5931 24508 5932 24548
rect 5972 24508 5973 24548
rect 5931 24499 5973 24508
rect 5643 24212 5685 24221
rect 5643 24172 5644 24212
rect 5684 24172 5685 24212
rect 5643 24163 5685 24172
rect 5644 23120 5684 24163
rect 6028 24137 6068 25432
rect 6220 25304 6260 25313
rect 6220 24800 6260 25264
rect 6316 25304 6356 26776
rect 6316 25061 6356 25264
rect 6411 25304 6453 25313
rect 6411 25264 6412 25304
rect 6452 25264 6453 25304
rect 6411 25255 6453 25264
rect 6315 25052 6357 25061
rect 6315 25012 6316 25052
rect 6356 25012 6357 25052
rect 6315 25003 6357 25012
rect 6316 24800 6356 24809
rect 6220 24760 6316 24800
rect 6316 24751 6356 24760
rect 6124 24632 6164 24641
rect 6124 24473 6164 24592
rect 6123 24464 6165 24473
rect 6123 24424 6124 24464
rect 6164 24424 6165 24464
rect 6123 24415 6165 24424
rect 6219 24380 6261 24389
rect 6219 24340 6220 24380
rect 6260 24340 6261 24380
rect 6219 24331 6261 24340
rect 6027 24128 6069 24137
rect 6027 24088 6028 24128
rect 6068 24088 6069 24128
rect 6027 24079 6069 24088
rect 5835 23876 5877 23885
rect 5835 23836 5836 23876
rect 5876 23836 5877 23876
rect 5835 23827 5877 23836
rect 5739 23792 5781 23801
rect 5739 23752 5740 23792
rect 5780 23752 5781 23792
rect 5739 23743 5781 23752
rect 5836 23792 5876 23827
rect 5740 23658 5780 23743
rect 5836 23741 5876 23752
rect 5644 23071 5684 23080
rect 6028 23045 6068 24079
rect 6220 23876 6260 24331
rect 6220 23827 6260 23836
rect 6315 23876 6357 23885
rect 6315 23836 6316 23876
rect 6356 23836 6357 23876
rect 6315 23827 6357 23836
rect 6316 23742 6356 23827
rect 6123 23708 6165 23717
rect 6123 23668 6124 23708
rect 6164 23668 6165 23708
rect 6123 23659 6165 23668
rect 6027 23036 6069 23045
rect 6027 22996 6028 23036
rect 6068 22996 6069 23036
rect 6027 22987 6069 22996
rect 6124 22448 6164 23659
rect 6412 23624 6452 25255
rect 6124 22399 6164 22408
rect 6316 23584 6452 23624
rect 5739 22280 5781 22289
rect 5739 22240 5740 22280
rect 5780 22240 5781 22280
rect 5739 22231 5781 22240
rect 6123 22280 6165 22289
rect 6123 22240 6124 22280
rect 6164 22240 6165 22280
rect 6123 22231 6165 22240
rect 6220 22280 6260 22291
rect 5740 22146 5780 22231
rect 6124 22146 6164 22231
rect 6220 22205 6260 22240
rect 6219 22196 6261 22205
rect 6219 22156 6220 22196
rect 6260 22156 6261 22196
rect 6219 22147 6261 22156
rect 5932 22112 5972 22121
rect 6316 22112 6356 23584
rect 6411 22364 6453 22373
rect 6411 22324 6412 22364
rect 6452 22324 6453 22364
rect 6411 22315 6453 22324
rect 6412 22280 6452 22315
rect 6412 22229 6452 22240
rect 6508 22112 6548 28288
rect 6699 28279 6741 28288
rect 6892 28328 6932 28447
rect 7084 28412 7124 29800
rect 6700 26816 6740 28279
rect 6795 28160 6837 28169
rect 6795 28120 6796 28160
rect 6836 28120 6837 28160
rect 6795 28111 6837 28120
rect 6796 27329 6836 28111
rect 6795 27320 6837 27329
rect 6795 27280 6796 27320
rect 6836 27280 6837 27320
rect 6795 27271 6837 27280
rect 6795 26900 6837 26909
rect 6795 26860 6796 26900
rect 6836 26860 6837 26900
rect 6795 26851 6837 26860
rect 6603 25724 6645 25733
rect 6603 25684 6604 25724
rect 6644 25684 6645 25724
rect 6603 25675 6645 25684
rect 6604 23885 6644 25675
rect 6700 25313 6740 26776
rect 6699 25304 6741 25313
rect 6699 25264 6700 25304
rect 6740 25264 6741 25304
rect 6699 25255 6741 25264
rect 6796 25304 6836 26851
rect 6892 26825 6932 28288
rect 6988 28372 7124 28412
rect 6891 26816 6933 26825
rect 6891 26776 6892 26816
rect 6932 26776 6933 26816
rect 6891 26767 6933 26776
rect 6988 25388 7028 28372
rect 7083 28244 7125 28253
rect 7083 28204 7084 28244
rect 7124 28204 7125 28244
rect 7083 28195 7125 28204
rect 7084 27656 7124 28195
rect 7180 27656 7220 27665
rect 7084 27616 7180 27656
rect 7084 26153 7124 27616
rect 7180 27607 7220 27616
rect 7276 27488 7316 31135
rect 7371 29168 7413 29177
rect 7371 29128 7372 29168
rect 7412 29128 7413 29168
rect 7371 29119 7413 29128
rect 7372 29034 7412 29119
rect 7468 29084 7508 29093
rect 7372 28333 7412 28342
rect 7372 27824 7412 28293
rect 7372 27775 7412 27784
rect 7468 28160 7508 29044
rect 7564 28160 7604 28169
rect 7468 28120 7564 28160
rect 7180 27448 7316 27488
rect 7083 26144 7125 26153
rect 7083 26104 7084 26144
rect 7124 26104 7125 26144
rect 7083 26095 7125 26104
rect 6988 25348 7124 25388
rect 6700 25170 6740 25255
rect 6796 25229 6836 25264
rect 6795 25220 6837 25229
rect 6795 25180 6796 25220
rect 6836 25180 6837 25220
rect 6795 25171 6837 25180
rect 6987 25220 7029 25229
rect 6987 25180 6988 25220
rect 7028 25180 7029 25220
rect 6987 25171 7029 25180
rect 6891 25052 6933 25061
rect 6891 25012 6892 25052
rect 6932 25012 6933 25052
rect 6891 25003 6933 25012
rect 6700 24632 6740 24641
rect 6603 23876 6645 23885
rect 6603 23836 6604 23876
rect 6644 23836 6645 23876
rect 6603 23827 6645 23836
rect 6700 23801 6740 24592
rect 6699 23792 6741 23801
rect 6699 23752 6700 23792
rect 6740 23752 6741 23792
rect 6699 23743 6741 23752
rect 6796 23792 6836 23801
rect 6603 22868 6645 22877
rect 6603 22828 6604 22868
rect 6644 22828 6645 22868
rect 6603 22819 6645 22828
rect 6604 22280 6644 22819
rect 6796 22289 6836 23752
rect 6892 23288 6932 25003
rect 6988 24809 7028 25171
rect 7084 24809 7124 25348
rect 6982 24800 7028 24809
rect 6982 24760 6983 24800
rect 7023 24760 7028 24800
rect 6982 24751 7028 24760
rect 7083 24800 7125 24809
rect 7083 24760 7084 24800
rect 7124 24760 7125 24800
rect 7083 24751 7125 24760
rect 6988 24632 7028 24751
rect 6988 24583 7028 24592
rect 7084 24632 7124 24641
rect 7084 24389 7124 24592
rect 7083 24380 7125 24389
rect 7083 24340 7084 24380
rect 7124 24340 7125 24380
rect 7083 24331 7125 24340
rect 7180 24305 7220 27448
rect 7275 26816 7317 26825
rect 7275 26776 7276 26816
rect 7316 26776 7317 26816
rect 7275 26767 7317 26776
rect 7276 25313 7316 26767
rect 7468 26321 7508 28120
rect 7564 28111 7604 28120
rect 7563 27992 7605 28001
rect 7563 27952 7564 27992
rect 7604 27952 7605 27992
rect 7563 27943 7605 27952
rect 7467 26312 7509 26321
rect 7467 26272 7468 26312
rect 7508 26272 7509 26312
rect 7467 26263 7509 26272
rect 7371 26144 7413 26153
rect 7564 26144 7604 27943
rect 7371 26104 7372 26144
rect 7412 26104 7413 26144
rect 7371 26095 7413 26104
rect 7468 26104 7604 26144
rect 7372 26010 7412 26095
rect 7275 25304 7317 25313
rect 7275 25264 7276 25304
rect 7316 25264 7317 25304
rect 7275 25255 7317 25264
rect 7276 25170 7316 25255
rect 7371 24464 7413 24473
rect 7371 24424 7372 24464
rect 7412 24424 7413 24464
rect 7371 24415 7413 24424
rect 7372 24330 7412 24415
rect 7179 24296 7221 24305
rect 7179 24256 7180 24296
rect 7220 24256 7221 24296
rect 7179 24247 7221 24256
rect 7468 24212 7508 26104
rect 7564 25901 7604 25986
rect 7563 25892 7605 25901
rect 7563 25852 7564 25892
rect 7604 25852 7605 25892
rect 7563 25843 7605 25852
rect 7660 25724 7700 32143
rect 7756 27077 7796 32479
rect 8140 32444 8180 33076
rect 8236 32857 8276 32866
rect 8236 32453 8276 32817
rect 7948 32404 8180 32444
rect 8235 32444 8277 32453
rect 8235 32404 8236 32444
rect 8276 32404 8277 32444
rect 8332 32444 8372 33151
rect 8523 33116 8565 33125
rect 8523 33076 8524 33116
rect 8564 33076 8565 33116
rect 8523 33067 8565 33076
rect 8427 32948 8469 32957
rect 8427 32908 8428 32948
rect 8468 32908 8469 32948
rect 8427 32899 8469 32908
rect 8428 32814 8468 32899
rect 8524 32864 8564 33067
rect 8524 32815 8564 32824
rect 8332 32404 8468 32444
rect 7851 32192 7893 32201
rect 7851 32152 7852 32192
rect 7892 32152 7893 32192
rect 7851 32143 7893 32152
rect 7852 28253 7892 32143
rect 7948 31520 7988 32404
rect 8235 32395 8277 32404
rect 8331 32276 8373 32285
rect 8331 32236 8332 32276
rect 8372 32236 8373 32276
rect 8331 32227 8373 32236
rect 8428 32276 8468 32404
rect 8428 32227 8468 32236
rect 8044 32192 8084 32201
rect 8044 31604 8084 32152
rect 8332 32192 8372 32227
rect 8332 32141 8372 32152
rect 8620 32108 8660 35176
rect 8812 34376 8852 35848
rect 8908 35888 8948 35897
rect 9100 35888 9140 38200
rect 9292 38156 9332 39292
rect 8948 35848 9140 35888
rect 9196 38116 9332 38156
rect 8908 35839 8948 35848
rect 9004 34385 9044 35848
rect 8908 34376 8948 34385
rect 8812 34336 8908 34376
rect 8811 34124 8853 34133
rect 8811 34084 8812 34124
rect 8852 34084 8853 34124
rect 8811 34075 8853 34084
rect 8715 33704 8757 33713
rect 8715 33664 8716 33704
rect 8756 33664 8757 33704
rect 8715 33655 8757 33664
rect 8716 32201 8756 33655
rect 8715 32192 8757 32201
rect 8715 32152 8716 32192
rect 8756 32152 8757 32192
rect 8715 32143 8757 32152
rect 8428 32068 8660 32108
rect 8332 31604 8372 31613
rect 8044 31564 8332 31604
rect 8332 31555 8372 31564
rect 7948 31480 8084 31520
rect 8044 31193 8084 31480
rect 8140 31445 8180 31476
rect 8139 31436 8181 31445
rect 8139 31396 8140 31436
rect 8180 31396 8181 31436
rect 8139 31387 8181 31396
rect 8331 31436 8373 31445
rect 8331 31396 8332 31436
rect 8372 31396 8373 31436
rect 8331 31387 8373 31396
rect 8140 31352 8180 31387
rect 8043 31184 8085 31193
rect 8043 31144 8044 31184
rect 8084 31144 8085 31184
rect 8043 31135 8085 31144
rect 7947 29336 7989 29345
rect 7947 29296 7948 29336
rect 7988 29296 7989 29336
rect 7947 29287 7989 29296
rect 7948 29168 7988 29287
rect 7851 28244 7893 28253
rect 7851 28204 7852 28244
rect 7892 28204 7893 28244
rect 7851 28195 7893 28204
rect 7755 27068 7797 27077
rect 7755 27028 7756 27068
rect 7796 27028 7797 27068
rect 7755 27019 7797 27028
rect 7948 26900 7988 29128
rect 8044 28328 8084 31135
rect 8044 28001 8084 28288
rect 8140 28169 8180 31312
rect 8235 31352 8277 31361
rect 8235 31312 8236 31352
rect 8276 31312 8277 31352
rect 8235 31303 8277 31312
rect 8139 28160 8181 28169
rect 8139 28120 8140 28160
rect 8180 28120 8181 28160
rect 8139 28111 8181 28120
rect 8043 27992 8085 28001
rect 8043 27952 8044 27992
rect 8084 27952 8085 27992
rect 8043 27943 8085 27952
rect 7947 26860 7988 26900
rect 7756 26821 7796 26830
rect 7756 26741 7796 26781
rect 7947 26741 7987 26860
rect 7755 26732 7797 26741
rect 7947 26732 7988 26741
rect 7755 26692 7756 26732
rect 7796 26692 7797 26732
rect 7755 26683 7797 26692
rect 7852 26692 7948 26732
rect 7755 26144 7797 26153
rect 7755 26104 7756 26144
rect 7796 26104 7797 26144
rect 7755 26095 7797 26104
rect 7756 26010 7796 26095
rect 7755 25892 7797 25901
rect 7755 25852 7756 25892
rect 7796 25852 7797 25892
rect 7755 25843 7797 25852
rect 7372 24172 7508 24212
rect 7564 25684 7700 25724
rect 7564 24632 7604 25684
rect 7659 25556 7701 25565
rect 7659 25516 7660 25556
rect 7700 25516 7701 25556
rect 7659 25507 7701 25516
rect 7275 23876 7317 23885
rect 7275 23836 7276 23876
rect 7316 23836 7317 23876
rect 7275 23827 7317 23836
rect 7276 23806 7316 23827
rect 7276 23741 7316 23766
rect 7083 23288 7125 23297
rect 6892 23248 7028 23288
rect 6892 23120 6932 23131
rect 6892 23045 6932 23080
rect 6891 23036 6933 23045
rect 6891 22996 6892 23036
rect 6932 22996 6933 23036
rect 6891 22987 6933 22996
rect 6988 22616 7028 23248
rect 7083 23248 7084 23288
rect 7124 23248 7125 23288
rect 7083 23239 7125 23248
rect 7084 23154 7124 23239
rect 7276 23120 7316 23129
rect 7372 23120 7412 24172
rect 7564 23969 7604 24592
rect 7563 23960 7605 23969
rect 7563 23920 7564 23960
rect 7604 23920 7605 23960
rect 7563 23911 7605 23920
rect 7467 23708 7509 23717
rect 7467 23668 7468 23708
rect 7508 23668 7509 23708
rect 7467 23659 7509 23668
rect 7468 23574 7508 23659
rect 7316 23080 7412 23120
rect 7083 22868 7125 22877
rect 7083 22828 7084 22868
rect 7124 22828 7125 22868
rect 7083 22819 7125 22828
rect 7084 22734 7124 22819
rect 6988 22576 7124 22616
rect 6604 22231 6644 22240
rect 6795 22280 6837 22289
rect 6795 22240 6796 22280
rect 6836 22240 6837 22280
rect 6795 22231 6837 22240
rect 6699 22196 6741 22205
rect 6699 22156 6700 22196
rect 6740 22156 6741 22196
rect 6699 22147 6741 22156
rect 6316 22072 6452 22112
rect 6508 22072 6644 22112
rect 5932 21869 5972 22072
rect 5547 21860 5589 21869
rect 5547 21820 5548 21860
rect 5588 21820 5589 21860
rect 5547 21811 5589 21820
rect 5931 21860 5973 21869
rect 5931 21820 5932 21860
rect 5972 21820 5973 21860
rect 5931 21811 5973 21820
rect 5932 21692 5972 21701
rect 5547 21608 5589 21617
rect 5547 21568 5548 21608
rect 5588 21568 5589 21608
rect 5547 21559 5589 21568
rect 5739 21608 5781 21617
rect 5739 21568 5740 21608
rect 5780 21568 5781 21608
rect 5739 21559 5781 21568
rect 5836 21608 5876 21617
rect 5356 21400 5492 21440
rect 5356 21197 5396 21400
rect 5355 21188 5397 21197
rect 5355 21148 5356 21188
rect 5396 21148 5397 21188
rect 5355 21139 5397 21148
rect 4876 21064 5204 21104
rect 4876 21020 4916 21064
rect 4876 20971 4916 20980
rect 5356 20945 5396 21139
rect 5548 21020 5588 21559
rect 5740 21474 5780 21559
rect 5452 20980 5588 21020
rect 5355 20936 5397 20945
rect 5355 20896 5356 20936
rect 5396 20896 5397 20936
rect 5355 20887 5397 20896
rect 5067 20852 5109 20861
rect 5067 20812 5068 20852
rect 5108 20812 5109 20852
rect 5067 20803 5109 20812
rect 5068 20768 5108 20803
rect 5068 20717 5108 20728
rect 5163 20768 5205 20777
rect 5163 20728 5164 20768
rect 5204 20728 5205 20768
rect 5163 20719 5205 20728
rect 5355 20768 5397 20777
rect 5355 20728 5356 20768
rect 5396 20728 5397 20768
rect 5355 20719 5397 20728
rect 5164 20634 5204 20719
rect 5356 20642 5396 20719
rect 5356 20593 5396 20602
rect 5452 20600 5492 20980
rect 5836 20777 5876 21568
rect 5932 21533 5972 21652
rect 6028 21608 6068 21617
rect 6220 21608 6260 21617
rect 5931 21524 5973 21533
rect 5931 21484 5932 21524
rect 5972 21484 5973 21524
rect 5931 21475 5973 21484
rect 6028 21449 6068 21568
rect 6124 21568 6220 21608
rect 6027 21440 6069 21449
rect 6027 21400 6028 21440
rect 6068 21400 6069 21440
rect 6027 21391 6069 21400
rect 6027 20936 6069 20945
rect 6027 20896 6028 20936
rect 6068 20896 6069 20936
rect 6027 20887 6069 20896
rect 5548 20768 5588 20777
rect 5835 20768 5877 20777
rect 5588 20728 5684 20768
rect 5548 20719 5588 20728
rect 5452 20560 5493 20600
rect 5453 20516 5493 20560
rect 5644 20525 5684 20728
rect 5835 20728 5836 20768
rect 5876 20728 5877 20768
rect 5835 20719 5877 20728
rect 5452 20476 5493 20516
rect 5643 20516 5685 20525
rect 5643 20476 5644 20516
rect 5684 20476 5685 20516
rect 4928 20432 5296 20441
rect 4968 20392 5010 20432
rect 5050 20392 5092 20432
rect 5132 20392 5174 20432
rect 5214 20392 5256 20432
rect 4928 20383 5296 20392
rect 5355 20432 5397 20441
rect 5355 20392 5356 20432
rect 5396 20392 5397 20432
rect 5355 20383 5397 20392
rect 5356 20264 5396 20383
rect 5164 20224 5396 20264
rect 4684 20140 4820 20180
rect 4875 20180 4917 20189
rect 4875 20140 4876 20180
rect 4916 20140 4917 20180
rect 4684 20096 4724 20140
rect 4875 20131 4917 20140
rect 5164 20180 5204 20224
rect 5164 20131 5204 20140
rect 4684 20047 4724 20056
rect 4683 19928 4725 19937
rect 4683 19888 4684 19928
rect 4724 19888 4725 19928
rect 4683 19879 4725 19888
rect 4876 19928 4916 20131
rect 5260 20096 5300 20105
rect 5260 20021 5300 20056
rect 5259 20012 5301 20021
rect 5259 19972 5260 20012
rect 5300 19972 5301 20012
rect 5259 19963 5301 19972
rect 4876 19879 4916 19888
rect 4396 19804 4628 19844
rect 3688 19676 4056 19685
rect 3728 19636 3770 19676
rect 3810 19636 3852 19676
rect 3892 19636 3934 19676
rect 3974 19636 4016 19676
rect 3688 19627 4056 19636
rect 4203 19340 4245 19349
rect 4203 19300 4204 19340
rect 4244 19300 4245 19340
rect 4203 19291 4245 19300
rect 4204 19256 4244 19291
rect 4204 19205 4244 19216
rect 4299 18584 4341 18593
rect 4299 18544 4300 18584
rect 4340 18544 4341 18584
rect 4299 18535 4341 18544
rect 4300 18450 4340 18535
rect 4107 18332 4149 18341
rect 4107 18292 4108 18332
rect 4148 18292 4149 18332
rect 4107 18283 4149 18292
rect 3531 18164 3573 18173
rect 3531 18124 3532 18164
rect 3572 18124 3573 18164
rect 3531 18115 3573 18124
rect 3688 18164 4056 18173
rect 3728 18124 3770 18164
rect 3810 18124 3852 18164
rect 3892 18124 3934 18164
rect 3974 18124 4016 18164
rect 3688 18115 4056 18124
rect 3532 17744 3572 18115
rect 3627 17996 3669 18005
rect 3627 17956 3628 17996
rect 3668 17956 3669 17996
rect 3627 17947 3669 17956
rect 3532 17695 3572 17704
rect 3628 17744 3668 17947
rect 4108 17828 4148 18283
rect 4108 17779 4148 17788
rect 3628 17695 3668 17704
rect 3723 17744 3765 17753
rect 3723 17704 3724 17744
rect 3764 17704 3765 17744
rect 3723 17695 3765 17704
rect 4012 17744 4052 17753
rect 3244 17023 3284 17032
rect 3340 17032 3345 17072
rect 3385 17032 3476 17072
rect 3724 17072 3764 17695
rect 3340 17023 3385 17032
rect 2860 16820 2900 16829
rect 2860 16409 2900 16780
rect 3340 16409 3380 17023
rect 3724 16829 3764 17032
rect 4012 16829 4052 17704
rect 3723 16820 3765 16829
rect 3723 16780 3724 16820
rect 3764 16780 3765 16820
rect 3723 16771 3765 16780
rect 4011 16820 4053 16829
rect 4011 16780 4012 16820
rect 4052 16780 4053 16820
rect 4011 16771 4053 16780
rect 4299 16820 4341 16829
rect 4299 16780 4300 16820
rect 4340 16780 4341 16820
rect 4299 16771 4341 16780
rect 3688 16652 4056 16661
rect 3728 16612 3770 16652
rect 3810 16612 3852 16652
rect 3892 16612 3934 16652
rect 3974 16612 4016 16652
rect 3688 16603 4056 16612
rect 4107 16484 4149 16493
rect 4107 16444 4108 16484
rect 4148 16444 4149 16484
rect 4107 16435 4149 16444
rect 2859 16400 2901 16409
rect 2859 16360 2860 16400
rect 2900 16360 2901 16400
rect 2859 16351 2901 16360
rect 3339 16400 3381 16409
rect 3339 16360 3340 16400
rect 3380 16360 3381 16400
rect 3339 16351 3381 16360
rect 3052 16303 3092 16312
rect 2476 15737 2516 16192
rect 2763 16232 2805 16241
rect 2763 16192 2764 16232
rect 2804 16192 2805 16232
rect 2763 16183 2805 16192
rect 2860 16064 2900 16073
rect 2475 15728 2517 15737
rect 2475 15688 2476 15728
rect 2516 15688 2517 15728
rect 2475 15679 2517 15688
rect 2763 15728 2805 15737
rect 2763 15688 2764 15728
rect 2804 15688 2805 15728
rect 2763 15679 2805 15688
rect 2380 15520 2612 15560
rect 1804 15436 1940 15476
rect 1804 14720 1844 15436
rect 1899 15308 1941 15317
rect 1899 15268 1900 15308
rect 1940 15268 1941 15308
rect 1899 15259 1941 15268
rect 1804 14671 1844 14680
rect 1612 14596 1748 14636
rect 1515 14300 1557 14309
rect 1515 14260 1516 14300
rect 1556 14260 1557 14300
rect 1515 14251 1557 14260
rect 1324 14167 1364 14176
rect 1516 13964 1556 14251
rect 1516 13915 1556 13924
rect 1227 13544 1269 13553
rect 1227 13504 1228 13544
rect 1268 13504 1269 13544
rect 1227 13495 1269 13504
rect 1612 13460 1652 14596
rect 1803 14216 1845 14225
rect 1803 14176 1804 14216
rect 1844 14176 1845 14216
rect 1803 14167 1845 14176
rect 1516 13420 1652 13460
rect 1708 13796 1748 13805
rect 1227 13292 1269 13301
rect 1227 13252 1228 13292
rect 1268 13252 1269 13292
rect 1227 13243 1269 13252
rect 1228 13208 1268 13243
rect 1228 13157 1268 13168
rect 1228 12536 1268 12545
rect 1323 12536 1365 12545
rect 1268 12496 1324 12536
rect 1364 12496 1365 12536
rect 1228 12487 1268 12496
rect 1323 12487 1365 12496
rect 1420 11528 1460 11537
rect 1420 11201 1460 11488
rect 1419 11192 1461 11201
rect 1419 11152 1420 11192
rect 1460 11152 1461 11192
rect 1419 11143 1461 11152
rect 1516 11024 1556 13420
rect 1611 13040 1653 13049
rect 1611 13000 1612 13040
rect 1652 13000 1653 13040
rect 1611 12991 1653 13000
rect 1612 11780 1652 12991
rect 1708 12881 1748 13756
rect 1707 12872 1749 12881
rect 1707 12832 1708 12872
rect 1748 12832 1749 12872
rect 1707 12823 1749 12832
rect 1804 11948 1844 14167
rect 1900 13964 1940 15259
rect 2091 14636 2133 14645
rect 2091 14596 2092 14636
rect 2132 14596 2133 14636
rect 2091 14587 2133 14596
rect 1995 14468 2037 14477
rect 1995 14428 1996 14468
rect 2036 14428 2037 14468
rect 1995 14419 2037 14428
rect 1900 13915 1940 13924
rect 1996 11957 2036 14419
rect 2092 14048 2132 14587
rect 2092 13999 2132 14008
rect 2283 14048 2325 14057
rect 2283 14008 2284 14048
rect 2324 14008 2325 14048
rect 2283 13999 2325 14008
rect 2380 14048 2420 14057
rect 2284 13914 2324 13999
rect 2188 13880 2228 13889
rect 2091 12788 2133 12797
rect 2091 12748 2092 12788
rect 2132 12748 2133 12788
rect 2091 12739 2133 12748
rect 1995 11948 2037 11957
rect 1804 11899 1844 11908
rect 1900 11908 1996 11948
rect 2036 11908 2037 11948
rect 1707 11864 1749 11873
rect 1707 11824 1708 11864
rect 1748 11824 1749 11864
rect 1707 11815 1749 11824
rect 1612 11731 1652 11740
rect 1708 11192 1748 11815
rect 1900 11780 1940 11908
rect 1995 11899 2037 11908
rect 1708 11143 1748 11152
rect 1804 11740 1940 11780
rect 1995 11780 2037 11789
rect 1995 11740 1996 11780
rect 2036 11740 2037 11780
rect 1420 10984 1556 11024
rect 1324 10772 1364 10781
rect 1324 9521 1364 10732
rect 1420 10436 1460 10984
rect 1611 10940 1653 10949
rect 1526 10929 1612 10940
rect 1566 10900 1612 10929
rect 1652 10900 1653 10940
rect 1611 10891 1653 10900
rect 1526 10880 1566 10889
rect 1420 10387 1460 10396
rect 1804 10352 1844 11740
rect 1995 11731 2037 11740
rect 1996 11646 2036 11731
rect 1899 11528 1941 11537
rect 1899 11488 1900 11528
rect 1940 11488 1941 11528
rect 1899 11479 1941 11488
rect 1900 10940 1940 11479
rect 2092 11360 2132 12739
rect 2188 12629 2228 13840
rect 2380 12713 2420 14008
rect 2572 14048 2612 15520
rect 2764 14384 2804 15679
rect 2860 14561 2900 16024
rect 3052 15896 3092 16263
rect 3147 16232 3189 16241
rect 3147 16192 3148 16232
rect 3188 16192 3189 16232
rect 3147 16183 3189 16192
rect 3244 16232 3284 16241
rect 2956 15856 3092 15896
rect 2956 14645 2996 15856
rect 3051 15728 3093 15737
rect 3051 15688 3052 15728
rect 3092 15688 3093 15728
rect 3051 15679 3093 15688
rect 3052 15560 3092 15679
rect 3148 15569 3188 16183
rect 3052 15511 3092 15520
rect 3147 15560 3189 15569
rect 3147 15520 3148 15560
rect 3188 15520 3189 15560
rect 3147 15511 3189 15520
rect 3148 15308 3188 15511
rect 3244 15476 3284 16192
rect 3339 16232 3381 16241
rect 3339 16192 3340 16232
rect 3380 16192 3381 16232
rect 3339 16183 3381 16192
rect 3531 16232 3573 16241
rect 3531 16192 3532 16232
rect 3572 16192 3573 16232
rect 3531 16183 3573 16192
rect 4108 16232 4148 16435
rect 4300 16241 4340 16771
rect 4108 16183 4148 16192
rect 4299 16232 4341 16241
rect 4299 16192 4300 16232
rect 4340 16192 4341 16232
rect 4299 16183 4341 16192
rect 3340 16098 3380 16183
rect 3532 16098 3572 16183
rect 3436 16064 3476 16073
rect 3436 15556 3476 16024
rect 4300 15821 4340 16183
rect 4299 15812 4341 15821
rect 4299 15772 4300 15812
rect 4340 15772 4341 15812
rect 4299 15763 4341 15772
rect 4396 15737 4436 19804
rect 4684 19794 4724 19879
rect 5260 19265 5300 19963
rect 5259 19256 5301 19265
rect 5259 19216 5260 19256
rect 5300 19216 5301 19256
rect 5259 19207 5301 19216
rect 5356 19088 5396 20224
rect 5452 20096 5492 20476
rect 5643 20467 5685 20476
rect 5547 20096 5589 20105
rect 5452 20056 5548 20096
rect 5588 20056 5589 20096
rect 5547 20047 5589 20056
rect 5548 19962 5588 20047
rect 5451 19760 5493 19769
rect 5451 19720 5452 19760
rect 5492 19720 5493 19760
rect 5451 19711 5493 19720
rect 5452 19256 5492 19711
rect 5644 19517 5684 20467
rect 5836 20096 5876 20105
rect 5740 20056 5836 20096
rect 5740 19685 5780 20056
rect 5836 20047 5876 20056
rect 5739 19676 5781 19685
rect 5739 19636 5740 19676
rect 5780 19636 5781 19676
rect 5739 19627 5781 19636
rect 5643 19508 5685 19517
rect 5643 19468 5644 19508
rect 5684 19468 5685 19508
rect 5643 19459 5685 19468
rect 5452 19207 5492 19216
rect 5644 19097 5684 19182
rect 5643 19088 5685 19097
rect 5356 19048 5492 19088
rect 4928 18920 5296 18929
rect 4968 18880 5010 18920
rect 5050 18880 5092 18920
rect 5132 18880 5174 18920
rect 5214 18880 5256 18920
rect 4928 18871 5296 18880
rect 4779 18836 4821 18845
rect 4779 18796 4780 18836
rect 4820 18796 4821 18836
rect 4779 18787 4821 18796
rect 4683 18080 4725 18089
rect 4683 18040 4684 18080
rect 4724 18040 4725 18080
rect 4683 18031 4725 18040
rect 4684 17912 4724 18031
rect 4599 17872 4724 17912
rect 4599 17828 4639 17872
rect 4588 17788 4639 17828
rect 4588 17786 4628 17788
rect 4780 17753 4820 18787
rect 5355 18584 5397 18593
rect 5355 18544 5356 18584
rect 5396 18544 5397 18584
rect 5355 18535 5397 18544
rect 4588 17737 4628 17746
rect 4684 17713 4820 17753
rect 5068 17749 5108 17758
rect 4684 17660 4724 17713
rect 4492 17620 4724 17660
rect 3974 15728 4016 15737
rect 3974 15688 3975 15728
rect 4015 15688 4016 15728
rect 3974 15679 4016 15688
rect 4395 15728 4437 15737
rect 4395 15688 4396 15728
rect 4436 15688 4437 15728
rect 4395 15679 4437 15688
rect 3436 15507 3476 15516
rect 3532 15560 3572 15571
rect 3532 15485 3572 15520
rect 3724 15560 3764 15569
rect 3339 15476 3381 15485
rect 3244 15436 3340 15476
rect 3380 15436 3381 15476
rect 3339 15427 3381 15436
rect 3531 15476 3573 15485
rect 3531 15436 3532 15476
rect 3572 15436 3573 15476
rect 3531 15427 3573 15436
rect 3244 15308 3284 15317
rect 3148 15268 3244 15308
rect 3052 14720 3092 14729
rect 3148 14720 3188 15268
rect 3244 15259 3284 15268
rect 3244 14972 3284 14981
rect 3340 14972 3380 15427
rect 3435 15308 3477 15317
rect 3724 15308 3764 15520
rect 3819 15560 3861 15569
rect 3819 15520 3820 15560
rect 3860 15520 3861 15560
rect 3819 15511 3861 15520
rect 3975 15560 4015 15679
rect 3975 15511 4015 15520
rect 3820 15426 3860 15511
rect 4395 15476 4437 15485
rect 4395 15436 4396 15476
rect 4436 15436 4437 15476
rect 4395 15427 4437 15436
rect 4396 15342 4436 15427
rect 3435 15268 3436 15308
rect 3476 15268 3477 15308
rect 3435 15259 3477 15268
rect 3532 15268 3764 15308
rect 4204 15308 4244 15317
rect 4244 15268 4340 15308
rect 3436 15174 3476 15259
rect 3284 14932 3380 14972
rect 3532 14972 3572 15268
rect 4204 15259 4244 15268
rect 3688 15140 4056 15149
rect 3728 15100 3770 15140
rect 3810 15100 3852 15140
rect 3892 15100 3934 15140
rect 3974 15100 4016 15140
rect 3688 15091 4056 15100
rect 3532 14932 3764 14972
rect 3244 14923 3284 14932
rect 3436 14720 3476 14729
rect 3148 14680 3436 14720
rect 2955 14636 2997 14645
rect 2955 14596 2956 14636
rect 2996 14596 2997 14636
rect 2955 14587 2997 14596
rect 2859 14552 2901 14561
rect 2859 14512 2860 14552
rect 2900 14512 2901 14552
rect 2859 14503 2901 14512
rect 3052 14384 3092 14680
rect 3436 14671 3476 14680
rect 3532 14720 3572 14729
rect 3532 14561 3572 14680
rect 3339 14552 3381 14561
rect 3339 14512 3340 14552
rect 3380 14512 3381 14552
rect 3339 14503 3381 14512
rect 3531 14552 3573 14561
rect 3531 14512 3532 14552
rect 3572 14512 3573 14552
rect 3531 14503 3573 14512
rect 3724 14552 3764 14932
rect 3724 14503 3764 14512
rect 4108 14720 4148 14729
rect 2764 14344 3092 14384
rect 2572 13553 2612 14008
rect 2667 14048 2709 14057
rect 2667 14008 2668 14048
rect 2708 14008 2709 14048
rect 2667 13999 2709 14008
rect 2571 13544 2613 13553
rect 2571 13504 2572 13544
rect 2612 13504 2613 13544
rect 2571 13495 2613 13504
rect 2668 13460 2708 13999
rect 2668 13411 2708 13420
rect 2764 13217 2804 14344
rect 3243 14048 3285 14057
rect 3243 14008 3244 14048
rect 3284 14008 3285 14048
rect 3243 13999 3285 14008
rect 2859 13544 2901 13553
rect 2859 13504 2860 13544
rect 2900 13504 2901 13544
rect 2859 13495 2901 13504
rect 2475 13208 2517 13217
rect 2475 13168 2476 13208
rect 2516 13168 2517 13208
rect 2475 13159 2517 13168
rect 2763 13208 2805 13217
rect 2763 13168 2764 13208
rect 2804 13168 2805 13208
rect 2763 13159 2805 13168
rect 2860 13208 2900 13495
rect 2900 13168 3092 13208
rect 2860 13159 2900 13168
rect 2379 12704 2421 12713
rect 2379 12664 2380 12704
rect 2420 12664 2421 12704
rect 2379 12655 2421 12664
rect 2187 12620 2229 12629
rect 2187 12580 2188 12620
rect 2228 12580 2229 12620
rect 2187 12571 2229 12580
rect 2476 12536 2516 13159
rect 2668 12713 2708 12798
rect 2667 12704 2709 12713
rect 2667 12664 2668 12704
rect 2708 12664 2709 12704
rect 2667 12655 2709 12664
rect 2955 12704 2997 12713
rect 2955 12664 2956 12704
rect 2996 12664 2997 12704
rect 2955 12655 2997 12664
rect 2763 12620 2805 12629
rect 2763 12580 2764 12620
rect 2804 12580 2900 12620
rect 2763 12571 2805 12580
rect 2187 11948 2229 11957
rect 2187 11908 2188 11948
rect 2228 11908 2229 11948
rect 2187 11899 2229 11908
rect 2188 11696 2228 11899
rect 2188 11647 2228 11656
rect 2379 11444 2421 11453
rect 2379 11404 2380 11444
rect 2420 11404 2421 11444
rect 2379 11395 2421 11404
rect 1900 10891 1940 10900
rect 1996 11320 2132 11360
rect 1708 10312 1844 10352
rect 1611 10268 1653 10277
rect 1611 10228 1612 10268
rect 1652 10228 1653 10268
rect 1611 10219 1653 10228
rect 1612 10134 1652 10219
rect 1708 9596 1748 10312
rect 1804 10184 1844 10193
rect 1804 10100 1844 10144
rect 1899 10100 1941 10109
rect 1804 10060 1900 10100
rect 1940 10060 1941 10100
rect 1899 10051 1941 10060
rect 1899 9848 1941 9857
rect 1899 9808 1900 9848
rect 1940 9808 1941 9848
rect 1899 9799 1941 9808
rect 1900 9680 1940 9799
rect 1900 9631 1940 9640
rect 1612 9556 1748 9596
rect 1323 9512 1365 9521
rect 1323 9472 1324 9512
rect 1364 9472 1365 9512
rect 1323 9463 1365 9472
rect 1323 9344 1365 9353
rect 1323 9304 1324 9344
rect 1364 9304 1365 9344
rect 1323 9295 1365 9304
rect 1227 8840 1269 8849
rect 1227 8800 1228 8840
rect 1268 8800 1269 8840
rect 1227 8791 1269 8800
rect 1228 8168 1268 8791
rect 1228 8119 1268 8128
rect 1324 7748 1364 9295
rect 1515 9260 1557 9269
rect 1515 9220 1516 9260
rect 1556 9220 1557 9260
rect 1515 9211 1557 9220
rect 1516 9126 1556 9211
rect 1419 8924 1461 8933
rect 1419 8884 1420 8924
rect 1460 8884 1461 8924
rect 1419 8875 1461 8884
rect 1420 7916 1460 8875
rect 1516 8504 1556 8513
rect 1516 8177 1556 8464
rect 1515 8168 1557 8177
rect 1515 8128 1516 8168
rect 1556 8128 1557 8168
rect 1612 8168 1652 9556
rect 1708 9428 1748 9437
rect 1996 9428 2036 11320
rect 2187 11108 2229 11117
rect 2187 11068 2188 11108
rect 2228 11068 2229 11108
rect 2187 11059 2229 11068
rect 2092 11024 2132 11033
rect 2092 9941 2132 10984
rect 2091 9932 2133 9941
rect 2091 9892 2092 9932
rect 2132 9892 2133 9932
rect 2091 9883 2133 9892
rect 1748 9388 2036 9428
rect 2091 9428 2133 9437
rect 2091 9388 2092 9428
rect 2132 9388 2133 9428
rect 1708 9379 1748 9388
rect 2091 9379 2133 9388
rect 2092 9294 2132 9379
rect 2188 9176 2228 11059
rect 2283 10184 2325 10193
rect 2283 10144 2284 10184
rect 2324 10144 2325 10184
rect 2283 10135 2325 10144
rect 2284 9680 2324 10135
rect 2284 9631 2324 9640
rect 1996 9136 2228 9176
rect 1707 8756 1749 8765
rect 1707 8716 1708 8756
rect 1748 8716 1749 8756
rect 1707 8707 1749 8716
rect 1708 8622 1748 8707
rect 1899 8504 1941 8513
rect 1899 8464 1900 8504
rect 1940 8464 1941 8504
rect 1899 8455 1941 8464
rect 1900 8370 1940 8455
rect 1803 8336 1845 8345
rect 1803 8296 1804 8336
rect 1844 8296 1845 8336
rect 1803 8287 1845 8296
rect 1612 8128 1748 8168
rect 1515 8119 1557 8128
rect 1515 8000 1557 8009
rect 1515 7960 1516 8000
rect 1556 7960 1557 8000
rect 1515 7951 1557 7960
rect 1612 8000 1652 8011
rect 1420 7867 1460 7876
rect 1324 7708 1460 7748
rect 1323 7496 1365 7505
rect 1323 7456 1324 7496
rect 1364 7456 1365 7496
rect 1323 7447 1365 7456
rect 1324 6656 1364 7447
rect 1324 6607 1364 6616
rect 1323 6152 1365 6161
rect 1323 6112 1324 6152
rect 1364 6112 1365 6152
rect 1323 6103 1365 6112
rect 1227 5396 1269 5405
rect 1227 5356 1228 5396
rect 1268 5356 1269 5396
rect 1227 5347 1269 5356
rect 1228 4724 1268 5347
rect 1324 4808 1364 6103
rect 1420 5648 1460 7708
rect 1516 7160 1556 7951
rect 1612 7925 1652 7960
rect 1611 7916 1653 7925
rect 1611 7876 1612 7916
rect 1652 7876 1653 7916
rect 1611 7867 1653 7876
rect 1708 7505 1748 8128
rect 1707 7496 1749 7505
rect 1707 7456 1708 7496
rect 1748 7456 1749 7496
rect 1707 7447 1749 7456
rect 1611 7412 1653 7421
rect 1611 7372 1612 7412
rect 1652 7372 1653 7412
rect 1611 7363 1653 7372
rect 1516 7111 1556 7120
rect 1516 6404 1556 6413
rect 1612 6404 1652 7363
rect 1707 6824 1749 6833
rect 1707 6784 1708 6824
rect 1748 6784 1749 6824
rect 1707 6775 1749 6784
rect 1708 6656 1748 6775
rect 1708 6607 1748 6616
rect 1556 6364 1652 6404
rect 1516 6355 1556 6364
rect 1420 5599 1460 5608
rect 1420 4976 1460 4985
rect 1804 4976 1844 8287
rect 1996 8252 2036 9136
rect 2380 8849 2420 11395
rect 2476 10613 2516 12496
rect 2860 12536 2900 12580
rect 2860 12487 2900 12496
rect 2956 12536 2996 12655
rect 3052 12629 3092 13168
rect 3244 12629 3284 13999
rect 3051 12620 3093 12629
rect 3051 12580 3052 12620
rect 3092 12580 3093 12620
rect 3051 12571 3093 12580
rect 3243 12620 3285 12629
rect 3243 12580 3244 12620
rect 3284 12580 3285 12620
rect 3243 12571 3285 12580
rect 2956 12487 2996 12496
rect 3147 12536 3189 12545
rect 3147 12496 3148 12536
rect 3188 12496 3189 12536
rect 3147 12487 3189 12496
rect 3244 12536 3284 12571
rect 3051 12452 3093 12461
rect 3051 12412 3052 12452
rect 3092 12412 3093 12452
rect 3051 12403 3093 12412
rect 2860 12284 2900 12293
rect 2475 10604 2517 10613
rect 2475 10564 2476 10604
rect 2516 10564 2517 10604
rect 2475 10555 2517 10564
rect 2475 10436 2517 10445
rect 2475 10396 2476 10436
rect 2516 10396 2517 10436
rect 2475 10387 2517 10396
rect 2476 9428 2516 10387
rect 2860 10025 2900 12244
rect 3052 11360 3092 12403
rect 3148 12402 3188 12487
rect 3244 12486 3284 12496
rect 3340 12545 3380 14503
rect 3819 14384 3861 14393
rect 3819 14344 3820 14384
rect 3860 14344 3861 14384
rect 3819 14335 3861 14344
rect 3820 14216 3860 14335
rect 3724 14176 3860 14216
rect 4012 14216 4052 14225
rect 4108 14216 4148 14680
rect 4203 14720 4245 14729
rect 4203 14680 4204 14720
rect 4244 14680 4245 14720
rect 4203 14671 4245 14680
rect 4204 14586 4244 14671
rect 4300 14393 4340 15268
rect 4299 14384 4341 14393
rect 4299 14344 4300 14384
rect 4340 14344 4341 14384
rect 4299 14335 4341 14344
rect 4052 14176 4148 14216
rect 3435 14048 3477 14057
rect 3435 14008 3436 14048
rect 3476 14008 3477 14048
rect 3435 13999 3477 14008
rect 3340 12536 3385 12545
rect 3340 12496 3345 12536
rect 3340 12487 3385 12496
rect 3340 11360 3380 12487
rect 2956 11320 3092 11360
rect 3148 11320 3380 11360
rect 3436 11696 3476 13999
rect 3724 13889 3764 14176
rect 4012 14167 4052 14176
rect 3819 14048 3861 14057
rect 4492 14048 4532 17620
rect 5068 17576 5108 17709
rect 5260 17585 5300 17670
rect 4780 17536 5108 17576
rect 5259 17576 5301 17585
rect 5259 17536 5260 17576
rect 5300 17536 5301 17576
rect 4780 17165 4820 17536
rect 5259 17527 5301 17536
rect 5356 17501 5396 18535
rect 5452 17660 5492 19048
rect 5643 19048 5644 19088
rect 5684 19048 5685 19088
rect 5643 19039 5685 19048
rect 5643 18920 5685 18929
rect 5643 18880 5644 18920
rect 5684 18880 5685 18920
rect 5643 18871 5685 18880
rect 5547 18752 5589 18761
rect 5547 18712 5548 18752
rect 5588 18712 5589 18752
rect 5547 18703 5589 18712
rect 5548 18593 5588 18703
rect 5547 18584 5589 18593
rect 5547 18544 5548 18584
rect 5588 18544 5589 18584
rect 5547 18535 5589 18544
rect 5548 18450 5588 18535
rect 5644 17753 5684 18871
rect 5740 18584 5780 19627
rect 5932 19256 5972 19265
rect 5932 19097 5972 19216
rect 6028 19256 6068 20887
rect 6124 20180 6164 21568
rect 6220 21559 6260 21568
rect 6315 21608 6357 21617
rect 6315 21568 6316 21608
rect 6356 21568 6357 21608
rect 6315 21559 6357 21568
rect 6316 21474 6356 21559
rect 6124 20140 6260 20180
rect 6220 19937 6260 20140
rect 6219 19928 6261 19937
rect 6219 19888 6220 19928
rect 6260 19888 6261 19928
rect 6219 19879 6261 19888
rect 6028 19181 6068 19216
rect 6123 19256 6165 19265
rect 6315 19256 6357 19265
rect 6123 19216 6124 19256
rect 6164 19216 6260 19256
rect 6123 19207 6165 19216
rect 6027 19172 6069 19181
rect 6027 19132 6028 19172
rect 6068 19132 6069 19172
rect 6027 19123 6069 19132
rect 5931 19088 5973 19097
rect 5931 19048 5932 19088
rect 5972 19048 5973 19088
rect 5931 19039 5973 19048
rect 6028 18584 6068 18595
rect 5740 18544 5876 18584
rect 5739 18416 5781 18425
rect 5739 18376 5740 18416
rect 5780 18376 5781 18416
rect 5739 18367 5781 18376
rect 5740 18282 5780 18367
rect 5643 17744 5685 17753
rect 5643 17704 5644 17744
rect 5684 17704 5685 17744
rect 5643 17695 5685 17704
rect 5452 17620 5588 17660
rect 5355 17492 5397 17501
rect 5355 17452 5356 17492
rect 5396 17452 5397 17492
rect 5355 17443 5397 17452
rect 4928 17408 5296 17417
rect 4968 17368 5010 17408
rect 5050 17368 5092 17408
rect 5132 17368 5174 17408
rect 5214 17368 5256 17408
rect 4928 17359 5296 17368
rect 4779 17156 4821 17165
rect 4779 17116 4780 17156
rect 4820 17116 4821 17156
rect 4779 17107 4821 17116
rect 5163 17156 5205 17165
rect 5163 17116 5164 17156
rect 5204 17116 5205 17156
rect 5163 17107 5205 17116
rect 4971 17072 5013 17081
rect 4971 17032 4972 17072
rect 5012 17032 5013 17072
rect 4971 17023 5013 17032
rect 4972 16938 5012 17023
rect 5164 17022 5204 17107
rect 5355 17072 5397 17081
rect 5355 17032 5356 17072
rect 5396 17032 5397 17072
rect 5355 17023 5397 17032
rect 4587 16652 4629 16661
rect 4587 16612 4588 16652
rect 4628 16612 4629 16652
rect 4587 16603 4629 16612
rect 3819 14008 3820 14048
rect 3860 14008 3861 14048
rect 3819 13999 3861 14008
rect 4204 14008 4532 14048
rect 4204 14006 4244 14008
rect 3820 13914 3860 13999
rect 4204 13957 4244 13966
rect 3723 13880 3765 13889
rect 3723 13840 3724 13880
rect 3764 13840 3765 13880
rect 3723 13831 3765 13840
rect 3688 13628 4056 13637
rect 3728 13588 3770 13628
rect 3810 13588 3852 13628
rect 3892 13588 3934 13628
rect 3974 13588 4016 13628
rect 3688 13579 4056 13588
rect 4492 13301 4532 14008
rect 4588 14804 4628 16603
rect 4779 16400 4821 16409
rect 4779 16360 4780 16400
rect 4820 16360 4821 16400
rect 4779 16351 4821 16360
rect 4588 13469 4628 14764
rect 4683 14804 4725 14813
rect 4683 14764 4684 14804
rect 4724 14764 4725 14804
rect 4683 14755 4725 14764
rect 4684 14670 4724 14755
rect 4587 13460 4629 13469
rect 4587 13420 4588 13460
rect 4628 13420 4629 13460
rect 4587 13411 4629 13420
rect 4683 13376 4725 13385
rect 4683 13336 4684 13376
rect 4724 13336 4725 13376
rect 4683 13327 4725 13336
rect 4491 13292 4533 13301
rect 4491 13252 4492 13292
rect 4532 13252 4533 13292
rect 4491 13243 4533 13252
rect 4107 13208 4149 13217
rect 4107 13168 4108 13208
rect 4148 13168 4149 13208
rect 4107 13159 4149 13168
rect 4108 13074 4148 13159
rect 4299 13124 4341 13133
rect 4299 13084 4300 13124
rect 4340 13084 4341 13124
rect 4299 13075 4341 13084
rect 4300 12990 4340 13075
rect 3916 12704 3956 12713
rect 3627 12620 3669 12629
rect 3627 12580 3628 12620
rect 3668 12580 3669 12620
rect 3627 12571 3669 12580
rect 3628 12536 3668 12571
rect 3628 12485 3668 12496
rect 3724 12536 3764 12547
rect 3916 12545 3956 12664
rect 3724 12461 3764 12496
rect 3915 12536 3957 12545
rect 3915 12496 3916 12536
rect 3956 12496 3957 12536
rect 4492 12536 4532 13243
rect 4588 13208 4628 13219
rect 4588 13133 4628 13168
rect 4684 13208 4724 13327
rect 4684 13159 4724 13168
rect 4587 13124 4629 13133
rect 4587 13084 4588 13124
rect 4628 13084 4629 13124
rect 4587 13075 4629 13084
rect 4588 12536 4628 12545
rect 4492 12496 4588 12536
rect 3915 12487 3957 12496
rect 4588 12487 4628 12496
rect 3723 12452 3765 12461
rect 3723 12412 3724 12452
rect 3764 12412 3765 12452
rect 3723 12403 3765 12412
rect 4395 12284 4437 12293
rect 4395 12244 4396 12284
rect 4436 12244 4437 12284
rect 4395 12235 4437 12244
rect 3688 12116 4056 12125
rect 3728 12076 3770 12116
rect 3810 12076 3852 12116
rect 3892 12076 3934 12116
rect 3974 12076 4016 12116
rect 3688 12067 4056 12076
rect 4396 11780 4436 12235
rect 4491 12032 4533 12041
rect 4491 11992 4492 12032
rect 4532 11992 4533 12032
rect 4491 11983 4533 11992
rect 4396 11731 4436 11740
rect 4492 11780 4532 11983
rect 4492 11731 4532 11740
rect 2859 10016 2901 10025
rect 2859 9976 2860 10016
rect 2900 9976 2901 10016
rect 2859 9967 2901 9976
rect 2956 9857 2996 11320
rect 3051 11192 3093 11201
rect 3051 11152 3052 11192
rect 3092 11152 3093 11192
rect 3051 11143 3093 11152
rect 3052 10184 3092 11143
rect 3052 10135 3092 10144
rect 2955 9848 2997 9857
rect 2955 9808 2956 9848
rect 2996 9808 2997 9848
rect 2955 9799 2997 9808
rect 2476 9379 2516 9388
rect 2764 9512 2804 9521
rect 2667 9176 2709 9185
rect 2667 9136 2668 9176
rect 2708 9136 2709 9176
rect 2667 9127 2709 9136
rect 2379 8840 2421 8849
rect 2379 8800 2380 8840
rect 2420 8800 2421 8840
rect 2379 8791 2421 8800
rect 1900 8212 2036 8252
rect 2092 8756 2132 8765
rect 1900 6404 1940 8212
rect 2092 7757 2132 8716
rect 2668 8672 2708 9127
rect 2764 9101 2804 9472
rect 2860 9512 2900 9521
rect 2763 9092 2805 9101
rect 2763 9052 2764 9092
rect 2804 9052 2805 9092
rect 2763 9043 2805 9052
rect 2860 8681 2900 9472
rect 3051 9512 3093 9521
rect 3051 9472 3052 9512
rect 3092 9472 3093 9512
rect 3051 9463 3093 9472
rect 3052 9378 3092 9463
rect 2956 9344 2996 9353
rect 2668 8623 2708 8632
rect 2764 8672 2804 8681
rect 2859 8672 2901 8681
rect 2804 8632 2860 8672
rect 2900 8632 2901 8672
rect 2764 8623 2804 8632
rect 2859 8623 2901 8632
rect 2956 8672 2996 9304
rect 3051 9092 3093 9101
rect 3051 9052 3052 9092
rect 3092 9052 3093 9092
rect 3051 9043 3093 9052
rect 2956 8623 2996 8632
rect 3052 8672 3092 9043
rect 2475 8504 2517 8513
rect 2475 8464 2476 8504
rect 2516 8464 2517 8504
rect 2475 8455 2517 8464
rect 2476 8370 2516 8455
rect 2667 8420 2709 8429
rect 2667 8380 2668 8420
rect 2708 8380 2709 8420
rect 2667 8371 2709 8380
rect 2668 8000 2708 8371
rect 2860 8177 2900 8623
rect 3052 8420 3092 8632
rect 2956 8380 3092 8420
rect 2859 8168 2901 8177
rect 2859 8128 2860 8168
rect 2900 8128 2901 8168
rect 2859 8119 2901 8128
rect 2860 8000 2900 8009
rect 2668 7960 2860 8000
rect 2091 7748 2133 7757
rect 2091 7708 2092 7748
rect 2132 7708 2133 7748
rect 2091 7699 2133 7708
rect 1995 7664 2037 7673
rect 1995 7624 1996 7664
rect 2036 7624 2037 7664
rect 1995 7615 2037 7624
rect 1900 6355 1940 6364
rect 1996 6320 2036 7615
rect 2764 7160 2804 7960
rect 2860 7951 2900 7960
rect 2859 7496 2901 7505
rect 2859 7456 2860 7496
rect 2900 7456 2901 7496
rect 2859 7447 2901 7456
rect 2764 7085 2804 7120
rect 2763 7076 2805 7085
rect 2763 7036 2764 7076
rect 2804 7036 2805 7076
rect 2763 7027 2805 7036
rect 2667 6992 2709 7001
rect 2764 6996 2804 7027
rect 2667 6952 2668 6992
rect 2708 6952 2709 6992
rect 2667 6943 2709 6952
rect 2668 6833 2708 6943
rect 2860 6833 2900 7447
rect 2956 7412 2996 8380
rect 3051 8168 3093 8177
rect 3051 8128 3052 8168
rect 3092 8128 3093 8168
rect 3051 8119 3093 8128
rect 3052 8034 3092 8119
rect 2956 7363 2996 7372
rect 3148 7160 3188 11320
rect 3339 11192 3381 11201
rect 3339 11152 3340 11192
rect 3380 11152 3381 11192
rect 3339 11143 3381 11152
rect 3340 11024 3380 11143
rect 3436 11033 3476 11656
rect 3916 11696 3956 11705
rect 3628 11612 3668 11621
rect 3916 11612 3956 11656
rect 3668 11572 3956 11612
rect 4012 11696 4052 11705
rect 3628 11563 3668 11572
rect 4012 11201 4052 11656
rect 4107 11528 4149 11537
rect 4780 11528 4820 16351
rect 5356 16232 5396 17023
rect 5548 16661 5588 17620
rect 5644 17610 5684 17695
rect 5836 16997 5876 18544
rect 6028 18509 6068 18544
rect 6123 18584 6165 18593
rect 6123 18544 6124 18584
rect 6164 18544 6165 18584
rect 6123 18535 6165 18544
rect 6027 18500 6069 18509
rect 6027 18460 6028 18500
rect 6068 18460 6069 18500
rect 6027 18451 6069 18460
rect 6124 18450 6164 18535
rect 5931 18416 5973 18425
rect 5931 18376 5932 18416
rect 5972 18376 5973 18416
rect 5931 18367 5973 18376
rect 5835 16988 5877 16997
rect 5835 16948 5836 16988
rect 5876 16948 5877 16988
rect 5835 16939 5877 16948
rect 5547 16652 5589 16661
rect 5547 16612 5548 16652
rect 5588 16612 5589 16652
rect 5547 16603 5589 16612
rect 5548 16400 5588 16409
rect 5932 16400 5972 18367
rect 6027 17324 6069 17333
rect 6027 17284 6028 17324
rect 6068 17284 6069 17324
rect 6027 17275 6069 17284
rect 6028 17072 6068 17275
rect 6028 16661 6068 17032
rect 6027 16652 6069 16661
rect 6027 16612 6028 16652
rect 6068 16612 6069 16652
rect 6027 16603 6069 16612
rect 5588 16360 5780 16400
rect 5932 16360 6068 16400
rect 5548 16351 5588 16360
rect 5740 16315 5780 16360
rect 5740 16275 5876 16315
rect 5836 16251 5876 16275
rect 5836 16202 5876 16211
rect 5931 16232 5973 16241
rect 4928 15896 5296 15905
rect 4968 15856 5010 15896
rect 5050 15856 5092 15896
rect 5132 15856 5174 15896
rect 5214 15856 5256 15896
rect 4928 15847 5296 15856
rect 5260 15560 5300 15569
rect 5260 15317 5300 15520
rect 5259 15308 5301 15317
rect 5259 15268 5260 15308
rect 5300 15268 5301 15308
rect 5259 15259 5301 15268
rect 5163 14972 5205 14981
rect 5163 14932 5164 14972
rect 5204 14932 5205 14972
rect 5163 14923 5205 14932
rect 5164 14720 5204 14923
rect 5164 14671 5204 14680
rect 4928 14384 5296 14393
rect 4968 14344 5010 14384
rect 5050 14344 5092 14384
rect 5132 14344 5174 14384
rect 5214 14344 5256 14384
rect 4928 14335 5296 14344
rect 4971 14132 5013 14141
rect 4971 14092 4972 14132
rect 5012 14092 5013 14132
rect 4971 14083 5013 14092
rect 4972 13124 5012 14083
rect 5356 14048 5396 16192
rect 5931 16192 5932 16232
rect 5972 16192 5973 16232
rect 5931 16183 5973 16192
rect 5932 15821 5972 16183
rect 5931 15812 5973 15821
rect 5931 15772 5932 15812
rect 5972 15772 5973 15812
rect 5931 15763 5973 15772
rect 5644 14725 5684 14734
rect 5644 14216 5684 14685
rect 5835 14636 5877 14645
rect 5835 14596 5836 14636
rect 5876 14596 5877 14636
rect 5835 14587 5877 14596
rect 5836 14502 5876 14587
rect 5644 14167 5684 14176
rect 5835 14216 5877 14225
rect 5835 14176 5836 14216
rect 5876 14176 5877 14216
rect 5835 14167 5877 14176
rect 5451 14048 5493 14057
rect 5356 14008 5452 14048
rect 5492 14008 5493 14048
rect 5451 13999 5493 14008
rect 5452 13914 5492 13999
rect 5067 13460 5109 13469
rect 5067 13420 5068 13460
rect 5108 13420 5109 13460
rect 5067 13411 5109 13420
rect 5068 13292 5108 13411
rect 5068 13243 5108 13252
rect 5643 13292 5685 13301
rect 5643 13252 5644 13292
rect 5684 13252 5685 13292
rect 5643 13243 5685 13252
rect 5164 13208 5204 13217
rect 5164 13124 5204 13168
rect 4972 13084 5204 13124
rect 5164 13040 5204 13084
rect 5644 13208 5684 13243
rect 5836 13217 5876 14167
rect 5164 13000 5396 13040
rect 4928 12872 5296 12881
rect 4968 12832 5010 12872
rect 5050 12832 5092 12872
rect 5132 12832 5174 12872
rect 5214 12832 5256 12872
rect 4928 12823 5296 12832
rect 5356 12041 5396 13000
rect 5355 12032 5397 12041
rect 5355 11992 5356 12032
rect 5396 11992 5397 12032
rect 5355 11983 5397 11992
rect 5644 11873 5684 13168
rect 5835 13208 5877 13217
rect 5835 13168 5836 13208
rect 5876 13168 5877 13208
rect 5835 13159 5877 13168
rect 5836 12536 5876 13159
rect 6028 12881 6068 16360
rect 6220 14813 6260 19216
rect 6315 19216 6316 19256
rect 6356 19216 6357 19256
rect 6315 19207 6357 19216
rect 6412 19256 6452 22072
rect 6507 21860 6549 21869
rect 6507 21820 6508 21860
rect 6548 21820 6549 21860
rect 6507 21811 6549 21820
rect 6508 21608 6548 21811
rect 6508 21559 6548 21568
rect 6604 19685 6644 22072
rect 6700 22062 6740 22147
rect 6796 22146 6836 22231
rect 6987 22028 7029 22037
rect 6987 21988 6988 22028
rect 7028 21988 7029 22028
rect 6987 21979 7029 21988
rect 6795 21944 6837 21953
rect 6795 21904 6796 21944
rect 6836 21904 6837 21944
rect 6795 21895 6837 21904
rect 6699 21776 6741 21785
rect 6699 21736 6700 21776
rect 6740 21736 6741 21776
rect 6699 21727 6741 21736
rect 6700 21608 6740 21727
rect 6700 21559 6740 21568
rect 6796 21608 6836 21895
rect 6988 21776 7028 21979
rect 6988 21727 7028 21736
rect 6796 21440 6836 21568
rect 6892 21608 6932 21617
rect 6932 21568 7028 21608
rect 6892 21559 6932 21568
rect 6796 21400 6932 21440
rect 6699 21356 6741 21365
rect 6699 21316 6700 21356
rect 6740 21316 6741 21356
rect 6699 21307 6741 21316
rect 6603 19676 6645 19685
rect 6603 19636 6604 19676
rect 6644 19636 6645 19676
rect 6603 19627 6645 19636
rect 6700 19349 6740 21307
rect 6796 20768 6836 20777
rect 6796 20441 6836 20728
rect 6795 20432 6837 20441
rect 6795 20392 6796 20432
rect 6836 20392 6837 20432
rect 6795 20383 6837 20392
rect 6796 19853 6836 20383
rect 6795 19844 6837 19853
rect 6795 19804 6796 19844
rect 6836 19804 6837 19844
rect 6795 19795 6837 19804
rect 6795 19676 6837 19685
rect 6795 19636 6796 19676
rect 6836 19636 6837 19676
rect 6795 19627 6837 19636
rect 6507 19340 6549 19349
rect 6507 19300 6508 19340
rect 6548 19300 6549 19340
rect 6507 19291 6549 19300
rect 6699 19340 6741 19349
rect 6699 19300 6700 19340
rect 6740 19300 6741 19340
rect 6699 19291 6741 19300
rect 6316 16829 6356 19207
rect 6412 18593 6452 19216
rect 6508 19206 6548 19291
rect 6603 19256 6645 19265
rect 6603 19216 6604 19256
rect 6644 19216 6645 19256
rect 6603 19207 6645 19216
rect 6604 19088 6644 19207
rect 6699 19172 6741 19181
rect 6699 19132 6700 19172
rect 6740 19132 6741 19172
rect 6699 19123 6741 19132
rect 6508 19048 6644 19088
rect 6411 18584 6453 18593
rect 6411 18544 6412 18584
rect 6452 18544 6453 18584
rect 6411 18535 6453 18544
rect 6508 18584 6548 19048
rect 6603 18836 6645 18845
rect 6603 18796 6604 18836
rect 6644 18796 6645 18836
rect 6603 18787 6645 18796
rect 6508 18535 6548 18544
rect 6604 18584 6644 18787
rect 6604 18500 6644 18544
rect 6599 18460 6644 18500
rect 6599 18416 6639 18460
rect 6508 18376 6639 18416
rect 6315 16820 6357 16829
rect 6315 16780 6316 16820
rect 6356 16780 6357 16820
rect 6315 16771 6357 16780
rect 6508 16325 6548 18376
rect 6700 18332 6740 19123
rect 6796 18761 6836 19627
rect 6795 18752 6837 18761
rect 6795 18712 6796 18752
rect 6836 18712 6837 18752
rect 6892 18752 6932 21400
rect 6988 20861 7028 21568
rect 7084 20945 7124 22576
rect 7179 21692 7221 21701
rect 7179 21652 7180 21692
rect 7220 21652 7221 21692
rect 7179 21643 7221 21652
rect 7180 21608 7220 21643
rect 7180 21557 7220 21568
rect 7179 21440 7221 21449
rect 7179 21400 7180 21440
rect 7220 21400 7221 21440
rect 7179 21391 7221 21400
rect 7180 21306 7220 21391
rect 7276 21188 7316 23080
rect 7564 21869 7604 23911
rect 7660 23549 7700 25507
rect 7756 25318 7796 25843
rect 7756 25269 7796 25278
rect 7852 24557 7892 26692
rect 7948 26683 7988 26692
rect 8139 26732 8181 26741
rect 8139 26692 8140 26732
rect 8180 26692 8181 26732
rect 8139 26683 8181 26692
rect 8140 26598 8180 26683
rect 8236 25472 8276 31303
rect 8332 30680 8372 31387
rect 8332 30631 8372 30640
rect 8332 29849 8372 29934
rect 8331 29840 8373 29849
rect 8331 29800 8332 29840
rect 8372 29800 8373 29840
rect 8331 29791 8373 29800
rect 8428 29672 8468 32068
rect 8716 31940 8756 31949
rect 8524 30764 8564 30775
rect 8524 30689 8564 30724
rect 8523 30680 8565 30689
rect 8523 30640 8524 30680
rect 8564 30640 8565 30680
rect 8523 30631 8565 30640
rect 8619 30512 8661 30521
rect 8619 30472 8620 30512
rect 8660 30472 8661 30512
rect 8619 30463 8661 30472
rect 8332 29632 8468 29672
rect 8524 29672 8564 29681
rect 8332 28337 8372 29632
rect 8524 29168 8564 29632
rect 8620 29588 8660 30463
rect 8716 29765 8756 31900
rect 8812 31025 8852 34075
rect 8908 33284 8948 34336
rect 9003 34376 9045 34385
rect 9003 34336 9004 34376
rect 9044 34336 9045 34376
rect 9003 34327 9045 34336
rect 9004 34242 9044 34327
rect 8908 33244 9044 33284
rect 8811 31016 8853 31025
rect 8811 30976 8812 31016
rect 8852 30976 8853 31016
rect 8811 30967 8853 30976
rect 8812 30689 8852 30774
rect 8811 30680 8853 30689
rect 8811 30640 8812 30680
rect 8852 30640 8853 30680
rect 8811 30631 8853 30640
rect 8908 30680 8948 30689
rect 8811 30512 8853 30521
rect 8908 30512 8948 30640
rect 8811 30472 8812 30512
rect 8852 30472 8948 30512
rect 8811 30463 8853 30472
rect 8907 30344 8949 30353
rect 8907 30304 8908 30344
rect 8948 30304 8949 30344
rect 8907 30295 8949 30304
rect 8715 29756 8757 29765
rect 8715 29716 8716 29756
rect 8756 29716 8757 29756
rect 8715 29707 8757 29716
rect 8620 29548 8756 29588
rect 8619 29252 8661 29261
rect 8619 29212 8620 29252
rect 8660 29212 8661 29252
rect 8619 29203 8661 29212
rect 8476 29158 8564 29168
rect 8516 29128 8564 29158
rect 8620 29118 8660 29203
rect 8476 29109 8516 29118
rect 8331 28328 8373 28337
rect 8331 28288 8332 28328
rect 8372 28288 8373 28328
rect 8331 28279 8373 28288
rect 8619 27656 8661 27665
rect 8619 27616 8620 27656
rect 8660 27616 8661 27656
rect 8619 27607 8661 27616
rect 8716 27656 8756 29548
rect 8811 29504 8853 29513
rect 8811 29464 8812 29504
rect 8852 29464 8853 29504
rect 8811 29455 8853 29464
rect 8620 27522 8660 27607
rect 8331 26984 8373 26993
rect 8331 26944 8332 26984
rect 8372 26944 8373 26984
rect 8331 26935 8373 26944
rect 8332 26816 8372 26935
rect 8332 26767 8372 26776
rect 8716 25640 8756 27616
rect 8812 26153 8852 29455
rect 8811 26144 8853 26153
rect 8811 26104 8812 26144
rect 8852 26104 8853 26144
rect 8811 26095 8853 26104
rect 8044 25432 8276 25472
rect 8524 25600 8756 25640
rect 7947 25220 7989 25229
rect 7947 25180 7948 25220
rect 7988 25180 7989 25220
rect 7947 25171 7989 25180
rect 7948 25086 7988 25171
rect 8044 24968 8084 25432
rect 7948 24928 8084 24968
rect 8140 25304 8180 25313
rect 7851 24548 7893 24557
rect 7851 24508 7852 24548
rect 7892 24508 7893 24548
rect 7851 24499 7893 24508
rect 7755 23792 7797 23801
rect 7755 23752 7756 23792
rect 7796 23752 7797 23792
rect 7755 23743 7797 23752
rect 7756 23658 7796 23743
rect 7659 23540 7701 23549
rect 7659 23500 7660 23540
rect 7700 23500 7796 23540
rect 7659 23491 7701 23500
rect 7659 22280 7701 22289
rect 7659 22240 7660 22280
rect 7700 22240 7701 22280
rect 7659 22231 7701 22240
rect 7371 21860 7413 21869
rect 7371 21820 7372 21860
rect 7412 21820 7413 21860
rect 7371 21811 7413 21820
rect 7563 21860 7605 21869
rect 7563 21820 7564 21860
rect 7604 21820 7605 21860
rect 7660 21860 7700 22231
rect 7756 21944 7796 23500
rect 7948 22028 7988 24928
rect 8043 23960 8085 23969
rect 8043 23920 8044 23960
rect 8084 23920 8085 23960
rect 8043 23911 8085 23920
rect 8044 23792 8084 23911
rect 8140 23885 8180 25264
rect 8236 25304 8276 25313
rect 8236 24473 8276 25264
rect 8428 25136 8468 25147
rect 8428 25061 8468 25096
rect 8427 25052 8469 25061
rect 8427 25012 8428 25052
rect 8468 25012 8469 25052
rect 8427 25003 8469 25012
rect 8235 24464 8277 24473
rect 8235 24424 8236 24464
rect 8276 24424 8277 24464
rect 8235 24415 8277 24424
rect 8428 23960 8468 23969
rect 8236 23920 8428 23960
rect 8139 23876 8181 23885
rect 8139 23836 8140 23876
rect 8180 23836 8181 23876
rect 8139 23827 8181 23836
rect 8044 23743 8084 23752
rect 8140 23708 8180 23717
rect 8140 23549 8180 23668
rect 8139 23540 8181 23549
rect 8139 23500 8140 23540
rect 8180 23500 8181 23540
rect 8139 23491 8181 23500
rect 8236 23120 8276 23920
rect 8428 23911 8468 23920
rect 8331 23792 8373 23801
rect 8331 23752 8332 23792
rect 8372 23752 8373 23792
rect 8331 23743 8373 23752
rect 8044 23080 8276 23120
rect 8044 22280 8084 23080
rect 8139 22868 8181 22877
rect 8139 22828 8140 22868
rect 8180 22828 8181 22868
rect 8139 22819 8181 22828
rect 8044 22231 8084 22240
rect 8140 22280 8180 22819
rect 8332 22532 8372 23743
rect 8427 23624 8469 23633
rect 8427 23584 8428 23624
rect 8468 23584 8469 23624
rect 8524 23624 8564 25600
rect 8715 25052 8757 25061
rect 8715 25012 8716 25052
rect 8756 25012 8757 25052
rect 8715 25003 8757 25012
rect 8620 23801 8660 23886
rect 8619 23792 8661 23801
rect 8619 23752 8620 23792
rect 8660 23752 8661 23792
rect 8619 23743 8661 23752
rect 8716 23792 8756 25003
rect 8812 24632 8852 26095
rect 8812 24305 8852 24592
rect 8811 24296 8853 24305
rect 8811 24256 8812 24296
rect 8852 24256 8853 24296
rect 8811 24247 8853 24256
rect 8908 24044 8948 30295
rect 9004 30269 9044 33244
rect 9100 31940 9140 31949
rect 9100 31352 9140 31900
rect 9196 31613 9236 38116
rect 9484 38072 9524 39796
rect 10635 39752 10677 39761
rect 10635 39712 10636 39752
rect 10676 39712 10677 39752
rect 10635 39703 10677 39712
rect 10444 39500 10484 39509
rect 10155 39080 10197 39089
rect 10155 39040 10156 39080
rect 10196 39040 10197 39080
rect 10155 39031 10197 39040
rect 10156 38926 10196 39031
rect 9676 38912 9716 38921
rect 10156 38877 10196 38886
rect 9676 38669 9716 38872
rect 10347 38744 10389 38753
rect 10347 38704 10348 38744
rect 10388 38704 10389 38744
rect 10347 38695 10389 38704
rect 9675 38660 9717 38669
rect 9675 38620 9676 38660
rect 9716 38620 9717 38660
rect 9675 38611 9717 38620
rect 9292 38032 9524 38072
rect 9580 38240 9620 38249
rect 9676 38240 9716 38611
rect 10348 38610 10388 38695
rect 9620 38200 9716 38240
rect 10252 38324 10292 38333
rect 10060 38226 10100 38235
rect 9292 32192 9332 38032
rect 9580 37820 9620 38200
rect 9388 37780 9620 37820
rect 9964 38186 10060 38226
rect 9388 35888 9428 37780
rect 9771 37736 9813 37745
rect 9771 37696 9772 37736
rect 9812 37696 9813 37736
rect 9771 37687 9813 37696
rect 9675 37652 9717 37661
rect 9675 37612 9676 37652
rect 9716 37612 9717 37652
rect 9675 37603 9717 37612
rect 9676 36737 9716 37603
rect 9772 37409 9812 37687
rect 9964 37493 10004 38186
rect 10060 38177 10100 38186
rect 10252 37913 10292 38284
rect 10251 37904 10293 37913
rect 10251 37864 10252 37904
rect 10292 37864 10293 37904
rect 10251 37855 10293 37864
rect 10444 37745 10484 39460
rect 10636 39257 10676 39703
rect 10635 39248 10677 39257
rect 10635 39208 10636 39248
rect 10676 39208 10677 39248
rect 10635 39199 10677 39208
rect 11116 37820 11156 40216
rect 11500 38912 11540 40459
rect 11404 38872 11500 38912
rect 11404 37988 11444 38872
rect 11500 38863 11540 38872
rect 11499 38240 11541 38249
rect 11499 38200 11500 38240
rect 11540 38200 11541 38240
rect 11499 38191 11541 38200
rect 11500 38106 11540 38191
rect 10732 37780 11156 37820
rect 11308 37948 11444 37988
rect 10347 37736 10389 37745
rect 10347 37696 10348 37736
rect 10388 37696 10389 37736
rect 10347 37687 10389 37696
rect 10443 37736 10485 37745
rect 10443 37696 10444 37736
rect 10484 37696 10485 37736
rect 10443 37687 10485 37696
rect 9963 37484 10005 37493
rect 9963 37444 9964 37484
rect 10004 37444 10005 37484
rect 9963 37435 10005 37444
rect 9771 37400 9813 37409
rect 10252 37400 10292 37409
rect 9771 37360 9772 37400
rect 9812 37360 9813 37400
rect 9771 37351 9813 37360
rect 10060 37360 10252 37400
rect 9675 36728 9717 36737
rect 9675 36688 9676 36728
rect 9716 36688 9717 36728
rect 9675 36679 9717 36688
rect 9579 36224 9621 36233
rect 9579 36184 9580 36224
rect 9620 36184 9621 36224
rect 9579 36175 9621 36184
rect 9580 35981 9620 36175
rect 9579 35972 9621 35981
rect 9579 35932 9580 35972
rect 9620 35932 9621 35972
rect 9579 35923 9621 35932
rect 9428 35848 9524 35888
rect 9388 35839 9428 35848
rect 9387 35552 9429 35561
rect 9387 35512 9388 35552
rect 9428 35512 9429 35552
rect 9387 35503 9429 35512
rect 9195 31604 9237 31613
rect 9195 31564 9196 31604
rect 9236 31564 9237 31604
rect 9195 31555 9237 31564
rect 9292 31445 9332 32152
rect 9291 31436 9333 31445
rect 9291 31396 9292 31436
rect 9332 31396 9333 31436
rect 9291 31387 9333 31396
rect 9003 30260 9045 30269
rect 9003 30220 9004 30260
rect 9044 30220 9045 30260
rect 9003 30211 9045 30220
rect 9004 29840 9044 29849
rect 9100 29840 9140 31312
rect 9388 31352 9428 35503
rect 9484 34376 9524 35848
rect 9484 33536 9524 34336
rect 9580 34133 9620 35923
rect 9676 35561 9716 36679
rect 9772 35804 9812 37351
rect 10060 36905 10100 37360
rect 10252 37351 10292 37360
rect 10155 36980 10197 36989
rect 10155 36940 10156 36980
rect 10196 36940 10197 36980
rect 10155 36931 10197 36940
rect 10059 36896 10101 36905
rect 10059 36856 10060 36896
rect 10100 36856 10101 36896
rect 10059 36847 10101 36856
rect 10060 36653 10100 36847
rect 10059 36644 10101 36653
rect 10059 36604 10060 36644
rect 10100 36604 10101 36644
rect 10059 36595 10101 36604
rect 10059 36392 10101 36401
rect 10059 36352 10060 36392
rect 10100 36352 10101 36392
rect 10059 36343 10101 36352
rect 9916 35897 9956 35906
rect 10060 35897 10100 36343
rect 10059 35888 10101 35897
rect 9956 35857 10004 35888
rect 9916 35848 10004 35857
rect 9772 35764 9908 35804
rect 9675 35552 9717 35561
rect 9675 35512 9676 35552
rect 9716 35512 9717 35552
rect 9675 35503 9717 35512
rect 9772 35216 9812 35225
rect 9676 35176 9772 35216
rect 9579 34124 9621 34133
rect 9579 34084 9580 34124
rect 9620 34084 9621 34124
rect 9579 34075 9621 34084
rect 9580 33713 9620 33798
rect 9579 33704 9621 33713
rect 9676 33704 9716 35176
rect 9772 35167 9812 35176
rect 9772 33881 9812 33966
rect 9771 33872 9813 33881
rect 9771 33832 9772 33872
rect 9812 33832 9813 33872
rect 9771 33823 9813 33832
rect 9868 33704 9908 35764
rect 9964 35384 10004 35848
rect 10059 35848 10060 35888
rect 10100 35848 10101 35888
rect 10059 35839 10101 35848
rect 9964 35335 10004 35344
rect 10060 35720 10100 35729
rect 10060 35057 10100 35680
rect 10059 35048 10101 35057
rect 10059 35008 10060 35048
rect 10100 35008 10101 35048
rect 10059 34999 10101 35008
rect 9964 34381 10004 34390
rect 9964 33881 10004 34341
rect 10059 34376 10101 34385
rect 10059 34336 10060 34376
rect 10100 34336 10101 34376
rect 10156 34376 10196 36931
rect 10348 36896 10388 37687
rect 10444 37568 10484 37579
rect 10444 37493 10484 37528
rect 10443 37484 10485 37493
rect 10443 37444 10444 37484
rect 10484 37444 10485 37484
rect 10443 37435 10485 37444
rect 10732 36989 10772 37780
rect 11308 37745 11348 37948
rect 11596 37829 11636 41467
rect 11691 39164 11733 39173
rect 11691 39124 11692 39164
rect 11732 39124 11733 39164
rect 11691 39115 11733 39124
rect 11692 38249 11732 39115
rect 11691 38240 11733 38249
rect 11691 38200 11692 38240
rect 11732 38200 11733 38240
rect 11691 38191 11733 38200
rect 11403 37820 11445 37829
rect 11403 37780 11404 37820
rect 11444 37780 11445 37820
rect 11403 37771 11445 37780
rect 11595 37820 11637 37829
rect 11788 37820 11828 43408
rect 12172 43373 12212 43408
rect 12171 43364 12213 43373
rect 12171 43324 12172 43364
rect 12212 43324 12213 43364
rect 12171 43315 12213 43324
rect 12364 42776 12404 42785
rect 12460 42776 12500 44407
rect 12404 42736 12500 42776
rect 12076 41945 12116 42030
rect 12075 41936 12117 41945
rect 12075 41896 12076 41936
rect 12116 41896 12117 41936
rect 12075 41887 12117 41896
rect 12268 41768 12308 41777
rect 12076 41728 12268 41768
rect 12076 41264 12116 41728
rect 12268 41719 12308 41728
rect 12028 41254 12116 41264
rect 12068 41224 12116 41254
rect 12172 41348 12212 41357
rect 12028 41205 12068 41214
rect 11883 39752 11925 39761
rect 11883 39712 11884 39752
rect 11924 39712 11925 39752
rect 11883 39703 11925 39712
rect 11884 39618 11924 39703
rect 11595 37780 11596 37820
rect 11636 37780 11637 37820
rect 11595 37771 11637 37780
rect 11692 37780 11828 37820
rect 11307 37736 11349 37745
rect 11307 37696 11308 37736
rect 11348 37696 11349 37736
rect 11307 37687 11349 37696
rect 11116 37400 11156 37409
rect 10923 37316 10965 37325
rect 10923 37276 10924 37316
rect 10964 37276 10965 37316
rect 10923 37267 10965 37276
rect 10731 36980 10773 36989
rect 10731 36940 10732 36980
rect 10772 36940 10773 36980
rect 10731 36931 10773 36940
rect 10251 36856 10388 36896
rect 10827 36896 10869 36905
rect 10827 36856 10828 36896
rect 10868 36856 10869 36896
rect 10251 36812 10291 36856
rect 10827 36847 10869 36856
rect 10251 36772 10292 36812
rect 10252 36728 10292 36772
rect 10828 36762 10868 36847
rect 10252 36065 10292 36688
rect 10347 36728 10389 36737
rect 10540 36728 10580 36737
rect 10347 36688 10348 36728
rect 10388 36688 10389 36728
rect 10347 36679 10389 36688
rect 10444 36688 10540 36728
rect 10348 36594 10388 36679
rect 10347 36392 10389 36401
rect 10347 36352 10348 36392
rect 10388 36352 10389 36392
rect 10347 36343 10389 36352
rect 10251 36056 10293 36065
rect 10251 36016 10252 36056
rect 10292 36016 10293 36056
rect 10251 36007 10293 36016
rect 10252 35888 10292 35897
rect 10252 34973 10292 35848
rect 10251 34964 10293 34973
rect 10251 34924 10252 34964
rect 10292 34924 10293 34964
rect 10251 34915 10293 34924
rect 10156 34336 10292 34376
rect 10059 34327 10101 34336
rect 9963 33872 10005 33881
rect 9963 33832 9964 33872
rect 10004 33832 10005 33872
rect 9963 33823 10005 33832
rect 9579 33664 9580 33704
rect 9620 33664 9716 33704
rect 9772 33664 9908 33704
rect 9964 33704 10004 33713
rect 9579 33655 9621 33664
rect 9484 33496 9620 33536
rect 9196 31184 9236 31193
rect 9196 31025 9236 31144
rect 9388 31109 9428 31312
rect 9387 31100 9429 31109
rect 9387 31060 9388 31100
rect 9428 31060 9429 31100
rect 9387 31051 9429 31060
rect 9195 31016 9237 31025
rect 9195 30976 9196 31016
rect 9236 30976 9237 31016
rect 9195 30967 9237 30976
rect 9387 30764 9429 30773
rect 9387 30724 9388 30764
rect 9428 30724 9429 30764
rect 9387 30715 9429 30724
rect 9292 30680 9332 30689
rect 9196 30640 9292 30666
rect 9196 30626 9332 30640
rect 9388 30638 9428 30715
rect 9196 30428 9236 30626
rect 9483 30680 9525 30689
rect 9483 30640 9484 30680
rect 9524 30640 9525 30680
rect 9483 30631 9525 30640
rect 9388 30589 9428 30598
rect 9196 30388 9332 30428
rect 9196 30017 9236 30102
rect 9195 30008 9237 30017
rect 9195 29968 9196 30008
rect 9236 29968 9237 30008
rect 9195 29959 9237 29968
rect 9044 29800 9140 29840
rect 9195 29840 9237 29849
rect 9195 29800 9196 29840
rect 9236 29800 9237 29840
rect 9004 29791 9044 29800
rect 9195 29791 9237 29800
rect 9196 29706 9236 29791
rect 9004 29168 9044 29177
rect 9004 28421 9044 29128
rect 9292 28664 9332 30388
rect 9387 30344 9429 30353
rect 9387 30304 9388 30344
rect 9428 30304 9429 30344
rect 9387 30295 9429 30304
rect 9100 28624 9332 28664
rect 9003 28412 9045 28421
rect 9003 28372 9004 28412
rect 9044 28372 9045 28412
rect 9003 28363 9045 28372
rect 9100 27749 9140 28624
rect 9292 28328 9332 28337
rect 9292 28169 9332 28288
rect 9291 28160 9333 28169
rect 9291 28120 9292 28160
rect 9332 28120 9333 28160
rect 9291 28111 9333 28120
rect 9291 27908 9333 27917
rect 9291 27868 9292 27908
rect 9332 27868 9333 27908
rect 9291 27859 9333 27868
rect 9099 27740 9141 27749
rect 9099 27700 9100 27740
rect 9140 27700 9141 27740
rect 9099 27691 9141 27700
rect 9100 27656 9140 27691
rect 9100 27606 9140 27616
rect 9196 27572 9236 27581
rect 9003 26144 9045 26153
rect 9003 26104 9004 26144
rect 9044 26104 9045 26144
rect 9003 26095 9045 26104
rect 9004 26010 9044 26095
rect 9196 26060 9236 27532
rect 9100 26020 9236 26060
rect 9100 25817 9140 26020
rect 9196 25892 9236 25901
rect 9099 25808 9141 25817
rect 9099 25768 9100 25808
rect 9140 25768 9141 25808
rect 9099 25759 9141 25768
rect 9196 25733 9236 25852
rect 9195 25724 9237 25733
rect 9195 25684 9196 25724
rect 9236 25684 9237 25724
rect 9195 25675 9237 25684
rect 9292 24809 9332 27859
rect 9291 24800 9333 24809
rect 9291 24760 9292 24800
rect 9332 24760 9333 24800
rect 9388 24800 9428 30295
rect 9484 29840 9524 30631
rect 9484 29791 9524 29800
rect 9483 29672 9525 29681
rect 9483 29632 9484 29672
rect 9524 29632 9525 29672
rect 9483 29623 9525 29632
rect 9484 29000 9524 29623
rect 9580 29177 9620 33496
rect 9675 30932 9717 30941
rect 9675 30892 9676 30932
rect 9716 30892 9717 30932
rect 9675 30883 9717 30892
rect 9676 30773 9716 30883
rect 9675 30764 9717 30773
rect 9675 30724 9676 30764
rect 9716 30724 9717 30764
rect 9675 30715 9717 30724
rect 9579 29168 9621 29177
rect 9579 29128 9580 29168
rect 9620 29128 9621 29168
rect 9579 29119 9621 29128
rect 9484 28960 9620 29000
rect 9484 28160 9524 28169
rect 9484 27665 9524 28120
rect 9483 27656 9525 27665
rect 9483 27616 9484 27656
rect 9524 27616 9525 27656
rect 9483 27607 9525 27616
rect 9580 27488 9620 28960
rect 9676 27656 9716 30715
rect 9676 27607 9716 27616
rect 9772 29840 9812 33664
rect 9964 33209 10004 33664
rect 9963 33200 10005 33209
rect 9963 33160 9964 33200
rect 10004 33160 10005 33200
rect 9963 33151 10005 33160
rect 9964 32369 10004 33151
rect 9963 32360 10005 32369
rect 9963 32320 9964 32360
rect 10004 32320 10005 32360
rect 9963 32311 10005 32320
rect 9867 31352 9909 31361
rect 9867 31312 9868 31352
rect 9908 31312 9909 31352
rect 9867 31303 9909 31312
rect 9868 30680 9908 31303
rect 9963 31016 10005 31025
rect 9963 30976 9964 31016
rect 10004 30976 10005 31016
rect 9963 30967 10005 30976
rect 9868 30631 9908 30640
rect 9580 27448 9716 27488
rect 9579 26816 9621 26825
rect 9579 26776 9580 26816
rect 9620 26776 9621 26816
rect 9579 26767 9621 26776
rect 9580 26682 9620 26767
rect 9484 26144 9524 26153
rect 9484 25733 9524 26104
rect 9580 26144 9620 26153
rect 9483 25724 9525 25733
rect 9483 25684 9484 25724
rect 9524 25684 9525 25724
rect 9483 25675 9525 25684
rect 9388 24760 9524 24800
rect 9291 24751 9333 24760
rect 9004 24716 9044 24725
rect 9044 24676 9236 24716
rect 9004 24667 9044 24676
rect 9196 24632 9236 24676
rect 9196 24613 9332 24632
rect 9196 24592 9292 24613
rect 9292 24564 9332 24573
rect 9388 24613 9428 24622
rect 9388 24389 9428 24573
rect 9387 24380 9429 24389
rect 9387 24340 9388 24380
rect 9428 24340 9429 24380
rect 9387 24331 9429 24340
rect 8812 24004 8948 24044
rect 8812 23801 8852 24004
rect 9100 23960 9140 23969
rect 9484 23960 9524 24760
rect 8908 23920 9100 23960
rect 8716 23743 8756 23752
rect 8811 23792 8853 23801
rect 8811 23752 8812 23792
rect 8852 23752 8853 23792
rect 8811 23743 8853 23752
rect 8908 23792 8948 23920
rect 9100 23911 9140 23920
rect 9388 23920 9524 23960
rect 8908 23743 8948 23752
rect 9100 23792 9140 23803
rect 9100 23717 9140 23752
rect 9292 23792 9332 23801
rect 9099 23708 9141 23717
rect 9099 23668 9100 23708
rect 9140 23668 9141 23708
rect 9099 23659 9141 23668
rect 8811 23624 8853 23633
rect 8524 23584 8660 23624
rect 8427 23575 8469 23584
rect 8428 22877 8468 23575
rect 8524 23120 8564 23131
rect 8524 23045 8564 23080
rect 8523 23036 8565 23045
rect 8523 22996 8524 23036
rect 8564 22996 8565 23036
rect 8523 22987 8565 22996
rect 8427 22868 8469 22877
rect 8427 22828 8428 22868
rect 8468 22828 8469 22868
rect 8427 22819 8469 22828
rect 8523 22616 8565 22625
rect 8523 22576 8524 22616
rect 8564 22576 8565 22616
rect 8523 22567 8565 22576
rect 8332 22483 8372 22492
rect 8140 22231 8180 22240
rect 8331 22280 8373 22289
rect 8331 22240 8332 22280
rect 8372 22240 8373 22280
rect 8331 22231 8373 22240
rect 8332 22146 8372 22231
rect 7948 21988 8468 22028
rect 7756 21904 8372 21944
rect 7660 21820 7892 21860
rect 7563 21811 7605 21820
rect 7372 21608 7412 21811
rect 7659 21692 7701 21701
rect 7372 21559 7412 21568
rect 7564 21652 7660 21692
rect 7700 21652 7701 21692
rect 7564 21608 7604 21652
rect 7659 21643 7701 21652
rect 7564 21559 7604 21568
rect 7852 21524 7892 21820
rect 7947 21692 7989 21701
rect 7947 21652 7948 21692
rect 7988 21652 7989 21692
rect 7947 21643 7989 21652
rect 7660 21484 7892 21524
rect 7563 21440 7605 21449
rect 7563 21400 7564 21440
rect 7604 21400 7605 21440
rect 7563 21391 7605 21400
rect 7180 21148 7316 21188
rect 7083 20936 7125 20945
rect 7083 20896 7084 20936
rect 7124 20896 7125 20936
rect 7083 20887 7125 20896
rect 6987 20852 7029 20861
rect 6987 20812 6988 20852
rect 7028 20812 7029 20852
rect 6987 20803 7029 20812
rect 6987 20600 7029 20609
rect 6987 20560 6988 20600
rect 7028 20560 7029 20600
rect 6987 20551 7029 20560
rect 6988 20466 7028 20551
rect 7084 20096 7124 20105
rect 7084 19769 7124 20056
rect 7083 19760 7125 19769
rect 7083 19720 7084 19760
rect 7124 19720 7125 19760
rect 7083 19711 7125 19720
rect 6987 19256 7029 19265
rect 6987 19216 6988 19256
rect 7028 19216 7029 19256
rect 6987 19207 7029 19216
rect 6988 19122 7028 19207
rect 7180 18929 7220 21148
rect 7371 21104 7413 21113
rect 7371 21064 7372 21104
rect 7412 21064 7413 21104
rect 7371 21055 7413 21064
rect 7276 20768 7316 20777
rect 7276 20609 7316 20728
rect 7372 20768 7412 21055
rect 7372 20719 7412 20728
rect 7275 20600 7317 20609
rect 7275 20560 7276 20600
rect 7316 20560 7317 20600
rect 7275 20551 7317 20560
rect 7564 20180 7604 21391
rect 7660 20684 7700 21484
rect 7755 21272 7797 21281
rect 7755 21232 7756 21272
rect 7796 21232 7797 21272
rect 7755 21223 7797 21232
rect 7756 20852 7796 21223
rect 7756 20803 7796 20812
rect 7851 20852 7893 20861
rect 7851 20812 7852 20852
rect 7892 20812 7893 20852
rect 7851 20803 7893 20812
rect 7852 20718 7892 20803
rect 7660 20644 7796 20684
rect 7564 20140 7700 20180
rect 7467 20096 7509 20105
rect 7467 20056 7468 20096
rect 7508 20056 7509 20096
rect 7467 20047 7509 20056
rect 7468 19962 7508 20047
rect 7563 20012 7605 20021
rect 7563 19972 7564 20012
rect 7604 19972 7605 20012
rect 7563 19963 7605 19972
rect 7276 19844 7316 19853
rect 7316 19804 7508 19844
rect 7276 19795 7316 19804
rect 7371 19340 7413 19349
rect 7371 19300 7372 19340
rect 7412 19300 7413 19340
rect 7371 19291 7413 19300
rect 7179 18920 7221 18929
rect 7179 18880 7180 18920
rect 7220 18880 7221 18920
rect 7179 18871 7221 18880
rect 6892 18712 7220 18752
rect 6795 18703 6837 18712
rect 6795 18584 6837 18593
rect 6795 18544 6796 18584
rect 6836 18544 6837 18584
rect 6795 18535 6837 18544
rect 7083 18584 7125 18593
rect 7083 18544 7084 18584
rect 7124 18544 7125 18584
rect 7083 18535 7125 18544
rect 6604 18292 6740 18332
rect 6412 16316 6452 16325
rect 6316 16232 6356 16241
rect 6316 16157 6356 16192
rect 6315 16148 6357 16157
rect 6315 16108 6316 16148
rect 6356 16108 6357 16148
rect 6315 16099 6357 16108
rect 6316 16097 6356 16099
rect 6412 15989 6452 16276
rect 6507 16316 6549 16325
rect 6507 16276 6508 16316
rect 6548 16276 6549 16316
rect 6507 16267 6549 16276
rect 6508 16157 6548 16267
rect 6507 16148 6549 16157
rect 6507 16108 6508 16148
rect 6548 16108 6549 16148
rect 6507 16099 6549 16108
rect 6411 15980 6453 15989
rect 6411 15940 6412 15980
rect 6452 15940 6453 15980
rect 6411 15931 6453 15940
rect 6508 15560 6548 15569
rect 6219 14804 6261 14813
rect 6219 14764 6220 14804
rect 6260 14764 6261 14804
rect 6219 14755 6261 14764
rect 6220 13301 6260 14755
rect 6508 14057 6548 15520
rect 6507 14048 6549 14057
rect 6507 14008 6508 14048
rect 6548 14008 6549 14048
rect 6507 13999 6549 14008
rect 6219 13292 6261 13301
rect 6219 13252 6220 13292
rect 6260 13252 6261 13292
rect 6219 13243 6261 13252
rect 6507 13292 6549 13301
rect 6507 13252 6508 13292
rect 6548 13252 6549 13292
rect 6507 13243 6549 13252
rect 6124 13213 6164 13222
rect 6027 12872 6069 12881
rect 6027 12832 6028 12872
rect 6068 12832 6069 12872
rect 6027 12823 6069 12832
rect 6028 12704 6068 12713
rect 6124 12704 6164 13173
rect 6316 13040 6356 13049
rect 6219 12872 6261 12881
rect 6219 12832 6220 12872
rect 6260 12832 6261 12872
rect 6219 12823 6261 12832
rect 6068 12664 6164 12704
rect 6028 12655 6068 12664
rect 5836 12487 5876 12496
rect 6220 12536 6260 12823
rect 6316 12797 6356 13000
rect 6315 12788 6357 12797
rect 6315 12748 6316 12788
rect 6356 12748 6357 12788
rect 6315 12739 6357 12748
rect 4971 11864 5013 11873
rect 4971 11824 4972 11864
rect 5012 11824 5013 11864
rect 4971 11815 5013 11824
rect 5643 11864 5685 11873
rect 5643 11824 5644 11864
rect 5684 11824 5685 11864
rect 5643 11815 5685 11824
rect 4972 11696 5012 11815
rect 5836 11738 5876 11747
rect 5500 11705 5540 11714
rect 5836 11696 5876 11698
rect 5540 11665 5588 11696
rect 5500 11656 5588 11665
rect 4972 11647 5012 11656
rect 4107 11488 4108 11528
rect 4148 11488 4149 11528
rect 4107 11479 4149 11488
rect 4300 11488 4820 11528
rect 4011 11192 4053 11201
rect 4011 11152 4012 11192
rect 4052 11152 4053 11192
rect 4011 11143 4053 11152
rect 3340 10975 3380 10984
rect 3435 11024 3477 11033
rect 3435 10984 3436 11024
rect 3476 10984 3477 11024
rect 3435 10975 3477 10984
rect 3532 10772 3572 10781
rect 3532 10436 3572 10732
rect 3688 10604 4056 10613
rect 3728 10564 3770 10604
rect 3810 10564 3852 10604
rect 3892 10564 3934 10604
rect 3974 10564 4016 10604
rect 3688 10555 4056 10564
rect 4108 10436 4148 11479
rect 4300 11024 4340 11488
rect 5548 11444 5588 11656
rect 5644 11621 5684 11665
rect 5836 11656 6068 11696
rect 5643 11612 5685 11621
rect 5643 11572 5644 11612
rect 5684 11572 5685 11612
rect 5643 11570 5685 11572
rect 5643 11563 5644 11570
rect 5684 11563 5685 11570
rect 5644 11521 5684 11530
rect 5931 11528 5973 11537
rect 5931 11488 5932 11528
rect 5972 11488 5973 11528
rect 5931 11479 5973 11488
rect 5548 11404 5684 11444
rect 4683 11360 4725 11369
rect 4683 11320 4684 11360
rect 4724 11320 4725 11360
rect 4683 11311 4725 11320
rect 4928 11360 5296 11369
rect 4968 11320 5010 11360
rect 5050 11320 5092 11360
rect 5132 11320 5174 11360
rect 5214 11320 5256 11360
rect 4928 11311 5296 11320
rect 4340 10984 4628 11024
rect 4300 10975 4340 10984
rect 3532 10396 3860 10436
rect 3244 10352 3284 10361
rect 3284 10312 3572 10352
rect 3244 10303 3284 10312
rect 3436 10184 3476 10193
rect 3243 9680 3285 9689
rect 3243 9640 3244 9680
rect 3284 9640 3285 9680
rect 3243 9631 3285 9640
rect 3340 9680 3380 9689
rect 3436 9680 3476 10144
rect 3380 9640 3476 9680
rect 3532 10184 3572 10312
rect 3820 10193 3860 10396
rect 3977 10396 4148 10436
rect 3977 10199 4017 10396
rect 4395 10352 4437 10361
rect 3340 9631 3380 9640
rect 3244 9521 3284 9631
rect 3243 9512 3285 9521
rect 3243 9472 3244 9512
rect 3284 9472 3285 9512
rect 3243 9463 3285 9472
rect 3435 9512 3477 9521
rect 3435 9472 3436 9512
rect 3476 9472 3477 9512
rect 3435 9463 3477 9472
rect 3532 9512 3572 10144
rect 3724 10184 3764 10193
rect 3724 10025 3764 10144
rect 3819 10184 3861 10193
rect 3819 10144 3820 10184
rect 3860 10144 3861 10184
rect 4300 10312 4396 10352
rect 4436 10312 4437 10352
rect 4203 10184 4245 10193
rect 4017 10159 4052 10184
rect 3977 10144 4052 10159
rect 3819 10135 3861 10144
rect 3532 9463 3572 9472
rect 3628 10016 3668 10025
rect 3244 9378 3284 9463
rect 3436 9378 3476 9463
rect 3628 9260 3668 9976
rect 3723 10016 3765 10025
rect 3723 9976 3724 10016
rect 3764 9976 3765 10016
rect 3723 9967 3765 9976
rect 3820 9521 3860 10135
rect 4012 9605 4052 10144
rect 4203 10144 4204 10184
rect 4244 10144 4245 10184
rect 4203 10135 4245 10144
rect 4300 10184 4340 10312
rect 4395 10303 4437 10312
rect 4204 10050 4244 10135
rect 4300 9932 4340 10144
rect 4491 10016 4533 10025
rect 4491 9976 4492 10016
rect 4532 9976 4533 10016
rect 4491 9967 4533 9976
rect 4204 9892 4340 9932
rect 4107 9764 4149 9773
rect 4107 9724 4108 9764
rect 4148 9724 4149 9764
rect 4107 9715 4149 9724
rect 4011 9596 4053 9605
rect 4011 9556 4012 9596
rect 4052 9556 4053 9596
rect 4011 9547 4053 9556
rect 3819 9512 3861 9521
rect 3819 9472 3820 9512
rect 3860 9472 3861 9512
rect 3819 9463 3861 9472
rect 3532 9220 3668 9260
rect 4012 9260 4052 9547
rect 4108 9512 4148 9715
rect 4108 9463 4148 9472
rect 4012 9220 4148 9260
rect 3532 8924 3572 9220
rect 3688 9092 4056 9101
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 3688 9043 4056 9052
rect 4108 8924 4148 9220
rect 4204 9185 4244 9892
rect 4492 9882 4532 9967
rect 4588 9857 4628 10984
rect 4684 10184 4724 11311
rect 5355 11276 5397 11285
rect 5355 11236 5356 11276
rect 5396 11236 5397 11276
rect 5355 11227 5397 11236
rect 4779 11192 4821 11201
rect 4779 11152 4780 11192
rect 4820 11152 4821 11192
rect 4779 11143 4821 11152
rect 4684 10109 4724 10144
rect 4683 10100 4725 10109
rect 4683 10060 4684 10100
rect 4724 10060 4725 10100
rect 4683 10051 4725 10060
rect 4587 9848 4629 9857
rect 4587 9808 4588 9848
rect 4628 9808 4629 9848
rect 4587 9799 4629 9808
rect 4780 9689 4820 11143
rect 4928 9848 5296 9857
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 4928 9799 5296 9808
rect 4779 9680 4821 9689
rect 4396 9640 4724 9680
rect 4299 9512 4341 9521
rect 4299 9472 4300 9512
rect 4340 9472 4341 9512
rect 4299 9463 4341 9472
rect 4396 9512 4436 9640
rect 4588 9512 4628 9521
rect 4396 9463 4436 9472
rect 4492 9472 4588 9512
rect 4300 9378 4340 9463
rect 4396 9344 4436 9353
rect 4492 9344 4532 9472
rect 4588 9463 4628 9472
rect 4684 9512 4724 9640
rect 4779 9640 4780 9680
rect 4820 9640 4821 9680
rect 4779 9631 4821 9640
rect 5072 9596 5114 9605
rect 5072 9556 5073 9596
rect 5113 9556 5114 9596
rect 5072 9547 5114 9556
rect 4876 9512 4916 9521
rect 4436 9304 4532 9344
rect 4396 9295 4436 9304
rect 4588 9260 4628 9269
rect 4203 9176 4245 9185
rect 4203 9136 4204 9176
rect 4244 9136 4245 9176
rect 4203 9127 4245 9136
rect 3532 8884 3668 8924
rect 3468 8681 3508 8766
rect 3244 8672 3284 8681
rect 3244 8513 3284 8632
rect 3339 8672 3381 8681
rect 3339 8632 3340 8672
rect 3380 8632 3381 8672
rect 3339 8623 3381 8632
rect 3467 8672 3509 8681
rect 3467 8632 3468 8672
rect 3508 8632 3509 8672
rect 3467 8623 3509 8632
rect 3340 8538 3380 8623
rect 3243 8504 3285 8513
rect 3243 8464 3244 8504
rect 3284 8464 3285 8504
rect 3243 8455 3285 8464
rect 3436 8504 3476 8513
rect 3436 8084 3476 8464
rect 3628 8168 3668 8884
rect 4012 8884 4148 8924
rect 3723 8840 3765 8849
rect 3723 8800 3724 8840
rect 3764 8800 3765 8840
rect 3723 8791 3765 8800
rect 3724 8706 3764 8791
rect 3916 8756 3956 8765
rect 3916 8429 3956 8716
rect 4012 8681 4052 8884
rect 4107 8756 4149 8765
rect 4107 8716 4108 8756
rect 4148 8716 4149 8756
rect 4107 8707 4149 8716
rect 4011 8672 4053 8681
rect 4011 8632 4012 8672
rect 4052 8632 4053 8672
rect 4011 8623 4053 8632
rect 4108 8672 4148 8707
rect 3915 8420 3957 8429
rect 3915 8380 3916 8420
rect 3956 8380 3957 8420
rect 3915 8371 3957 8380
rect 3340 8044 3476 8084
rect 3532 8128 3668 8168
rect 3243 7832 3285 7841
rect 3243 7792 3244 7832
rect 3284 7792 3285 7832
rect 3243 7783 3285 7792
rect 3244 7698 3284 7783
rect 3340 7412 3380 8044
rect 3435 7916 3477 7925
rect 3435 7876 3436 7916
rect 3476 7876 3477 7916
rect 3435 7867 3477 7876
rect 3436 7782 3476 7867
rect 3052 7120 3188 7160
rect 3244 7372 3380 7412
rect 3052 6859 3092 7120
rect 3148 6992 3188 7001
rect 2091 6824 2133 6833
rect 2091 6784 2092 6824
rect 2132 6784 2133 6824
rect 2091 6775 2133 6784
rect 2667 6824 2709 6833
rect 2667 6784 2668 6824
rect 2708 6784 2709 6824
rect 2667 6775 2709 6784
rect 2859 6824 2901 6833
rect 2859 6784 2860 6824
rect 2900 6784 2901 6824
rect 2859 6775 2901 6784
rect 2092 6488 2132 6775
rect 3052 6749 3097 6859
rect 2283 6740 2325 6749
rect 2283 6700 2284 6740
rect 2324 6700 2325 6740
rect 2283 6691 2325 6700
rect 2955 6740 2997 6749
rect 2955 6700 2956 6740
rect 2996 6700 2997 6740
rect 2955 6691 2997 6700
rect 3052 6740 3098 6749
rect 3052 6700 3057 6740
rect 3097 6700 3098 6740
rect 3052 6691 3098 6700
rect 2187 6572 2229 6581
rect 2187 6532 2188 6572
rect 2228 6532 2229 6572
rect 2187 6523 2229 6532
rect 2092 6439 2132 6448
rect 2188 6438 2228 6523
rect 2284 6488 2324 6691
rect 2284 6439 2324 6448
rect 2380 6488 2420 6499
rect 2572 6497 2612 6582
rect 2380 6413 2420 6448
rect 2571 6488 2613 6497
rect 2571 6448 2572 6488
rect 2612 6448 2613 6488
rect 2571 6439 2613 6448
rect 2668 6488 2708 6497
rect 2860 6488 2900 6497
rect 2668 6413 2708 6448
rect 2764 6448 2860 6488
rect 2379 6404 2421 6413
rect 2379 6364 2380 6404
rect 2420 6364 2421 6404
rect 2379 6355 2421 6364
rect 2667 6404 2709 6413
rect 2667 6364 2668 6404
rect 2708 6364 2709 6404
rect 2667 6355 2709 6364
rect 1996 6280 2132 6320
rect 1899 5480 1941 5489
rect 1899 5440 1900 5480
rect 1940 5440 1941 5480
rect 1899 5431 1941 5440
rect 1460 4936 1844 4976
rect 1420 4927 1460 4936
rect 1803 4808 1845 4817
rect 1324 4768 1556 4808
rect 1228 4684 1364 4724
rect 1131 1196 1173 1205
rect 1131 1156 1132 1196
rect 1172 1156 1173 1196
rect 1131 1147 1173 1156
rect 1324 701 1364 4684
rect 1419 4472 1461 4481
rect 1419 4432 1420 4472
rect 1460 4432 1461 4472
rect 1419 4423 1461 4432
rect 1420 3632 1460 4423
rect 1516 4388 1556 4768
rect 1803 4768 1804 4808
rect 1844 4768 1845 4808
rect 1803 4759 1845 4768
rect 1707 4640 1749 4649
rect 1707 4600 1708 4640
rect 1748 4600 1749 4640
rect 1707 4591 1749 4600
rect 1516 4339 1556 4348
rect 1708 4220 1748 4591
rect 1708 4171 1748 4180
rect 1516 3632 1556 3641
rect 1420 3592 1516 3632
rect 1804 3632 1844 4759
rect 1900 4388 1940 5431
rect 1900 4339 1940 4348
rect 1995 4388 2037 4397
rect 1995 4348 1996 4388
rect 2036 4348 2037 4388
rect 1995 4339 2037 4348
rect 1900 3632 1940 3641
rect 1804 3592 1900 3632
rect 1516 3583 1556 3592
rect 1900 3583 1940 3592
rect 1419 3464 1461 3473
rect 1419 3424 1420 3464
rect 1460 3424 1461 3464
rect 1419 3415 1461 3424
rect 1420 2876 1460 3415
rect 1708 3380 1748 3389
rect 1611 3296 1653 3305
rect 1611 3256 1612 3296
rect 1652 3256 1653 3296
rect 1611 3247 1653 3256
rect 1516 2876 1556 2885
rect 1420 2836 1516 2876
rect 1516 2827 1556 2836
rect 1612 2708 1652 3247
rect 1708 3221 1748 3340
rect 1707 3212 1749 3221
rect 1707 3172 1708 3212
rect 1748 3172 1749 3212
rect 1707 3163 1749 3172
rect 1899 3044 1941 3053
rect 1899 3004 1900 3044
rect 1940 3004 1941 3044
rect 1899 2995 1941 3004
rect 1803 2960 1845 2969
rect 1803 2920 1804 2960
rect 1844 2920 1845 2960
rect 1803 2911 1845 2920
rect 1708 2708 1748 2717
rect 1612 2668 1708 2708
rect 1708 2659 1748 2668
rect 1611 2540 1653 2549
rect 1611 2500 1612 2540
rect 1652 2500 1653 2540
rect 1611 2491 1653 2500
rect 1515 1784 1557 1793
rect 1515 1744 1516 1784
rect 1556 1744 1557 1784
rect 1515 1735 1557 1744
rect 1516 1650 1556 1735
rect 1612 1196 1652 2491
rect 1708 1868 1748 1877
rect 1804 1868 1844 2911
rect 1900 2876 1940 2995
rect 1900 2827 1940 2836
rect 1996 2708 2036 4339
rect 2092 4220 2132 6280
rect 2572 6236 2612 6245
rect 2380 6196 2572 6236
rect 2187 5900 2229 5909
rect 2187 5860 2188 5900
rect 2228 5860 2229 5900
rect 2187 5851 2229 5860
rect 2092 4171 2132 4180
rect 2188 4052 2228 5851
rect 2283 5816 2325 5825
rect 2283 5776 2284 5816
rect 2324 5776 2325 5816
rect 2283 5767 2325 5776
rect 2284 4388 2324 5767
rect 2284 4339 2324 4348
rect 2283 4136 2325 4145
rect 2283 4096 2284 4136
rect 2324 4096 2325 4136
rect 2283 4087 2325 4096
rect 2092 4012 2228 4052
rect 2092 3380 2132 4012
rect 2284 3632 2324 4087
rect 2284 3583 2324 3592
rect 2283 3464 2325 3473
rect 2283 3424 2284 3464
rect 2324 3424 2325 3464
rect 2283 3415 2325 3424
rect 2092 3331 2132 3340
rect 2187 3380 2229 3389
rect 2187 3340 2188 3380
rect 2228 3340 2229 3380
rect 2187 3331 2229 3340
rect 2092 2708 2132 2717
rect 1996 2668 2092 2708
rect 2092 2659 2132 2668
rect 2091 2204 2133 2213
rect 2091 2164 2092 2204
rect 2132 2164 2133 2204
rect 2091 2155 2133 2164
rect 1899 2120 1941 2129
rect 1899 2080 1900 2120
rect 1940 2080 1941 2120
rect 1899 2071 1941 2080
rect 1900 1986 1940 2071
rect 1748 1828 1844 1868
rect 2092 1868 2132 2155
rect 1708 1819 1748 1828
rect 2092 1819 2132 1828
rect 1995 1784 2037 1793
rect 1995 1744 1996 1784
rect 2036 1744 2037 1784
rect 1995 1735 2037 1744
rect 1708 1196 1748 1205
rect 1612 1156 1708 1196
rect 1708 1147 1748 1156
rect 1515 1112 1557 1121
rect 1515 1072 1516 1112
rect 1556 1072 1557 1112
rect 1515 1063 1557 1072
rect 1516 944 1556 1063
rect 1803 1028 1845 1037
rect 1803 988 1804 1028
rect 1844 988 1845 1028
rect 1803 979 1845 988
rect 1516 895 1556 904
rect 1323 692 1365 701
rect 1323 652 1324 692
rect 1364 652 1365 692
rect 1323 643 1365 652
rect 1804 80 1844 979
rect 1900 944 1940 953
rect 1900 197 1940 904
rect 1899 188 1941 197
rect 1899 148 1900 188
rect 1940 148 1941 188
rect 1899 139 1941 148
rect 1996 80 2036 1735
rect 2092 1196 2132 1205
rect 2092 869 2132 1156
rect 2188 1112 2228 3331
rect 2284 2204 2324 3415
rect 2380 3380 2420 6196
rect 2572 6187 2612 6196
rect 2668 5900 2708 6355
rect 2572 5860 2708 5900
rect 2572 5321 2612 5860
rect 2668 5648 2708 5657
rect 2571 5312 2613 5321
rect 2571 5272 2572 5312
rect 2612 5272 2613 5312
rect 2571 5263 2613 5272
rect 2668 4976 2708 5608
rect 2668 4901 2708 4936
rect 2667 4892 2709 4901
rect 2667 4852 2668 4892
rect 2708 4852 2709 4892
rect 2667 4843 2709 4852
rect 2475 4220 2517 4229
rect 2475 4180 2476 4220
rect 2516 4180 2517 4220
rect 2475 4171 2517 4180
rect 2476 4086 2516 4171
rect 2475 3968 2517 3977
rect 2475 3928 2476 3968
rect 2516 3928 2517 3968
rect 2764 3968 2804 6448
rect 2860 6439 2900 6448
rect 2956 6488 2996 6691
rect 3052 6497 3092 6691
rect 3148 6665 3188 6952
rect 3147 6656 3189 6665
rect 3147 6616 3148 6656
rect 3188 6616 3189 6656
rect 3147 6607 3189 6616
rect 3244 6497 3284 7372
rect 3532 7328 3572 8128
rect 4108 8093 4148 8632
rect 4107 8084 4149 8093
rect 4107 8044 4108 8084
rect 4148 8044 4149 8084
rect 4107 8035 4149 8044
rect 3627 8000 3669 8009
rect 3627 7960 3628 8000
rect 3668 7960 3669 8000
rect 3627 7951 3669 7960
rect 3628 7866 3668 7951
rect 4588 7673 4628 9220
rect 4587 7664 4629 7673
rect 4587 7624 4588 7664
rect 4628 7624 4629 7664
rect 4587 7615 4629 7624
rect 3688 7580 4056 7589
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 3688 7531 4056 7540
rect 3436 7288 3572 7328
rect 3723 7328 3765 7337
rect 3723 7288 3724 7328
rect 3764 7288 3765 7328
rect 3339 7244 3381 7253
rect 3339 7204 3340 7244
rect 3380 7204 3381 7244
rect 3339 7195 3381 7204
rect 3340 7110 3380 7195
rect 3339 6824 3381 6833
rect 3339 6784 3340 6824
rect 3380 6784 3381 6824
rect 3339 6775 3381 6784
rect 3340 6581 3380 6775
rect 3339 6572 3381 6581
rect 3339 6532 3340 6572
rect 3380 6532 3381 6572
rect 3339 6523 3381 6532
rect 3052 6488 3097 6497
rect 3052 6448 3057 6488
rect 2956 6320 2996 6448
rect 3057 6439 3097 6448
rect 3243 6488 3285 6497
rect 3243 6448 3244 6488
rect 3284 6448 3285 6488
rect 3243 6439 3285 6448
rect 3340 6320 3380 6523
rect 2956 6280 3092 6320
rect 2860 5816 2900 5825
rect 3052 5816 3092 6280
rect 2900 5776 3092 5816
rect 2860 5767 2900 5776
rect 2955 5648 2997 5657
rect 2955 5608 2956 5648
rect 2996 5608 2997 5648
rect 2955 5599 2997 5608
rect 2859 5312 2901 5321
rect 2859 5272 2860 5312
rect 2900 5272 2901 5312
rect 2859 5263 2901 5272
rect 2860 5144 2900 5263
rect 2860 5095 2900 5104
rect 2860 3968 2900 3977
rect 2764 3928 2860 3968
rect 2475 3919 2517 3928
rect 2860 3919 2900 3928
rect 2476 3557 2516 3919
rect 2571 3884 2613 3893
rect 2571 3844 2572 3884
rect 2612 3844 2613 3884
rect 2571 3835 2613 3844
rect 2475 3548 2517 3557
rect 2475 3508 2476 3548
rect 2516 3508 2517 3548
rect 2475 3499 2517 3508
rect 2572 3464 2612 3835
rect 2667 3800 2709 3809
rect 2667 3760 2668 3800
rect 2708 3760 2709 3800
rect 2667 3751 2709 3760
rect 2668 3632 2708 3751
rect 2668 3583 2708 3592
rect 2572 3424 2708 3464
rect 2476 3380 2516 3389
rect 2380 3340 2476 3380
rect 2476 3331 2516 3340
rect 2571 3044 2613 3053
rect 2571 3004 2572 3044
rect 2612 3004 2613 3044
rect 2571 2995 2613 3004
rect 2572 2708 2612 2995
rect 2572 2659 2612 2668
rect 2668 2540 2708 3424
rect 2860 3380 2900 3389
rect 2956 3380 2996 5599
rect 3052 5480 3092 5776
rect 3148 6280 3380 6320
rect 3148 5648 3188 6280
rect 3436 6236 3476 7288
rect 3723 7279 3765 7288
rect 3531 7160 3573 7169
rect 3531 7120 3532 7160
rect 3572 7120 3573 7160
rect 3531 7111 3573 7120
rect 3532 7026 3572 7111
rect 3531 6488 3573 6497
rect 3531 6448 3532 6488
rect 3572 6448 3573 6488
rect 3531 6439 3573 6448
rect 3628 6488 3668 6497
rect 3724 6488 3764 7279
rect 4299 7244 4341 7253
rect 4299 7204 4300 7244
rect 4340 7204 4341 7244
rect 4299 7195 4341 7204
rect 4300 6656 4340 7195
rect 4684 6992 4724 9472
rect 4780 9472 4876 9512
rect 4780 7589 4820 9472
rect 4876 9463 4916 9472
rect 4971 9512 5013 9521
rect 4971 9472 4972 9512
rect 5012 9472 5013 9512
rect 4971 9463 5013 9472
rect 5073 9512 5113 9547
rect 4972 9378 5012 9463
rect 5073 9461 5113 9472
rect 5259 9512 5301 9521
rect 5259 9472 5260 9512
rect 5300 9472 5301 9512
rect 5259 9463 5301 9472
rect 5260 8504 5300 9463
rect 5356 8681 5396 11227
rect 5644 11192 5684 11404
rect 5740 11192 5780 11201
rect 5644 11152 5740 11192
rect 5740 11143 5780 11152
rect 5547 11024 5589 11033
rect 5547 10984 5548 11024
rect 5588 10984 5589 11024
rect 5547 10975 5589 10984
rect 5451 10352 5493 10361
rect 5451 10312 5452 10352
rect 5492 10312 5493 10352
rect 5451 10303 5493 10312
rect 5355 8672 5397 8681
rect 5355 8632 5356 8672
rect 5396 8632 5397 8672
rect 5355 8623 5397 8632
rect 5260 8464 5396 8504
rect 4928 8336 5296 8345
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 4928 8287 5296 8296
rect 5068 8168 5108 8177
rect 5356 8168 5396 8464
rect 5108 8128 5396 8168
rect 5068 8119 5108 8128
rect 4875 8084 4917 8093
rect 4875 8044 4876 8084
rect 4916 8044 4917 8084
rect 4875 8035 4917 8044
rect 4876 8000 4916 8035
rect 4779 7580 4821 7589
rect 4779 7540 4780 7580
rect 4820 7540 4821 7580
rect 4779 7531 4821 7540
rect 4780 7160 4820 7169
rect 4876 7160 4916 7960
rect 4820 7120 4916 7160
rect 5164 7160 5204 8128
rect 5260 8000 5300 8009
rect 5260 7841 5300 7960
rect 5259 7832 5301 7841
rect 5259 7792 5260 7832
rect 5300 7792 5301 7832
rect 5259 7783 5301 7792
rect 5452 7748 5492 10303
rect 5548 10193 5588 10975
rect 5932 10352 5972 11479
rect 6028 11453 6068 11656
rect 6220 11537 6260 12496
rect 6315 12032 6357 12041
rect 6315 11992 6316 12032
rect 6356 11992 6357 12032
rect 6315 11983 6357 11992
rect 6219 11528 6261 11537
rect 6219 11488 6220 11528
rect 6260 11488 6261 11528
rect 6219 11479 6261 11488
rect 6027 11444 6069 11453
rect 6027 11404 6028 11444
rect 6068 11404 6069 11444
rect 6027 11395 6069 11404
rect 6123 11276 6165 11285
rect 6123 11236 6124 11276
rect 6164 11236 6165 11276
rect 6123 11227 6165 11236
rect 6028 11024 6068 11033
rect 6028 10436 6068 10984
rect 6124 11024 6164 11227
rect 6124 10697 6164 10984
rect 6316 10781 6356 11983
rect 6411 11276 6453 11285
rect 6411 11236 6412 11276
rect 6452 11236 6453 11276
rect 6411 11227 6453 11236
rect 6315 10772 6357 10781
rect 6315 10732 6316 10772
rect 6356 10732 6357 10772
rect 6315 10723 6357 10732
rect 6123 10688 6165 10697
rect 6123 10648 6124 10688
rect 6164 10648 6165 10688
rect 6123 10639 6165 10648
rect 6124 10436 6164 10445
rect 6028 10396 6124 10436
rect 6124 10387 6164 10396
rect 6412 10361 6452 11227
rect 6508 11024 6548 13243
rect 6604 11108 6644 18292
rect 6796 16064 6836 18535
rect 7084 18341 7124 18535
rect 7083 18332 7125 18341
rect 7083 18292 7084 18332
rect 7124 18292 7125 18332
rect 7083 18283 7125 18292
rect 6891 17996 6933 18005
rect 7083 17996 7125 18005
rect 6891 17956 6892 17996
rect 6932 17956 7028 17996
rect 6891 17947 6933 17956
rect 6892 17744 6932 17755
rect 6892 17081 6932 17704
rect 6891 17072 6933 17081
rect 6891 17032 6892 17072
rect 6932 17032 6933 17072
rect 6891 17023 6933 17032
rect 6891 16820 6933 16829
rect 6891 16780 6892 16820
rect 6932 16780 6933 16820
rect 6891 16771 6933 16780
rect 6892 16232 6932 16771
rect 6988 16316 7028 17956
rect 7083 17956 7084 17996
rect 7124 17956 7125 17996
rect 7083 17947 7125 17956
rect 7084 17862 7124 17947
rect 6988 16276 7124 16316
rect 6892 16183 6932 16192
rect 7084 16157 7124 16276
rect 7083 16148 7125 16157
rect 7083 16108 7084 16148
rect 7124 16108 7125 16148
rect 7083 16099 7125 16108
rect 6796 16024 6932 16064
rect 6699 15392 6741 15401
rect 6699 15352 6700 15392
rect 6740 15352 6741 15392
rect 6699 15343 6741 15352
rect 6700 15258 6740 15343
rect 6795 15224 6837 15233
rect 6795 15184 6796 15224
rect 6836 15184 6837 15224
rect 6795 15175 6837 15184
rect 6699 14552 6741 14561
rect 6699 14512 6700 14552
rect 6740 14512 6741 14552
rect 6699 14503 6741 14512
rect 6700 11285 6740 14503
rect 6796 13124 6836 15175
rect 6796 13075 6836 13084
rect 6892 11360 6932 16024
rect 6988 15560 7028 15569
rect 6988 15401 7028 15520
rect 7084 15560 7124 16099
rect 7084 15511 7124 15520
rect 6987 15392 7029 15401
rect 6987 15352 6988 15392
rect 7028 15352 7029 15392
rect 6987 15343 7029 15352
rect 7083 13880 7125 13889
rect 7083 13840 7084 13880
rect 7124 13840 7125 13880
rect 7083 13831 7125 13840
rect 6988 13213 7028 13222
rect 6988 12629 7028 13173
rect 6987 12620 7029 12629
rect 6987 12580 6988 12620
rect 7028 12580 7029 12620
rect 6987 12571 7029 12580
rect 7084 12461 7124 13831
rect 7083 12452 7125 12461
rect 6988 12412 7084 12452
rect 7124 12412 7125 12452
rect 6988 11621 7028 12412
rect 7083 12403 7125 12412
rect 7083 11948 7125 11957
rect 7083 11908 7084 11948
rect 7124 11908 7125 11948
rect 7083 11899 7125 11908
rect 7084 11696 7124 11899
rect 7084 11647 7124 11656
rect 6987 11612 7029 11621
rect 6987 11572 6988 11612
rect 7028 11572 7029 11612
rect 6987 11563 7029 11572
rect 6796 11320 6932 11360
rect 6699 11276 6741 11285
rect 6699 11236 6700 11276
rect 6740 11236 6741 11276
rect 6699 11227 6741 11236
rect 6604 11068 6740 11108
rect 6508 10975 6548 10984
rect 6604 10940 6644 10949
rect 6604 10781 6644 10900
rect 6603 10772 6645 10781
rect 6603 10732 6604 10772
rect 6644 10732 6645 10772
rect 6603 10723 6645 10732
rect 6507 10604 6549 10613
rect 6507 10564 6508 10604
rect 6548 10564 6549 10604
rect 6507 10555 6549 10564
rect 6411 10352 6453 10361
rect 5932 10312 6068 10352
rect 5547 10184 5589 10193
rect 5547 10144 5548 10184
rect 5588 10144 5589 10184
rect 5547 10135 5589 10144
rect 5931 10184 5973 10193
rect 5931 10144 5932 10184
rect 5972 10144 5973 10184
rect 5931 10135 5973 10144
rect 5932 10050 5972 10135
rect 6028 9941 6068 10312
rect 6411 10312 6412 10352
rect 6452 10312 6453 10352
rect 6411 10303 6453 10312
rect 6027 9932 6069 9941
rect 6027 9892 6028 9932
rect 6068 9892 6069 9932
rect 6027 9883 6069 9892
rect 6315 9932 6357 9941
rect 6315 9892 6316 9932
rect 6356 9892 6357 9932
rect 6315 9883 6357 9892
rect 5835 9680 5877 9689
rect 5835 9640 5836 9680
rect 5876 9640 5877 9680
rect 5835 9631 5877 9640
rect 5547 8588 5589 8597
rect 5547 8548 5548 8588
rect 5588 8548 5589 8588
rect 5547 8539 5589 8548
rect 5548 8454 5588 8539
rect 5740 8504 5780 8513
rect 5740 7925 5780 8464
rect 5739 7916 5781 7925
rect 5739 7876 5740 7916
rect 5780 7876 5781 7916
rect 5739 7867 5781 7876
rect 5356 7708 5492 7748
rect 4780 7111 4820 7120
rect 5164 7111 5204 7120
rect 5260 7160 5300 7169
rect 5356 7160 5396 7708
rect 5451 7580 5493 7589
rect 5451 7540 5452 7580
rect 5492 7540 5493 7580
rect 5451 7531 5493 7540
rect 5300 7120 5396 7160
rect 5260 7111 5300 7120
rect 4972 6992 5012 7001
rect 4684 6952 4972 6992
rect 4972 6943 5012 6952
rect 5452 6992 5492 7531
rect 5739 7160 5781 7169
rect 5836 7160 5876 9631
rect 6316 9512 6356 9883
rect 6316 9463 6356 9472
rect 5932 8677 5972 8686
rect 5932 8177 5972 8637
rect 6412 8672 6452 10303
rect 6412 8623 6452 8632
rect 5931 8168 5973 8177
rect 6508 8168 6548 10555
rect 6604 8681 6644 10723
rect 6603 8672 6645 8681
rect 6603 8632 6604 8672
rect 6644 8632 6645 8672
rect 6603 8623 6645 8632
rect 5931 8128 5932 8168
rect 5972 8128 5973 8168
rect 5931 8119 5973 8128
rect 6412 8128 6548 8168
rect 6027 7832 6069 7841
rect 6027 7792 6028 7832
rect 6068 7792 6069 7832
rect 6027 7783 6069 7792
rect 5739 7120 5740 7160
rect 5780 7120 5876 7160
rect 5739 7111 5781 7120
rect 5547 7076 5589 7085
rect 5547 7036 5548 7076
rect 5588 7036 5589 7076
rect 5547 7027 5589 7036
rect 5452 6943 5492 6952
rect 4928 6824 5296 6833
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 4928 6775 5296 6784
rect 4592 6740 4634 6749
rect 4592 6700 4593 6740
rect 4633 6700 4634 6740
rect 4592 6691 4634 6700
rect 3916 6616 4244 6656
rect 3668 6448 3764 6488
rect 3819 6488 3861 6497
rect 3819 6448 3820 6488
rect 3860 6448 3861 6488
rect 3628 6439 3668 6448
rect 3819 6439 3861 6448
rect 3916 6488 3956 6616
rect 4108 6488 4148 6497
rect 3916 6439 3956 6448
rect 4012 6448 4108 6488
rect 3148 5599 3188 5608
rect 3244 6196 3476 6236
rect 3052 5440 3188 5480
rect 3051 5144 3093 5153
rect 3051 5104 3052 5144
rect 3092 5104 3093 5144
rect 3051 5095 3093 5104
rect 3052 4808 3092 5095
rect 3052 4759 3092 4768
rect 3051 4640 3093 4649
rect 3051 4600 3052 4640
rect 3092 4600 3093 4640
rect 3051 4591 3093 4600
rect 3052 4136 3092 4591
rect 3052 4087 3092 4096
rect 3148 4136 3188 5440
rect 3244 4892 3284 6196
rect 3244 4843 3284 4852
rect 3436 4976 3476 4985
rect 3436 4817 3476 4936
rect 3435 4808 3477 4817
rect 3435 4768 3436 4808
rect 3476 4768 3477 4808
rect 3435 4759 3477 4768
rect 3243 4640 3285 4649
rect 3243 4600 3244 4640
rect 3284 4600 3285 4640
rect 3243 4591 3285 4600
rect 3148 4087 3188 4096
rect 3147 3968 3189 3977
rect 3147 3928 3148 3968
rect 3188 3928 3189 3968
rect 3147 3919 3189 3928
rect 2900 3340 2996 3380
rect 2860 3331 2900 3340
rect 3052 3212 3092 3221
rect 2955 3128 2997 3137
rect 2955 3088 2956 3128
rect 2996 3088 2997 3128
rect 2955 3079 2997 3088
rect 2859 2624 2901 2633
rect 2859 2584 2860 2624
rect 2900 2584 2901 2624
rect 2859 2575 2901 2584
rect 2572 2500 2708 2540
rect 2379 2456 2421 2465
rect 2379 2416 2380 2456
rect 2420 2416 2421 2456
rect 2379 2407 2421 2416
rect 2380 2322 2420 2407
rect 2284 2164 2420 2204
rect 2284 1700 2324 1709
rect 2284 1457 2324 1660
rect 2283 1448 2325 1457
rect 2283 1408 2284 1448
rect 2324 1408 2325 1448
rect 2283 1399 2325 1408
rect 2380 1196 2420 2164
rect 2475 1868 2517 1877
rect 2475 1828 2476 1868
rect 2516 1828 2517 1868
rect 2475 1819 2517 1828
rect 2476 1734 2516 1819
rect 2476 1196 2516 1205
rect 2380 1156 2476 1196
rect 2476 1147 2516 1156
rect 2188 1072 2420 1112
rect 2284 944 2324 953
rect 2091 860 2133 869
rect 2091 820 2092 860
rect 2132 820 2133 860
rect 2091 811 2133 820
rect 2284 785 2324 904
rect 2283 776 2325 785
rect 2283 736 2284 776
rect 2324 736 2325 776
rect 2283 727 2325 736
rect 2187 692 2229 701
rect 2187 652 2188 692
rect 2228 652 2229 692
rect 2187 643 2229 652
rect 2188 80 2228 643
rect 2380 80 2420 1072
rect 2572 80 2612 2500
rect 2860 2036 2900 2575
rect 2764 1996 2900 2036
rect 2668 1700 2708 1709
rect 2668 449 2708 1660
rect 2667 440 2709 449
rect 2667 400 2668 440
rect 2708 400 2709 440
rect 2667 391 2709 400
rect 2764 80 2804 1996
rect 2860 1868 2900 1877
rect 2956 1868 2996 3079
rect 3052 2801 3092 3172
rect 3051 2792 3093 2801
rect 3051 2752 3052 2792
rect 3092 2752 3093 2792
rect 3051 2743 3093 2752
rect 2900 1828 2996 1868
rect 3148 1868 3188 3919
rect 3244 3380 3284 4591
rect 3435 4136 3477 4145
rect 3435 4096 3436 4136
rect 3476 4096 3477 4136
rect 3435 4087 3477 4096
rect 3244 3331 3284 3340
rect 3243 2876 3285 2885
rect 3243 2836 3244 2876
rect 3284 2836 3285 2876
rect 3243 2827 3285 2836
rect 2860 1819 2900 1828
rect 3148 1819 3188 1828
rect 3147 1280 3189 1289
rect 3147 1240 3148 1280
rect 3188 1240 3189 1280
rect 3244 1280 3284 2827
rect 3436 1952 3476 4087
rect 3532 3053 3572 6439
rect 3820 6354 3860 6439
rect 3916 6320 3956 6329
rect 4012 6320 4052 6448
rect 4108 6439 4148 6448
rect 4204 6488 4244 6616
rect 4300 6607 4340 6616
rect 3956 6280 4052 6320
rect 3916 6271 3956 6280
rect 3688 6068 4056 6077
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 3688 6019 4056 6028
rect 4204 5900 4244 6448
rect 4396 6488 4436 6497
rect 4396 6077 4436 6448
rect 4491 6488 4533 6497
rect 4491 6448 4492 6488
rect 4532 6448 4533 6488
rect 4491 6439 4533 6448
rect 4593 6488 4633 6691
rect 4875 6572 4917 6581
rect 4875 6532 4876 6572
rect 4916 6532 4917 6572
rect 4875 6523 4917 6532
rect 4593 6439 4633 6448
rect 4876 6488 4916 6523
rect 4395 6068 4437 6077
rect 4395 6028 4396 6068
rect 4436 6028 4437 6068
rect 4492 6068 4532 6439
rect 4876 6437 4916 6448
rect 5355 6068 5397 6077
rect 4492 6028 4724 6068
rect 4395 6019 4437 6028
rect 4588 5900 4628 5909
rect 4204 5860 4588 5900
rect 4588 5851 4628 5860
rect 4395 5732 4437 5741
rect 4395 5692 4396 5732
rect 4436 5692 4437 5732
rect 4395 5683 4437 5692
rect 4587 5732 4629 5741
rect 4587 5692 4588 5732
rect 4628 5692 4629 5732
rect 4587 5683 4629 5692
rect 4396 5648 4436 5683
rect 4396 5597 4436 5608
rect 4588 4901 4628 5683
rect 4684 5228 4724 6028
rect 5355 6028 5356 6068
rect 5396 6028 5397 6068
rect 5355 6019 5397 6028
rect 4779 5648 4821 5657
rect 4779 5608 4780 5648
rect 4820 5608 4821 5648
rect 4779 5599 4821 5608
rect 4780 5514 4820 5599
rect 4928 5312 5296 5321
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 4928 5263 5296 5272
rect 4684 5188 4820 5228
rect 4780 5060 4820 5188
rect 5356 5144 5396 6019
rect 5356 5095 5396 5104
rect 4876 5060 4916 5069
rect 4780 5020 4876 5060
rect 4916 5020 5108 5060
rect 4876 5011 4916 5020
rect 5068 4976 5108 5020
rect 4684 4934 4724 4943
rect 4587 4892 4629 4901
rect 5068 4927 5108 4936
rect 5163 4976 5205 4985
rect 5163 4936 5164 4976
rect 5204 4936 5205 4976
rect 5163 4927 5205 4936
rect 4684 4892 4724 4894
rect 4875 4892 4917 4901
rect 4587 4852 4588 4892
rect 4628 4852 4820 4892
rect 4587 4843 4629 4852
rect 4588 4758 4628 4843
rect 3688 4556 4056 4565
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 3688 4507 4056 4516
rect 3627 4304 3669 4313
rect 3627 4264 3628 4304
rect 3668 4264 3669 4304
rect 3627 4255 3669 4264
rect 3628 4136 3668 4255
rect 3628 4087 3668 4096
rect 4587 3968 4629 3977
rect 4587 3928 4588 3968
rect 4628 3928 4629 3968
rect 4587 3919 4629 3928
rect 3627 3716 3669 3725
rect 3627 3676 3628 3716
rect 3668 3676 3669 3716
rect 3627 3667 3669 3676
rect 3628 3464 3668 3667
rect 3628 3415 3668 3424
rect 3531 3044 3573 3053
rect 3531 3004 3532 3044
rect 3572 3004 3573 3044
rect 3531 2995 3573 3004
rect 3688 3044 4056 3053
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 3688 2995 4056 3004
rect 4203 3044 4245 3053
rect 4203 3004 4204 3044
rect 4244 3004 4245 3044
rect 4203 2995 4245 3004
rect 3531 2876 3573 2885
rect 3531 2836 3532 2876
rect 3572 2836 3573 2876
rect 3531 2827 3573 2836
rect 3532 2624 3572 2827
rect 4204 2633 4244 2995
rect 3532 2575 3572 2584
rect 4203 2624 4245 2633
rect 4203 2584 4204 2624
rect 4244 2584 4245 2624
rect 4203 2575 4245 2584
rect 4395 2372 4437 2381
rect 4395 2332 4396 2372
rect 4436 2332 4437 2372
rect 4395 2323 4437 2332
rect 3532 1952 3572 1961
rect 3436 1912 3532 1952
rect 3532 1903 3572 1912
rect 4203 1952 4245 1961
rect 4203 1912 4204 1952
rect 4244 1912 4245 1952
rect 4203 1903 4245 1912
rect 3339 1700 3381 1709
rect 3339 1660 3340 1700
rect 3380 1660 3381 1700
rect 3339 1651 3381 1660
rect 3340 1566 3380 1651
rect 3688 1532 4056 1541
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 3688 1483 4056 1492
rect 3915 1280 3957 1289
rect 3244 1240 3380 1280
rect 3147 1231 3189 1240
rect 2955 272 2997 281
rect 2955 232 2956 272
rect 2996 232 2997 272
rect 2955 223 2997 232
rect 2956 80 2996 223
rect 3148 80 3188 1231
rect 3340 80 3380 1240
rect 3915 1240 3916 1280
rect 3956 1240 3957 1280
rect 3915 1231 3957 1240
rect 3723 356 3765 365
rect 3723 316 3724 356
rect 3764 316 3765 356
rect 3723 307 3765 316
rect 3531 272 3573 281
rect 3531 232 3532 272
rect 3572 232 3573 272
rect 3531 223 3573 232
rect 3532 80 3572 223
rect 3724 80 3764 307
rect 3916 80 3956 1231
rect 4107 1196 4149 1205
rect 4107 1156 4108 1196
rect 4148 1156 4149 1196
rect 4107 1147 4149 1156
rect 4108 80 4148 1147
rect 4204 617 4244 1903
rect 4299 1868 4341 1877
rect 4299 1828 4300 1868
rect 4340 1828 4341 1868
rect 4299 1819 4341 1828
rect 4203 608 4245 617
rect 4203 568 4204 608
rect 4244 568 4245 608
rect 4203 559 4245 568
rect 4300 80 4340 1819
rect 4396 1541 4436 2323
rect 4491 2288 4533 2297
rect 4491 2248 4492 2288
rect 4532 2248 4533 2288
rect 4491 2239 4533 2248
rect 4492 1709 4532 2239
rect 4588 1952 4628 3919
rect 4780 3464 4820 4852
rect 4875 4852 4876 4892
rect 4916 4852 4917 4892
rect 4875 4843 4917 4852
rect 4876 4136 4916 4843
rect 5164 4842 5204 4927
rect 5548 4901 5588 7027
rect 5740 7026 5780 7111
rect 6028 5741 6068 7783
rect 6123 7076 6165 7085
rect 6123 7036 6124 7076
rect 6164 7036 6165 7076
rect 6123 7027 6165 7036
rect 6124 6488 6164 7027
rect 6412 6656 6452 8128
rect 6508 8000 6548 8009
rect 6508 7841 6548 7960
rect 6604 7925 6644 8623
rect 6700 8345 6740 11068
rect 6796 8504 6836 11320
rect 7083 11276 7125 11285
rect 7083 11236 7084 11276
rect 7124 11236 7125 11276
rect 7083 11227 7125 11236
rect 7084 11024 7124 11227
rect 7084 10975 7124 10984
rect 7084 10184 7124 10193
rect 7084 10109 7124 10144
rect 7083 10100 7125 10109
rect 7083 10060 7084 10100
rect 7124 10060 7125 10100
rect 7083 10051 7125 10060
rect 7084 9269 7124 10051
rect 7083 9260 7125 9269
rect 7083 9220 7084 9260
rect 7124 9220 7125 9260
rect 7083 9211 7125 9220
rect 6892 8681 6932 8766
rect 6988 8756 7028 8765
rect 7180 8756 7220 18712
rect 7275 18164 7317 18173
rect 7275 18124 7276 18164
rect 7316 18124 7317 18164
rect 7275 18115 7317 18124
rect 7276 17744 7316 18115
rect 7276 17695 7316 17704
rect 7275 17072 7317 17081
rect 7275 17032 7276 17072
rect 7316 17032 7317 17072
rect 7275 17023 7317 17032
rect 7276 16938 7316 17023
rect 7372 16400 7412 19291
rect 7468 19270 7508 19804
rect 7468 19221 7508 19230
rect 7564 18668 7604 19963
rect 7660 19265 7700 20140
rect 7659 19256 7701 19265
rect 7659 19216 7660 19256
rect 7700 19216 7701 19256
rect 7659 19207 7701 19216
rect 7660 19088 7700 19097
rect 7660 18836 7700 19048
rect 7756 18836 7796 20644
rect 7948 18920 7988 21643
rect 8332 20768 8372 21904
rect 8332 20180 8372 20728
rect 8236 20140 8372 20180
rect 7948 18880 8084 18920
rect 7660 18796 7988 18836
rect 7756 18668 7796 18677
rect 7564 18628 7700 18668
rect 7564 18570 7604 18579
rect 7564 18005 7604 18530
rect 7563 17996 7605 18005
rect 7563 17956 7564 17996
rect 7604 17956 7605 17996
rect 7563 17947 7605 17956
rect 7660 17240 7700 18628
rect 7564 17200 7700 17240
rect 7276 16360 7412 16400
rect 7468 16820 7508 16829
rect 7276 14048 7316 16360
rect 7468 16316 7508 16780
rect 7420 16276 7508 16316
rect 7420 16274 7460 16276
rect 7420 16225 7460 16234
rect 7564 16232 7604 17200
rect 7659 17072 7701 17081
rect 7659 17032 7660 17072
rect 7700 17032 7701 17072
rect 7659 17023 7701 17032
rect 7660 16938 7700 17023
rect 7564 16192 7700 16232
rect 7564 16064 7604 16073
rect 7467 15980 7509 15989
rect 7467 15940 7468 15980
rect 7508 15940 7509 15980
rect 7467 15931 7509 15940
rect 7371 15896 7413 15905
rect 7371 15856 7372 15896
rect 7412 15856 7413 15896
rect 7371 15847 7413 15856
rect 7372 14561 7412 15847
rect 7468 15560 7508 15931
rect 7564 15653 7604 16024
rect 7563 15644 7605 15653
rect 7563 15604 7564 15644
rect 7604 15604 7605 15644
rect 7563 15595 7605 15604
rect 7468 15511 7508 15520
rect 7564 15476 7604 15485
rect 7660 15476 7700 16192
rect 7604 15436 7700 15476
rect 7564 15427 7604 15436
rect 7660 15233 7700 15436
rect 7659 15224 7701 15233
rect 7659 15184 7660 15224
rect 7700 15184 7701 15224
rect 7659 15175 7701 15184
rect 7563 15140 7605 15149
rect 7563 15100 7564 15140
rect 7604 15100 7605 15140
rect 7563 15091 7605 15100
rect 7371 14552 7413 14561
rect 7371 14512 7372 14552
rect 7412 14512 7413 14552
rect 7371 14503 7413 14512
rect 7372 14048 7412 14057
rect 7276 14008 7372 14048
rect 7275 13208 7317 13217
rect 7275 13168 7276 13208
rect 7316 13168 7317 13208
rect 7275 13159 7317 13168
rect 7276 11948 7316 13159
rect 7276 11899 7316 11908
rect 7275 11696 7317 11705
rect 7275 11656 7276 11696
rect 7316 11656 7317 11696
rect 7275 11647 7317 11656
rect 7028 8716 7220 8756
rect 6988 8707 7028 8716
rect 6891 8672 6933 8681
rect 6891 8632 6892 8672
rect 6932 8632 6933 8672
rect 6891 8623 6933 8632
rect 7179 8504 7221 8513
rect 6796 8464 6932 8504
rect 6699 8336 6741 8345
rect 6699 8296 6700 8336
rect 6740 8296 6741 8336
rect 6699 8287 6741 8296
rect 6699 8168 6741 8177
rect 6699 8128 6700 8168
rect 6740 8128 6741 8168
rect 6699 8119 6741 8128
rect 6700 8034 6740 8119
rect 6603 7916 6645 7925
rect 6603 7876 6604 7916
rect 6644 7876 6645 7916
rect 6603 7867 6645 7876
rect 6507 7832 6549 7841
rect 6507 7792 6508 7832
rect 6548 7792 6549 7832
rect 6507 7783 6549 7792
rect 6604 7337 6644 7867
rect 6603 7328 6645 7337
rect 6603 7288 6604 7328
rect 6644 7288 6645 7328
rect 6603 7279 6645 7288
rect 6796 6656 6836 6665
rect 6412 6616 6644 6656
rect 6124 6439 6164 6448
rect 6508 6488 6548 6497
rect 6508 6404 6548 6448
rect 6220 6364 6548 6404
rect 6604 6488 6644 6616
rect 6220 5900 6260 6364
rect 6604 6320 6644 6448
rect 6412 6280 6644 6320
rect 6220 5851 6260 5860
rect 6316 6236 6356 6245
rect 6316 5741 6356 6196
rect 6027 5732 6069 5741
rect 6027 5692 6028 5732
rect 6068 5692 6069 5732
rect 6027 5683 6069 5692
rect 6315 5732 6357 5741
rect 6315 5692 6316 5732
rect 6356 5692 6357 5732
rect 6315 5683 6357 5692
rect 6028 5648 6068 5683
rect 6028 5237 6068 5608
rect 6220 5480 6260 5489
rect 6123 5312 6165 5321
rect 6123 5272 6124 5312
rect 6164 5272 6165 5312
rect 6123 5263 6165 5272
rect 6027 5228 6069 5237
rect 6027 5188 6028 5228
rect 6068 5188 6069 5228
rect 6027 5179 6069 5188
rect 5740 4976 5780 4985
rect 5547 4892 5589 4901
rect 5547 4852 5548 4892
rect 5588 4852 5589 4892
rect 5547 4843 5589 4852
rect 5740 4817 5780 4936
rect 5739 4808 5781 4817
rect 5739 4768 5740 4808
rect 5780 4768 5781 4808
rect 5739 4759 5781 4768
rect 5931 4640 5973 4649
rect 5931 4600 5932 4640
rect 5972 4600 5973 4640
rect 5931 4591 5973 4600
rect 4876 3977 4916 4096
rect 5740 4136 5780 4145
rect 4875 3968 4917 3977
rect 4875 3928 4876 3968
rect 4916 3928 4917 3968
rect 4875 3919 4917 3928
rect 5068 3968 5108 3977
rect 5548 3968 5588 3977
rect 5108 3928 5492 3968
rect 5068 3919 5108 3928
rect 4928 3800 5296 3809
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 4928 3751 5296 3760
rect 4971 3632 5013 3641
rect 5355 3632 5397 3641
rect 4971 3592 4972 3632
rect 5012 3592 5013 3632
rect 4971 3583 5013 3592
rect 5164 3592 5300 3632
rect 4876 3464 4916 3473
rect 4780 3424 4876 3464
rect 4683 2624 4725 2633
rect 4683 2584 4684 2624
rect 4724 2584 4725 2624
rect 4683 2575 4725 2584
rect 4780 2624 4820 3424
rect 4876 3415 4916 3424
rect 4972 2876 5012 3583
rect 5067 3464 5109 3473
rect 5067 3424 5068 3464
rect 5108 3424 5109 3464
rect 5067 3415 5109 3424
rect 4972 2633 5012 2836
rect 5068 3212 5108 3415
rect 5164 3221 5204 3592
rect 5260 3548 5300 3592
rect 5355 3592 5356 3632
rect 5396 3592 5397 3632
rect 5355 3583 5397 3592
rect 5260 3499 5300 3508
rect 5356 3464 5396 3583
rect 5260 3441 5300 3450
rect 5356 3415 5396 3424
rect 5068 2717 5108 3172
rect 5163 3212 5205 3221
rect 5163 3172 5164 3212
rect 5204 3172 5205 3212
rect 5163 3163 5205 3172
rect 5163 2960 5205 2969
rect 5163 2920 5164 2960
rect 5204 2920 5205 2960
rect 5163 2911 5205 2920
rect 5164 2876 5204 2911
rect 5260 2876 5300 3401
rect 5452 3044 5492 3928
rect 5548 3464 5588 3928
rect 5740 3809 5780 4096
rect 5836 4136 5876 4145
rect 5739 3800 5781 3809
rect 5739 3760 5740 3800
rect 5780 3760 5781 3800
rect 5739 3751 5781 3760
rect 5836 3632 5876 4096
rect 5644 3592 5876 3632
rect 5644 3473 5684 3592
rect 5932 3548 5972 4591
rect 6124 4061 6164 5263
rect 6220 5069 6260 5440
rect 6219 5060 6261 5069
rect 6412 5060 6452 6280
rect 6507 5732 6549 5741
rect 6507 5692 6508 5732
rect 6548 5692 6549 5732
rect 6507 5683 6549 5692
rect 6508 5648 6548 5683
rect 6604 5657 6644 5742
rect 6508 5597 6548 5608
rect 6603 5648 6645 5657
rect 6603 5608 6604 5648
rect 6644 5608 6645 5648
rect 6603 5599 6645 5608
rect 6699 5144 6741 5153
rect 6699 5104 6700 5144
rect 6740 5104 6741 5144
rect 6699 5095 6741 5104
rect 6219 5020 6220 5060
rect 6260 5020 6261 5060
rect 6219 5011 6261 5020
rect 6316 5020 6452 5060
rect 6123 4052 6165 4061
rect 6123 4012 6124 4052
rect 6164 4012 6165 4052
rect 6123 4003 6165 4012
rect 6316 3968 6356 5020
rect 6411 4892 6453 4901
rect 6411 4852 6412 4892
rect 6452 4852 6453 4892
rect 6411 4843 6453 4852
rect 6220 3928 6356 3968
rect 6124 3809 6164 3828
rect 6123 3800 6165 3809
rect 6220 3800 6260 3928
rect 6123 3760 6124 3800
rect 6164 3760 6260 3800
rect 6123 3751 6165 3760
rect 5772 3508 5972 3548
rect 5548 3415 5588 3424
rect 5643 3464 5685 3473
rect 5643 3424 5644 3464
rect 5684 3424 5685 3464
rect 5643 3415 5685 3424
rect 5772 3461 5812 3508
rect 6220 3473 6260 3760
rect 6315 3800 6357 3809
rect 6315 3760 6316 3800
rect 6356 3760 6357 3800
rect 6315 3751 6357 3760
rect 5644 3330 5684 3415
rect 5772 3380 5812 3421
rect 6219 3464 6261 3473
rect 6219 3424 6220 3464
rect 6260 3424 6261 3464
rect 6219 3415 6261 3424
rect 5740 3340 5812 3380
rect 5452 3004 5588 3044
rect 5260 2836 5396 2876
rect 5164 2825 5204 2836
rect 5067 2708 5109 2717
rect 5067 2668 5068 2708
rect 5108 2668 5109 2708
rect 5067 2659 5109 2668
rect 5164 2647 5204 2656
rect 4780 2575 4820 2584
rect 4971 2624 5013 2633
rect 4971 2584 4972 2624
rect 5012 2584 5013 2624
rect 4971 2575 5013 2584
rect 5260 2633 5300 2718
rect 4684 2120 4724 2575
rect 5164 2465 5204 2607
rect 5259 2624 5301 2633
rect 5259 2584 5260 2624
rect 5300 2584 5301 2624
rect 5259 2575 5301 2584
rect 5163 2456 5205 2465
rect 5163 2416 5164 2456
rect 5204 2416 5205 2456
rect 5163 2407 5205 2416
rect 4928 2288 5296 2297
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 4928 2239 5296 2248
rect 5259 2120 5301 2129
rect 4684 2080 5108 2120
rect 4780 1952 4820 1961
rect 4588 1912 4780 1952
rect 4780 1903 4820 1912
rect 4971 1952 5013 1961
rect 4971 1912 4972 1952
rect 5012 1912 5013 1952
rect 5068 1952 5108 2080
rect 5259 2080 5260 2120
rect 5300 2080 5301 2120
rect 5259 2071 5301 2080
rect 5356 2120 5396 2836
rect 5452 2633 5492 2718
rect 5451 2624 5493 2633
rect 5451 2584 5452 2624
rect 5492 2584 5493 2624
rect 5451 2575 5493 2584
rect 5548 2624 5588 3004
rect 5740 2648 5780 3340
rect 5705 2639 5780 2648
rect 5745 2599 5780 2639
rect 5931 2624 5973 2633
rect 5705 2590 5745 2599
rect 5548 2540 5588 2584
rect 5931 2584 5932 2624
rect 5972 2584 5973 2624
rect 5931 2575 5973 2584
rect 6316 2624 6356 3751
rect 6412 3464 6452 4843
rect 6412 3415 6452 3424
rect 6316 2575 6356 2584
rect 5548 2500 5684 2540
rect 5547 2372 5589 2381
rect 5547 2332 5548 2372
rect 5588 2332 5589 2372
rect 5547 2323 5589 2332
rect 5451 2288 5493 2297
rect 5451 2248 5452 2288
rect 5492 2248 5493 2288
rect 5451 2239 5493 2248
rect 5356 2071 5396 2080
rect 5164 1952 5204 1961
rect 5068 1912 5164 1952
rect 4971 1903 5013 1912
rect 5164 1903 5204 1912
rect 5260 1952 5300 2071
rect 5260 1903 5300 1912
rect 5452 1952 5492 2239
rect 4972 1784 5012 1903
rect 5012 1744 5204 1784
rect 4972 1735 5012 1744
rect 4491 1700 4533 1709
rect 4491 1660 4492 1700
rect 4532 1660 4533 1700
rect 4491 1651 4533 1660
rect 4395 1532 4437 1541
rect 4395 1492 4396 1532
rect 4436 1492 4437 1532
rect 4395 1483 4437 1492
rect 4683 1448 4725 1457
rect 4683 1408 4684 1448
rect 4724 1408 4725 1448
rect 4683 1399 4725 1408
rect 4491 104 4533 113
rect 4491 80 4492 104
rect 1784 0 1864 80
rect 1976 0 2056 80
rect 2168 0 2248 80
rect 2360 0 2440 80
rect 2552 0 2632 80
rect 2744 0 2824 80
rect 2936 0 3016 80
rect 3128 0 3208 80
rect 3320 0 3400 80
rect 3512 0 3592 80
rect 3704 0 3784 80
rect 3896 0 3976 80
rect 4088 0 4168 80
rect 4280 0 4360 80
rect 4472 64 4492 80
rect 4532 80 4533 104
rect 4684 80 4724 1399
rect 5164 1112 5204 1744
rect 5355 1448 5397 1457
rect 5355 1408 5356 1448
rect 5396 1408 5397 1448
rect 5355 1399 5397 1408
rect 5356 1280 5396 1399
rect 5452 1280 5492 1912
rect 5548 1457 5588 2323
rect 5644 1952 5684 2500
rect 5739 2288 5781 2297
rect 5739 2248 5740 2288
rect 5780 2248 5781 2288
rect 5739 2239 5781 2248
rect 5547 1448 5589 1457
rect 5547 1408 5548 1448
rect 5588 1408 5589 1448
rect 5547 1399 5589 1408
rect 5356 1231 5396 1240
rect 5445 1240 5492 1280
rect 5445 1196 5485 1240
rect 5445 1156 5492 1196
rect 5164 1063 5204 1072
rect 5260 1112 5300 1121
rect 5452 1112 5492 1156
rect 5300 1072 5396 1112
rect 5260 1063 5300 1072
rect 5356 944 5396 1072
rect 5452 1063 5492 1072
rect 5644 944 5684 1912
rect 5740 1952 5780 2239
rect 5932 2120 5972 2575
rect 6700 2381 6740 5095
rect 6796 5069 6836 6616
rect 6795 5060 6837 5069
rect 6795 5020 6796 5060
rect 6836 5020 6837 5060
rect 6795 5011 6837 5020
rect 6892 4640 6932 8464
rect 7179 8464 7180 8504
rect 7220 8464 7221 8504
rect 7179 8455 7221 8464
rect 7083 8336 7125 8345
rect 7083 8296 7084 8336
rect 7124 8296 7125 8336
rect 7083 8287 7125 8296
rect 6988 8000 7028 8009
rect 6988 7412 7028 7960
rect 7084 8000 7124 8287
rect 7084 7673 7124 7960
rect 7180 7841 7220 8455
rect 7276 8009 7316 11647
rect 7372 10109 7412 14008
rect 7467 13880 7509 13889
rect 7467 13840 7468 13880
rect 7508 13840 7509 13880
rect 7467 13831 7509 13840
rect 7468 13208 7508 13831
rect 7468 13159 7508 13168
rect 7468 12536 7508 12547
rect 7468 12461 7508 12496
rect 7467 12452 7509 12461
rect 7467 12412 7468 12452
rect 7508 12412 7509 12452
rect 7467 12403 7509 12412
rect 7467 12200 7509 12209
rect 7467 12160 7468 12200
rect 7508 12160 7509 12200
rect 7467 12151 7509 12160
rect 7468 11948 7508 12151
rect 7468 11899 7508 11908
rect 7564 11108 7604 15091
rect 7659 14888 7701 14897
rect 7659 14848 7660 14888
rect 7700 14848 7701 14888
rect 7659 14839 7701 14848
rect 7660 14754 7700 14839
rect 7659 12620 7701 12629
rect 7659 12580 7660 12620
rect 7700 12580 7701 12620
rect 7659 12571 7701 12580
rect 7660 12486 7700 12571
rect 7660 11780 7700 11789
rect 7756 11780 7796 18628
rect 7851 14804 7893 14813
rect 7851 14764 7852 14804
rect 7892 14764 7893 14804
rect 7851 14755 7893 14764
rect 7852 14670 7892 14755
rect 7948 13208 7988 18796
rect 8044 16409 8084 18880
rect 8139 17996 8181 18005
rect 8139 17956 8140 17996
rect 8180 17956 8181 17996
rect 8139 17947 8181 17956
rect 8043 16400 8085 16409
rect 8043 16360 8044 16400
rect 8084 16360 8085 16400
rect 8043 16351 8085 16360
rect 8043 15896 8085 15905
rect 8043 15856 8044 15896
rect 8084 15856 8085 15896
rect 8043 15847 8085 15856
rect 8044 15560 8084 15847
rect 8140 15728 8180 17947
rect 8236 15905 8276 20140
rect 8428 20021 8468 21988
rect 8427 20012 8469 20021
rect 8427 19972 8428 20012
rect 8468 19972 8469 20012
rect 8427 19963 8469 19972
rect 8331 19256 8373 19265
rect 8331 19216 8332 19256
rect 8372 19216 8373 19256
rect 8331 19207 8373 19216
rect 8235 15896 8277 15905
rect 8235 15856 8236 15896
rect 8276 15856 8277 15896
rect 8235 15847 8277 15856
rect 8140 15688 8276 15728
rect 8044 15511 8084 15520
rect 8043 15056 8085 15065
rect 8043 15016 8044 15056
rect 8084 15016 8085 15056
rect 8043 15007 8085 15016
rect 8044 14720 8084 15007
rect 8139 14888 8181 14897
rect 8139 14848 8140 14888
rect 8180 14848 8181 14888
rect 8139 14839 8181 14848
rect 8044 14671 8084 14680
rect 8043 13292 8085 13301
rect 8043 13252 8044 13292
rect 8084 13252 8085 13292
rect 8043 13243 8085 13252
rect 7948 13040 7988 13168
rect 8044 13158 8084 13243
rect 7948 13000 8084 13040
rect 7851 12956 7893 12965
rect 7851 12916 7852 12956
rect 7892 12916 7893 12956
rect 7851 12907 7893 12916
rect 7700 11740 7796 11780
rect 7852 12536 7892 12907
rect 7660 11731 7700 11740
rect 7852 11705 7892 12496
rect 7947 12452 7989 12461
rect 7947 12412 7948 12452
rect 7988 12412 7989 12452
rect 7947 12403 7989 12412
rect 7948 11957 7988 12403
rect 8044 12293 8084 13000
rect 8043 12284 8085 12293
rect 8043 12244 8044 12284
rect 8084 12244 8085 12284
rect 8043 12235 8085 12244
rect 7947 11948 7989 11957
rect 7947 11908 7948 11948
rect 7988 11908 7989 11948
rect 7947 11899 7989 11908
rect 7851 11696 7893 11705
rect 7851 11656 7852 11696
rect 7892 11656 7893 11696
rect 7851 11647 7893 11656
rect 8140 11537 8180 14839
rect 8139 11528 8181 11537
rect 8139 11488 8140 11528
rect 8180 11488 8181 11528
rect 8139 11479 8181 11488
rect 7468 11068 7604 11108
rect 7756 11108 7796 11117
rect 7796 11068 8180 11108
rect 7468 10856 7508 11068
rect 7756 11059 7796 11068
rect 7612 10982 7652 10991
rect 7612 10940 7652 10942
rect 8140 10940 8180 11068
rect 7612 10900 7796 10940
rect 7468 10816 7604 10856
rect 7467 10688 7509 10697
rect 7467 10648 7468 10688
rect 7508 10648 7509 10688
rect 7467 10639 7509 10648
rect 7371 10100 7413 10109
rect 7371 10060 7372 10100
rect 7412 10060 7413 10100
rect 7371 10051 7413 10060
rect 7468 9932 7508 10639
rect 7372 9892 7508 9932
rect 7372 9353 7412 9892
rect 7564 9680 7604 10816
rect 7659 10184 7701 10193
rect 7659 10144 7660 10184
rect 7700 10144 7701 10184
rect 7659 10135 7701 10144
rect 7468 9640 7604 9680
rect 7371 9344 7413 9353
rect 7371 9304 7372 9344
rect 7412 9304 7413 9344
rect 7468 9344 7508 9640
rect 7564 9512 7604 9521
rect 7660 9512 7700 10135
rect 7756 9680 7796 10900
rect 8140 10891 8180 10900
rect 7948 10772 7988 10781
rect 7948 10529 7988 10732
rect 7947 10520 7989 10529
rect 7947 10480 7948 10520
rect 7988 10480 7989 10520
rect 7947 10471 7989 10480
rect 8236 9680 8276 15688
rect 8332 12881 8372 19207
rect 8524 18005 8564 22567
rect 8620 19424 8660 23584
rect 8811 23584 8812 23624
rect 8852 23584 8853 23624
rect 8811 23575 8853 23584
rect 8812 23490 8852 23575
rect 9292 23372 9332 23752
rect 9004 23332 9332 23372
rect 8716 23204 8756 23213
rect 8716 23120 8756 23164
rect 9004 23120 9044 23332
rect 8716 23080 9004 23120
rect 9004 23071 9044 23080
rect 8715 22952 8757 22961
rect 8715 22912 8716 22952
rect 8756 22912 8757 22952
rect 8715 22903 8757 22912
rect 8716 21608 8756 22903
rect 8908 22868 8948 22877
rect 8908 22289 8948 22828
rect 8907 22280 8949 22289
rect 8907 22240 8908 22280
rect 8948 22240 8949 22280
rect 8907 22231 8949 22240
rect 9388 22121 9428 23920
rect 9483 23792 9525 23801
rect 9483 23752 9484 23792
rect 9524 23752 9525 23792
rect 9483 23743 9525 23752
rect 9484 23213 9524 23743
rect 9483 23204 9525 23213
rect 9483 23164 9484 23204
rect 9524 23164 9525 23204
rect 9483 23155 9525 23164
rect 9580 23036 9620 26104
rect 9484 22996 9620 23036
rect 8907 22112 8949 22121
rect 8907 22072 8908 22112
rect 8948 22072 8949 22112
rect 8907 22063 8949 22072
rect 9387 22112 9429 22121
rect 9387 22072 9388 22112
rect 9428 22072 9429 22112
rect 9387 22063 9429 22072
rect 8800 21617 8840 21636
rect 8800 21608 8852 21617
rect 8716 21568 8812 21608
rect 8812 21281 8852 21568
rect 8811 21272 8853 21281
rect 8811 21232 8812 21272
rect 8852 21232 8853 21272
rect 8811 21223 8853 21232
rect 8908 20936 8948 22063
rect 9004 21692 9044 21701
rect 9044 21652 9332 21692
rect 9004 21643 9044 21652
rect 9292 21608 9332 21652
rect 9292 21559 9332 21568
rect 9387 21608 9429 21617
rect 9387 21568 9388 21608
rect 9428 21568 9429 21608
rect 9387 21559 9429 21568
rect 9195 21524 9237 21533
rect 9195 21484 9196 21524
rect 9236 21484 9237 21524
rect 9195 21475 9237 21484
rect 8716 20896 8948 20936
rect 8716 20684 8756 20896
rect 8860 20777 8900 20786
rect 8900 20737 8948 20768
rect 8860 20728 8948 20737
rect 8716 20644 8852 20684
rect 8715 20432 8757 20441
rect 8715 20392 8716 20432
rect 8756 20392 8757 20432
rect 8715 20383 8757 20392
rect 8716 20096 8756 20383
rect 8716 20021 8756 20056
rect 8715 20012 8757 20021
rect 8715 19972 8716 20012
rect 8756 19972 8757 20012
rect 8715 19963 8757 19972
rect 8620 19384 8756 19424
rect 8620 19256 8660 19265
rect 8523 17996 8565 18005
rect 8523 17956 8524 17996
rect 8564 17956 8565 17996
rect 8620 17996 8660 19216
rect 8716 19256 8756 19384
rect 8716 18164 8756 19216
rect 8812 18845 8852 20644
rect 8908 20264 8948 20728
rect 8908 20215 8948 20224
rect 9004 20600 9044 20609
rect 8811 18836 8853 18845
rect 8811 18796 8812 18836
rect 8852 18796 8853 18836
rect 8811 18787 8853 18796
rect 8812 18425 8852 18787
rect 8811 18416 8853 18425
rect 8811 18376 8812 18416
rect 8852 18376 8853 18416
rect 8811 18367 8853 18376
rect 8716 18124 8852 18164
rect 8716 17996 8756 18005
rect 8620 17956 8716 17996
rect 8523 17947 8565 17956
rect 8716 17947 8756 17956
rect 8524 17753 8564 17838
rect 8812 17828 8852 18124
rect 8716 17788 8852 17828
rect 8907 17828 8949 17837
rect 8907 17788 8908 17828
rect 8948 17788 8949 17828
rect 8523 17744 8565 17753
rect 8523 17704 8524 17744
rect 8564 17704 8565 17744
rect 8523 17695 8565 17704
rect 8716 17249 8756 17788
rect 8907 17779 8949 17788
rect 8908 17744 8948 17779
rect 8908 17693 8948 17704
rect 8811 17660 8853 17669
rect 8811 17620 8812 17660
rect 8852 17620 8853 17660
rect 8811 17611 8853 17620
rect 8715 17240 8757 17249
rect 8715 17200 8716 17240
rect 8756 17200 8757 17240
rect 8715 17191 8757 17200
rect 8427 17156 8469 17165
rect 8427 17116 8428 17156
rect 8468 17116 8469 17156
rect 8427 17107 8469 17116
rect 8428 16661 8468 17107
rect 8812 17072 8852 17611
rect 8908 17072 8948 17081
rect 8812 17032 8908 17072
rect 8908 17023 8948 17032
rect 8427 16652 8469 16661
rect 8427 16612 8428 16652
rect 8468 16612 8469 16652
rect 8427 16603 8469 16612
rect 8907 15980 8949 15989
rect 8907 15940 8908 15980
rect 8948 15940 8949 15980
rect 8907 15931 8949 15940
rect 8716 15644 8756 15653
rect 8572 15518 8612 15527
rect 8572 15476 8612 15478
rect 8572 15436 8660 15476
rect 8427 15308 8469 15317
rect 8427 15268 8428 15308
rect 8468 15268 8469 15308
rect 8427 15259 8469 15268
rect 8428 14897 8468 15259
rect 8427 14888 8469 14897
rect 8427 14848 8428 14888
rect 8468 14848 8469 14888
rect 8427 14839 8469 14848
rect 8620 14216 8660 15436
rect 8716 14813 8756 15604
rect 8715 14804 8757 14813
rect 8715 14764 8716 14804
rect 8756 14764 8757 14804
rect 8715 14755 8757 14764
rect 8812 14216 8852 14225
rect 8620 14176 8812 14216
rect 8812 14167 8852 14176
rect 8619 14048 8661 14057
rect 8619 14008 8620 14048
rect 8660 14008 8661 14048
rect 8619 13999 8661 14008
rect 8427 13376 8469 13385
rect 8427 13336 8428 13376
rect 8468 13336 8469 13376
rect 8427 13327 8469 13336
rect 8428 13208 8468 13327
rect 8428 13159 8468 13168
rect 8523 13208 8565 13217
rect 8523 13168 8524 13208
rect 8564 13168 8565 13208
rect 8523 13159 8565 13168
rect 8524 13074 8564 13159
rect 8331 12872 8373 12881
rect 8331 12832 8332 12872
rect 8372 12832 8373 12872
rect 8331 12823 8373 12832
rect 8620 11957 8660 13999
rect 8715 13964 8757 13973
rect 8715 13924 8716 13964
rect 8756 13924 8757 13964
rect 8715 13915 8757 13924
rect 8619 11948 8661 11957
rect 8619 11908 8620 11948
rect 8660 11908 8661 11948
rect 8619 11899 8661 11908
rect 8332 11696 8372 11705
rect 8332 11360 8372 11656
rect 8428 11696 8468 11705
rect 8716 11696 8756 13915
rect 8811 11864 8853 11873
rect 8811 11824 8812 11864
rect 8852 11824 8853 11864
rect 8811 11815 8853 11824
rect 8468 11656 8756 11696
rect 8812 11780 8852 11815
rect 8428 11647 8468 11656
rect 8332 11320 8564 11360
rect 8524 10436 8564 11320
rect 8524 10387 8564 10396
rect 8331 10184 8373 10193
rect 8331 10144 8332 10184
rect 8372 10144 8373 10184
rect 8331 10135 8373 10144
rect 8332 10050 8372 10135
rect 8620 9689 8660 11656
rect 8715 11528 8757 11537
rect 8715 11488 8716 11528
rect 8756 11488 8757 11528
rect 8715 11479 8757 11488
rect 8716 11024 8756 11479
rect 7756 9631 7796 9640
rect 8044 9640 8276 9680
rect 8619 9680 8661 9689
rect 8619 9640 8620 9680
rect 8660 9640 8661 9680
rect 7604 9472 7700 9512
rect 7948 9512 7988 9521
rect 7564 9463 7604 9472
rect 7468 9304 7604 9344
rect 7371 9295 7413 9304
rect 7372 8672 7412 9295
rect 7372 8623 7412 8632
rect 7468 8672 7508 8683
rect 7468 8597 7508 8632
rect 7467 8588 7509 8597
rect 7467 8548 7468 8588
rect 7508 8548 7509 8588
rect 7467 8539 7509 8548
rect 7275 8000 7317 8009
rect 7275 7960 7276 8000
rect 7316 7960 7317 8000
rect 7275 7951 7317 7960
rect 7467 8000 7509 8009
rect 7467 7960 7468 8000
rect 7508 7960 7509 8000
rect 7467 7951 7509 7960
rect 7564 8000 7604 9304
rect 7659 9260 7701 9269
rect 7659 9220 7660 9260
rect 7700 9220 7701 9260
rect 7659 9211 7701 9220
rect 7564 7951 7604 7960
rect 7179 7832 7221 7841
rect 7179 7792 7180 7832
rect 7220 7792 7221 7832
rect 7179 7783 7221 7792
rect 7083 7664 7125 7673
rect 7083 7624 7084 7664
rect 7124 7624 7125 7664
rect 7083 7615 7125 7624
rect 7180 7412 7220 7421
rect 6988 7372 7180 7412
rect 7180 7363 7220 7372
rect 6988 7160 7028 7171
rect 7276 7160 7316 7951
rect 7468 7866 7508 7951
rect 7372 7160 7412 7169
rect 7276 7120 7372 7160
rect 6988 7085 7028 7120
rect 7372 7111 7412 7120
rect 6987 7076 7029 7085
rect 6987 7036 6988 7076
rect 7028 7036 7029 7076
rect 6987 7027 7029 7036
rect 7467 6992 7509 7001
rect 7467 6952 7468 6992
rect 7508 6952 7509 6992
rect 7467 6943 7509 6952
rect 6987 6488 7029 6497
rect 6987 6448 6988 6488
rect 7028 6448 7029 6488
rect 6987 6439 7029 6448
rect 6988 6354 7028 6439
rect 6987 5816 7029 5825
rect 6987 5776 6988 5816
rect 7028 5776 7029 5816
rect 6987 5767 7029 5776
rect 6988 5732 7028 5767
rect 6988 5405 7028 5692
rect 7083 5732 7125 5741
rect 7083 5692 7084 5732
rect 7124 5692 7125 5732
rect 7083 5683 7125 5692
rect 7084 5598 7124 5683
rect 6987 5396 7029 5405
rect 6987 5356 6988 5396
rect 7028 5356 7029 5396
rect 6987 5347 7029 5356
rect 6987 5228 7029 5237
rect 6987 5188 6988 5228
rect 7028 5188 7029 5228
rect 7468 5228 7508 6943
rect 7564 5648 7604 5657
rect 7660 5648 7700 9211
rect 7948 8252 7988 9472
rect 7852 8212 7988 8252
rect 7852 8009 7892 8212
rect 8044 8177 8084 9640
rect 8619 9631 8661 9640
rect 8140 9512 8180 9521
rect 8140 9185 8180 9472
rect 8236 9512 8276 9521
rect 8620 9512 8660 9521
rect 8276 9472 8372 9512
rect 8236 9463 8276 9472
rect 8236 9344 8276 9353
rect 8139 9176 8181 9185
rect 8139 9136 8140 9176
rect 8180 9136 8181 9176
rect 8139 9127 8181 9136
rect 8236 8681 8276 9304
rect 8332 8849 8372 9472
rect 8524 9472 8620 9512
rect 8428 9260 8468 9271
rect 8428 9185 8468 9220
rect 8427 9176 8469 9185
rect 8427 9136 8428 9176
rect 8468 9136 8469 9176
rect 8427 9127 8469 9136
rect 8331 8840 8373 8849
rect 8331 8800 8332 8840
rect 8372 8800 8373 8840
rect 8331 8791 8373 8800
rect 8332 8706 8372 8791
rect 8235 8672 8277 8681
rect 8235 8632 8236 8672
rect 8276 8632 8277 8672
rect 8235 8623 8277 8632
rect 8524 8672 8564 9472
rect 8620 9463 8660 9472
rect 8619 9260 8661 9269
rect 8619 9220 8620 9260
rect 8660 9220 8661 9260
rect 8619 9211 8661 9220
rect 8524 8513 8564 8632
rect 8523 8504 8565 8513
rect 8523 8464 8524 8504
rect 8564 8464 8565 8504
rect 8523 8455 8565 8464
rect 8620 8336 8660 9211
rect 8332 8296 8660 8336
rect 8043 8168 8085 8177
rect 8043 8128 8044 8168
rect 8084 8128 8085 8168
rect 8043 8119 8085 8128
rect 7851 8000 7893 8009
rect 7851 7960 7852 8000
rect 7892 7960 7893 8000
rect 7851 7951 7893 7960
rect 8044 8000 8084 8011
rect 8044 7925 8084 7960
rect 8043 7916 8085 7925
rect 8043 7876 8044 7916
rect 8084 7876 8085 7916
rect 8043 7867 8085 7876
rect 8235 7076 8277 7085
rect 8235 7036 8236 7076
rect 8276 7036 8277 7076
rect 8235 7027 8277 7036
rect 8236 6488 8276 7027
rect 8332 6833 8372 8296
rect 8716 8261 8756 10984
rect 8812 9941 8852 11740
rect 8908 11780 8948 15931
rect 8908 11731 8948 11740
rect 8811 9932 8853 9941
rect 8811 9892 8812 9932
rect 8852 9892 8853 9932
rect 8811 9883 8853 9892
rect 8715 8252 8757 8261
rect 8715 8212 8716 8252
rect 8756 8212 8757 8252
rect 8715 8203 8757 8212
rect 8716 8084 8756 8093
rect 8428 8044 8716 8084
rect 8331 6824 8373 6833
rect 8331 6784 8332 6824
rect 8372 6784 8373 6824
rect 8331 6775 8373 6784
rect 8236 6439 8276 6448
rect 8428 6404 8468 8044
rect 8716 8035 8756 8044
rect 8572 7958 8612 7967
rect 8572 7916 8612 7918
rect 8907 7916 8949 7925
rect 8572 7876 8756 7916
rect 8523 7580 8565 7589
rect 8523 7540 8524 7580
rect 8564 7540 8565 7580
rect 8523 7531 8565 7540
rect 8524 6908 8564 7531
rect 8716 7412 8756 7876
rect 8907 7876 8908 7916
rect 8948 7876 8949 7916
rect 8907 7867 8949 7876
rect 8812 7412 8852 7421
rect 8716 7372 8812 7412
rect 8812 7363 8852 7372
rect 8908 7244 8948 7867
rect 9004 7589 9044 20560
rect 9099 20096 9141 20105
rect 9099 20056 9100 20096
rect 9140 20056 9141 20096
rect 9099 20047 9141 20056
rect 9100 19962 9140 20047
rect 9099 19424 9141 19433
rect 9099 19384 9100 19424
rect 9140 19384 9141 19424
rect 9099 19375 9141 19384
rect 9100 19340 9140 19375
rect 9100 19289 9140 19300
rect 9196 19256 9236 21475
rect 9388 19601 9428 21559
rect 9387 19592 9429 19601
rect 9387 19552 9388 19592
rect 9428 19552 9429 19592
rect 9387 19543 9429 19552
rect 9196 19088 9236 19216
rect 9100 19048 9236 19088
rect 9100 17585 9140 19048
rect 9195 18920 9237 18929
rect 9195 18880 9196 18920
rect 9236 18880 9237 18920
rect 9195 18871 9237 18880
rect 9099 17576 9141 17585
rect 9099 17536 9100 17576
rect 9140 17536 9141 17576
rect 9099 17527 9141 17536
rect 9099 17156 9141 17165
rect 9099 17116 9100 17156
rect 9140 17116 9141 17156
rect 9099 17107 9141 17116
rect 9100 17022 9140 17107
rect 9099 12620 9141 12629
rect 9099 12580 9100 12620
rect 9140 12580 9141 12620
rect 9099 12571 9141 12580
rect 9100 12536 9140 12571
rect 9100 12485 9140 12496
rect 9100 10184 9140 10193
rect 9100 9521 9140 10144
rect 9099 9512 9141 9521
rect 9099 9472 9100 9512
rect 9140 9472 9141 9512
rect 9099 9463 9141 9472
rect 9196 8168 9236 18871
rect 9292 18584 9332 18593
rect 9292 17669 9332 18544
rect 9484 18257 9524 22996
rect 9580 20777 9620 20862
rect 9579 20768 9621 20777
rect 9579 20728 9580 20768
rect 9620 20728 9621 20768
rect 9579 20719 9621 20728
rect 9579 20600 9621 20609
rect 9579 20560 9580 20600
rect 9620 20560 9621 20600
rect 9579 20551 9621 20560
rect 9580 18593 9620 20551
rect 9676 20180 9716 27448
rect 9772 26909 9812 29800
rect 9868 29756 9908 29767
rect 9868 29681 9908 29716
rect 9867 29672 9909 29681
rect 9867 29632 9868 29672
rect 9908 29632 9909 29672
rect 9867 29623 9909 29632
rect 9964 29345 10004 30967
rect 9963 29336 10005 29345
rect 9963 29296 9964 29336
rect 10004 29296 10005 29336
rect 9963 29287 10005 29296
rect 9867 28328 9909 28337
rect 9867 28288 9868 28328
rect 9908 28288 9909 28328
rect 9867 28279 9909 28288
rect 9868 28194 9908 28279
rect 10060 27740 10100 34327
rect 10155 34208 10197 34217
rect 10155 34168 10156 34208
rect 10196 34168 10197 34208
rect 10155 34159 10197 34168
rect 10156 34074 10196 34159
rect 10156 30008 10196 30017
rect 10156 29177 10196 29968
rect 10252 29429 10292 34336
rect 10348 33629 10388 36343
rect 10444 35972 10484 36688
rect 10540 36679 10580 36688
rect 10732 36728 10772 36737
rect 10539 36560 10581 36569
rect 10539 36520 10540 36560
rect 10580 36520 10581 36560
rect 10539 36511 10581 36520
rect 10540 36426 10580 36511
rect 10732 36065 10772 36688
rect 10924 36728 10964 37267
rect 10924 36679 10964 36688
rect 11019 36728 11061 36737
rect 11019 36688 11020 36728
rect 11060 36688 11061 36728
rect 11019 36679 11061 36688
rect 10827 36644 10869 36653
rect 10827 36604 10828 36644
rect 10868 36604 10869 36644
rect 10827 36595 10869 36604
rect 10539 36056 10581 36065
rect 10539 36016 10540 36056
rect 10580 36016 10581 36056
rect 10539 36007 10581 36016
rect 10731 36056 10773 36065
rect 10731 36016 10732 36056
rect 10772 36016 10773 36056
rect 10731 36007 10773 36016
rect 10444 35923 10484 35932
rect 10540 35888 10580 36007
rect 10540 35729 10580 35848
rect 10635 35888 10677 35897
rect 10635 35848 10636 35888
rect 10676 35848 10677 35888
rect 10635 35839 10677 35848
rect 10732 35888 10772 35899
rect 10539 35720 10581 35729
rect 10444 35680 10540 35720
rect 10580 35680 10581 35720
rect 10444 35216 10484 35680
rect 10539 35671 10581 35680
rect 10636 35384 10676 35839
rect 10732 35813 10772 35848
rect 10731 35804 10773 35813
rect 10731 35764 10732 35804
rect 10772 35764 10773 35804
rect 10731 35755 10773 35764
rect 10540 35344 10676 35384
rect 10540 35300 10580 35344
rect 10732 35300 10772 35755
rect 10828 35561 10868 36595
rect 11020 36594 11060 36679
rect 11020 36140 11060 36149
rect 11116 36140 11156 37360
rect 11308 37400 11348 37409
rect 11212 37232 11252 37241
rect 11212 37073 11252 37192
rect 11211 37064 11253 37073
rect 11211 37024 11212 37064
rect 11252 37024 11253 37064
rect 11211 37015 11253 37024
rect 11308 36896 11348 37360
rect 11224 36856 11348 36896
rect 11404 37400 11444 37771
rect 11224 36644 11264 36856
rect 11404 36812 11444 37360
rect 11595 37400 11637 37409
rect 11595 37360 11596 37400
rect 11636 37360 11637 37400
rect 11595 37351 11637 37360
rect 11596 37266 11636 37351
rect 11692 36896 11732 37780
rect 11884 37568 11924 37577
rect 11924 37528 12020 37568
rect 11884 37519 11924 37528
rect 11788 37400 11828 37409
rect 11788 37241 11828 37360
rect 11884 37400 11924 37409
rect 11787 37232 11829 37241
rect 11787 37192 11788 37232
rect 11828 37192 11829 37232
rect 11787 37183 11829 37192
rect 11308 36772 11444 36812
rect 11500 36856 11732 36896
rect 11308 36743 11348 36772
rect 11308 36694 11348 36703
rect 11500 36644 11540 36856
rect 11596 36728 11636 36739
rect 11788 36737 11828 37183
rect 11596 36653 11636 36688
rect 11692 36728 11732 36737
rect 11212 36604 11264 36644
rect 11404 36604 11540 36644
rect 11595 36644 11637 36653
rect 11595 36604 11596 36644
rect 11636 36604 11637 36644
rect 11212 36224 11252 36604
rect 11307 36476 11349 36485
rect 11307 36436 11308 36476
rect 11348 36436 11349 36476
rect 11307 36427 11349 36436
rect 11308 36233 11348 36427
rect 11060 36100 11156 36140
rect 11209 36184 11252 36224
rect 11307 36224 11349 36233
rect 11307 36184 11308 36224
rect 11348 36184 11349 36224
rect 11209 36140 11249 36184
rect 11307 36175 11349 36184
rect 11209 36100 11252 36140
rect 11020 36091 11060 36100
rect 10923 36056 10965 36065
rect 11212 36056 11252 36100
rect 10923 36016 10924 36056
rect 10964 36016 10965 36056
rect 10923 36007 10965 36016
rect 11209 36016 11252 36056
rect 10827 35552 10869 35561
rect 10827 35512 10828 35552
rect 10868 35512 10869 35552
rect 10827 35503 10869 35512
rect 10732 35260 10868 35300
rect 10540 35251 10580 35260
rect 10444 35167 10484 35176
rect 10636 35216 10676 35225
rect 10828 35216 10868 35260
rect 10676 35176 10772 35216
rect 10636 35167 10676 35176
rect 10539 35132 10581 35141
rect 10539 35092 10540 35132
rect 10580 35092 10581 35132
rect 10539 35083 10581 35092
rect 10443 35048 10485 35057
rect 10443 35008 10444 35048
rect 10484 35008 10485 35048
rect 10443 34999 10485 35008
rect 10347 33620 10389 33629
rect 10347 33580 10348 33620
rect 10388 33580 10389 33620
rect 10347 33571 10389 33580
rect 10348 30941 10388 33571
rect 10444 33125 10484 34999
rect 10540 34376 10580 35083
rect 10635 34964 10677 34973
rect 10635 34924 10636 34964
rect 10676 34924 10677 34964
rect 10635 34915 10677 34924
rect 10540 34327 10580 34336
rect 10636 34376 10676 34915
rect 10732 34385 10772 35176
rect 10828 35167 10868 35176
rect 10827 35048 10869 35057
rect 10827 35008 10828 35048
rect 10868 35008 10869 35048
rect 10827 34999 10869 35008
rect 10636 34327 10676 34336
rect 10731 34376 10773 34385
rect 10731 34336 10732 34376
rect 10772 34336 10773 34376
rect 10731 34327 10773 34336
rect 10828 34208 10868 34999
rect 10924 34553 10964 36007
rect 11020 35981 11060 35983
rect 11019 35972 11061 35981
rect 11019 35932 11020 35972
rect 11060 35932 11061 35972
rect 11209 35972 11249 36016
rect 11209 35932 11252 35972
rect 11019 35923 11061 35932
rect 11020 35888 11060 35923
rect 11020 35839 11060 35848
rect 11019 35720 11061 35729
rect 11019 35680 11020 35720
rect 11060 35680 11061 35720
rect 11019 35671 11061 35680
rect 10923 34544 10965 34553
rect 10923 34504 10924 34544
rect 10964 34504 10965 34544
rect 10923 34495 10965 34504
rect 10636 34168 10868 34208
rect 10443 33116 10485 33125
rect 10443 33076 10444 33116
rect 10484 33076 10485 33116
rect 10443 33067 10485 33076
rect 10347 30932 10389 30941
rect 10347 30892 10348 30932
rect 10388 30892 10389 30932
rect 10347 30883 10389 30892
rect 10444 30773 10484 33067
rect 10540 32192 10580 32201
rect 10636 32192 10676 34168
rect 10924 34133 10964 34495
rect 11020 34376 11060 35671
rect 11115 35216 11157 35225
rect 11115 35176 11116 35216
rect 11156 35176 11157 35216
rect 11115 35167 11157 35176
rect 11116 35082 11156 35167
rect 11115 34964 11157 34973
rect 11115 34924 11116 34964
rect 11156 34924 11157 34964
rect 11115 34915 11157 34924
rect 11116 34830 11156 34915
rect 11115 34628 11157 34637
rect 11115 34588 11116 34628
rect 11156 34588 11157 34628
rect 11115 34579 11157 34588
rect 11116 34460 11156 34579
rect 11116 34411 11156 34420
rect 10923 34124 10965 34133
rect 10923 34084 10924 34124
rect 10964 34084 10965 34124
rect 10923 34075 10965 34084
rect 11020 33116 11060 34336
rect 11212 33881 11252 35932
rect 11308 35888 11348 35897
rect 11308 35729 11348 35848
rect 11307 35720 11349 35729
rect 11307 35680 11308 35720
rect 11348 35680 11349 35720
rect 11307 35671 11349 35680
rect 11307 35552 11349 35561
rect 11307 35512 11308 35552
rect 11348 35512 11349 35552
rect 11404 35552 11444 36604
rect 11595 36595 11637 36604
rect 11596 35888 11636 35899
rect 11500 35729 11540 35814
rect 11596 35813 11636 35848
rect 11595 35804 11637 35813
rect 11595 35764 11596 35804
rect 11636 35764 11637 35804
rect 11595 35755 11637 35764
rect 11499 35720 11541 35729
rect 11499 35680 11500 35720
rect 11540 35680 11541 35720
rect 11499 35671 11541 35680
rect 11692 35636 11732 36688
rect 11787 36728 11829 36737
rect 11787 36688 11788 36728
rect 11828 36688 11829 36728
rect 11787 36679 11829 36688
rect 11788 36476 11828 36679
rect 11884 36560 11924 37360
rect 11980 36728 12020 37528
rect 12172 37493 12212 41308
rect 12364 41273 12404 42736
rect 12556 41777 12596 44584
rect 12844 44456 12884 48616
rect 12940 45968 12980 48700
rect 13131 48700 13132 48740
rect 13172 48700 13173 48740
rect 13131 48691 13173 48700
rect 13132 46556 13172 48691
rect 13227 48572 13269 48581
rect 13227 48532 13228 48572
rect 13268 48532 13269 48572
rect 13227 48523 13269 48532
rect 13132 46507 13172 46516
rect 13035 46472 13077 46481
rect 13035 46432 13036 46472
rect 13076 46432 13077 46472
rect 13035 46423 13077 46432
rect 13036 46338 13076 46423
rect 12940 45919 12980 45928
rect 13132 45716 13172 45725
rect 12844 44416 12980 44456
rect 12844 44288 12884 44297
rect 12844 44129 12884 44248
rect 12843 44120 12885 44129
rect 12843 44080 12844 44120
rect 12884 44080 12885 44120
rect 12843 44071 12885 44080
rect 12748 43448 12788 43457
rect 12844 43448 12884 44071
rect 12788 43408 12884 43448
rect 12748 43399 12788 43408
rect 12940 41945 12980 44416
rect 13132 43280 13172 45676
rect 13228 45128 13268 48523
rect 13324 46313 13364 48784
rect 13419 48824 13461 48833
rect 13419 48784 13420 48824
rect 13460 48784 13461 48824
rect 13419 48775 13461 48784
rect 13420 47909 13460 48775
rect 13516 47984 13556 49111
rect 13612 48581 13652 51883
rect 13708 51008 13748 52219
rect 13708 48740 13748 50968
rect 13804 51008 13844 52303
rect 13804 48749 13844 50968
rect 13708 48665 13748 48700
rect 13803 48740 13845 48749
rect 13803 48700 13804 48740
rect 13844 48700 13845 48740
rect 13803 48691 13845 48700
rect 13707 48656 13749 48665
rect 13707 48616 13708 48656
rect 13748 48616 13749 48656
rect 13707 48607 13749 48616
rect 13804 48606 13844 48691
rect 13611 48572 13653 48581
rect 13611 48532 13612 48572
rect 13652 48532 13653 48572
rect 13611 48523 13653 48532
rect 13612 47984 13652 47993
rect 13516 47944 13612 47984
rect 13419 47900 13461 47909
rect 13419 47860 13420 47900
rect 13460 47860 13461 47900
rect 13419 47851 13461 47860
rect 13323 46304 13365 46313
rect 13323 46264 13324 46304
rect 13364 46264 13365 46304
rect 13323 46255 13365 46264
rect 13324 45389 13364 46255
rect 13420 45800 13460 47851
rect 13516 47321 13556 47944
rect 13612 47935 13652 47944
rect 13515 47312 13557 47321
rect 13515 47272 13516 47312
rect 13556 47272 13557 47312
rect 13515 47263 13557 47272
rect 13900 47060 13940 56923
rect 13996 53873 14036 59872
rect 14379 59576 14421 59585
rect 14379 59536 14380 59576
rect 14420 59536 14421 59576
rect 14379 59527 14421 59536
rect 14380 59442 14420 59527
rect 14187 59408 14229 59417
rect 14187 59368 14188 59408
rect 14228 59368 14229 59408
rect 14187 59359 14229 59368
rect 14091 58904 14133 58913
rect 14091 58864 14092 58904
rect 14132 58864 14133 58904
rect 14091 58855 14133 58864
rect 14092 58568 14132 58855
rect 14092 57989 14132 58528
rect 14091 57980 14133 57989
rect 14091 57940 14092 57980
rect 14132 57940 14133 57980
rect 14091 57931 14133 57940
rect 14091 55376 14133 55385
rect 14091 55336 14092 55376
rect 14132 55336 14133 55376
rect 14091 55327 14133 55336
rect 14092 54881 14132 55327
rect 14091 54872 14133 54881
rect 14091 54832 14092 54872
rect 14132 54832 14133 54872
rect 14091 54823 14133 54832
rect 14092 54738 14132 54823
rect 13995 53864 14037 53873
rect 13995 53824 13996 53864
rect 14036 53824 14037 53864
rect 13995 53815 14037 53824
rect 13995 53528 14037 53537
rect 13995 53488 13996 53528
rect 14036 53488 14037 53528
rect 13995 53479 14037 53488
rect 13996 53360 14036 53479
rect 14188 53355 14228 59359
rect 14476 57980 14516 60712
rect 14572 59576 14612 60871
rect 14668 60005 14708 61552
rect 14764 61543 14804 61552
rect 14860 61592 14900 61601
rect 14860 61433 14900 61552
rect 14859 61424 14901 61433
rect 14859 61384 14860 61424
rect 14900 61384 14901 61424
rect 14859 61375 14901 61384
rect 14956 61349 14996 61627
rect 15052 61424 15092 62215
rect 15052 61375 15092 61384
rect 14955 61340 14997 61349
rect 14955 61300 14956 61340
rect 14996 61300 14997 61340
rect 14955 61291 14997 61300
rect 14763 61256 14805 61265
rect 14763 61216 14764 61256
rect 14804 61216 14805 61256
rect 14763 61207 14805 61216
rect 14764 60089 14804 61207
rect 14955 61172 14997 61181
rect 14955 61132 14956 61172
rect 14996 61132 14997 61172
rect 14955 61123 14997 61132
rect 14956 60920 14996 61123
rect 14860 60880 14956 60920
rect 14763 60080 14805 60089
rect 14763 60040 14764 60080
rect 14804 60040 14805 60080
rect 14763 60031 14805 60040
rect 14667 59996 14709 60005
rect 14667 59956 14668 59996
rect 14708 59956 14709 59996
rect 14667 59947 14709 59956
rect 14572 59527 14612 59536
rect 14764 59408 14804 60031
rect 14764 59359 14804 59368
rect 14476 57940 14612 57980
rect 14475 57812 14517 57821
rect 14475 57772 14476 57812
rect 14516 57772 14517 57812
rect 14475 57763 14517 57772
rect 14283 57308 14325 57317
rect 14283 57268 14284 57308
rect 14324 57268 14325 57308
rect 14283 57259 14325 57268
rect 14284 57149 14324 57259
rect 14379 57224 14421 57233
rect 14379 57184 14380 57224
rect 14420 57184 14421 57224
rect 14379 57175 14421 57184
rect 14283 57140 14325 57149
rect 14283 57100 14284 57140
rect 14324 57100 14325 57140
rect 14283 57091 14325 57100
rect 14380 57140 14420 57175
rect 14284 57006 14324 57091
rect 14283 56636 14325 56645
rect 14283 56596 14284 56636
rect 14324 56596 14325 56636
rect 14283 56587 14325 56596
rect 13996 53311 14036 53320
rect 14087 53315 14228 53355
rect 13995 53192 14037 53201
rect 13995 53152 13996 53192
rect 14036 53152 14037 53192
rect 14087 53192 14127 53315
rect 14188 53192 14228 53201
rect 14087 53152 14132 53192
rect 13995 53143 14037 53152
rect 13996 52697 14036 53143
rect 13995 52688 14037 52697
rect 13995 52648 13996 52688
rect 14036 52648 14037 52688
rect 13995 52639 14037 52648
rect 13996 51017 14036 52639
rect 14092 52016 14132 53152
rect 14188 52534 14228 53152
rect 14188 52485 14228 52494
rect 14284 52436 14324 56587
rect 14380 55973 14420 57100
rect 14476 56393 14516 57763
rect 14572 56645 14612 57940
rect 14764 57896 14804 57905
rect 14764 57569 14804 57856
rect 14763 57560 14805 57569
rect 14763 57520 14764 57560
rect 14804 57520 14805 57560
rect 14763 57511 14805 57520
rect 14860 57233 14900 60880
rect 14956 60871 14996 60880
rect 14955 59324 14997 59333
rect 14955 59284 14956 59324
rect 14996 59284 14997 59324
rect 14955 59275 14997 59284
rect 14859 57224 14901 57233
rect 14859 57184 14860 57224
rect 14900 57184 14901 57224
rect 14859 57175 14901 57184
rect 14859 57056 14901 57065
rect 14859 57016 14860 57056
rect 14900 57016 14901 57056
rect 14859 57007 14901 57016
rect 14860 56922 14900 57007
rect 14667 56720 14709 56729
rect 14667 56680 14668 56720
rect 14708 56680 14709 56720
rect 14667 56671 14709 56680
rect 14571 56636 14613 56645
rect 14571 56596 14572 56636
rect 14612 56596 14613 56636
rect 14571 56587 14613 56596
rect 14475 56384 14517 56393
rect 14475 56344 14476 56384
rect 14516 56344 14517 56384
rect 14475 56335 14517 56344
rect 14476 56250 14516 56335
rect 14668 56300 14708 56671
rect 14572 56260 14708 56300
rect 14379 55964 14421 55973
rect 14379 55924 14380 55964
rect 14420 55924 14421 55964
rect 14379 55915 14421 55924
rect 14380 55721 14420 55915
rect 14379 55712 14421 55721
rect 14379 55672 14380 55712
rect 14420 55672 14421 55712
rect 14379 55663 14421 55672
rect 14380 55544 14420 55553
rect 14572 55544 14612 56260
rect 14668 56132 14708 56141
rect 14860 56132 14900 56141
rect 14708 56092 14804 56132
rect 14668 56083 14708 56092
rect 14667 55964 14709 55973
rect 14667 55924 14668 55964
rect 14708 55924 14709 55964
rect 14667 55915 14709 55924
rect 14420 55504 14612 55544
rect 14380 54965 14420 55504
rect 14572 55376 14612 55385
rect 14379 54956 14421 54965
rect 14379 54916 14380 54956
rect 14420 54916 14421 54956
rect 14379 54907 14421 54916
rect 14380 53537 14420 54907
rect 14572 54867 14612 55336
rect 14572 54818 14612 54827
rect 14668 53696 14708 55915
rect 14764 55460 14804 56092
rect 14860 55889 14900 56092
rect 14859 55880 14901 55889
rect 14859 55840 14860 55880
rect 14900 55840 14901 55880
rect 14859 55831 14901 55840
rect 14956 55460 14996 59275
rect 15148 58577 15188 64240
rect 15340 64028 15380 64240
rect 15628 64112 15668 64576
rect 15724 64567 15764 64576
rect 15723 64364 15765 64373
rect 15723 64324 15724 64364
rect 15764 64324 15765 64364
rect 15723 64315 15765 64324
rect 15724 64121 15764 64315
rect 15244 63988 15380 64028
rect 15532 64072 15668 64112
rect 15723 64112 15765 64121
rect 15723 64072 15724 64112
rect 15764 64072 15765 64112
rect 15532 64070 15572 64072
rect 15723 64063 15765 64072
rect 15532 64021 15572 64030
rect 15244 62777 15284 63988
rect 15723 63944 15765 63953
rect 15340 63930 15380 63939
rect 15723 63904 15724 63944
rect 15764 63904 15765 63944
rect 15723 63895 15765 63904
rect 15340 63869 15380 63890
rect 15339 63860 15381 63869
rect 15339 63820 15340 63860
rect 15380 63820 15381 63860
rect 15339 63811 15381 63820
rect 15340 63795 15380 63811
rect 15724 63810 15764 63895
rect 15243 62768 15285 62777
rect 15243 62728 15244 62768
rect 15284 62728 15285 62768
rect 15243 62719 15285 62728
rect 15724 62600 15764 62609
rect 15820 62600 15860 65164
rect 16012 64616 16052 64625
rect 16108 64616 16148 65248
rect 16204 64616 16244 64625
rect 16108 64576 16204 64616
rect 15916 64448 15956 64457
rect 15916 64121 15956 64408
rect 16012 64205 16052 64576
rect 16204 64567 16244 64576
rect 16203 64448 16245 64457
rect 16203 64408 16204 64448
rect 16244 64408 16245 64448
rect 16203 64399 16245 64408
rect 16011 64196 16053 64205
rect 16011 64156 16012 64196
rect 16052 64156 16053 64196
rect 16011 64147 16053 64156
rect 15915 64112 15957 64121
rect 15915 64072 15916 64112
rect 15956 64072 15957 64112
rect 15915 64063 15957 64072
rect 15915 63944 15957 63953
rect 15915 63904 15916 63944
rect 15956 63904 15957 63944
rect 15915 63895 15957 63904
rect 16012 63944 16052 63953
rect 15916 63810 15956 63895
rect 15820 62560 15956 62600
rect 15244 62432 15284 62441
rect 15244 61853 15284 62392
rect 15340 62432 15380 62441
rect 15340 62273 15380 62392
rect 15436 62432 15476 62441
rect 15339 62264 15381 62273
rect 15339 62224 15340 62264
rect 15380 62224 15381 62264
rect 15339 62215 15381 62224
rect 15243 61844 15285 61853
rect 15243 61804 15244 61844
rect 15284 61804 15285 61844
rect 15436 61844 15476 62392
rect 15531 62432 15573 62441
rect 15531 62392 15532 62432
rect 15572 62392 15573 62432
rect 15531 62383 15573 62392
rect 15532 62298 15572 62383
rect 15436 61804 15572 61844
rect 15243 61795 15285 61804
rect 15244 61571 15284 61580
rect 15244 61349 15284 61531
rect 15340 61571 15380 61580
rect 15243 61340 15285 61349
rect 15243 61300 15244 61340
rect 15284 61300 15285 61340
rect 15243 61291 15285 61300
rect 15340 61181 15380 61531
rect 15436 61571 15476 61580
rect 15532 61571 15572 61804
rect 15724 61685 15764 62560
rect 15820 62432 15860 62441
rect 15820 61769 15860 62392
rect 15916 61928 15956 62560
rect 16012 62441 16052 63904
rect 16204 63944 16244 64399
rect 16204 63869 16244 63904
rect 16203 63860 16245 63869
rect 16203 63820 16204 63860
rect 16244 63820 16245 63860
rect 16203 63811 16245 63820
rect 16204 63780 16244 63811
rect 16300 63524 16340 65416
rect 16396 65297 16436 65920
rect 16684 65456 16724 65995
rect 16684 65407 16724 65416
rect 16779 65372 16821 65381
rect 16779 65332 16780 65372
rect 16820 65332 16821 65372
rect 16779 65323 16821 65332
rect 16395 65288 16437 65297
rect 16395 65248 16396 65288
rect 16436 65248 16437 65288
rect 16395 65239 16437 65248
rect 16780 65238 16820 65323
rect 16683 65120 16725 65129
rect 16683 65080 16684 65120
rect 16724 65080 16725 65120
rect 16683 65071 16725 65080
rect 16684 64280 16724 65071
rect 17164 64280 17204 69784
rect 17452 67136 17492 70204
rect 17836 70204 18164 70244
rect 17644 69992 17684 70001
rect 17547 69740 17589 69749
rect 17547 69700 17548 69740
rect 17588 69700 17589 69740
rect 17547 69691 17589 69700
rect 17548 68984 17588 69691
rect 17644 69413 17684 69952
rect 17740 69992 17780 70001
rect 17740 69749 17780 69952
rect 17739 69740 17781 69749
rect 17739 69700 17740 69740
rect 17780 69700 17781 69740
rect 17739 69691 17781 69700
rect 17836 69572 17876 70204
rect 18027 70076 18069 70085
rect 18027 70036 18028 70076
rect 18068 70036 18069 70076
rect 18027 70027 18069 70036
rect 17931 69908 17973 69917
rect 17931 69868 17932 69908
rect 17972 69868 17973 69908
rect 17931 69859 17973 69868
rect 17740 69532 17876 69572
rect 17643 69404 17685 69413
rect 17643 69364 17644 69404
rect 17684 69364 17685 69404
rect 17643 69355 17685 69364
rect 17643 69236 17685 69245
rect 17643 69196 17644 69236
rect 17684 69196 17685 69236
rect 17643 69187 17685 69196
rect 17644 69152 17684 69187
rect 17644 69101 17684 69112
rect 17548 68944 17684 68984
rect 17547 68228 17589 68237
rect 17547 68188 17548 68228
rect 17588 68188 17589 68228
rect 17547 68179 17589 68188
rect 17548 67640 17588 68179
rect 17548 67591 17588 67600
rect 17644 67640 17684 68944
rect 17740 67649 17780 69532
rect 17835 69404 17877 69413
rect 17835 69364 17836 69404
rect 17876 69364 17877 69404
rect 17835 69355 17877 69364
rect 17836 69270 17876 69355
rect 17644 67565 17684 67600
rect 17739 67640 17781 67649
rect 17739 67600 17740 67640
rect 17780 67600 17781 67640
rect 17739 67591 17781 67600
rect 17643 67556 17685 67565
rect 17643 67516 17644 67556
rect 17684 67516 17685 67556
rect 17643 67507 17685 67516
rect 17452 67096 17684 67136
rect 17260 66968 17300 66977
rect 17260 66137 17300 66928
rect 17356 66968 17396 66977
rect 17548 66968 17588 66977
rect 17356 66725 17396 66928
rect 17452 66928 17548 66968
rect 17355 66716 17397 66725
rect 17355 66676 17356 66716
rect 17396 66676 17397 66716
rect 17355 66667 17397 66676
rect 17452 66221 17492 66928
rect 17548 66919 17588 66928
rect 17547 66800 17589 66809
rect 17547 66760 17548 66800
rect 17588 66760 17589 66800
rect 17547 66751 17589 66760
rect 17548 66666 17588 66751
rect 17644 66548 17684 67096
rect 17932 66809 17972 69859
rect 18028 68153 18068 70027
rect 18124 69992 18164 70204
rect 18124 69943 18164 69952
rect 18220 69908 18260 69917
rect 18220 69833 18260 69868
rect 18219 69824 18261 69833
rect 18219 69784 18220 69824
rect 18260 69784 18261 69824
rect 18219 69775 18261 69784
rect 18220 69320 18260 69775
rect 18124 69280 18260 69320
rect 18027 68144 18069 68153
rect 18027 68104 18028 68144
rect 18068 68104 18069 68144
rect 18027 68095 18069 68104
rect 18027 67976 18069 67985
rect 18027 67936 18028 67976
rect 18068 67936 18069 67976
rect 18027 67927 18069 67936
rect 18028 67724 18068 67927
rect 18028 67675 18068 67684
rect 18124 67640 18164 69280
rect 18316 69236 18356 71875
rect 18603 71672 18645 71681
rect 18603 71632 18604 71672
rect 18644 71632 18645 71672
rect 18603 71623 18645 71632
rect 18604 70673 18644 71623
rect 18603 70664 18645 70673
rect 18603 70624 18604 70664
rect 18644 70624 18645 70664
rect 18603 70615 18645 70624
rect 18411 69320 18453 69329
rect 18411 69280 18412 69320
rect 18452 69280 18453 69320
rect 18411 69271 18453 69280
rect 18220 69196 18356 69236
rect 18220 69152 18260 69196
rect 18412 69152 18452 69271
rect 18604 69245 18644 70615
rect 18700 70169 18740 82039
rect 18796 82013 18836 82804
rect 19180 82844 19220 82853
rect 19180 82256 19220 82804
rect 20044 82601 20084 82686
rect 19180 82207 19220 82216
rect 19660 82592 19700 82601
rect 19660 82097 19700 82552
rect 20043 82592 20085 82601
rect 20043 82552 20044 82592
rect 20084 82552 20085 82592
rect 20043 82543 20085 82552
rect 20048 82424 20416 82433
rect 20088 82384 20130 82424
rect 20170 82384 20212 82424
rect 20252 82384 20294 82424
rect 20334 82384 20376 82424
rect 20048 82375 20416 82384
rect 19659 82088 19701 82097
rect 19659 82048 19660 82088
rect 19700 82048 19701 82088
rect 19659 82039 19701 82048
rect 18795 82004 18837 82013
rect 18795 81964 18796 82004
rect 18836 81964 18837 82004
rect 18795 81955 18837 81964
rect 18796 81870 18836 81955
rect 19275 81920 19317 81929
rect 19275 81880 19276 81920
rect 19316 81880 19317 81920
rect 19275 81871 19317 81880
rect 19276 81786 19316 81871
rect 18808 81668 19176 81677
rect 18848 81628 18890 81668
rect 18930 81628 18972 81668
rect 19012 81628 19054 81668
rect 19094 81628 19136 81668
rect 18808 81619 19176 81628
rect 20048 80912 20416 80921
rect 20088 80872 20130 80912
rect 20170 80872 20212 80912
rect 20252 80872 20294 80912
rect 20334 80872 20376 80912
rect 20048 80863 20416 80872
rect 18808 80156 19176 80165
rect 18848 80116 18890 80156
rect 18930 80116 18972 80156
rect 19012 80116 19054 80156
rect 19094 80116 19136 80156
rect 18808 80107 19176 80116
rect 20048 79400 20416 79409
rect 20088 79360 20130 79400
rect 20170 79360 20212 79400
rect 20252 79360 20294 79400
rect 20334 79360 20376 79400
rect 20048 79351 20416 79360
rect 18808 78644 19176 78653
rect 18848 78604 18890 78644
rect 18930 78604 18972 78644
rect 19012 78604 19054 78644
rect 19094 78604 19136 78644
rect 18808 78595 19176 78604
rect 20811 78560 20853 78569
rect 20811 78520 20812 78560
rect 20852 78520 20853 78560
rect 20811 78511 20853 78520
rect 20048 77888 20416 77897
rect 20088 77848 20130 77888
rect 20170 77848 20212 77888
rect 20252 77848 20294 77888
rect 20334 77848 20376 77888
rect 20048 77839 20416 77848
rect 18808 77132 19176 77141
rect 18848 77092 18890 77132
rect 18930 77092 18972 77132
rect 19012 77092 19054 77132
rect 19094 77092 19136 77132
rect 18808 77083 19176 77092
rect 20523 76544 20565 76553
rect 20523 76504 20524 76544
rect 20564 76504 20565 76544
rect 20523 76495 20565 76504
rect 20048 76376 20416 76385
rect 20088 76336 20130 76376
rect 20170 76336 20212 76376
rect 20252 76336 20294 76376
rect 20334 76336 20376 76376
rect 20048 76327 20416 76336
rect 18808 75620 19176 75629
rect 18848 75580 18890 75620
rect 18930 75580 18972 75620
rect 19012 75580 19054 75620
rect 19094 75580 19136 75620
rect 18808 75571 19176 75580
rect 20048 74864 20416 74873
rect 20088 74824 20130 74864
rect 20170 74824 20212 74864
rect 20252 74824 20294 74864
rect 20334 74824 20376 74864
rect 20048 74815 20416 74824
rect 18808 74108 19176 74117
rect 18848 74068 18890 74108
rect 18930 74068 18972 74108
rect 19012 74068 19054 74108
rect 19094 74068 19136 74108
rect 18808 74059 19176 74068
rect 20048 73352 20416 73361
rect 20088 73312 20130 73352
rect 20170 73312 20212 73352
rect 20252 73312 20294 73352
rect 20334 73312 20376 73352
rect 20048 73303 20416 73312
rect 18808 72596 19176 72605
rect 18848 72556 18890 72596
rect 18930 72556 18972 72596
rect 19012 72556 19054 72596
rect 19094 72556 19136 72596
rect 18808 72547 19176 72556
rect 20048 71840 20416 71849
rect 20088 71800 20130 71840
rect 20170 71800 20212 71840
rect 20252 71800 20294 71840
rect 20334 71800 20376 71840
rect 20048 71791 20416 71800
rect 18795 71672 18837 71681
rect 18795 71632 18796 71672
rect 18836 71632 18837 71672
rect 18795 71623 18837 71632
rect 18796 71504 18836 71623
rect 19372 71513 19412 71598
rect 18796 71455 18836 71464
rect 19371 71504 19413 71513
rect 19371 71464 19372 71504
rect 19412 71464 19413 71504
rect 19371 71455 19413 71464
rect 18988 71252 19028 71261
rect 19468 71252 19508 71261
rect 19028 71212 19316 71252
rect 18988 71203 19028 71212
rect 18808 71084 19176 71093
rect 18848 71044 18890 71084
rect 18930 71044 18972 71084
rect 19012 71044 19054 71084
rect 19094 71044 19136 71084
rect 18808 71035 19176 71044
rect 18891 70664 18933 70673
rect 19276 70664 19316 71212
rect 19468 70916 19508 71212
rect 19468 70876 19700 70916
rect 19371 70832 19413 70841
rect 19371 70792 19372 70832
rect 19412 70792 19413 70832
rect 19371 70783 19413 70792
rect 18891 70624 18892 70664
rect 18932 70624 18933 70664
rect 18891 70615 18933 70624
rect 19180 70624 19276 70664
rect 18892 70530 18932 70615
rect 18795 70496 18837 70505
rect 18795 70456 18796 70496
rect 18836 70456 18837 70496
rect 18795 70447 18837 70456
rect 19084 70496 19124 70505
rect 18699 70160 18741 70169
rect 18699 70120 18700 70160
rect 18740 70120 18741 70160
rect 18699 70111 18741 70120
rect 18699 69992 18741 70001
rect 18699 69952 18700 69992
rect 18740 69952 18741 69992
rect 18699 69943 18741 69952
rect 18700 69858 18740 69943
rect 18796 69740 18836 70447
rect 18987 70076 19029 70085
rect 18987 70036 18988 70076
rect 19028 70036 19029 70076
rect 18987 70027 19029 70036
rect 18988 69833 19028 70027
rect 19084 70001 19124 70456
rect 19083 69992 19125 70001
rect 19083 69952 19084 69992
rect 19124 69952 19125 69992
rect 19083 69943 19125 69952
rect 19180 69987 19220 70624
rect 19276 70615 19316 70624
rect 19372 70664 19412 70783
rect 19372 70615 19412 70624
rect 19467 70664 19509 70673
rect 19467 70624 19468 70664
rect 19508 70624 19509 70664
rect 19467 70615 19509 70624
rect 19468 70530 19508 70615
rect 19564 70496 19604 70505
rect 19371 70076 19413 70085
rect 19371 70036 19372 70076
rect 19412 70036 19413 70076
rect 19371 70027 19413 70036
rect 18987 69824 19029 69833
rect 18987 69784 18988 69824
rect 19028 69784 19029 69824
rect 18987 69775 19029 69784
rect 19084 69749 19124 69943
rect 19180 69824 19220 69947
rect 19372 69942 19412 70027
rect 19564 69992 19604 70456
rect 19564 69943 19604 69952
rect 19660 69992 19700 70876
rect 19852 70664 19892 70673
rect 19755 70496 19797 70505
rect 19755 70456 19756 70496
rect 19796 70456 19797 70496
rect 19755 70447 19797 70456
rect 19756 70362 19796 70447
rect 19852 70160 19892 70624
rect 20043 70580 20085 70589
rect 20043 70540 20044 70580
rect 20084 70540 20085 70580
rect 20043 70531 20085 70540
rect 20044 70446 20084 70531
rect 20048 70328 20416 70337
rect 20088 70288 20130 70328
rect 20170 70288 20212 70328
rect 20252 70288 20294 70328
rect 20334 70288 20376 70328
rect 20048 70279 20416 70288
rect 19660 69943 19700 69952
rect 19756 70120 19892 70160
rect 19756 69824 19796 70120
rect 20043 70076 20085 70085
rect 20043 70036 20044 70076
rect 20084 70036 20085 70076
rect 20043 70027 20085 70036
rect 19852 69992 19892 70001
rect 20044 69992 20084 70027
rect 19892 69952 19988 69992
rect 19852 69943 19892 69952
rect 19180 69784 19412 69824
rect 18700 69700 18836 69740
rect 19083 69740 19125 69749
rect 19083 69700 19084 69740
rect 19124 69700 19125 69740
rect 18700 69413 18740 69700
rect 19083 69691 19125 69700
rect 19275 69656 19317 69665
rect 19275 69616 19276 69656
rect 19316 69616 19317 69656
rect 19275 69607 19317 69616
rect 18808 69572 19176 69581
rect 18848 69532 18890 69572
rect 18930 69532 18972 69572
rect 19012 69532 19054 69572
rect 19094 69532 19136 69572
rect 18808 69523 19176 69532
rect 19276 69413 19316 69607
rect 18699 69404 18741 69413
rect 18699 69364 18700 69404
rect 18740 69364 18741 69404
rect 18699 69355 18741 69364
rect 18891 69404 18933 69413
rect 18891 69364 18892 69404
rect 18932 69364 18933 69404
rect 18891 69355 18933 69364
rect 19275 69404 19317 69413
rect 19275 69364 19276 69404
rect 19316 69364 19317 69404
rect 19275 69355 19317 69364
rect 18603 69236 18645 69245
rect 18603 69196 18604 69236
rect 18644 69196 18645 69236
rect 18603 69187 18645 69196
rect 18220 68816 18260 69112
rect 18316 69131 18356 69140
rect 18412 69103 18452 69112
rect 18700 69152 18740 69355
rect 18700 69103 18740 69112
rect 18796 69152 18836 69161
rect 18316 68993 18356 69091
rect 18315 68984 18357 68993
rect 18315 68944 18316 68984
rect 18356 68944 18357 68984
rect 18315 68935 18357 68944
rect 18508 68984 18548 68993
rect 18796 68984 18836 69112
rect 18892 69152 18932 69355
rect 18987 69236 19029 69245
rect 18987 69196 18988 69236
rect 19028 69196 19029 69236
rect 18987 69187 19029 69196
rect 18892 69103 18932 69112
rect 18988 69152 19028 69187
rect 18988 69101 19028 69112
rect 19180 69152 19220 69163
rect 19372 69161 19412 69784
rect 19468 69784 19796 69824
rect 19948 69824 19988 69952
rect 20044 69941 20084 69952
rect 20235 69992 20277 70001
rect 20235 69952 20236 69992
rect 20276 69952 20277 69992
rect 20235 69943 20277 69952
rect 20236 69858 20276 69943
rect 20044 69824 20084 69833
rect 19948 69784 20044 69824
rect 19180 69077 19220 69112
rect 19276 69152 19316 69161
rect 19371 69152 19413 69161
rect 19316 69112 19372 69152
rect 19412 69112 19413 69152
rect 19179 69068 19221 69077
rect 19179 69028 19180 69068
rect 19220 69028 19221 69068
rect 19179 69019 19221 69028
rect 19276 68993 19316 69112
rect 19371 69103 19413 69112
rect 19372 69018 19412 69103
rect 18548 68944 18836 68984
rect 19275 68984 19317 68993
rect 19275 68944 19276 68984
rect 19316 68944 19317 68984
rect 18508 68935 18548 68944
rect 19275 68935 19317 68944
rect 19468 68984 19508 69784
rect 20044 69775 20084 69784
rect 19852 69740 19892 69749
rect 19659 69656 19701 69665
rect 19659 69616 19660 69656
rect 19700 69616 19701 69656
rect 19659 69607 19701 69616
rect 19660 69152 19700 69607
rect 19852 69497 19892 69700
rect 19851 69488 19893 69497
rect 19851 69448 19852 69488
rect 19892 69448 19893 69488
rect 19851 69439 19893 69448
rect 19947 69320 19989 69329
rect 19947 69280 19948 69320
rect 19988 69280 19989 69320
rect 19947 69271 19989 69280
rect 19660 69103 19700 69112
rect 19755 69152 19797 69161
rect 19755 69112 19756 69152
rect 19796 69112 19797 69152
rect 19755 69103 19797 69112
rect 19756 69018 19796 69103
rect 19468 68935 19508 68944
rect 19948 68984 19988 69271
rect 19948 68935 19988 68944
rect 18795 68816 18837 68825
rect 18220 68776 18644 68816
rect 18220 68480 18260 68489
rect 18220 68069 18260 68440
rect 18604 68480 18644 68776
rect 18795 68776 18796 68816
rect 18836 68776 18837 68816
rect 18795 68767 18837 68776
rect 20048 68816 20416 68825
rect 20088 68776 20130 68816
rect 20170 68776 20212 68816
rect 20252 68776 20294 68816
rect 20334 68776 20376 68816
rect 20048 68767 20416 68776
rect 18604 68431 18644 68440
rect 18699 68480 18741 68489
rect 18699 68440 18700 68480
rect 18740 68440 18741 68480
rect 18699 68431 18741 68440
rect 18700 68346 18740 68431
rect 18411 68228 18453 68237
rect 18796 68228 18836 68767
rect 18892 68480 18932 68489
rect 18892 68237 18932 68440
rect 19084 68480 19124 68489
rect 18411 68188 18412 68228
rect 18452 68188 18453 68228
rect 18411 68179 18453 68188
rect 18700 68188 18836 68228
rect 18891 68228 18933 68237
rect 18891 68188 18892 68228
rect 18932 68188 18933 68228
rect 19084 68228 19124 68440
rect 19275 68480 19317 68489
rect 19275 68440 19276 68480
rect 19316 68440 19317 68480
rect 19275 68431 19317 68440
rect 19372 68480 19412 68489
rect 19412 68440 19796 68480
rect 19372 68431 19412 68440
rect 19276 68346 19316 68431
rect 19372 68312 19412 68321
rect 19084 68188 19316 68228
rect 18412 68094 18452 68179
rect 18603 68144 18645 68153
rect 18603 68104 18604 68144
rect 18644 68104 18645 68144
rect 18603 68095 18645 68104
rect 18219 68060 18261 68069
rect 18219 68020 18220 68060
rect 18260 68020 18261 68060
rect 18219 68011 18261 68020
rect 18124 67556 18164 67600
rect 18604 67640 18644 68095
rect 18124 67516 18356 67556
rect 18028 66968 18068 66977
rect 17931 66800 17973 66809
rect 17931 66760 17932 66800
rect 17972 66760 17973 66800
rect 17931 66751 17973 66760
rect 17548 66508 17684 66548
rect 17451 66212 17493 66221
rect 17451 66172 17452 66212
rect 17492 66172 17493 66212
rect 17451 66163 17493 66172
rect 17259 66128 17301 66137
rect 17259 66088 17260 66128
rect 17300 66088 17301 66128
rect 17259 66079 17301 66088
rect 17548 65960 17588 66508
rect 17260 65920 17588 65960
rect 17260 65456 17300 65920
rect 17451 65540 17493 65549
rect 17451 65500 17452 65540
rect 17492 65500 17493 65540
rect 17451 65491 17493 65500
rect 17931 65540 17973 65549
rect 17931 65500 17932 65540
rect 17972 65500 17973 65540
rect 17931 65491 17973 65500
rect 17300 65416 17396 65456
rect 17260 65407 17300 65416
rect 16684 64240 16916 64280
rect 16779 64112 16821 64121
rect 16779 64072 16780 64112
rect 16820 64072 16821 64112
rect 16779 64063 16821 64072
rect 16395 63944 16437 63953
rect 16395 63904 16396 63944
rect 16436 63904 16437 63944
rect 16395 63895 16437 63904
rect 16492 63944 16532 63953
rect 16780 63944 16820 64063
rect 16532 63904 16628 63944
rect 16492 63895 16532 63904
rect 16396 63810 16436 63895
rect 16491 63776 16533 63785
rect 16491 63736 16492 63776
rect 16532 63736 16533 63776
rect 16491 63727 16533 63736
rect 16492 63642 16532 63727
rect 16204 63484 16340 63524
rect 16011 62432 16053 62441
rect 16011 62392 16012 62432
rect 16052 62392 16053 62432
rect 16011 62383 16053 62392
rect 16011 62180 16053 62189
rect 16011 62140 16012 62180
rect 16052 62140 16053 62180
rect 16011 62131 16053 62140
rect 16012 62046 16052 62131
rect 15916 61888 16052 61928
rect 15819 61760 15861 61769
rect 15819 61720 15820 61760
rect 15860 61720 15861 61760
rect 15819 61711 15861 61720
rect 15723 61676 15765 61685
rect 15723 61636 15724 61676
rect 15764 61636 15765 61676
rect 15723 61627 15765 61636
rect 15819 61592 15861 61601
rect 15532 61531 15764 61571
rect 15819 61552 15820 61592
rect 15860 61552 15861 61592
rect 15819 61543 15861 61552
rect 15916 61592 15956 61601
rect 15436 61517 15476 61531
rect 15435 61508 15477 61517
rect 15435 61468 15436 61508
rect 15476 61468 15477 61508
rect 15435 61459 15477 61468
rect 15436 61436 15476 61459
rect 15724 61433 15764 61531
rect 15532 61424 15572 61433
rect 15435 61340 15477 61349
rect 15435 61300 15436 61340
rect 15476 61300 15477 61340
rect 15532 61340 15572 61384
rect 15723 61424 15765 61433
rect 15723 61384 15724 61424
rect 15764 61384 15765 61424
rect 15723 61375 15765 61384
rect 15627 61340 15669 61349
rect 15532 61300 15628 61340
rect 15668 61300 15669 61340
rect 15435 61291 15477 61300
rect 15627 61291 15669 61300
rect 15339 61172 15381 61181
rect 15339 61132 15340 61172
rect 15380 61132 15381 61172
rect 15339 61123 15381 61132
rect 15436 60906 15476 61291
rect 15724 61290 15764 61375
rect 15820 61172 15860 61543
rect 15916 61265 15956 61552
rect 15915 61256 15957 61265
rect 15915 61216 15916 61256
rect 15956 61216 15957 61256
rect 15915 61207 15957 61216
rect 15724 61132 15860 61172
rect 15627 61088 15669 61097
rect 15627 61048 15628 61088
rect 15668 61048 15669 61088
rect 15627 61039 15669 61048
rect 15628 60954 15668 61039
rect 15243 59240 15285 59249
rect 15243 59200 15244 59240
rect 15284 59200 15285 59240
rect 15243 59191 15285 59200
rect 15147 58568 15189 58577
rect 15147 58528 15148 58568
rect 15188 58528 15189 58568
rect 15147 58519 15189 58528
rect 15244 56972 15284 59191
rect 15436 58661 15476 60866
rect 15627 60584 15669 60593
rect 15627 60544 15628 60584
rect 15668 60544 15669 60584
rect 15627 60535 15669 60544
rect 15628 60080 15668 60535
rect 15628 60031 15668 60040
rect 15531 58736 15573 58745
rect 15531 58696 15532 58736
rect 15572 58696 15573 58736
rect 15531 58687 15573 58696
rect 15435 58652 15477 58661
rect 15435 58612 15436 58652
rect 15476 58612 15477 58652
rect 15435 58603 15477 58612
rect 15532 58602 15572 58687
rect 15340 58568 15380 58577
rect 15340 57821 15380 58528
rect 15724 58400 15764 61132
rect 16012 61097 16052 61888
rect 16011 61088 16053 61097
rect 16011 61048 16012 61088
rect 16052 61048 16053 61088
rect 16011 61039 16053 61048
rect 15820 60929 15860 61014
rect 16204 61004 16244 63484
rect 16299 63356 16341 63365
rect 16299 63316 16300 63356
rect 16340 63316 16341 63356
rect 16299 63307 16341 63316
rect 16300 63104 16340 63307
rect 16300 63055 16340 63064
rect 16491 63104 16533 63113
rect 16491 63064 16492 63104
rect 16532 63064 16533 63104
rect 16491 63055 16533 63064
rect 16492 62970 16532 63055
rect 16395 62768 16437 62777
rect 16395 62728 16396 62768
rect 16436 62728 16437 62768
rect 16395 62719 16437 62728
rect 16204 60964 16340 61004
rect 15819 60920 15861 60929
rect 16012 60920 16052 60929
rect 15819 60880 15820 60920
rect 15860 60880 15861 60920
rect 15819 60871 15861 60880
rect 15916 60880 16012 60920
rect 15819 60668 15861 60677
rect 15819 60628 15820 60668
rect 15860 60628 15861 60668
rect 15819 60619 15861 60628
rect 15820 60534 15860 60619
rect 15820 60080 15860 60089
rect 15820 59921 15860 60040
rect 15819 59912 15861 59921
rect 15819 59872 15820 59912
rect 15860 59872 15861 59912
rect 15819 59863 15861 59872
rect 15820 58400 15860 58409
rect 15724 58360 15820 58400
rect 15820 58351 15860 58360
rect 15916 58064 15956 60880
rect 16012 60871 16052 60880
rect 16108 60920 16148 60929
rect 16012 59408 16052 59417
rect 16012 58997 16052 59368
rect 16011 58988 16053 58997
rect 16011 58948 16012 58988
rect 16052 58948 16053 58988
rect 16011 58939 16053 58948
rect 16108 58829 16148 60880
rect 16300 60257 16340 60964
rect 16396 60929 16436 62719
rect 16588 62609 16628 63904
rect 16780 63895 16820 63904
rect 16779 63776 16821 63785
rect 16779 63736 16780 63776
rect 16820 63736 16821 63776
rect 16779 63727 16821 63736
rect 16780 63642 16820 63727
rect 16587 62600 16629 62609
rect 16587 62560 16588 62600
rect 16628 62560 16629 62600
rect 16587 62551 16629 62560
rect 16492 62432 16532 62441
rect 16532 62392 16820 62432
rect 16492 62383 16532 62392
rect 16491 62180 16533 62189
rect 16491 62140 16492 62180
rect 16532 62140 16533 62180
rect 16491 62131 16533 62140
rect 16395 60920 16437 60929
rect 16395 60880 16396 60920
rect 16436 60880 16437 60920
rect 16395 60871 16437 60880
rect 16396 60786 16436 60871
rect 16299 60248 16341 60257
rect 16299 60208 16300 60248
rect 16340 60208 16341 60248
rect 16299 60199 16341 60208
rect 16299 59408 16341 59417
rect 16299 59368 16300 59408
rect 16340 59368 16341 59408
rect 16299 59359 16341 59368
rect 16300 59274 16340 59359
rect 16107 58820 16149 58829
rect 16107 58780 16108 58820
rect 16148 58780 16149 58820
rect 16107 58771 16149 58780
rect 16011 58652 16053 58661
rect 16011 58612 16012 58652
rect 16052 58612 16053 58652
rect 16011 58603 16053 58612
rect 16012 58568 16052 58603
rect 16108 58577 16148 58662
rect 16012 58517 16052 58528
rect 16107 58568 16149 58577
rect 16107 58528 16108 58568
rect 16148 58528 16149 58568
rect 16107 58519 16149 58528
rect 16299 58568 16341 58577
rect 16299 58528 16300 58568
rect 16340 58528 16341 58568
rect 16299 58519 16341 58528
rect 16396 58568 16436 58577
rect 15916 58024 16052 58064
rect 16012 57905 16052 58024
rect 15916 57896 15956 57905
rect 15339 57812 15381 57821
rect 15339 57772 15340 57812
rect 15380 57772 15381 57812
rect 15339 57763 15381 57772
rect 15916 57569 15956 57856
rect 16011 57896 16053 57905
rect 16011 57856 16012 57896
rect 16052 57856 16053 57896
rect 16011 57847 16053 57856
rect 15915 57560 15957 57569
rect 15915 57520 15916 57560
rect 15956 57520 15957 57560
rect 15915 57511 15957 57520
rect 15339 57392 15381 57401
rect 15339 57352 15340 57392
rect 15380 57352 15381 57392
rect 15339 57343 15381 57352
rect 15340 57070 15380 57343
rect 15340 57021 15380 57030
rect 16012 57140 16052 57149
rect 15244 56932 15380 56972
rect 15244 56384 15284 56393
rect 15051 56300 15093 56309
rect 15051 56260 15052 56300
rect 15092 56260 15093 56300
rect 15051 56251 15093 56260
rect 15052 56166 15092 56251
rect 15244 56225 15284 56344
rect 15243 56216 15285 56225
rect 15243 56176 15244 56216
rect 15284 56176 15285 56216
rect 15243 56167 15285 56176
rect 15052 55544 15092 55553
rect 15052 55460 15092 55504
rect 14764 55420 14900 55460
rect 14956 55420 15092 55460
rect 14763 54956 14805 54965
rect 14763 54916 14764 54956
rect 14804 54916 14805 54956
rect 14763 54907 14805 54916
rect 14764 54822 14804 54907
rect 14860 54872 14900 55420
rect 15052 55133 15092 55420
rect 15051 55124 15093 55133
rect 15051 55084 15052 55124
rect 15092 55084 15093 55124
rect 15051 55075 15093 55084
rect 15052 54872 15092 54881
rect 14860 54832 15052 54872
rect 15052 54823 15092 54832
rect 15148 54872 15188 54883
rect 15148 54797 15188 54832
rect 15147 54788 15189 54797
rect 15147 54748 15148 54788
rect 15188 54748 15189 54788
rect 15147 54739 15189 54748
rect 15051 54536 15093 54545
rect 15051 54496 15052 54536
rect 15092 54496 15093 54536
rect 15051 54487 15093 54496
rect 15052 54209 15092 54487
rect 15051 54200 15093 54209
rect 15051 54160 15052 54200
rect 15092 54160 15093 54200
rect 15051 54151 15093 54160
rect 15052 54032 15092 54151
rect 15052 53983 15092 53992
rect 14763 53864 14805 53873
rect 15244 53864 15284 53873
rect 14763 53824 14764 53864
rect 14804 53824 14805 53864
rect 14763 53815 14805 53824
rect 15148 53824 15244 53864
rect 14476 53656 14708 53696
rect 14379 53528 14421 53537
rect 14379 53488 14380 53528
rect 14420 53488 14421 53528
rect 14379 53479 14421 53488
rect 14380 52436 14420 52445
rect 14284 52396 14380 52436
rect 14380 52387 14420 52396
rect 14092 51976 14420 52016
rect 14187 51848 14229 51857
rect 14187 51808 14188 51848
rect 14228 51808 14229 51848
rect 14187 51799 14229 51808
rect 13995 51008 14037 51017
rect 13995 50968 13996 51008
rect 14036 50968 14037 51008
rect 13995 50959 14037 50968
rect 13995 50420 14037 50429
rect 13995 50380 13996 50420
rect 14036 50380 14037 50420
rect 13995 50371 14037 50380
rect 13996 50336 14036 50371
rect 13996 50285 14036 50296
rect 13995 49664 14037 49673
rect 13995 49624 13996 49664
rect 14036 49624 14037 49664
rect 13995 49615 14037 49624
rect 13996 48833 14036 49615
rect 13995 48824 14037 48833
rect 13995 48784 13996 48824
rect 14036 48784 14037 48824
rect 13995 48775 14037 48784
rect 14188 47825 14228 51799
rect 14283 51008 14325 51017
rect 14283 50968 14284 51008
rect 14324 50968 14325 51008
rect 14283 50959 14325 50968
rect 14284 48824 14324 50959
rect 14284 48775 14324 48784
rect 14187 47816 14229 47825
rect 14187 47776 14188 47816
rect 14228 47776 14229 47816
rect 14187 47767 14229 47776
rect 13996 47312 14036 47323
rect 13996 47237 14036 47272
rect 13995 47228 14037 47237
rect 13995 47188 13996 47228
rect 14036 47188 14037 47228
rect 13995 47179 14037 47188
rect 14188 47060 14228 47069
rect 13900 47020 14036 47060
rect 13611 46556 13653 46565
rect 13611 46516 13612 46556
rect 13652 46516 13653 46556
rect 13611 46507 13653 46516
rect 13612 46472 13652 46507
rect 13612 46421 13652 46432
rect 13707 46388 13749 46397
rect 13707 46348 13708 46388
rect 13748 46348 13749 46388
rect 13707 46339 13749 46348
rect 13420 45751 13460 45760
rect 13323 45380 13365 45389
rect 13323 45340 13324 45380
rect 13364 45340 13365 45380
rect 13323 45331 13365 45340
rect 13708 45212 13748 46339
rect 13708 45163 13748 45172
rect 13228 45088 13652 45128
rect 13323 44960 13365 44969
rect 13323 44920 13324 44960
rect 13364 44920 13365 44960
rect 13323 44911 13365 44920
rect 13324 44826 13364 44911
rect 13516 44792 13556 44801
rect 13420 44752 13516 44792
rect 13324 44274 13364 44283
rect 13324 43625 13364 44234
rect 13323 43616 13365 43625
rect 13323 43576 13324 43616
rect 13364 43576 13365 43616
rect 13323 43567 13365 43576
rect 13276 43457 13316 43466
rect 13420 43448 13460 44752
rect 13516 44743 13556 44752
rect 13515 44624 13557 44633
rect 13515 44584 13516 44624
rect 13556 44584 13557 44624
rect 13515 44575 13557 44584
rect 13516 44456 13556 44575
rect 13516 44407 13556 44416
rect 13316 43417 13460 43448
rect 13276 43408 13460 43417
rect 13420 43280 13460 43289
rect 13132 43240 13420 43280
rect 13420 43231 13460 43240
rect 13612 42944 13652 45088
rect 13900 45044 13940 45053
rect 13803 44960 13845 44969
rect 13803 44920 13804 44960
rect 13844 44920 13845 44960
rect 13803 44911 13845 44920
rect 13707 44624 13749 44633
rect 13707 44584 13708 44624
rect 13748 44584 13749 44624
rect 13707 44575 13749 44584
rect 13708 44297 13748 44575
rect 13707 44288 13749 44297
rect 13707 44248 13708 44288
rect 13748 44248 13749 44288
rect 13707 44239 13749 44248
rect 13804 43784 13844 44911
rect 13900 44717 13940 45004
rect 13899 44708 13941 44717
rect 13899 44668 13900 44708
rect 13940 44668 13941 44708
rect 13899 44659 13941 44668
rect 13996 44540 14036 47020
rect 14188 46556 14228 47020
rect 14140 46516 14228 46556
rect 14140 46514 14180 46516
rect 14140 46465 14180 46474
rect 14284 46304 14324 46313
rect 13900 44500 14036 44540
rect 14092 46264 14284 46304
rect 13900 44372 13940 44500
rect 13899 44332 13940 44372
rect 13899 44204 13939 44332
rect 13996 44330 14036 44383
rect 13995 44290 13996 44297
rect 14036 44290 14037 44297
rect 13995 44288 14037 44290
rect 13995 44248 13996 44288
rect 14036 44248 14037 44288
rect 13995 44239 14037 44248
rect 13899 44164 13940 44204
rect 13900 44120 13940 44164
rect 13900 44080 14036 44120
rect 13516 42904 13652 42944
rect 13708 43744 13844 43784
rect 12939 41936 12981 41945
rect 12939 41896 12940 41936
rect 12980 41896 12981 41936
rect 12939 41887 12981 41896
rect 12555 41768 12597 41777
rect 12555 41728 12556 41768
rect 12596 41728 12597 41768
rect 12555 41719 12597 41728
rect 12939 41432 12981 41441
rect 12939 41392 12940 41432
rect 12980 41392 12981 41432
rect 12939 41383 12981 41392
rect 12940 41298 12980 41383
rect 12363 41264 12405 41273
rect 12363 41224 12364 41264
rect 12404 41224 12405 41264
rect 12363 41215 12405 41224
rect 12748 41180 12788 41189
rect 12748 40349 12788 41140
rect 13227 40676 13269 40685
rect 13227 40636 13228 40676
rect 13268 40636 13269 40676
rect 13227 40627 13269 40636
rect 13228 40542 13268 40627
rect 13035 40508 13077 40517
rect 13035 40468 13036 40508
rect 13076 40468 13077 40508
rect 13035 40459 13077 40468
rect 13036 40374 13076 40459
rect 12747 40340 12789 40349
rect 12747 40300 12748 40340
rect 12788 40300 12789 40340
rect 12747 40291 12789 40300
rect 12844 39880 13076 39920
rect 12652 39752 12692 39761
rect 12652 37745 12692 39712
rect 12844 39752 12884 39880
rect 12844 39703 12884 39712
rect 12940 39752 12980 39761
rect 12843 39584 12885 39593
rect 12843 39544 12844 39584
rect 12884 39544 12885 39584
rect 12843 39535 12885 39544
rect 12844 39450 12884 39535
rect 12747 39248 12789 39257
rect 12747 39208 12748 39248
rect 12788 39208 12789 39248
rect 12747 39199 12789 39208
rect 12748 38954 12788 39199
rect 12940 39164 12980 39712
rect 12940 39005 12980 39124
rect 12939 38996 12981 39005
rect 12748 38240 12788 38914
rect 12748 38191 12788 38200
rect 12844 38956 12940 38996
rect 12980 38956 12981 38996
rect 12747 37988 12789 37997
rect 12747 37948 12748 37988
rect 12788 37948 12789 37988
rect 12747 37939 12789 37948
rect 12651 37736 12693 37745
rect 12651 37696 12652 37736
rect 12692 37696 12693 37736
rect 12651 37687 12693 37696
rect 12556 37568 12596 37577
rect 12364 37528 12556 37568
rect 12171 37484 12213 37493
rect 12171 37444 12172 37484
rect 12212 37444 12213 37484
rect 12171 37435 12213 37444
rect 12076 37400 12116 37409
rect 12076 36989 12116 37360
rect 12268 37400 12308 37409
rect 12171 37316 12213 37325
rect 12171 37276 12172 37316
rect 12212 37276 12213 37316
rect 12171 37267 12213 37276
rect 12172 37182 12212 37267
rect 12075 36980 12117 36989
rect 12075 36940 12076 36980
rect 12116 36940 12117 36980
rect 12075 36931 12117 36940
rect 12268 36905 12308 37360
rect 12364 37400 12404 37528
rect 12364 37351 12404 37360
rect 12460 37148 12500 37528
rect 12556 37519 12596 37528
rect 12555 37400 12597 37409
rect 12748 37400 12788 37939
rect 12555 37360 12556 37400
rect 12596 37360 12788 37400
rect 12555 37351 12597 37360
rect 12556 37266 12596 37351
rect 12460 37108 12596 37148
rect 12267 36896 12309 36905
rect 12267 36856 12268 36896
rect 12308 36856 12309 36896
rect 12267 36847 12309 36856
rect 12364 36896 12404 36905
rect 12172 36728 12212 36737
rect 11980 36688 12172 36728
rect 12172 36679 12212 36688
rect 12268 36728 12308 36737
rect 11980 36560 12020 36569
rect 11884 36520 11980 36560
rect 11980 36511 12020 36520
rect 11788 36436 11924 36476
rect 11884 36140 11924 36436
rect 12268 36149 12308 36688
rect 12267 36140 12309 36149
rect 11884 36100 12212 36140
rect 11787 35888 11829 35897
rect 11787 35848 11788 35888
rect 11828 35848 11829 35888
rect 11787 35839 11829 35848
rect 11884 35888 11924 36100
rect 12172 36056 12212 36100
rect 12267 36100 12268 36140
rect 12308 36100 12309 36140
rect 12267 36091 12309 36100
rect 12172 36016 12217 36056
rect 12076 35897 12116 35982
rect 12177 35905 12217 36016
rect 12268 36006 12308 36091
rect 11884 35839 11924 35848
rect 12075 35888 12117 35897
rect 12075 35848 12076 35888
rect 12116 35848 12117 35888
rect 12177 35888 12308 35905
rect 12177 35865 12268 35888
rect 12075 35839 12117 35848
rect 12364 35888 12404 36856
rect 12460 36728 12500 36737
rect 12460 36569 12500 36688
rect 12556 36728 12596 37108
rect 12651 37064 12693 37073
rect 12651 37024 12652 37064
rect 12692 37024 12693 37064
rect 12651 37015 12693 37024
rect 12652 36737 12692 37015
rect 12652 36728 12697 36737
rect 12652 36688 12657 36728
rect 12556 36679 12596 36688
rect 12657 36679 12697 36688
rect 12748 36653 12788 37360
rect 12844 37400 12884 38956
rect 12939 38947 12981 38956
rect 12940 38408 12980 38417
rect 13036 38408 13076 39880
rect 13227 39584 13269 39593
rect 13227 39544 13228 39584
rect 13268 39544 13269 39584
rect 13227 39535 13269 39544
rect 13131 38996 13173 39005
rect 13131 38956 13132 38996
rect 13172 38956 13173 38996
rect 13131 38947 13173 38956
rect 13132 38912 13172 38947
rect 13132 38861 13172 38872
rect 12980 38368 13076 38408
rect 12940 38359 12980 38368
rect 13035 38240 13077 38249
rect 13035 38200 13036 38240
rect 13076 38200 13077 38240
rect 13035 38191 13077 38200
rect 13132 38240 13172 38249
rect 13228 38240 13268 39535
rect 13420 38921 13460 39006
rect 13419 38912 13461 38921
rect 13419 38872 13420 38912
rect 13460 38872 13461 38912
rect 13419 38863 13461 38872
rect 13324 38744 13364 38753
rect 13364 38704 13460 38744
rect 13324 38695 13364 38704
rect 13324 38240 13364 38249
rect 13228 38200 13324 38240
rect 12940 37997 12980 38082
rect 12939 37988 12981 37997
rect 12939 37948 12940 37988
rect 12980 37948 12981 37988
rect 12939 37939 12981 37948
rect 13036 37568 13076 38191
rect 13132 37913 13172 38200
rect 13324 38191 13364 38200
rect 13420 38240 13460 38704
rect 13516 38249 13556 42904
rect 13612 42776 13652 42785
rect 13708 42776 13748 43744
rect 13803 43616 13845 43625
rect 13803 43576 13804 43616
rect 13844 43576 13845 43616
rect 13803 43567 13845 43576
rect 13804 42860 13844 43567
rect 13899 43448 13941 43457
rect 13899 43408 13900 43448
rect 13940 43408 13941 43448
rect 13899 43399 13941 43408
rect 13900 43280 13940 43399
rect 13900 43231 13940 43240
rect 13804 42811 13844 42820
rect 13652 42736 13748 42776
rect 13612 42727 13652 42736
rect 13804 38324 13844 38333
rect 13420 38191 13460 38200
rect 13515 38240 13557 38249
rect 13515 38200 13516 38240
rect 13556 38200 13557 38240
rect 13515 38191 13557 38200
rect 13612 38240 13652 38249
rect 13420 38072 13460 38081
rect 13612 38072 13652 38200
rect 13460 38032 13652 38072
rect 13708 38240 13748 38249
rect 13420 38023 13460 38032
rect 13131 37904 13173 37913
rect 13131 37864 13132 37904
rect 13172 37864 13173 37904
rect 13131 37855 13173 37864
rect 13323 37904 13365 37913
rect 13323 37864 13324 37904
rect 13364 37864 13365 37904
rect 13323 37855 13365 37864
rect 13515 37904 13557 37913
rect 13515 37864 13516 37904
rect 13556 37864 13557 37904
rect 13515 37855 13557 37864
rect 13036 37528 13268 37568
rect 12844 37241 12884 37360
rect 13036 37400 13076 37411
rect 13036 37325 13076 37360
rect 13132 37400 13172 37409
rect 13035 37316 13077 37325
rect 13035 37276 13036 37316
rect 13076 37276 13077 37316
rect 13035 37267 13077 37276
rect 12843 37232 12885 37241
rect 12843 37192 12844 37232
rect 12884 37192 12885 37232
rect 12843 37183 12885 37192
rect 12844 36821 12884 37183
rect 13035 36896 13077 36905
rect 13035 36856 13036 36896
rect 13076 36856 13077 36896
rect 13035 36847 13077 36856
rect 12843 36812 12885 36821
rect 12843 36772 12844 36812
rect 12884 36772 12885 36812
rect 12843 36763 12885 36772
rect 13036 36762 13076 36847
rect 12939 36728 12981 36737
rect 12939 36688 12940 36728
rect 12980 36688 12981 36728
rect 12939 36679 12981 36688
rect 12747 36644 12789 36653
rect 12747 36604 12748 36644
rect 12788 36604 12789 36644
rect 12747 36595 12789 36604
rect 12459 36560 12501 36569
rect 12459 36520 12460 36560
rect 12500 36520 12501 36560
rect 12459 36511 12501 36520
rect 12748 36224 12788 36595
rect 12940 36594 12980 36679
rect 12556 36184 12788 36224
rect 12556 35897 12596 36184
rect 12843 36140 12885 36149
rect 12843 36100 12844 36140
rect 12884 36100 12885 36140
rect 12843 36091 12885 36100
rect 12651 36056 12693 36065
rect 12651 36016 12652 36056
rect 12692 36016 12693 36056
rect 12651 36007 12693 36016
rect 12555 35888 12597 35897
rect 12364 35848 12500 35888
rect 12268 35839 12308 35848
rect 11788 35754 11828 35839
rect 12076 35720 12116 35729
rect 12116 35680 12308 35720
rect 12076 35671 12116 35680
rect 11596 35596 11732 35636
rect 11787 35636 11829 35645
rect 11787 35596 11788 35636
rect 11828 35596 12020 35636
rect 11404 35512 11540 35552
rect 11307 35503 11349 35512
rect 11211 33872 11253 33881
rect 11211 33832 11212 33872
rect 11252 33832 11253 33872
rect 11211 33823 11253 33832
rect 11211 33704 11253 33713
rect 11211 33664 11212 33704
rect 11252 33664 11253 33704
rect 11211 33655 11253 33664
rect 11212 33570 11252 33655
rect 11308 33536 11348 35503
rect 11404 35225 11444 35310
rect 11403 35216 11445 35225
rect 11403 35176 11404 35216
rect 11444 35176 11445 35216
rect 11403 35167 11445 35176
rect 11500 35141 11540 35512
rect 11499 35132 11541 35141
rect 11499 35092 11500 35132
rect 11540 35092 11541 35132
rect 11499 35083 11541 35092
rect 11403 35048 11445 35057
rect 11403 35008 11404 35048
rect 11444 35008 11445 35048
rect 11403 34999 11445 35008
rect 11404 33872 11444 34999
rect 11499 34964 11541 34973
rect 11499 34924 11500 34964
rect 11540 34924 11541 34964
rect 11499 34915 11541 34924
rect 11404 33713 11444 33832
rect 11403 33704 11445 33713
rect 11403 33664 11404 33704
rect 11444 33664 11445 33704
rect 11500 33704 11540 34915
rect 11596 34553 11636 35596
rect 11787 35587 11829 35596
rect 11980 35384 12020 35596
rect 12268 35468 12308 35680
rect 12268 35428 12404 35468
rect 11980 35344 12308 35384
rect 11883 35300 11925 35309
rect 11883 35260 11884 35300
rect 11924 35260 11925 35300
rect 11883 35251 11925 35260
rect 11692 35216 11732 35225
rect 11595 34544 11637 34553
rect 11595 34504 11596 34544
rect 11636 34504 11637 34544
rect 11595 34495 11637 34504
rect 11595 34376 11637 34385
rect 11595 34336 11596 34376
rect 11636 34336 11637 34376
rect 11595 34327 11637 34336
rect 11596 34242 11636 34327
rect 11692 34133 11732 35176
rect 11787 35216 11829 35225
rect 11787 35176 11788 35216
rect 11828 35176 11829 35216
rect 11787 35167 11829 35176
rect 11788 35082 11828 35167
rect 11884 34133 11924 35251
rect 12075 35216 12117 35225
rect 12075 35176 12076 35216
rect 12116 35176 12117 35216
rect 12075 35167 12117 35176
rect 12268 35216 12308 35344
rect 12268 35167 12308 35176
rect 12364 35216 12404 35428
rect 12364 35167 12404 35176
rect 12460 35216 12500 35848
rect 12555 35848 12556 35888
rect 12596 35848 12597 35888
rect 12555 35839 12597 35848
rect 12556 35754 12596 35839
rect 12556 35300 12596 35309
rect 12652 35300 12692 36007
rect 12748 35888 12788 35897
rect 12748 35729 12788 35848
rect 12844 35888 12884 36091
rect 12939 35972 12981 35981
rect 12939 35932 12940 35972
rect 12980 35932 12981 35972
rect 12939 35923 12981 35932
rect 12844 35839 12884 35848
rect 12747 35720 12789 35729
rect 12747 35680 12748 35720
rect 12788 35680 12789 35720
rect 12747 35671 12789 35680
rect 12940 35384 12980 35923
rect 13036 35720 13076 35729
rect 13132 35720 13172 37360
rect 13228 36905 13268 37528
rect 13324 37400 13364 37855
rect 13324 37351 13364 37360
rect 13324 37232 13364 37241
rect 13516 37232 13556 37855
rect 13611 37652 13653 37661
rect 13611 37612 13612 37652
rect 13652 37612 13653 37652
rect 13611 37603 13653 37612
rect 13612 37400 13652 37603
rect 13612 37351 13652 37360
rect 13364 37192 13460 37232
rect 13516 37192 13652 37232
rect 13324 37183 13364 37192
rect 13323 37064 13365 37073
rect 13323 37024 13324 37064
rect 13364 37024 13365 37064
rect 13323 37015 13365 37024
rect 13227 36896 13269 36905
rect 13227 36856 13228 36896
rect 13268 36856 13269 36896
rect 13227 36847 13269 36856
rect 13228 36728 13268 36737
rect 13228 36065 13268 36688
rect 13324 36644 13364 37015
rect 13420 36896 13460 37192
rect 13420 36856 13556 36896
rect 13324 36595 13364 36604
rect 13516 36644 13556 36856
rect 13612 36728 13652 37192
rect 13708 36896 13748 38200
rect 13804 37073 13844 38284
rect 13899 38240 13941 38249
rect 13899 38200 13900 38240
rect 13940 38200 13941 38240
rect 13899 38191 13941 38200
rect 13900 37913 13940 38191
rect 13899 37904 13941 37913
rect 13899 37864 13900 37904
rect 13940 37864 13941 37904
rect 13899 37855 13941 37864
rect 13803 37064 13845 37073
rect 13803 37024 13804 37064
rect 13844 37024 13845 37064
rect 13803 37015 13845 37024
rect 13804 36896 13844 36905
rect 13708 36856 13804 36896
rect 13996 36896 14036 44080
rect 14092 43532 14132 46264
rect 14284 46255 14324 46264
rect 14187 45128 14229 45137
rect 14187 45088 14188 45128
rect 14228 45088 14229 45128
rect 14187 45079 14229 45088
rect 14188 44297 14228 45079
rect 14187 44288 14229 44297
rect 14187 44248 14188 44288
rect 14228 44248 14229 44288
rect 14187 44239 14229 44248
rect 14092 43483 14132 43492
rect 14380 39089 14420 51976
rect 14476 50849 14516 53656
rect 14764 53612 14804 53815
rect 14668 53572 14804 53612
rect 14571 53444 14613 53453
rect 14571 53404 14572 53444
rect 14612 53404 14613 53444
rect 14571 53395 14613 53404
rect 14572 52520 14612 53395
rect 14475 50840 14517 50849
rect 14475 50800 14476 50840
rect 14516 50800 14517 50840
rect 14475 50791 14517 50800
rect 14475 50336 14517 50345
rect 14475 50296 14476 50336
rect 14516 50296 14517 50336
rect 14475 50287 14517 50296
rect 14476 47993 14516 50287
rect 14572 49673 14612 52480
rect 14571 49664 14613 49673
rect 14571 49624 14572 49664
rect 14612 49624 14613 49664
rect 14571 49615 14613 49624
rect 14572 49169 14612 49615
rect 14571 49160 14613 49169
rect 14571 49120 14572 49160
rect 14612 49120 14613 49160
rect 14571 49111 14613 49120
rect 14571 48572 14613 48581
rect 14571 48532 14572 48572
rect 14612 48532 14613 48572
rect 14571 48523 14613 48532
rect 14475 47984 14517 47993
rect 14475 47944 14476 47984
rect 14516 47944 14517 47984
rect 14475 47935 14517 47944
rect 14475 47816 14517 47825
rect 14475 47776 14476 47816
rect 14516 47776 14517 47816
rect 14475 47767 14517 47776
rect 14476 39257 14516 47767
rect 14572 40685 14612 48523
rect 14668 46640 14708 53572
rect 15148 53360 15188 53824
rect 15244 53815 15284 53824
rect 15148 53311 15188 53320
rect 15244 53360 15284 53369
rect 15147 53024 15189 53033
rect 15147 52984 15148 53024
rect 15188 52984 15189 53024
rect 15147 52975 15189 52984
rect 14763 51848 14805 51857
rect 14763 51808 14764 51848
rect 14804 51808 14805 51848
rect 14763 51799 14805 51808
rect 14764 51714 14804 51799
rect 14956 51596 14996 51605
rect 14860 51556 14956 51596
rect 14860 51092 14900 51556
rect 14956 51547 14996 51556
rect 15148 51101 15188 52975
rect 15244 51857 15284 53320
rect 15243 51848 15285 51857
rect 15243 51808 15244 51848
rect 15284 51808 15285 51848
rect 15243 51799 15285 51808
rect 14812 51052 14900 51092
rect 15147 51092 15189 51101
rect 15147 51052 15148 51092
rect 15188 51052 15189 51092
rect 14812 51050 14852 51052
rect 15147 51043 15189 51052
rect 14812 51001 14852 51010
rect 15243 51008 15285 51017
rect 15243 50968 15244 51008
rect 15284 50968 15285 51008
rect 15243 50959 15285 50968
rect 14955 50840 14997 50849
rect 14955 50800 14956 50840
rect 14996 50800 14997 50840
rect 14955 50791 14997 50800
rect 14956 50706 14996 50791
rect 15244 50336 15284 50959
rect 15244 50287 15284 50296
rect 14763 49748 14805 49757
rect 14763 49708 14764 49748
rect 14804 49708 14805 49748
rect 14763 49699 14805 49708
rect 14764 49496 14804 49699
rect 15340 49664 15380 56932
rect 15532 56888 15572 56897
rect 15532 56309 15572 56848
rect 15820 56888 15860 56897
rect 15627 56468 15669 56477
rect 15627 56428 15628 56468
rect 15668 56428 15669 56468
rect 15627 56419 15669 56428
rect 15531 56300 15573 56309
rect 15531 56260 15532 56300
rect 15572 56260 15573 56300
rect 15531 56251 15573 56260
rect 15531 54872 15573 54881
rect 15531 54832 15532 54872
rect 15572 54832 15573 54872
rect 15531 54823 15573 54832
rect 15628 54872 15668 56419
rect 15820 55553 15860 56848
rect 15915 56300 15957 56309
rect 15915 56260 15916 56300
rect 15956 56260 15957 56300
rect 15915 56251 15957 56260
rect 15819 55544 15861 55553
rect 15819 55504 15820 55544
rect 15860 55504 15861 55544
rect 15819 55495 15861 55504
rect 15532 54738 15572 54823
rect 15531 54452 15573 54461
rect 15531 54412 15532 54452
rect 15572 54412 15573 54452
rect 15531 54403 15573 54412
rect 15532 54032 15572 54403
rect 15436 53992 15532 54032
rect 15436 50429 15476 53992
rect 15532 53983 15572 53992
rect 15628 53864 15668 54832
rect 15819 54032 15861 54041
rect 15819 53992 15820 54032
rect 15860 53992 15861 54032
rect 15819 53983 15861 53992
rect 15532 53824 15668 53864
rect 15435 50420 15477 50429
rect 15435 50380 15436 50420
rect 15476 50380 15477 50420
rect 15435 50371 15477 50380
rect 15244 49624 15380 49664
rect 15436 50084 15476 50093
rect 15051 49580 15093 49589
rect 15051 49540 15052 49580
rect 15092 49540 15093 49580
rect 15051 49531 15093 49540
rect 14764 49447 14804 49456
rect 14956 49328 14996 49337
rect 14860 49288 14956 49328
rect 14860 48824 14900 49288
rect 14956 49279 14996 49288
rect 14956 48992 14996 49001
rect 15052 48992 15092 49531
rect 15147 49412 15189 49421
rect 15147 49372 15148 49412
rect 15188 49372 15189 49412
rect 15147 49363 15189 49372
rect 14996 48952 15092 48992
rect 14956 48943 14996 48952
rect 14812 48814 14900 48824
rect 14852 48784 14900 48814
rect 14812 48765 14852 48774
rect 14859 47984 14901 47993
rect 14859 47944 14860 47984
rect 14900 47944 14901 47984
rect 14859 47935 14901 47944
rect 14668 46600 14804 46640
rect 14667 46304 14709 46313
rect 14667 46264 14668 46304
rect 14708 46264 14709 46304
rect 14667 46255 14709 46264
rect 14668 45800 14708 46255
rect 14668 44969 14708 45760
rect 14667 44960 14709 44969
rect 14667 44920 14668 44960
rect 14708 44920 14709 44960
rect 14667 44911 14709 44920
rect 14571 40676 14613 40685
rect 14571 40636 14572 40676
rect 14612 40636 14613 40676
rect 14571 40627 14613 40636
rect 14571 39584 14613 39593
rect 14571 39544 14572 39584
rect 14612 39544 14613 39584
rect 14571 39535 14613 39544
rect 14475 39248 14517 39257
rect 14475 39208 14476 39248
rect 14516 39208 14517 39248
rect 14475 39199 14517 39208
rect 14379 39080 14421 39089
rect 14379 39040 14380 39080
rect 14420 39040 14421 39080
rect 14379 39031 14421 39040
rect 14476 38996 14516 39005
rect 14091 38240 14133 38249
rect 14091 38200 14092 38240
rect 14132 38200 14133 38240
rect 14091 38191 14133 38200
rect 14188 38240 14228 38249
rect 14092 38106 14132 38191
rect 14188 37997 14228 38200
rect 14380 38156 14420 38165
rect 14187 37988 14229 37997
rect 14187 37948 14188 37988
rect 14228 37948 14229 37988
rect 14187 37939 14229 37948
rect 14380 37577 14420 38116
rect 14476 37829 14516 38956
rect 14572 38408 14612 39535
rect 14667 38744 14709 38753
rect 14667 38704 14668 38744
rect 14708 38704 14709 38744
rect 14667 38695 14709 38704
rect 14668 38610 14708 38695
rect 14572 38359 14612 38368
rect 14475 37820 14517 37829
rect 14764 37820 14804 46600
rect 14860 46313 14900 47935
rect 15052 47816 15092 47825
rect 15052 47312 15092 47776
rect 15052 47263 15092 47272
rect 15148 47312 15188 49363
rect 15244 49328 15284 49624
rect 15436 49580 15476 50044
rect 15532 49589 15572 53824
rect 15723 53360 15765 53369
rect 15723 53320 15724 53360
rect 15764 53320 15765 53360
rect 15723 53311 15765 53320
rect 15627 53276 15669 53285
rect 15627 53236 15628 53276
rect 15668 53236 15669 53276
rect 15627 53227 15669 53236
rect 15628 53142 15668 53227
rect 15724 53226 15764 53311
rect 15820 53117 15860 53983
rect 15819 53108 15861 53117
rect 15819 53068 15820 53108
rect 15860 53068 15861 53108
rect 15819 53059 15861 53068
rect 15820 52520 15860 53059
rect 15916 52520 15956 56251
rect 16012 55469 16052 57100
rect 16011 55460 16053 55469
rect 16011 55420 16012 55460
rect 16052 55420 16053 55460
rect 16108 55460 16148 58519
rect 16300 58434 16340 58519
rect 16396 57653 16436 58528
rect 16492 58568 16532 62131
rect 16587 61088 16629 61097
rect 16587 61048 16588 61088
rect 16628 61048 16629 61088
rect 16587 61039 16629 61048
rect 16588 59501 16628 61039
rect 16683 60920 16725 60929
rect 16683 60880 16684 60920
rect 16724 60880 16725 60920
rect 16683 60871 16725 60880
rect 16587 59492 16629 59501
rect 16587 59452 16588 59492
rect 16628 59452 16629 59492
rect 16587 59443 16629 59452
rect 16587 58820 16629 58829
rect 16587 58780 16588 58820
rect 16628 58780 16629 58820
rect 16587 58771 16629 58780
rect 16492 58519 16532 58528
rect 16588 58568 16628 58771
rect 16588 58519 16628 58528
rect 16395 57644 16437 57653
rect 16395 57604 16396 57644
rect 16436 57604 16437 57644
rect 16395 57595 16437 57604
rect 16299 57308 16341 57317
rect 16299 57268 16300 57308
rect 16340 57268 16341 57308
rect 16299 57259 16341 57268
rect 16300 57174 16340 57259
rect 16492 57140 16532 57149
rect 16396 57100 16492 57140
rect 16299 56384 16341 56393
rect 16396 56384 16436 57100
rect 16492 57091 16532 57100
rect 16684 56720 16724 60871
rect 16780 59072 16820 62392
rect 16876 59249 16916 64240
rect 17068 64240 17204 64280
rect 16971 63692 17013 63701
rect 16971 63652 16972 63692
rect 17012 63652 17013 63692
rect 16971 63643 17013 63652
rect 16972 63558 17012 63643
rect 16971 60920 17013 60929
rect 16971 60880 16972 60920
rect 17012 60880 17013 60920
rect 16971 60871 17013 60880
rect 16972 60080 17012 60871
rect 17068 60248 17108 64240
rect 17356 64112 17396 65416
rect 17452 64616 17492 65491
rect 17740 65442 17780 65451
rect 17932 65406 17972 65491
rect 17644 64868 17684 64877
rect 17740 64868 17780 65402
rect 17835 65288 17877 65297
rect 17835 65248 17836 65288
rect 17876 65248 17877 65288
rect 17835 65239 17877 65248
rect 17684 64828 17780 64868
rect 17644 64819 17684 64828
rect 17452 64567 17492 64576
rect 17836 64616 17876 65239
rect 17836 64567 17876 64576
rect 17451 64448 17493 64457
rect 17451 64408 17452 64448
rect 17492 64408 17493 64448
rect 17451 64399 17493 64408
rect 17931 64448 17973 64457
rect 17931 64408 17932 64448
rect 17972 64408 17973 64448
rect 17931 64399 17973 64408
rect 17356 64063 17396 64072
rect 17350 63944 17392 63953
rect 17350 63904 17351 63944
rect 17391 63904 17392 63944
rect 17350 63895 17392 63904
rect 17452 63944 17492 64399
rect 17932 64314 17972 64399
rect 18028 64373 18068 66928
rect 18219 65456 18261 65465
rect 18219 65416 18220 65456
rect 18260 65416 18261 65456
rect 18219 65407 18261 65416
rect 18027 64364 18069 64373
rect 18027 64324 18028 64364
rect 18068 64324 18069 64364
rect 18027 64315 18069 64324
rect 18028 64112 18068 64121
rect 17740 64072 18028 64112
rect 17643 64028 17685 64037
rect 17643 63988 17644 64028
rect 17684 63988 17685 64028
rect 17643 63979 17685 63988
rect 17452 63895 17492 63904
rect 17548 63944 17588 63953
rect 17351 63810 17391 63895
rect 17548 63365 17588 63904
rect 17644 63776 17684 63979
rect 17740 63944 17780 64072
rect 18028 64063 18068 64072
rect 17740 63895 17780 63904
rect 17836 63944 17876 63953
rect 18220 63944 18260 65407
rect 18316 64280 18356 67516
rect 18412 66128 18452 66137
rect 18412 64961 18452 66088
rect 18604 65381 18644 67600
rect 18603 65372 18645 65381
rect 18603 65332 18604 65372
rect 18644 65332 18645 65372
rect 18603 65323 18645 65332
rect 18411 64952 18453 64961
rect 18411 64912 18412 64952
rect 18452 64912 18453 64952
rect 18411 64903 18453 64912
rect 18604 64280 18644 65323
rect 18316 64240 18452 64280
rect 17876 63904 18164 63944
rect 17836 63895 17876 63904
rect 18027 63776 18069 63785
rect 17644 63736 17876 63776
rect 17547 63356 17589 63365
rect 17547 63316 17548 63356
rect 17588 63316 17589 63356
rect 17547 63307 17589 63316
rect 17740 63104 17780 63113
rect 17740 62432 17780 63064
rect 17836 62432 17876 63736
rect 18027 63736 18028 63776
rect 18068 63736 18069 63776
rect 18027 63727 18069 63736
rect 17931 63356 17973 63365
rect 17931 63316 17932 63356
rect 17972 63316 17973 63356
rect 17931 63307 17973 63316
rect 17932 63222 17972 63307
rect 17931 63104 17973 63113
rect 17931 63064 17932 63104
rect 17972 63064 17973 63104
rect 17931 63055 17973 63064
rect 17932 62600 17972 63055
rect 17932 62551 17972 62560
rect 17836 62392 17972 62432
rect 17164 61592 17204 61601
rect 17164 61349 17204 61552
rect 17451 61424 17493 61433
rect 17451 61384 17452 61424
rect 17492 61384 17493 61424
rect 17451 61375 17493 61384
rect 17163 61340 17205 61349
rect 17163 61300 17164 61340
rect 17204 61300 17205 61340
rect 17163 61291 17205 61300
rect 17068 60208 17204 60248
rect 17068 60080 17108 60089
rect 16972 60040 17068 60080
rect 16875 59240 16917 59249
rect 16875 59200 16876 59240
rect 16916 59200 16917 59240
rect 16875 59191 16917 59200
rect 16972 59156 17012 59165
rect 16780 59032 16916 59072
rect 16780 58568 16820 58577
rect 16780 58241 16820 58528
rect 16779 58232 16821 58241
rect 16779 58192 16780 58232
rect 16820 58192 16821 58232
rect 16779 58183 16821 58192
rect 16876 57569 16916 59032
rect 16875 57560 16917 57569
rect 16875 57520 16876 57560
rect 16916 57520 16917 57560
rect 16875 57511 16917 57520
rect 16588 56680 16724 56720
rect 16780 57056 16820 57065
rect 16299 56344 16300 56384
rect 16340 56344 16436 56384
rect 16491 56384 16533 56393
rect 16491 56344 16492 56384
rect 16532 56344 16533 56384
rect 16299 56335 16341 56344
rect 16491 56335 16533 56344
rect 16300 55637 16340 56335
rect 16299 55628 16341 55637
rect 16299 55588 16300 55628
rect 16340 55588 16341 55628
rect 16492 55628 16532 56335
rect 16588 55973 16628 56680
rect 16684 56552 16724 56561
rect 16780 56552 16820 57016
rect 16875 57056 16917 57065
rect 16875 57016 16876 57056
rect 16916 57016 16917 57056
rect 16875 57007 16917 57016
rect 16876 56922 16916 57007
rect 16724 56512 16820 56552
rect 16875 56552 16917 56561
rect 16875 56512 16876 56552
rect 16916 56512 16917 56552
rect 16684 56503 16724 56512
rect 16875 56503 16917 56512
rect 16876 56418 16916 56503
rect 16972 56132 17012 59116
rect 17068 57896 17108 60040
rect 17164 59492 17204 60208
rect 17164 59443 17204 59452
rect 17260 59912 17300 59921
rect 17260 59417 17300 59872
rect 17259 59408 17301 59417
rect 17259 59368 17260 59408
rect 17300 59368 17301 59408
rect 17259 59359 17301 59368
rect 17355 59156 17397 59165
rect 17355 59116 17356 59156
rect 17396 59116 17397 59156
rect 17355 59107 17397 59116
rect 17164 57896 17204 57905
rect 17068 57856 17164 57896
rect 17068 56729 17108 57856
rect 17164 57847 17204 57856
rect 17356 57812 17396 59107
rect 17452 57896 17492 61375
rect 17643 60920 17685 60929
rect 17643 60880 17644 60920
rect 17684 60880 17685 60920
rect 17643 60871 17685 60880
rect 17644 60786 17684 60871
rect 17547 60584 17589 60593
rect 17547 60544 17548 60584
rect 17588 60544 17589 60584
rect 17547 60535 17589 60544
rect 17548 60080 17588 60535
rect 17643 60500 17685 60509
rect 17643 60460 17644 60500
rect 17684 60460 17685 60500
rect 17643 60451 17685 60460
rect 17548 60031 17588 60040
rect 17644 60080 17684 60451
rect 17740 60425 17780 62392
rect 17836 60677 17876 60762
rect 17835 60668 17877 60677
rect 17835 60628 17836 60668
rect 17876 60628 17877 60668
rect 17835 60619 17877 60628
rect 17932 60500 17972 62392
rect 17836 60460 17972 60500
rect 17739 60416 17781 60425
rect 17739 60376 17740 60416
rect 17780 60376 17781 60416
rect 17739 60367 17781 60376
rect 17548 59417 17588 59502
rect 17547 59408 17589 59417
rect 17547 59368 17548 59408
rect 17588 59368 17589 59408
rect 17547 59359 17589 59368
rect 17644 59408 17684 60040
rect 17644 59249 17684 59368
rect 17739 59324 17781 59333
rect 17739 59284 17740 59324
rect 17780 59284 17781 59324
rect 17739 59275 17781 59284
rect 17643 59240 17685 59249
rect 17643 59200 17644 59240
rect 17684 59200 17685 59240
rect 17643 59191 17685 59200
rect 17548 57896 17588 57905
rect 17452 57856 17548 57896
rect 17548 57847 17588 57856
rect 17643 57896 17685 57905
rect 17643 57856 17644 57896
rect 17684 57856 17685 57896
rect 17643 57847 17685 57856
rect 17356 57772 17492 57812
rect 17452 57728 17492 57772
rect 17644 57762 17684 57847
rect 17452 57688 17588 57728
rect 17163 57644 17205 57653
rect 17163 57604 17164 57644
rect 17204 57604 17205 57644
rect 17163 57595 17205 57604
rect 17356 57644 17396 57653
rect 17396 57604 17492 57644
rect 17356 57595 17396 57604
rect 17164 56804 17204 57595
rect 17260 57056 17300 57067
rect 17260 56981 17300 57016
rect 17356 57056 17396 57065
rect 17259 56972 17301 56981
rect 17259 56932 17260 56972
rect 17300 56932 17301 56972
rect 17259 56923 17301 56932
rect 17164 56764 17300 56804
rect 17067 56720 17109 56729
rect 17067 56680 17068 56720
rect 17108 56680 17109 56720
rect 17067 56671 17109 56680
rect 17068 56300 17108 56309
rect 17108 56260 17204 56300
rect 17068 56251 17108 56260
rect 16972 56092 17108 56132
rect 16587 55964 16629 55973
rect 16587 55924 16588 55964
rect 16628 55924 16629 55964
rect 16587 55915 16629 55924
rect 16971 55964 17013 55973
rect 16971 55924 16972 55964
rect 17012 55924 17013 55964
rect 16971 55915 17013 55924
rect 16875 55628 16917 55637
rect 16492 55588 16628 55628
rect 16299 55579 16341 55588
rect 16300 55544 16340 55579
rect 16300 55494 16340 55504
rect 16108 55420 16244 55460
rect 16011 55411 16053 55420
rect 16108 54872 16148 54883
rect 16108 54797 16148 54832
rect 16107 54788 16149 54797
rect 16107 54748 16108 54788
rect 16148 54748 16149 54788
rect 16107 54739 16149 54748
rect 16204 53360 16244 55420
rect 16492 55376 16532 55385
rect 16395 55208 16437 55217
rect 16395 55168 16396 55208
rect 16436 55168 16437 55208
rect 16395 55159 16437 55168
rect 16299 55040 16341 55049
rect 16299 55000 16300 55040
rect 16340 55000 16341 55040
rect 16299 54991 16341 55000
rect 16300 53369 16340 54991
rect 16204 52613 16244 53320
rect 16299 53360 16341 53369
rect 16299 53320 16300 53360
rect 16340 53320 16341 53360
rect 16299 53311 16341 53320
rect 16203 52604 16245 52613
rect 16203 52564 16204 52604
rect 16244 52564 16245 52604
rect 16203 52555 16245 52564
rect 15916 52480 16148 52520
rect 15723 52352 15765 52361
rect 15723 52312 15724 52352
rect 15764 52312 15765 52352
rect 15723 52303 15765 52312
rect 15724 51848 15764 52303
rect 15820 52016 15860 52480
rect 16011 52352 16053 52361
rect 16011 52312 16012 52352
rect 16052 52312 16053 52352
rect 16011 52303 16053 52312
rect 16012 52218 16052 52303
rect 16011 52016 16053 52025
rect 15820 51976 15956 52016
rect 15724 51799 15764 51808
rect 15819 51848 15861 51857
rect 15819 51808 15820 51848
rect 15860 51808 15861 51848
rect 15819 51799 15861 51808
rect 15627 51764 15669 51773
rect 15627 51724 15628 51764
rect 15668 51724 15669 51764
rect 15627 51715 15669 51724
rect 15340 49540 15476 49580
rect 15531 49580 15573 49589
rect 15531 49540 15532 49580
rect 15572 49540 15573 49580
rect 15340 49496 15380 49540
rect 15531 49531 15573 49540
rect 15340 49447 15380 49456
rect 15436 49476 15476 49485
rect 15436 49421 15476 49436
rect 15435 49412 15477 49421
rect 15435 49372 15436 49412
rect 15476 49372 15477 49412
rect 15435 49363 15477 49372
rect 15436 49341 15476 49363
rect 15628 49328 15668 51715
rect 15820 51714 15860 51799
rect 15819 51092 15861 51101
rect 15819 51052 15820 51092
rect 15860 51052 15861 51092
rect 15819 51043 15861 51052
rect 15820 50252 15860 51043
rect 15916 51017 15956 51976
rect 16011 51976 16012 52016
rect 16052 51976 16053 52016
rect 16011 51967 16053 51976
rect 15915 51008 15957 51017
rect 15915 50968 15916 51008
rect 15956 50968 15957 51008
rect 15915 50959 15957 50968
rect 16012 50756 16052 51967
rect 16108 51596 16148 52480
rect 16204 52025 16244 52555
rect 16203 52016 16245 52025
rect 16203 51976 16204 52016
rect 16244 51976 16245 52016
rect 16203 51967 16245 51976
rect 16204 51773 16244 51858
rect 16300 51848 16340 53311
rect 16300 51799 16340 51808
rect 16203 51764 16245 51773
rect 16203 51724 16204 51764
rect 16244 51724 16245 51764
rect 16203 51715 16245 51724
rect 16108 51556 16340 51596
rect 16203 51092 16245 51101
rect 16203 51052 16204 51092
rect 16244 51052 16245 51092
rect 16203 51043 16245 51052
rect 16204 51008 16244 51043
rect 16012 50716 16148 50756
rect 16011 50252 16053 50261
rect 15820 50212 15956 50252
rect 15819 50084 15861 50093
rect 15819 50044 15820 50084
rect 15860 50044 15861 50084
rect 15819 50035 15861 50044
rect 15820 49950 15860 50035
rect 15916 49748 15956 50212
rect 16011 50212 16012 50252
rect 16052 50212 16053 50252
rect 16011 50203 16053 50212
rect 16012 50118 16052 50203
rect 15916 49708 16052 49748
rect 15915 49580 15957 49589
rect 15915 49540 15916 49580
rect 15956 49540 15957 49580
rect 15915 49531 15957 49540
rect 15723 49496 15765 49505
rect 15723 49456 15724 49496
rect 15764 49456 15765 49496
rect 15723 49447 15765 49456
rect 15820 49496 15860 49505
rect 15244 49288 15380 49328
rect 14859 46304 14901 46313
rect 14859 46264 14860 46304
rect 14900 46264 14901 46304
rect 14859 46255 14901 46264
rect 15148 45968 15188 47272
rect 15243 46808 15285 46817
rect 15243 46768 15244 46808
rect 15284 46768 15285 46808
rect 15243 46759 15285 46768
rect 15244 46472 15284 46759
rect 15244 46423 15284 46432
rect 15148 45928 15284 45968
rect 14860 45884 14900 45893
rect 14900 45844 15188 45884
rect 14860 45835 14900 45844
rect 15148 45800 15188 45844
rect 15244 45809 15284 45928
rect 15148 45751 15188 45760
rect 15243 45800 15285 45809
rect 15243 45760 15244 45800
rect 15284 45760 15285 45800
rect 15243 45751 15285 45760
rect 15244 45666 15284 45751
rect 15243 44960 15285 44969
rect 15148 44920 15244 44960
rect 15284 44920 15285 44960
rect 15051 43868 15093 43877
rect 15051 43828 15052 43868
rect 15092 43828 15093 43868
rect 15051 43819 15093 43828
rect 15052 43700 15092 43819
rect 15052 43651 15092 43660
rect 14860 43532 14900 43541
rect 14860 42365 14900 43492
rect 14859 42356 14901 42365
rect 14859 42316 14860 42356
rect 14900 42316 14901 42356
rect 14859 42307 14901 42316
rect 15148 39509 15188 44920
rect 15243 44911 15285 44920
rect 15244 44826 15284 44911
rect 15243 44288 15285 44297
rect 15243 44248 15244 44288
rect 15284 44248 15285 44288
rect 15243 44239 15285 44248
rect 15244 44154 15284 44239
rect 15147 39500 15189 39509
rect 15147 39460 15148 39500
rect 15188 39460 15189 39500
rect 15147 39451 15189 39460
rect 14859 39248 14901 39257
rect 14859 39208 14860 39248
rect 14900 39208 14901 39248
rect 14859 39199 14901 39208
rect 14475 37780 14476 37820
rect 14516 37780 14517 37820
rect 14475 37771 14517 37780
rect 14668 37780 14804 37820
rect 14379 37568 14421 37577
rect 14379 37528 14380 37568
rect 14420 37528 14421 37568
rect 14379 37519 14421 37528
rect 13996 36856 14612 36896
rect 13804 36847 13844 36856
rect 13612 36679 13652 36688
rect 13900 36728 13940 36739
rect 13900 36653 13940 36688
rect 13995 36728 14037 36737
rect 13995 36688 13996 36728
rect 14036 36688 14037 36728
rect 13995 36679 14037 36688
rect 14092 36728 14132 36737
rect 13516 36595 13556 36604
rect 13899 36644 13941 36653
rect 13899 36604 13900 36644
rect 13940 36604 13941 36644
rect 13899 36595 13941 36604
rect 13996 36594 14036 36679
rect 13420 36560 13460 36569
rect 14092 36560 14132 36688
rect 14284 36728 14324 36737
rect 14324 36688 14516 36728
rect 14284 36679 14324 36688
rect 14380 36560 14420 36569
rect 14092 36520 14380 36560
rect 13323 36308 13365 36317
rect 13323 36268 13324 36308
rect 13364 36268 13365 36308
rect 13323 36259 13365 36268
rect 13227 36056 13269 36065
rect 13227 36016 13228 36056
rect 13268 36016 13269 36056
rect 13227 36007 13269 36016
rect 13324 36056 13364 36259
rect 13324 36007 13364 36016
rect 13420 35897 13460 36520
rect 14380 36511 14420 36520
rect 13707 36308 13749 36317
rect 13707 36268 13708 36308
rect 13748 36268 13749 36308
rect 13707 36259 13749 36268
rect 13228 35888 13268 35897
rect 13228 35729 13268 35848
rect 13324 35888 13364 35897
rect 13076 35680 13172 35720
rect 13227 35720 13269 35729
rect 13227 35680 13228 35720
rect 13268 35680 13269 35720
rect 13036 35671 13076 35680
rect 13227 35671 13269 35680
rect 13227 35468 13269 35477
rect 13227 35428 13228 35468
rect 13268 35428 13269 35468
rect 13227 35419 13269 35428
rect 12844 35344 12980 35384
rect 13228 35384 13268 35419
rect 13324 35393 13364 35848
rect 13419 35888 13461 35897
rect 13419 35848 13420 35888
rect 13460 35848 13461 35888
rect 13419 35839 13461 35848
rect 13516 35888 13556 35897
rect 13708 35888 13748 36259
rect 13996 36100 14420 36140
rect 13556 35848 13652 35888
rect 13516 35839 13556 35848
rect 12596 35260 12692 35300
rect 12747 35300 12789 35309
rect 12747 35260 12748 35300
rect 12788 35260 12789 35300
rect 12556 35251 12596 35260
rect 12747 35251 12789 35260
rect 12460 35167 12500 35176
rect 12076 35048 12116 35167
rect 12171 35132 12213 35141
rect 12171 35092 12172 35132
rect 12212 35092 12213 35132
rect 12171 35083 12213 35092
rect 12555 35132 12597 35141
rect 12555 35092 12556 35132
rect 12596 35092 12597 35132
rect 12555 35083 12597 35092
rect 12076 34999 12116 35008
rect 11979 34544 12021 34553
rect 11979 34504 11980 34544
rect 12020 34504 12021 34544
rect 11979 34495 12021 34504
rect 11691 34124 11733 34133
rect 11691 34084 11692 34124
rect 11732 34084 11733 34124
rect 11691 34075 11733 34084
rect 11883 34124 11925 34133
rect 11883 34084 11884 34124
rect 11924 34084 11925 34124
rect 11883 34075 11925 34084
rect 11691 33956 11733 33965
rect 11691 33916 11692 33956
rect 11732 33916 11733 33956
rect 11691 33907 11733 33916
rect 11692 33872 11732 33907
rect 11692 33821 11732 33832
rect 11787 33872 11829 33881
rect 11787 33832 11788 33872
rect 11828 33832 11829 33872
rect 11787 33823 11829 33832
rect 11596 33704 11636 33713
rect 11500 33664 11596 33704
rect 11403 33655 11445 33664
rect 11596 33655 11636 33664
rect 11788 33704 11828 33823
rect 11308 33496 11444 33536
rect 11020 33076 11156 33116
rect 10580 32152 10676 32192
rect 10732 32360 10772 32369
rect 10540 31025 10580 32152
rect 10635 31436 10677 31445
rect 10635 31396 10636 31436
rect 10676 31396 10677 31436
rect 10635 31387 10677 31396
rect 10636 31352 10676 31387
rect 10636 31277 10676 31312
rect 10635 31268 10677 31277
rect 10635 31228 10636 31268
rect 10676 31228 10677 31268
rect 10635 31219 10677 31228
rect 10636 31188 10676 31219
rect 10732 31100 10772 32320
rect 10828 32320 11060 32360
rect 10828 31604 10868 32320
rect 10828 31555 10868 31564
rect 10924 32192 10964 32201
rect 10636 31060 10772 31100
rect 10828 31184 10868 31193
rect 10539 31016 10581 31025
rect 10539 30976 10540 31016
rect 10580 30976 10581 31016
rect 10539 30967 10581 30976
rect 10443 30764 10485 30773
rect 10443 30724 10444 30764
rect 10484 30724 10485 30764
rect 10443 30715 10485 30724
rect 10540 30764 10580 30773
rect 10348 30666 10388 30691
rect 10348 30605 10388 30626
rect 10347 30596 10389 30605
rect 10347 30556 10348 30596
rect 10388 30556 10389 30596
rect 10347 30547 10389 30556
rect 10443 30008 10485 30017
rect 10443 29968 10444 30008
rect 10484 29968 10485 30008
rect 10443 29959 10485 29968
rect 10444 29840 10484 29959
rect 10540 29849 10580 30724
rect 10444 29791 10484 29800
rect 10539 29840 10581 29849
rect 10539 29800 10540 29840
rect 10580 29800 10581 29840
rect 10539 29791 10581 29800
rect 10636 29840 10676 31060
rect 10828 31016 10868 31144
rect 10732 30976 10868 31016
rect 10732 30605 10772 30976
rect 10827 30680 10869 30689
rect 10827 30640 10828 30680
rect 10868 30640 10869 30680
rect 10827 30631 10869 30640
rect 10731 30596 10773 30605
rect 10731 30556 10732 30596
rect 10772 30556 10773 30596
rect 10731 30547 10773 30556
rect 10732 30428 10772 30547
rect 10828 30546 10868 30631
rect 10924 30521 10964 32152
rect 11020 32192 11060 32320
rect 11020 32143 11060 32152
rect 11019 32024 11061 32033
rect 11019 31984 11020 32024
rect 11060 31984 11061 32024
rect 11019 31975 11061 31984
rect 11020 31184 11060 31975
rect 11020 31135 11060 31144
rect 11116 31016 11156 33076
rect 11211 32360 11253 32369
rect 11211 32320 11212 32360
rect 11252 32320 11253 32360
rect 11211 32311 11253 32320
rect 11212 32226 11252 32311
rect 11404 32192 11444 33496
rect 11691 33368 11733 33377
rect 11691 33328 11692 33368
rect 11732 33328 11733 33368
rect 11691 33319 11733 33328
rect 11212 31940 11252 31949
rect 11212 31520 11252 31900
rect 11404 31529 11444 32152
rect 11499 31604 11541 31613
rect 11499 31564 11500 31604
rect 11540 31564 11541 31604
rect 11499 31555 11541 31564
rect 11403 31520 11445 31529
rect 11212 31480 11348 31520
rect 11211 31352 11253 31361
rect 11211 31312 11212 31352
rect 11252 31312 11253 31352
rect 11211 31303 11253 31312
rect 11308 31352 11348 31480
rect 11403 31480 11404 31520
rect 11444 31480 11445 31520
rect 11403 31471 11445 31480
rect 11308 31303 11348 31312
rect 11500 31352 11540 31555
rect 11500 31303 11540 31312
rect 11212 31218 11252 31303
rect 11307 31184 11349 31193
rect 11307 31144 11308 31184
rect 11348 31144 11349 31184
rect 11307 31135 11349 31144
rect 11020 30976 11156 31016
rect 10923 30512 10965 30521
rect 10923 30472 10924 30512
rect 10964 30472 10965 30512
rect 10923 30463 10965 30472
rect 10732 30388 10868 30428
rect 10636 29791 10676 29800
rect 10732 29840 10772 29849
rect 10539 29672 10581 29681
rect 10539 29632 10540 29672
rect 10580 29632 10581 29672
rect 10539 29623 10581 29632
rect 10540 29538 10580 29623
rect 10251 29420 10293 29429
rect 10251 29380 10252 29420
rect 10292 29380 10293 29420
rect 10251 29371 10293 29380
rect 10539 29420 10581 29429
rect 10539 29380 10540 29420
rect 10580 29380 10581 29420
rect 10539 29371 10581 29380
rect 10155 29168 10197 29177
rect 10155 29128 10156 29168
rect 10196 29128 10197 29168
rect 10155 29119 10197 29128
rect 10252 29168 10292 29177
rect 10252 29000 10292 29128
rect 10156 28960 10292 29000
rect 10156 28169 10196 28960
rect 10444 28916 10484 28925
rect 10252 28876 10444 28916
rect 10155 28160 10197 28169
rect 10155 28120 10156 28160
rect 10196 28120 10197 28160
rect 10155 28111 10197 28120
rect 9964 27700 10100 27740
rect 9964 27656 10004 27700
rect 10252 27656 10292 28876
rect 10444 28867 10484 28876
rect 10347 28580 10389 28589
rect 10347 28540 10348 28580
rect 10388 28540 10389 28580
rect 10347 28531 10389 28540
rect 10348 27740 10388 28531
rect 10540 27824 10580 29371
rect 10635 29336 10677 29345
rect 10635 29296 10636 29336
rect 10676 29296 10677 29336
rect 10635 29287 10677 29296
rect 10732 29336 10772 29800
rect 10732 29287 10772 29296
rect 10636 29168 10676 29287
rect 10636 29119 10676 29128
rect 10828 29168 10868 30388
rect 10923 30176 10965 30185
rect 10923 30136 10924 30176
rect 10964 30136 10965 30176
rect 10923 30127 10965 30136
rect 10924 29849 10964 30127
rect 10923 29840 10965 29849
rect 10923 29800 10924 29840
rect 10964 29800 10965 29840
rect 10923 29791 10965 29800
rect 10924 29705 10964 29791
rect 11020 29261 11060 30976
rect 11211 30932 11253 30941
rect 11116 30892 11212 30932
rect 11252 30892 11253 30932
rect 11116 30680 11156 30892
rect 11211 30883 11253 30892
rect 11211 30764 11253 30773
rect 11211 30724 11212 30764
rect 11252 30724 11253 30764
rect 11211 30715 11253 30724
rect 11116 30176 11156 30640
rect 11212 30630 11252 30715
rect 11308 30605 11348 31135
rect 11307 30596 11349 30605
rect 11307 30556 11308 30596
rect 11348 30556 11349 30596
rect 11307 30547 11349 30556
rect 11499 30512 11541 30521
rect 11499 30472 11500 30512
rect 11540 30472 11541 30512
rect 11499 30463 11541 30472
rect 11500 30378 11540 30463
rect 11116 30136 11348 30176
rect 11115 30008 11157 30017
rect 11115 29968 11116 30008
rect 11156 29968 11157 30008
rect 11115 29959 11157 29968
rect 11116 29513 11156 29959
rect 11115 29504 11157 29513
rect 11115 29464 11116 29504
rect 11156 29464 11157 29504
rect 11115 29455 11157 29464
rect 11019 29252 11061 29261
rect 11019 29212 11020 29252
rect 11060 29212 11061 29252
rect 11019 29203 11061 29212
rect 10828 29119 10868 29128
rect 10923 29168 10965 29177
rect 10923 29128 10924 29168
rect 10964 29128 10965 29168
rect 10923 29119 10965 29128
rect 11116 29168 11156 29177
rect 10924 29034 10964 29119
rect 10827 29000 10869 29009
rect 11116 29000 11156 29128
rect 10732 28960 10828 29000
rect 10868 28960 10869 29000
rect 10635 28916 10677 28925
rect 10635 28876 10636 28916
rect 10676 28876 10677 28916
rect 10635 28867 10677 28876
rect 10348 27691 10388 27700
rect 10444 27784 10580 27824
rect 9868 27616 10004 27656
rect 10060 27646 10292 27656
rect 10060 27616 10204 27646
rect 9771 26900 9813 26909
rect 9771 26860 9772 26900
rect 9812 26860 9813 26900
rect 9771 26851 9813 26860
rect 9868 25976 9908 27616
rect 9963 27152 10005 27161
rect 9963 27112 9964 27152
rect 10004 27112 10005 27152
rect 9963 27103 10005 27112
rect 9964 26321 10004 27103
rect 10060 26909 10100 27616
rect 10244 27616 10292 27646
rect 10204 27597 10244 27606
rect 10155 27488 10197 27497
rect 10155 27448 10156 27488
rect 10196 27448 10197 27488
rect 10155 27439 10197 27448
rect 10059 26900 10101 26909
rect 10059 26860 10060 26900
rect 10100 26860 10101 26900
rect 10059 26851 10101 26860
rect 10060 26816 10100 26851
rect 10060 26766 10100 26776
rect 10156 26816 10196 27439
rect 10251 27236 10293 27245
rect 10251 27196 10252 27236
rect 10292 27196 10293 27236
rect 10251 27187 10293 27196
rect 9963 26312 10005 26321
rect 9963 26272 9964 26312
rect 10004 26272 10005 26312
rect 9963 26263 10005 26272
rect 9964 26060 10004 26069
rect 9964 25976 10004 26020
rect 10059 26060 10101 26069
rect 10059 26020 10060 26060
rect 10100 26020 10101 26060
rect 10059 26011 10101 26020
rect 9868 25936 10004 25976
rect 9771 25304 9813 25313
rect 9771 25264 9772 25304
rect 9812 25264 9813 25304
rect 9771 25255 9813 25264
rect 9772 25170 9812 25255
rect 9868 24809 9908 25936
rect 10060 25926 10100 26011
rect 9963 25808 10005 25817
rect 9963 25768 9964 25808
rect 10004 25768 10005 25808
rect 9963 25759 10005 25768
rect 9867 24800 9909 24809
rect 9867 24760 9868 24800
rect 9908 24760 9909 24800
rect 9867 24751 9909 24760
rect 9867 24632 9909 24641
rect 9867 24592 9868 24632
rect 9908 24592 9909 24632
rect 9867 24583 9909 24592
rect 9772 24548 9812 24557
rect 9772 22457 9812 24508
rect 9868 24498 9908 24583
rect 9867 22952 9909 22961
rect 9867 22912 9868 22952
rect 9908 22912 9909 22952
rect 9867 22903 9909 22912
rect 9771 22448 9813 22457
rect 9771 22408 9772 22448
rect 9812 22408 9813 22448
rect 9771 22399 9813 22408
rect 9772 21608 9812 22399
rect 9772 21559 9812 21568
rect 9868 21608 9908 22903
rect 9868 21559 9908 21568
rect 9867 21356 9909 21365
rect 9867 21316 9868 21356
rect 9908 21316 9909 21356
rect 9867 21307 9909 21316
rect 9868 20357 9908 21307
rect 9964 20609 10004 25759
rect 10059 23120 10101 23129
rect 10059 23080 10060 23120
rect 10100 23080 10101 23120
rect 10059 23071 10101 23080
rect 10060 22986 10100 23071
rect 10156 22868 10196 26776
rect 10252 26816 10292 27187
rect 10252 26767 10292 26776
rect 10347 26732 10389 26741
rect 10347 26692 10348 26732
rect 10388 26692 10389 26732
rect 10347 26683 10389 26692
rect 10348 26598 10388 26683
rect 10251 26564 10293 26573
rect 10251 26524 10252 26564
rect 10292 26524 10293 26564
rect 10251 26515 10293 26524
rect 10252 25817 10292 26515
rect 10444 26144 10484 27784
rect 10539 27656 10581 27665
rect 10539 27616 10540 27656
rect 10580 27616 10581 27656
rect 10539 27607 10581 27616
rect 10540 26816 10580 27607
rect 10636 26984 10676 28867
rect 10732 27497 10772 28960
rect 10827 28951 10869 28960
rect 11020 28960 11156 29000
rect 11212 29168 11252 29177
rect 11020 27992 11060 28960
rect 11212 28589 11252 29128
rect 11308 29093 11348 30136
rect 11595 30008 11637 30017
rect 11595 29968 11596 30008
rect 11636 29968 11637 30008
rect 11595 29959 11637 29968
rect 11596 29513 11636 29959
rect 11595 29504 11637 29513
rect 11595 29464 11596 29504
rect 11636 29464 11637 29504
rect 11595 29455 11637 29464
rect 11404 29336 11444 29345
rect 11307 29084 11349 29093
rect 11307 29044 11308 29084
rect 11348 29044 11349 29084
rect 11307 29035 11349 29044
rect 11404 29000 11444 29296
rect 11692 29177 11732 33319
rect 11691 29168 11733 29177
rect 11691 29128 11692 29168
rect 11732 29128 11733 29168
rect 11691 29119 11733 29128
rect 11404 28960 11732 29000
rect 11499 28664 11541 28673
rect 11404 28624 11500 28664
rect 11540 28624 11541 28664
rect 11211 28580 11253 28589
rect 11211 28540 11212 28580
rect 11252 28540 11253 28580
rect 11211 28531 11253 28540
rect 11116 28328 11156 28337
rect 11116 28169 11156 28288
rect 11115 28160 11157 28169
rect 11115 28120 11116 28160
rect 11156 28120 11157 28160
rect 11115 28111 11157 28120
rect 11308 28160 11348 28169
rect 11308 27992 11348 28120
rect 10828 27952 11348 27992
rect 10731 27488 10773 27497
rect 10731 27448 10732 27488
rect 10772 27448 10773 27488
rect 10731 27439 10773 27448
rect 10636 26944 10772 26984
rect 10540 26767 10580 26776
rect 10635 26816 10677 26825
rect 10635 26776 10636 26816
rect 10676 26776 10677 26816
rect 10635 26767 10677 26776
rect 10636 26682 10676 26767
rect 10540 26144 10580 26153
rect 10444 26104 10540 26144
rect 10251 25808 10293 25817
rect 10251 25768 10252 25808
rect 10292 25768 10293 25808
rect 10251 25759 10293 25768
rect 10251 25304 10293 25313
rect 10251 25264 10252 25304
rect 10292 25264 10293 25304
rect 10251 25255 10293 25264
rect 10060 22828 10196 22868
rect 9963 20600 10005 20609
rect 9963 20560 9964 20600
rect 10004 20560 10005 20600
rect 9963 20551 10005 20560
rect 9867 20348 9909 20357
rect 9867 20308 9868 20348
rect 9908 20308 9909 20348
rect 9867 20299 9909 20308
rect 9676 20140 9812 20180
rect 9676 19256 9716 19265
rect 9772 19256 9812 20140
rect 9716 19216 9812 19256
rect 9579 18584 9621 18593
rect 9579 18544 9580 18584
rect 9620 18544 9621 18584
rect 9579 18535 9621 18544
rect 9483 18248 9525 18257
rect 9483 18208 9484 18248
rect 9524 18208 9525 18248
rect 9483 18199 9525 18208
rect 9676 18089 9716 19216
rect 9675 18080 9717 18089
rect 9675 18040 9676 18080
rect 9716 18040 9717 18080
rect 9675 18031 9717 18040
rect 9291 17660 9333 17669
rect 9291 17620 9292 17660
rect 9332 17620 9333 17660
rect 9291 17611 9333 17620
rect 9675 17660 9717 17669
rect 9675 17620 9676 17660
rect 9716 17620 9717 17660
rect 9675 17611 9717 17620
rect 9387 17156 9429 17165
rect 9387 17116 9388 17156
rect 9428 17116 9429 17156
rect 9387 17107 9429 17116
rect 9388 17072 9428 17107
rect 9388 17021 9428 17032
rect 9483 17072 9525 17081
rect 9483 17032 9484 17072
rect 9524 17032 9525 17072
rect 9483 17023 9525 17032
rect 9484 16577 9524 17023
rect 9483 16568 9525 16577
rect 9483 16528 9484 16568
rect 9524 16528 9525 16568
rect 9483 16519 9525 16528
rect 9676 16493 9716 17611
rect 9868 17072 9908 20299
rect 10060 19172 10100 22828
rect 10252 22784 10292 25255
rect 10156 22744 10292 22784
rect 10348 24632 10388 24641
rect 10156 19853 10196 22744
rect 10348 21608 10388 24592
rect 10540 24389 10580 26104
rect 10539 24380 10581 24389
rect 10539 24340 10540 24380
rect 10580 24340 10581 24380
rect 10539 24331 10581 24340
rect 10732 23960 10772 26944
rect 10828 26825 10868 27952
rect 11019 27740 11061 27749
rect 11019 27700 11020 27740
rect 11060 27700 11061 27740
rect 11019 27691 11061 27700
rect 10924 27656 10964 27667
rect 10924 27581 10964 27616
rect 10923 27572 10965 27581
rect 10923 27532 10924 27572
rect 10964 27532 10965 27572
rect 10923 27523 10965 27532
rect 10924 27329 10964 27523
rect 10923 27320 10965 27329
rect 10923 27280 10924 27320
rect 10964 27280 10965 27320
rect 10923 27271 10965 27280
rect 11020 26984 11060 27691
rect 11307 27236 11349 27245
rect 11307 27196 11308 27236
rect 11348 27196 11349 27236
rect 11307 27187 11349 27196
rect 10924 26944 11060 26984
rect 10827 26816 10869 26825
rect 10827 26776 10828 26816
rect 10868 26776 10869 26816
rect 10827 26767 10869 26776
rect 10827 26648 10869 26657
rect 10827 26608 10828 26648
rect 10868 26608 10869 26648
rect 10827 26599 10869 26608
rect 10828 26514 10868 26599
rect 10924 25313 10964 26944
rect 11115 26900 11157 26909
rect 11115 26860 11116 26900
rect 11156 26860 11157 26900
rect 11115 26851 11157 26860
rect 11020 26816 11060 26825
rect 11020 26573 11060 26776
rect 11116 26816 11156 26851
rect 11116 26765 11156 26776
rect 11308 26648 11348 27187
rect 11404 26732 11444 28624
rect 11499 28615 11541 28624
rect 11500 28328 11540 28337
rect 11500 26993 11540 28288
rect 11596 28328 11636 28337
rect 11499 26984 11541 26993
rect 11499 26944 11500 26984
rect 11540 26944 11541 26984
rect 11499 26935 11541 26944
rect 11596 26825 11636 28288
rect 11692 28328 11732 28960
rect 11788 28328 11828 33664
rect 11883 33704 11925 33713
rect 11883 33664 11884 33704
rect 11924 33664 11925 33704
rect 11883 33655 11925 33664
rect 11884 33570 11924 33655
rect 11883 31604 11925 31613
rect 11883 31564 11884 31604
rect 11924 31564 11925 31604
rect 11883 31555 11925 31564
rect 11884 29840 11924 31555
rect 11980 30773 12020 34495
rect 12076 34469 12116 34505
rect 12075 34460 12117 34469
rect 12075 34420 12076 34460
rect 12116 34420 12117 34460
rect 12075 34411 12117 34420
rect 12076 34381 12116 34411
rect 12076 33713 12116 34341
rect 12075 33704 12117 33713
rect 12075 33664 12076 33704
rect 12116 33664 12117 33704
rect 12075 33655 12117 33664
rect 12076 32873 12116 33655
rect 12172 33461 12212 35083
rect 12556 34469 12596 35083
rect 12651 35048 12693 35057
rect 12651 35008 12652 35048
rect 12692 35008 12693 35048
rect 12651 34999 12693 35008
rect 12555 34460 12597 34469
rect 12555 34420 12556 34460
rect 12596 34420 12597 34460
rect 12555 34411 12597 34420
rect 12459 34376 12501 34385
rect 12459 34336 12460 34376
rect 12500 34336 12501 34376
rect 12459 34327 12501 34336
rect 12556 34376 12596 34411
rect 12268 34208 12308 34217
rect 12308 34168 12404 34208
rect 12268 34159 12308 34168
rect 12267 34040 12309 34049
rect 12267 34000 12268 34040
rect 12308 34000 12309 34040
rect 12267 33991 12309 34000
rect 12171 33452 12213 33461
rect 12171 33412 12172 33452
rect 12212 33412 12213 33452
rect 12171 33403 12213 33412
rect 12171 33284 12213 33293
rect 12171 33244 12172 33284
rect 12212 33244 12213 33284
rect 12171 33235 12213 33244
rect 12075 32864 12117 32873
rect 12075 32824 12076 32864
rect 12116 32824 12117 32864
rect 12075 32815 12117 32824
rect 12075 32360 12117 32369
rect 12075 32320 12076 32360
rect 12116 32320 12117 32360
rect 12075 32311 12117 32320
rect 11979 30764 12021 30773
rect 11979 30724 11980 30764
rect 12020 30724 12021 30764
rect 11979 30715 12021 30724
rect 12076 30680 12116 32311
rect 12172 30941 12212 33235
rect 12268 32864 12308 33991
rect 12364 33704 12404 34168
rect 12460 33872 12500 34327
rect 12556 34325 12596 34336
rect 12460 33823 12500 33832
rect 12364 33655 12404 33664
rect 12652 33704 12692 34999
rect 12748 34049 12788 35251
rect 12844 34712 12884 35344
rect 13228 35333 13268 35344
rect 13323 35384 13365 35393
rect 13323 35344 13324 35384
rect 13364 35344 13365 35384
rect 13323 35335 13365 35344
rect 13515 35384 13557 35393
rect 13515 35344 13516 35384
rect 13556 35344 13557 35384
rect 13515 35335 13557 35344
rect 13419 35300 13461 35309
rect 13419 35260 13420 35300
rect 13460 35260 13461 35300
rect 13419 35251 13461 35260
rect 12940 35216 12980 35225
rect 12940 35057 12980 35176
rect 13035 35216 13077 35225
rect 13035 35176 13036 35216
rect 13076 35176 13077 35216
rect 13035 35167 13077 35176
rect 13132 35216 13172 35227
rect 13036 35082 13076 35167
rect 13132 35141 13172 35176
rect 13420 35216 13460 35251
rect 13420 35165 13460 35176
rect 13516 35216 13556 35335
rect 13516 35167 13556 35176
rect 13131 35132 13173 35141
rect 13131 35092 13132 35132
rect 13172 35092 13173 35132
rect 13131 35083 13173 35092
rect 12939 35048 12981 35057
rect 12939 35008 12940 35048
rect 12980 35008 12981 35048
rect 12939 34999 12981 35008
rect 13515 35048 13557 35057
rect 13515 35008 13516 35048
rect 13556 35008 13557 35048
rect 13515 34999 13557 35008
rect 13419 34964 13461 34973
rect 13419 34924 13420 34964
rect 13460 34924 13461 34964
rect 13419 34915 13461 34924
rect 13323 34880 13365 34889
rect 13323 34840 13324 34880
rect 13364 34840 13365 34880
rect 13323 34831 13365 34840
rect 12844 34672 13172 34712
rect 12939 34544 12981 34553
rect 12939 34504 12940 34544
rect 12980 34504 12981 34544
rect 12939 34495 12981 34504
rect 12844 34376 12884 34385
rect 12844 34217 12884 34336
rect 12940 34376 12980 34495
rect 13035 34460 13077 34469
rect 13035 34420 13036 34460
rect 13076 34420 13077 34460
rect 13035 34411 13077 34420
rect 12940 34327 12980 34336
rect 12843 34208 12885 34217
rect 12843 34168 12844 34208
rect 12884 34168 12885 34208
rect 12843 34159 12885 34168
rect 12939 34124 12981 34133
rect 12939 34084 12940 34124
rect 12980 34084 12981 34124
rect 12939 34075 12981 34084
rect 12747 34040 12789 34049
rect 12747 34000 12748 34040
rect 12788 34000 12789 34040
rect 12747 33991 12789 34000
rect 12940 33956 12980 34075
rect 12844 33916 12980 33956
rect 12747 33872 12789 33881
rect 12747 33832 12748 33872
rect 12788 33832 12789 33872
rect 12747 33823 12789 33832
rect 12748 33738 12788 33823
rect 12652 33655 12692 33664
rect 12844 33704 12884 33916
rect 12555 33452 12597 33461
rect 12555 33412 12556 33452
rect 12596 33412 12597 33452
rect 12555 33403 12597 33412
rect 12268 32815 12308 32824
rect 12460 32864 12500 32873
rect 12364 32780 12404 32789
rect 12267 32696 12309 32705
rect 12267 32656 12268 32696
rect 12308 32656 12309 32696
rect 12267 32647 12309 32656
rect 12171 30932 12213 30941
rect 12171 30892 12172 30932
rect 12212 30892 12213 30932
rect 12171 30883 12213 30892
rect 12076 30631 12116 30640
rect 12172 30008 12212 30883
rect 12076 29968 12212 30008
rect 11884 29800 12020 29840
rect 11883 29672 11925 29681
rect 11883 29632 11884 29672
rect 11924 29632 11925 29672
rect 11883 29623 11925 29632
rect 11884 29188 11924 29623
rect 11980 29345 12020 29800
rect 11979 29336 12021 29345
rect 11979 29296 11980 29336
rect 12020 29296 12021 29336
rect 11979 29287 12021 29296
rect 12076 29177 12116 29968
rect 12172 29840 12212 29849
rect 12172 29513 12212 29800
rect 12171 29504 12213 29513
rect 12171 29464 12172 29504
rect 12212 29464 12213 29504
rect 12171 29455 12213 29464
rect 12171 29336 12213 29345
rect 12171 29296 12172 29336
rect 12212 29296 12213 29336
rect 12171 29287 12213 29296
rect 11884 29139 11924 29148
rect 11980 29168 12020 29177
rect 11980 29084 12020 29128
rect 12075 29168 12117 29177
rect 12075 29128 12076 29168
rect 12116 29128 12117 29168
rect 12075 29119 12117 29128
rect 11884 29044 12020 29084
rect 11884 28589 11924 29044
rect 12172 29000 12212 29287
rect 12268 29168 12308 32647
rect 12364 32201 12404 32740
rect 12460 32369 12500 32824
rect 12459 32360 12501 32369
rect 12459 32320 12460 32360
rect 12500 32320 12501 32360
rect 12459 32311 12501 32320
rect 12363 32192 12405 32201
rect 12363 32152 12364 32192
rect 12404 32152 12405 32192
rect 12363 32143 12405 32152
rect 12459 30764 12501 30773
rect 12459 30724 12460 30764
rect 12500 30724 12501 30764
rect 12459 30715 12501 30724
rect 12363 30680 12405 30689
rect 12363 30640 12364 30680
rect 12404 30640 12405 30680
rect 12363 30631 12405 30640
rect 12364 30546 12404 30631
rect 12460 30630 12500 30715
rect 12459 29924 12501 29933
rect 12459 29884 12460 29924
rect 12500 29884 12501 29924
rect 12459 29875 12501 29884
rect 12363 29672 12405 29681
rect 12363 29632 12364 29672
rect 12404 29632 12405 29672
rect 12363 29623 12405 29632
rect 12364 29538 12404 29623
rect 12364 29168 12404 29177
rect 12268 29128 12364 29168
rect 12076 28960 12212 29000
rect 12267 29000 12309 29009
rect 12267 28960 12268 29000
rect 12308 28960 12309 29000
rect 11979 28916 12021 28925
rect 11979 28876 11980 28916
rect 12020 28876 12021 28916
rect 11979 28867 12021 28876
rect 11883 28580 11925 28589
rect 11883 28540 11884 28580
rect 11924 28540 11925 28580
rect 11883 28531 11925 28540
rect 11788 28288 11924 28328
rect 11692 28279 11732 28288
rect 11787 28160 11829 28169
rect 11787 28120 11788 28160
rect 11828 28120 11829 28160
rect 11787 28111 11829 28120
rect 11788 28026 11828 28111
rect 11884 27917 11924 28288
rect 11883 27908 11925 27917
rect 11883 27868 11884 27908
rect 11924 27868 11925 27908
rect 11883 27859 11925 27868
rect 11691 27488 11733 27497
rect 11691 27448 11692 27488
rect 11732 27448 11733 27488
rect 11691 27439 11733 27448
rect 11595 26816 11637 26825
rect 11595 26776 11596 26816
rect 11636 26776 11637 26816
rect 11595 26767 11637 26776
rect 11404 26692 11540 26732
rect 11308 26599 11348 26608
rect 11019 26564 11061 26573
rect 11019 26524 11020 26564
rect 11060 26524 11061 26564
rect 11019 26515 11061 26524
rect 11403 26564 11445 26573
rect 11403 26524 11404 26564
rect 11444 26524 11445 26564
rect 11500 26564 11540 26692
rect 11500 26524 11636 26564
rect 11403 26515 11445 26524
rect 11211 26312 11253 26321
rect 11211 26272 11212 26312
rect 11252 26272 11253 26312
rect 11211 26263 11253 26272
rect 11212 26178 11252 26263
rect 11068 26134 11108 26143
rect 11108 26094 11252 26134
rect 11068 26085 11108 26094
rect 11212 25556 11252 26094
rect 11212 25507 11252 25516
rect 11404 25481 11444 26515
rect 11499 26228 11541 26237
rect 11499 26188 11500 26228
rect 11540 26188 11541 26228
rect 11499 26179 11541 26188
rect 11403 25472 11445 25481
rect 11403 25432 11404 25472
rect 11444 25432 11445 25472
rect 11403 25423 11445 25432
rect 10923 25304 10965 25313
rect 10923 25264 10924 25304
rect 10964 25264 10965 25304
rect 10923 25255 10965 25264
rect 11020 25304 11060 25313
rect 11060 25264 11348 25304
rect 11020 25255 11060 25264
rect 11020 24842 11060 24851
rect 11020 24800 11060 24802
rect 11115 24800 11157 24809
rect 11020 24760 11116 24800
rect 11156 24760 11157 24800
rect 11115 24751 11157 24760
rect 11308 24632 11348 25264
rect 11404 24632 11444 24641
rect 10828 24618 10868 24627
rect 10828 24044 10868 24578
rect 11308 24592 11404 24632
rect 11115 24380 11157 24389
rect 11115 24340 11116 24380
rect 11156 24340 11157 24380
rect 11115 24331 11157 24340
rect 11212 24380 11252 24389
rect 10924 24044 10964 24053
rect 10828 24004 10924 24044
rect 10924 23995 10964 24004
rect 10636 23920 10772 23960
rect 10443 23204 10485 23213
rect 10443 23164 10444 23204
rect 10484 23164 10485 23204
rect 10443 23155 10485 23164
rect 10444 22709 10484 23155
rect 10443 22700 10485 22709
rect 10443 22660 10444 22700
rect 10484 22660 10485 22700
rect 10443 22651 10485 22660
rect 10443 21692 10485 21701
rect 10443 21652 10444 21692
rect 10484 21652 10485 21692
rect 10443 21643 10485 21652
rect 10252 21568 10348 21608
rect 10155 19844 10197 19853
rect 10155 19804 10156 19844
rect 10196 19804 10197 19844
rect 10155 19795 10197 19804
rect 10252 19685 10292 21568
rect 10348 21559 10388 21568
rect 10444 21440 10484 21643
rect 10348 21400 10484 21440
rect 10348 21197 10388 21400
rect 10347 21188 10389 21197
rect 10347 21148 10348 21188
rect 10388 21148 10389 21188
rect 10347 21139 10389 21148
rect 10348 20096 10388 21139
rect 10636 21113 10676 23920
rect 10732 23792 10772 23803
rect 10732 23717 10772 23752
rect 10731 23708 10773 23717
rect 10731 23668 10732 23708
rect 10772 23668 10773 23708
rect 10731 23659 10773 23668
rect 11020 21692 11060 21701
rect 10732 21652 11020 21692
rect 10635 21104 10677 21113
rect 10635 21064 10636 21104
rect 10676 21064 10677 21104
rect 10635 21055 10677 21064
rect 10636 20525 10676 21055
rect 10635 20516 10677 20525
rect 10635 20476 10636 20516
rect 10676 20476 10677 20516
rect 10635 20467 10677 20476
rect 10732 20348 10772 21652
rect 11020 21643 11060 21652
rect 10876 21598 10916 21607
rect 10916 21558 11060 21594
rect 10876 21554 11060 21558
rect 10876 21549 10916 21554
rect 10827 21272 10869 21281
rect 10827 21232 10828 21272
rect 10868 21232 10869 21272
rect 10827 21223 10869 21232
rect 10828 20768 10868 21223
rect 11020 21020 11060 21554
rect 11020 20971 11060 20980
rect 11116 20852 11156 24331
rect 11212 23801 11252 24340
rect 11308 24305 11348 24592
rect 11404 24583 11444 24592
rect 11500 24464 11540 26179
rect 11596 24725 11636 26524
rect 11595 24716 11637 24725
rect 11595 24676 11596 24716
rect 11636 24676 11637 24716
rect 11595 24667 11637 24676
rect 11404 24424 11540 24464
rect 11307 24296 11349 24305
rect 11307 24256 11308 24296
rect 11348 24256 11349 24296
rect 11307 24247 11349 24256
rect 11211 23792 11253 23801
rect 11211 23752 11212 23792
rect 11252 23752 11253 23792
rect 11211 23743 11253 23752
rect 11308 23717 11348 24247
rect 11307 23708 11349 23717
rect 11307 23668 11308 23708
rect 11348 23668 11349 23708
rect 11307 23659 11349 23668
rect 11308 23120 11348 23659
rect 11308 21701 11348 23080
rect 11404 21944 11444 24424
rect 11692 24221 11732 27439
rect 11787 27404 11829 27413
rect 11787 27364 11788 27404
rect 11828 27364 11829 27404
rect 11787 27355 11829 27364
rect 11788 26816 11828 27355
rect 11980 26993 12020 28867
rect 12076 28673 12116 28960
rect 12267 28951 12309 28960
rect 12075 28664 12117 28673
rect 12075 28624 12076 28664
rect 12116 28624 12117 28664
rect 12075 28615 12117 28624
rect 12076 28328 12116 28615
rect 12171 28580 12213 28589
rect 12171 28540 12172 28580
rect 12212 28540 12213 28580
rect 12171 28531 12213 28540
rect 12076 28279 12116 28288
rect 12172 28160 12212 28531
rect 12076 28120 12212 28160
rect 11979 26984 12021 26993
rect 11979 26944 11980 26984
rect 12020 26944 12021 26984
rect 11979 26935 12021 26944
rect 11788 26767 11828 26776
rect 11884 26816 11924 26825
rect 11884 26732 11924 26776
rect 12076 26732 12116 28120
rect 12171 27656 12213 27665
rect 12171 27616 12172 27656
rect 12212 27616 12213 27656
rect 12171 27607 12213 27616
rect 12172 27522 12212 27607
rect 12268 27497 12308 28951
rect 12364 27656 12404 29128
rect 12460 29168 12500 29875
rect 12460 27917 12500 29128
rect 12459 27908 12501 27917
rect 12459 27868 12460 27908
rect 12500 27868 12501 27908
rect 12459 27859 12501 27868
rect 12364 27616 12500 27656
rect 12267 27488 12309 27497
rect 12267 27448 12268 27488
rect 12308 27448 12309 27488
rect 12267 27439 12309 27448
rect 12364 27413 12404 27498
rect 12363 27404 12405 27413
rect 12363 27364 12364 27404
rect 12404 27364 12405 27404
rect 12363 27355 12405 27364
rect 12460 27236 12500 27616
rect 12268 27196 12500 27236
rect 12171 26984 12213 26993
rect 12171 26944 12172 26984
rect 12212 26944 12213 26984
rect 12171 26935 12213 26944
rect 11884 26692 12116 26732
rect 11884 24977 11924 26692
rect 11980 26144 12020 26153
rect 11980 25985 12020 26104
rect 11979 25976 12021 25985
rect 11979 25936 11980 25976
rect 12020 25936 12021 25976
rect 11979 25927 12021 25936
rect 11883 24968 11925 24977
rect 11883 24928 11884 24968
rect 11924 24928 11925 24968
rect 11883 24919 11925 24928
rect 11691 24212 11733 24221
rect 11691 24172 11692 24212
rect 11732 24172 11733 24212
rect 11691 24163 11733 24172
rect 11692 23969 11732 24054
rect 11691 23960 11733 23969
rect 11691 23920 11692 23960
rect 11732 23920 11733 23960
rect 12172 23960 12212 26935
rect 12268 26816 12308 27196
rect 12459 26984 12501 26993
rect 12459 26944 12460 26984
rect 12500 26944 12501 26984
rect 12459 26935 12501 26944
rect 12268 26489 12308 26776
rect 12364 26816 12404 26825
rect 12267 26480 12309 26489
rect 12267 26440 12268 26480
rect 12308 26440 12309 26480
rect 12267 26431 12309 26440
rect 12364 26237 12404 26776
rect 12363 26228 12405 26237
rect 12363 26188 12364 26228
rect 12404 26188 12405 26228
rect 12363 26179 12405 26188
rect 12363 24380 12405 24389
rect 12363 24340 12364 24380
rect 12404 24340 12405 24380
rect 12363 24331 12405 24340
rect 12364 24044 12404 24331
rect 12460 24137 12500 26935
rect 12459 24128 12501 24137
rect 12459 24088 12460 24128
rect 12500 24088 12501 24128
rect 12459 24079 12501 24088
rect 12364 23995 12404 24004
rect 12556 23960 12596 33403
rect 12844 32444 12884 33664
rect 12940 33704 12980 33713
rect 13036 33704 13076 34411
rect 12980 33664 13076 33704
rect 13132 33704 13172 34672
rect 13228 34553 13268 34638
rect 13227 34544 13269 34553
rect 13227 34504 13228 34544
rect 13268 34504 13269 34544
rect 13227 34495 13269 34504
rect 13324 34376 13364 34831
rect 13420 34628 13460 34915
rect 13420 34579 13460 34588
rect 12940 33655 12980 33664
rect 13132 32789 13172 33664
rect 13228 34336 13364 34376
rect 13420 34376 13460 34385
rect 13228 33620 13268 34336
rect 13420 33881 13460 34336
rect 13516 34376 13556 34999
rect 13516 34217 13556 34336
rect 13515 34208 13557 34217
rect 13515 34168 13516 34208
rect 13556 34168 13557 34208
rect 13515 34159 13557 34168
rect 13419 33872 13461 33881
rect 13419 33832 13420 33872
rect 13460 33832 13461 33872
rect 13419 33823 13461 33832
rect 13612 33713 13652 35848
rect 13708 35839 13748 35848
rect 13804 35888 13844 35897
rect 13804 35477 13844 35848
rect 13900 35888 13940 35897
rect 13803 35468 13845 35477
rect 13803 35428 13804 35468
rect 13844 35428 13845 35468
rect 13803 35419 13845 35428
rect 13708 35384 13748 35393
rect 13708 34889 13748 35344
rect 13707 34880 13749 34889
rect 13707 34840 13708 34880
rect 13748 34840 13749 34880
rect 13707 34831 13749 34840
rect 13900 34796 13940 35848
rect 13996 35888 14036 36100
rect 14188 35897 14228 35982
rect 13996 35839 14036 35848
rect 14187 35888 14229 35897
rect 14187 35848 14188 35888
rect 14228 35848 14229 35888
rect 14187 35839 14229 35848
rect 14284 35888 14324 35897
rect 14284 35384 14324 35848
rect 14380 35888 14420 36100
rect 14476 35981 14516 36688
rect 14475 35972 14517 35981
rect 14475 35932 14476 35972
rect 14516 35932 14517 35972
rect 14475 35923 14517 35932
rect 14380 35839 14420 35848
rect 14476 35720 14516 35729
rect 14188 35344 14324 35384
rect 14380 35680 14476 35720
rect 14091 35048 14133 35057
rect 14091 35008 14092 35048
rect 14132 35008 14133 35048
rect 14091 34999 14133 35008
rect 14092 34914 14132 34999
rect 14188 34973 14228 35344
rect 14283 35216 14325 35225
rect 14283 35176 14284 35216
rect 14324 35176 14325 35216
rect 14283 35167 14325 35176
rect 14284 35082 14324 35167
rect 14187 34964 14229 34973
rect 14187 34924 14188 34964
rect 14228 34924 14229 34964
rect 14187 34915 14229 34924
rect 13900 34756 14324 34796
rect 14188 34553 14228 34638
rect 13803 34544 13845 34553
rect 13803 34504 13804 34544
rect 13844 34504 13845 34544
rect 13803 34495 13845 34504
rect 14187 34544 14229 34553
rect 14187 34504 14188 34544
rect 14228 34504 14229 34544
rect 14187 34495 14229 34504
rect 13707 34376 13749 34385
rect 13707 34336 13708 34376
rect 13748 34336 13749 34376
rect 13707 34327 13749 34336
rect 13804 34376 13844 34495
rect 13804 34327 13844 34336
rect 13959 34376 13999 34385
rect 14188 34376 14228 34385
rect 13999 34336 14036 34376
rect 13959 34327 14036 34336
rect 13708 34242 13748 34327
rect 13803 34208 13845 34217
rect 13803 34168 13804 34208
rect 13844 34168 13845 34208
rect 13803 34159 13845 34168
rect 13707 34040 13749 34049
rect 13707 34000 13708 34040
rect 13748 34000 13749 34040
rect 13707 33991 13749 34000
rect 13419 33704 13461 33713
rect 13419 33664 13420 33704
rect 13460 33664 13461 33704
rect 13419 33655 13461 33664
rect 13516 33704 13556 33713
rect 13228 33571 13268 33580
rect 13420 33620 13460 33655
rect 13420 33569 13460 33580
rect 13324 33536 13364 33545
rect 13227 32864 13269 32873
rect 13227 32824 13228 32864
rect 13268 32824 13269 32864
rect 13324 32864 13364 33496
rect 13516 33461 13556 33664
rect 13611 33704 13653 33713
rect 13611 33664 13612 33704
rect 13652 33664 13653 33704
rect 13611 33655 13653 33664
rect 13708 33704 13748 33991
rect 13804 33704 13844 34159
rect 13996 34049 14036 34327
rect 14092 34336 14188 34376
rect 13899 34040 13941 34049
rect 13899 34000 13900 34040
rect 13940 34000 13941 34040
rect 13996 34040 14044 34049
rect 13996 34000 14003 34040
rect 14043 34000 14044 34040
rect 13899 33991 13941 34000
rect 14002 33991 14044 34000
rect 13900 33872 13940 33991
rect 13900 33832 14036 33872
rect 13900 33704 13940 33713
rect 13804 33664 13900 33704
rect 13708 33655 13748 33664
rect 13515 33452 13557 33461
rect 13515 33412 13516 33452
rect 13556 33412 13557 33452
rect 13515 33403 13557 33412
rect 13515 33284 13557 33293
rect 13515 33244 13516 33284
rect 13556 33244 13557 33284
rect 13515 33235 13557 33244
rect 13420 33041 13460 33126
rect 13419 33032 13461 33041
rect 13419 32992 13420 33032
rect 13460 32992 13461 33032
rect 13419 32983 13461 32992
rect 13420 32864 13460 32873
rect 13324 32824 13420 32864
rect 13227 32815 13269 32824
rect 13420 32815 13460 32824
rect 13516 32864 13556 33235
rect 13612 33116 13652 33655
rect 13809 33452 13849 33664
rect 13900 33655 13940 33664
rect 13996 33704 14036 33832
rect 13996 33655 14036 33664
rect 13996 33536 14036 33545
rect 13804 33412 13849 33452
rect 13899 33452 13941 33461
rect 13899 33412 13900 33452
rect 13940 33412 13941 33452
rect 13708 33116 13748 33125
rect 13612 33076 13708 33116
rect 13708 33067 13748 33076
rect 13516 32815 13556 32824
rect 13804 32864 13844 33412
rect 13899 33403 13941 33412
rect 13804 32815 13844 32824
rect 13131 32780 13173 32789
rect 13131 32740 13132 32780
rect 13172 32740 13173 32780
rect 13131 32731 13173 32740
rect 13228 32730 13268 32815
rect 13900 32696 13940 33403
rect 13996 33293 14036 33496
rect 14092 33461 14132 34336
rect 14188 34327 14228 34336
rect 14284 33872 14324 34756
rect 14380 34637 14420 35680
rect 14476 35671 14516 35680
rect 14475 35048 14517 35057
rect 14475 35008 14476 35048
rect 14516 35008 14517 35048
rect 14475 34999 14517 35008
rect 14379 34628 14421 34637
rect 14379 34588 14380 34628
rect 14420 34588 14421 34628
rect 14379 34579 14421 34588
rect 14476 34460 14516 34999
rect 14572 34469 14612 36856
rect 14380 34420 14516 34460
rect 14571 34460 14613 34469
rect 14571 34420 14572 34460
rect 14612 34420 14613 34460
rect 14380 34373 14420 34420
rect 14571 34411 14613 34420
rect 14380 34324 14420 34333
rect 14572 34217 14612 34302
rect 14379 34208 14421 34217
rect 14379 34168 14380 34208
rect 14420 34168 14421 34208
rect 14379 34159 14421 34168
rect 14571 34208 14613 34217
rect 14571 34168 14572 34208
rect 14612 34168 14613 34208
rect 14571 34159 14613 34168
rect 14284 33823 14324 33832
rect 14188 33704 14228 33713
rect 14091 33452 14133 33461
rect 14091 33412 14092 33452
rect 14132 33412 14133 33452
rect 14091 33403 14133 33412
rect 13995 33284 14037 33293
rect 13995 33244 13996 33284
rect 14036 33244 14037 33284
rect 13995 33235 14037 33244
rect 13995 33116 14037 33125
rect 13995 33076 13996 33116
rect 14036 33076 14037 33116
rect 13995 33067 14037 33076
rect 13996 32873 14036 33067
rect 14188 33041 14228 33664
rect 14187 33032 14229 33041
rect 14187 32992 14188 33032
rect 14228 32992 14229 33032
rect 14187 32983 14229 32992
rect 13995 32864 14037 32873
rect 14380 32864 14420 34159
rect 14668 34040 14708 37780
rect 14860 37400 14900 39199
rect 15243 39080 15285 39089
rect 15243 39040 15244 39080
rect 15284 39040 15285 39080
rect 15243 39031 15285 39040
rect 15051 37988 15093 37997
rect 15051 37948 15052 37988
rect 15092 37948 15093 37988
rect 15051 37939 15093 37948
rect 15052 37652 15092 37939
rect 15052 37603 15092 37612
rect 14764 37360 14860 37400
rect 14764 35225 14804 37360
rect 14860 37351 14900 37360
rect 14859 35888 14901 35897
rect 14859 35848 14860 35888
rect 14900 35848 14901 35888
rect 14859 35839 14901 35848
rect 14763 35216 14805 35225
rect 14763 35176 14764 35216
rect 14804 35176 14805 35216
rect 14763 35167 14805 35176
rect 14764 34376 14804 35167
rect 14764 34049 14804 34336
rect 14572 34000 14708 34040
rect 14763 34040 14805 34049
rect 14763 34000 14764 34040
rect 14804 34000 14805 34040
rect 14475 33704 14517 33713
rect 14475 33664 14476 33704
rect 14516 33664 14517 33704
rect 14475 33655 14517 33664
rect 14476 33570 14516 33655
rect 13995 32824 13996 32864
rect 14036 32824 14037 32864
rect 13995 32815 14037 32824
rect 14092 32824 14420 32864
rect 13996 32730 14036 32815
rect 13708 32656 13940 32696
rect 12844 32404 13652 32444
rect 12651 32276 12693 32285
rect 12651 32236 12652 32276
rect 12692 32236 12693 32276
rect 12651 32227 12693 32236
rect 13515 32276 13557 32285
rect 13515 32236 13516 32276
rect 13556 32236 13557 32276
rect 13515 32227 13557 32236
rect 12652 32192 12692 32227
rect 12652 32141 12692 32152
rect 12843 32192 12885 32201
rect 12843 32152 12844 32192
rect 12884 32152 12885 32192
rect 12843 32143 12885 32152
rect 12940 32192 12980 32201
rect 13035 32192 13077 32201
rect 12980 32152 13036 32192
rect 13076 32152 13077 32192
rect 12940 32143 12980 32152
rect 13035 32143 13077 32152
rect 13132 32192 13172 32201
rect 13419 32192 13461 32201
rect 13172 32152 13268 32192
rect 13132 32143 13172 32152
rect 12844 32058 12884 32143
rect 12940 31940 12980 31949
rect 12980 31900 13076 31940
rect 12940 31891 12980 31900
rect 12939 31604 12981 31613
rect 12939 31564 12940 31604
rect 12980 31564 12981 31604
rect 12939 31555 12981 31564
rect 12747 31520 12789 31529
rect 12747 31480 12748 31520
rect 12788 31480 12789 31520
rect 12747 31471 12789 31480
rect 12748 31352 12788 31471
rect 12940 31470 12980 31555
rect 12748 31109 12788 31312
rect 12939 31184 12981 31193
rect 12939 31144 12940 31184
rect 12980 31144 12981 31184
rect 12939 31135 12981 31144
rect 12747 31100 12789 31109
rect 12747 31060 12748 31100
rect 12788 31060 12789 31100
rect 12747 31051 12789 31060
rect 12940 30680 12980 31135
rect 12652 30640 12940 30680
rect 12652 29840 12692 30640
rect 12940 30631 12980 30640
rect 13036 30680 13076 31900
rect 13228 31613 13268 32152
rect 13419 32152 13420 32192
rect 13460 32152 13461 32192
rect 13419 32143 13461 32152
rect 13227 31604 13269 31613
rect 13227 31564 13228 31604
rect 13268 31564 13269 31604
rect 13227 31555 13269 31564
rect 12747 30512 12789 30521
rect 12747 30472 12748 30512
rect 12788 30472 12789 30512
rect 12747 30463 12789 30472
rect 12748 30378 12788 30463
rect 12652 29791 12692 29800
rect 12940 29840 12980 29849
rect 13036 29840 13076 30640
rect 13132 31352 13172 31361
rect 13228 31352 13268 31555
rect 13324 31352 13364 31361
rect 13228 31312 13324 31352
rect 13132 30521 13172 31312
rect 13324 31303 13364 31312
rect 13227 31184 13269 31193
rect 13227 31144 13228 31184
rect 13268 31144 13269 31184
rect 13227 31135 13269 31144
rect 13228 31050 13268 31135
rect 13323 31100 13365 31109
rect 13323 31060 13324 31100
rect 13364 31060 13365 31100
rect 13323 31051 13365 31060
rect 13228 30848 13268 30859
rect 13228 30773 13268 30808
rect 13227 30764 13269 30773
rect 13227 30724 13228 30764
rect 13268 30724 13269 30764
rect 13227 30715 13269 30724
rect 13131 30512 13173 30521
rect 13131 30472 13132 30512
rect 13172 30472 13173 30512
rect 13131 30463 13173 30472
rect 12980 29800 13076 29840
rect 13228 29840 13268 29849
rect 12940 29791 12980 29800
rect 13131 29756 13173 29765
rect 13131 29716 13132 29756
rect 13172 29716 13173 29756
rect 13131 29707 13173 29716
rect 12748 29672 12788 29681
rect 13035 29672 13077 29681
rect 12788 29632 12980 29672
rect 12748 29623 12788 29632
rect 12940 29168 12980 29632
rect 13035 29632 13036 29672
rect 13076 29632 13077 29672
rect 13035 29623 13077 29632
rect 12747 28580 12789 28589
rect 12747 28540 12748 28580
rect 12788 28540 12789 28580
rect 12747 28531 12789 28540
rect 12651 28412 12693 28421
rect 12651 28372 12652 28412
rect 12692 28372 12693 28412
rect 12651 28363 12693 28372
rect 12652 24641 12692 28363
rect 12748 28337 12788 28531
rect 12747 28328 12789 28337
rect 12747 28288 12748 28328
rect 12788 28288 12789 28328
rect 12747 28279 12789 28288
rect 12651 24632 12693 24641
rect 12651 24592 12652 24632
rect 12692 24592 12693 24632
rect 12651 24583 12693 24592
rect 12652 24498 12692 24583
rect 12748 23969 12788 28279
rect 12844 26816 12884 26825
rect 12940 26816 12980 29128
rect 13036 27656 13076 29623
rect 13132 29513 13172 29707
rect 13131 29504 13173 29513
rect 13131 29464 13132 29504
rect 13172 29464 13173 29504
rect 13131 29455 13173 29464
rect 13132 28328 13172 29455
rect 13228 28589 13268 29800
rect 13324 29000 13364 31051
rect 13420 30773 13460 32143
rect 13516 31940 13556 32227
rect 13612 32192 13652 32404
rect 13708 32360 13748 32656
rect 13708 32311 13748 32320
rect 13804 32192 13844 32201
rect 13612 32152 13804 32192
rect 13804 32143 13844 32152
rect 13516 31900 13844 31940
rect 13515 31352 13557 31361
rect 13515 31312 13516 31352
rect 13556 31312 13557 31352
rect 13515 31303 13557 31312
rect 13516 31218 13556 31303
rect 13804 30848 13844 31900
rect 13804 30808 13940 30848
rect 13419 30764 13461 30773
rect 13419 30724 13420 30764
rect 13460 30724 13652 30764
rect 13419 30715 13461 30724
rect 13612 29924 13652 30724
rect 13708 30680 13748 30689
rect 13708 30101 13748 30640
rect 13803 30680 13845 30689
rect 13803 30640 13804 30680
rect 13844 30640 13845 30680
rect 13803 30631 13845 30640
rect 13804 30546 13844 30631
rect 13707 30092 13749 30101
rect 13707 30052 13708 30092
rect 13748 30052 13749 30092
rect 13707 30043 13749 30052
rect 13612 29884 13748 29924
rect 13611 29336 13653 29345
rect 13611 29296 13612 29336
rect 13652 29296 13653 29336
rect 13611 29287 13653 29296
rect 13612 29202 13652 29287
rect 13468 29126 13508 29135
rect 13468 29084 13508 29086
rect 13468 29044 13604 29084
rect 13564 29000 13604 29044
rect 13324 28960 13460 29000
rect 13227 28580 13269 28589
rect 13227 28540 13228 28580
rect 13268 28540 13269 28580
rect 13227 28531 13269 28540
rect 13324 28328 13364 28337
rect 13132 28288 13324 28328
rect 13324 28279 13364 28288
rect 13036 27607 13076 27616
rect 13227 27656 13269 27665
rect 13227 27616 13228 27656
rect 13268 27616 13269 27656
rect 13227 27607 13269 27616
rect 12884 26776 12980 26816
rect 12844 26767 12884 26776
rect 12172 23920 12308 23960
rect 11691 23911 11733 23920
rect 11499 23792 11541 23801
rect 11499 23752 11500 23792
rect 11540 23752 11541 23792
rect 11499 23743 11541 23752
rect 11692 23792 11732 23801
rect 11500 23658 11540 23743
rect 11692 23288 11732 23752
rect 11883 23792 11925 23801
rect 11883 23752 11884 23792
rect 11924 23752 11925 23792
rect 11883 23743 11925 23752
rect 12075 23792 12117 23801
rect 12075 23752 12076 23792
rect 12116 23752 12117 23792
rect 12075 23743 12117 23752
rect 12172 23792 12212 23801
rect 11884 23658 11924 23743
rect 12076 23658 12116 23743
rect 11692 23239 11732 23248
rect 12075 23288 12117 23297
rect 12075 23248 12076 23288
rect 12116 23248 12117 23288
rect 12075 23239 12117 23248
rect 11499 23204 11541 23213
rect 11499 23164 11500 23204
rect 11540 23164 11541 23204
rect 11499 23155 11541 23164
rect 11500 23070 11540 23155
rect 11691 23120 11733 23129
rect 11691 23080 11692 23120
rect 11732 23080 11733 23120
rect 11691 23071 11733 23080
rect 11884 23106 11924 23115
rect 11595 22280 11637 22289
rect 11595 22240 11596 22280
rect 11636 22240 11637 22280
rect 11595 22231 11637 22240
rect 11692 22280 11732 23071
rect 11787 22532 11829 22541
rect 11787 22492 11788 22532
rect 11828 22492 11829 22532
rect 11787 22483 11829 22492
rect 11692 22231 11732 22240
rect 11788 22280 11828 22483
rect 11884 22373 11924 23066
rect 12076 22961 12116 23239
rect 12075 22952 12117 22961
rect 12075 22912 12076 22952
rect 12116 22912 12117 22952
rect 12075 22903 12117 22912
rect 11979 22700 12021 22709
rect 11979 22660 11980 22700
rect 12020 22660 12021 22700
rect 11979 22651 12021 22660
rect 11883 22364 11925 22373
rect 11883 22324 11884 22364
rect 11924 22324 11925 22364
rect 11883 22315 11925 22324
rect 11788 22231 11828 22240
rect 11884 22280 11924 22315
rect 11596 22146 11636 22231
rect 11884 22230 11924 22240
rect 11980 22112 12020 22651
rect 12172 22457 12212 23752
rect 12171 22448 12213 22457
rect 12171 22408 12172 22448
rect 12212 22408 12213 22448
rect 12171 22399 12213 22408
rect 12075 22364 12117 22373
rect 12075 22324 12076 22364
rect 12116 22324 12117 22364
rect 12075 22315 12117 22324
rect 12076 22196 12116 22315
rect 12172 22280 12212 22289
rect 12172 22205 12212 22240
rect 12171 22196 12213 22205
rect 12076 22156 12172 22196
rect 12212 22156 12213 22196
rect 12171 22147 12213 22156
rect 11788 22072 12020 22112
rect 11404 21904 11732 21944
rect 11307 21692 11349 21701
rect 11307 21652 11308 21692
rect 11348 21652 11349 21692
rect 11307 21643 11349 21652
rect 11404 21608 11444 21619
rect 11404 21533 11444 21568
rect 11403 21524 11445 21533
rect 11403 21484 11404 21524
rect 11444 21484 11445 21524
rect 11403 21475 11445 21484
rect 11307 21104 11349 21113
rect 11307 21064 11308 21104
rect 11348 21064 11349 21104
rect 11307 21055 11349 21064
rect 10828 20609 10868 20728
rect 11020 20812 11156 20852
rect 10827 20600 10869 20609
rect 10827 20560 10828 20600
rect 10868 20560 10869 20600
rect 10827 20551 10869 20560
rect 10348 20047 10388 20056
rect 10444 20308 10772 20348
rect 10251 19676 10293 19685
rect 10251 19636 10252 19676
rect 10292 19636 10293 19676
rect 10251 19627 10293 19636
rect 10204 19265 10244 19274
rect 10244 19225 10292 19256
rect 10204 19216 10292 19225
rect 10060 19132 10196 19172
rect 10059 18500 10101 18509
rect 10059 18460 10060 18500
rect 10100 18460 10101 18500
rect 10059 18451 10101 18460
rect 9963 18248 10005 18257
rect 9963 18208 9964 18248
rect 10004 18208 10005 18248
rect 9963 18199 10005 18208
rect 9868 17023 9908 17032
rect 9964 17072 10004 18199
rect 10060 17921 10100 18451
rect 10156 18005 10196 19132
rect 10155 17996 10197 18005
rect 10155 17956 10156 17996
rect 10196 17956 10197 17996
rect 10252 17996 10292 19216
rect 10347 19088 10389 19097
rect 10347 19048 10348 19088
rect 10388 19048 10389 19088
rect 10347 19039 10389 19048
rect 10348 18954 10388 19039
rect 10348 17996 10388 18005
rect 10252 17956 10348 17996
rect 10155 17947 10197 17956
rect 10348 17947 10388 17956
rect 10059 17912 10101 17921
rect 10059 17872 10060 17912
rect 10100 17872 10101 17912
rect 10059 17863 10101 17872
rect 10156 17753 10196 17838
rect 10251 17828 10293 17837
rect 10251 17788 10252 17828
rect 10292 17788 10293 17828
rect 10251 17779 10293 17788
rect 10155 17744 10197 17753
rect 10155 17704 10156 17744
rect 10196 17704 10197 17744
rect 10155 17695 10197 17704
rect 10252 17324 10292 17779
rect 9964 17023 10004 17032
rect 10156 17284 10292 17324
rect 9675 16484 9717 16493
rect 9675 16444 9676 16484
rect 9716 16444 9717 16484
rect 9675 16435 9717 16444
rect 9292 16232 9332 16241
rect 9292 14972 9332 16192
rect 9388 16232 9428 16243
rect 9388 16157 9428 16192
rect 9387 16148 9429 16157
rect 9387 16108 9388 16148
rect 9428 16108 9429 16148
rect 9387 16099 9429 16108
rect 9484 14972 9524 14981
rect 9292 14932 9484 14972
rect 9484 14923 9524 14932
rect 9291 14720 9333 14729
rect 9291 14680 9292 14720
rect 9332 14680 9333 14720
rect 9676 14720 9716 16435
rect 9867 16316 9909 16325
rect 9867 16276 9868 16316
rect 9908 16276 9909 16316
rect 9867 16267 9909 16276
rect 9771 16232 9813 16241
rect 9771 16192 9772 16232
rect 9812 16192 9813 16232
rect 9771 16183 9813 16192
rect 9772 14888 9812 16183
rect 9868 16182 9908 16267
rect 10059 16232 10101 16241
rect 10059 16192 10060 16232
rect 10100 16192 10101 16232
rect 10059 16183 10101 16192
rect 9963 15224 10005 15233
rect 9963 15184 9964 15224
rect 10004 15184 10005 15224
rect 9963 15175 10005 15184
rect 9772 14848 9908 14888
rect 9772 14720 9812 14729
rect 9676 14680 9772 14720
rect 9291 14671 9333 14680
rect 9772 14671 9812 14680
rect 9292 14225 9332 14671
rect 9291 14216 9333 14225
rect 9291 14176 9292 14216
rect 9332 14176 9333 14216
rect 9291 14167 9333 14176
rect 9484 14141 9524 14143
rect 9483 14132 9525 14141
rect 9483 14092 9484 14132
rect 9524 14092 9525 14132
rect 9483 14083 9525 14092
rect 9388 14048 9428 14057
rect 9292 14008 9388 14048
rect 9292 12620 9332 14008
rect 9388 13999 9428 14008
rect 9484 14048 9524 14083
rect 9484 13999 9524 14008
rect 9868 14048 9908 14848
rect 9579 13880 9621 13889
rect 9579 13840 9580 13880
rect 9620 13840 9621 13880
rect 9579 13831 9621 13840
rect 9387 13796 9429 13805
rect 9387 13756 9388 13796
rect 9428 13756 9429 13796
rect 9387 13747 9429 13756
rect 9292 12571 9332 12580
rect 9388 12452 9428 13747
rect 9100 8128 9236 8168
rect 9292 12412 9428 12452
rect 9484 12536 9524 12545
rect 9003 7580 9045 7589
rect 9003 7540 9004 7580
rect 9044 7540 9045 7580
rect 9003 7531 9045 7540
rect 8812 7204 8948 7244
rect 8620 7160 8660 7171
rect 8620 7085 8660 7120
rect 8619 7076 8661 7085
rect 8619 7036 8620 7076
rect 8660 7036 8661 7076
rect 8619 7027 8661 7036
rect 8524 6868 8660 6908
rect 8620 6473 8660 6868
rect 8715 6656 8757 6665
rect 8715 6616 8716 6656
rect 8756 6616 8757 6656
rect 8715 6607 8757 6616
rect 8716 6522 8756 6607
rect 8620 6433 8756 6473
rect 8428 6364 8564 6404
rect 8043 6236 8085 6245
rect 8043 6196 8044 6236
rect 8084 6196 8085 6236
rect 8043 6187 8085 6196
rect 8427 6236 8469 6245
rect 8427 6196 8428 6236
rect 8468 6196 8469 6236
rect 8427 6187 8469 6196
rect 7604 5608 7700 5648
rect 8044 5662 8084 6187
rect 8428 6102 8468 6187
rect 8524 6152 8564 6364
rect 8524 6112 8660 6152
rect 8523 5984 8565 5993
rect 8523 5944 8524 5984
rect 8564 5944 8565 5984
rect 8523 5935 8565 5944
rect 8044 5613 8084 5622
rect 8524 5648 8564 5935
rect 7564 5599 7604 5608
rect 8524 5599 8564 5608
rect 8236 5480 8276 5489
rect 8276 5440 8372 5480
rect 8236 5431 8276 5440
rect 7468 5188 7604 5228
rect 6987 5179 7029 5188
rect 6988 4976 7028 5179
rect 7276 5104 7508 5144
rect 6988 4927 7028 4936
rect 7180 5060 7220 5069
rect 7276 5060 7316 5104
rect 7220 5020 7316 5060
rect 6796 4600 6932 4640
rect 6699 2372 6741 2381
rect 6699 2332 6700 2372
rect 6740 2332 6741 2372
rect 6699 2323 6741 2332
rect 6603 2204 6645 2213
rect 6603 2164 6604 2204
rect 6644 2164 6645 2204
rect 6603 2155 6645 2164
rect 5932 2071 5972 2080
rect 6604 2120 6644 2155
rect 6604 2069 6644 2080
rect 6796 1952 6836 4600
rect 7083 4556 7125 4565
rect 7083 4516 7084 4556
rect 7124 4516 7125 4556
rect 7083 4507 7125 4516
rect 6891 4472 6933 4481
rect 6891 4432 6892 4472
rect 6932 4432 6933 4472
rect 6891 4423 6933 4432
rect 6892 4136 6932 4423
rect 6892 2540 6932 4096
rect 7084 4136 7124 4507
rect 7084 4087 7124 4096
rect 7180 4136 7220 5020
rect 7372 4976 7412 4985
rect 7180 4087 7220 4096
rect 7276 4936 7372 4976
rect 6988 3968 7028 3977
rect 7276 3968 7316 4936
rect 7372 4927 7412 4936
rect 7468 4976 7508 5104
rect 7468 4927 7508 4936
rect 7564 4808 7604 5188
rect 7659 5060 7701 5069
rect 7659 5020 7660 5060
rect 7700 5020 7701 5060
rect 7659 5011 7701 5020
rect 7660 4976 7700 5011
rect 7660 4925 7700 4936
rect 7755 4976 7797 4985
rect 7857 4976 7897 4985
rect 7755 4936 7756 4976
rect 7796 4936 7797 4976
rect 7755 4927 7797 4936
rect 7852 4936 7857 4976
rect 7852 4927 7897 4936
rect 7468 4768 7604 4808
rect 7371 4724 7413 4733
rect 7371 4684 7372 4724
rect 7412 4684 7413 4724
rect 7371 4675 7413 4684
rect 7372 4590 7412 4675
rect 7468 4481 7508 4768
rect 7756 4565 7796 4927
rect 7852 4649 7892 4927
rect 7851 4640 7893 4649
rect 7851 4600 7852 4640
rect 7892 4600 7893 4640
rect 7851 4591 7893 4600
rect 7755 4556 7797 4565
rect 7755 4516 7756 4556
rect 7796 4516 7797 4556
rect 7755 4507 7797 4516
rect 7467 4472 7509 4481
rect 7467 4432 7468 4472
rect 7508 4432 7509 4472
rect 7467 4423 7509 4432
rect 7852 4220 7892 4591
rect 7852 4180 7897 4220
rect 7857 4145 7897 4180
rect 7028 3928 7316 3968
rect 7372 4136 7412 4145
rect 6988 3919 7028 3928
rect 7372 3296 7412 4096
rect 7468 4136 7508 4145
rect 7468 3557 7508 4096
rect 7660 4136 7700 4145
rect 7660 3977 7700 4096
rect 7756 4136 7796 4145
rect 7857 4136 7924 4145
rect 7857 4096 7884 4136
rect 7564 3968 7604 3977
rect 7467 3548 7509 3557
rect 7467 3508 7468 3548
rect 7508 3508 7509 3548
rect 7467 3499 7509 3508
rect 7564 3305 7604 3928
rect 7659 3968 7701 3977
rect 7659 3928 7660 3968
rect 7700 3928 7701 3968
rect 7659 3919 7701 3928
rect 7756 3716 7796 4096
rect 7884 4087 7924 4096
rect 8235 3968 8277 3977
rect 8235 3928 8236 3968
rect 8276 3928 8277 3968
rect 8332 3968 8372 5440
rect 8620 5312 8660 6112
rect 8524 5272 8660 5312
rect 8427 5228 8469 5237
rect 8427 5188 8428 5228
rect 8468 5188 8469 5228
rect 8427 5179 8469 5188
rect 8428 4976 8468 5179
rect 8428 4927 8468 4936
rect 8332 3928 8468 3968
rect 8235 3919 8277 3928
rect 8236 3800 8276 3919
rect 8236 3760 8372 3800
rect 7756 3676 7892 3716
rect 7852 3632 7892 3676
rect 7852 3583 7892 3592
rect 8235 3632 8277 3641
rect 8235 3592 8236 3632
rect 8276 3592 8277 3632
rect 8235 3583 8277 3592
rect 8332 3632 8372 3760
rect 8332 3583 8372 3592
rect 7755 3548 7797 3557
rect 7755 3508 7756 3548
rect 7796 3508 7797 3548
rect 7755 3499 7797 3508
rect 7660 3464 7700 3475
rect 7660 3389 7700 3424
rect 7659 3380 7701 3389
rect 7659 3340 7660 3380
rect 7700 3340 7701 3380
rect 7659 3331 7701 3340
rect 7563 3296 7605 3305
rect 7372 3256 7508 3296
rect 6892 2500 7412 2540
rect 6987 2120 7029 2129
rect 6987 2080 6988 2120
rect 7028 2080 7029 2120
rect 6987 2071 7029 2080
rect 6988 1986 7028 2071
rect 5740 1903 5780 1912
rect 6604 1912 6836 1952
rect 7372 1952 7412 2500
rect 7468 2120 7508 3256
rect 7563 3256 7564 3296
rect 7604 3256 7605 3296
rect 7563 3247 7605 3256
rect 7660 3128 7700 3331
rect 7564 3088 7700 3128
rect 7564 2624 7604 3088
rect 7756 2876 7796 3499
rect 8044 3464 8084 3473
rect 8044 3221 8084 3424
rect 8139 3464 8181 3473
rect 8139 3424 8140 3464
rect 8180 3424 8181 3464
rect 8139 3415 8181 3424
rect 8140 3330 8180 3415
rect 7851 3212 7893 3221
rect 7851 3172 7852 3212
rect 7892 3172 7893 3212
rect 7851 3163 7893 3172
rect 8043 3212 8085 3221
rect 8043 3172 8044 3212
rect 8084 3172 8085 3212
rect 8043 3163 8085 3172
rect 7564 2575 7604 2584
rect 7660 2836 7756 2876
rect 7468 2071 7508 2080
rect 6412 1868 6452 1877
rect 6220 1700 6260 1709
rect 6220 1373 6260 1660
rect 6219 1364 6261 1373
rect 6219 1324 6220 1364
rect 6260 1324 6261 1364
rect 6219 1315 6261 1324
rect 6123 1196 6165 1205
rect 6123 1156 6124 1196
rect 6164 1156 6165 1196
rect 6123 1147 6165 1156
rect 6124 1062 6164 1147
rect 6219 1112 6261 1121
rect 6219 1072 6220 1112
rect 6260 1072 6261 1112
rect 6219 1063 6261 1072
rect 5356 904 5684 944
rect 5931 944 5973 953
rect 5931 904 5932 944
rect 5972 904 5973 944
rect 5931 895 5973 904
rect 5835 860 5877 869
rect 5835 820 5836 860
rect 5876 820 5877 860
rect 5835 811 5877 820
rect 4928 776 5296 785
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 4928 727 5296 736
rect 4875 608 4917 617
rect 4875 568 4876 608
rect 4916 568 4917 608
rect 4875 559 4917 568
rect 5067 608 5109 617
rect 5067 568 5068 608
rect 5108 568 5109 608
rect 5067 559 5109 568
rect 4876 80 4916 559
rect 5068 80 5108 559
rect 5451 524 5493 533
rect 5451 484 5452 524
rect 5492 484 5493 524
rect 5451 475 5493 484
rect 5259 188 5301 197
rect 5259 148 5260 188
rect 5300 148 5301 188
rect 5259 139 5301 148
rect 5260 80 5300 139
rect 5452 80 5492 475
rect 5643 440 5685 449
rect 5643 400 5644 440
rect 5684 400 5685 440
rect 5643 391 5685 400
rect 5644 80 5684 391
rect 5836 80 5876 811
rect 5932 810 5972 895
rect 6027 272 6069 281
rect 6027 232 6028 272
rect 6068 232 6069 272
rect 6027 223 6069 232
rect 6028 80 6068 223
rect 6220 80 6260 1063
rect 6412 1037 6452 1828
rect 6508 1196 6548 1205
rect 6411 1028 6453 1037
rect 6411 988 6412 1028
rect 6452 988 6453 1028
rect 6411 979 6453 988
rect 6315 944 6357 953
rect 6315 904 6316 944
rect 6356 904 6357 944
rect 6315 895 6357 904
rect 6316 810 6356 895
rect 6411 776 6453 785
rect 6411 736 6412 776
rect 6452 736 6453 776
rect 6411 727 6453 736
rect 6412 80 6452 727
rect 6508 617 6548 1156
rect 6507 608 6549 617
rect 6507 568 6508 608
rect 6548 568 6549 608
rect 6507 559 6549 568
rect 6604 449 6644 1912
rect 7372 1903 7412 1912
rect 7564 1952 7604 1961
rect 7180 1868 7220 1877
rect 6796 1857 6836 1866
rect 6796 1457 6836 1817
rect 6795 1448 6837 1457
rect 6795 1408 6796 1448
rect 6836 1408 6837 1448
rect 6795 1399 6837 1408
rect 7180 1373 7220 1828
rect 7564 1784 7604 1912
rect 7660 1952 7700 2836
rect 7756 2827 7796 2836
rect 7852 2540 7892 3163
rect 8140 2624 8180 2633
rect 8236 2624 8276 3583
rect 8428 2801 8468 3928
rect 8427 2792 8469 2801
rect 8427 2752 8428 2792
rect 8468 2752 8469 2792
rect 8427 2743 8469 2752
rect 8180 2584 8276 2624
rect 8140 2575 8180 2584
rect 7660 1903 7700 1912
rect 7756 2500 7892 2540
rect 7756 1784 7796 2500
rect 7851 1868 7893 1877
rect 7851 1828 7852 1868
rect 7892 1828 7893 1868
rect 7851 1819 7893 1828
rect 8235 1868 8277 1877
rect 8235 1828 8236 1868
rect 8276 1828 8277 1868
rect 8235 1819 8277 1828
rect 7564 1744 7796 1784
rect 7852 1734 7892 1819
rect 8236 1734 8276 1819
rect 8044 1700 8084 1709
rect 8428 1700 8468 1709
rect 8084 1660 8180 1700
rect 8044 1651 8084 1660
rect 7851 1448 7893 1457
rect 7851 1408 7852 1448
rect 7892 1408 7893 1448
rect 7851 1399 7893 1408
rect 7179 1364 7221 1373
rect 7179 1324 7180 1364
rect 7220 1324 7221 1364
rect 7179 1315 7221 1324
rect 6699 1280 6741 1289
rect 6699 1240 6700 1280
rect 6740 1240 6741 1280
rect 6699 1231 6741 1240
rect 7371 1280 7413 1289
rect 7371 1240 7372 1280
rect 7412 1240 7413 1280
rect 7371 1231 7413 1240
rect 7755 1280 7797 1289
rect 7755 1240 7756 1280
rect 7796 1240 7797 1280
rect 7755 1231 7797 1240
rect 6700 1146 6740 1231
rect 6892 1196 6932 1205
rect 6795 944 6837 953
rect 6795 904 6796 944
rect 6836 904 6837 944
rect 6795 895 6837 904
rect 6603 440 6645 449
rect 6603 400 6604 440
rect 6644 400 6645 440
rect 6603 391 6645 400
rect 6603 188 6645 197
rect 6603 148 6604 188
rect 6644 148 6645 188
rect 6603 139 6645 148
rect 6604 80 6644 139
rect 6796 80 6836 895
rect 6892 449 6932 1156
rect 7179 1196 7221 1205
rect 7179 1156 7180 1196
rect 7220 1156 7221 1196
rect 7179 1147 7221 1156
rect 6987 776 7029 785
rect 6987 736 6988 776
rect 7028 736 7029 776
rect 6987 727 7029 736
rect 6891 440 6933 449
rect 6891 400 6892 440
rect 6932 400 6933 440
rect 6891 391 6933 400
rect 6988 80 7028 727
rect 7180 80 7220 1147
rect 7372 1146 7412 1231
rect 7564 1196 7604 1205
rect 7564 617 7604 1156
rect 7756 1146 7796 1231
rect 7755 1028 7797 1037
rect 7755 988 7756 1028
rect 7796 988 7797 1028
rect 7755 979 7797 988
rect 7371 608 7413 617
rect 7371 568 7372 608
rect 7412 568 7413 608
rect 7371 559 7413 568
rect 7563 608 7605 617
rect 7563 568 7564 608
rect 7604 568 7605 608
rect 7563 559 7605 568
rect 7372 80 7412 559
rect 7563 440 7605 449
rect 7563 400 7564 440
rect 7604 400 7605 440
rect 7563 391 7605 400
rect 7564 80 7604 391
rect 7756 80 7796 979
rect 7852 944 7892 1399
rect 8043 1364 8085 1373
rect 8043 1324 8044 1364
rect 8084 1324 8085 1364
rect 8043 1315 8085 1324
rect 7947 1196 7989 1205
rect 7947 1156 7948 1196
rect 7988 1156 7989 1196
rect 7947 1147 7989 1156
rect 7948 1062 7988 1147
rect 8044 1028 8084 1315
rect 8140 1289 8180 1660
rect 8428 1541 8468 1660
rect 8427 1532 8469 1541
rect 8427 1492 8428 1532
rect 8468 1492 8469 1532
rect 8427 1483 8469 1492
rect 8524 1448 8564 5272
rect 8619 4640 8661 4649
rect 8619 4600 8620 4640
rect 8660 4600 8661 4640
rect 8619 4591 8661 4600
rect 8620 4061 8660 4591
rect 8619 4052 8661 4061
rect 8619 4012 8620 4052
rect 8660 4012 8661 4052
rect 8619 4003 8661 4012
rect 8619 3464 8661 3473
rect 8619 3424 8620 3464
rect 8660 3424 8661 3464
rect 8619 3415 8661 3424
rect 8620 3330 8660 3415
rect 8716 2540 8756 6433
rect 8812 4901 8852 7204
rect 8907 6908 8949 6917
rect 8907 6868 8908 6908
rect 8948 6868 8949 6908
rect 8907 6859 8949 6868
rect 8908 6488 8948 6859
rect 9003 6572 9045 6581
rect 9003 6532 9004 6572
rect 9044 6532 9045 6572
rect 9003 6523 9045 6532
rect 8908 6439 8948 6448
rect 9004 6488 9044 6523
rect 9004 6437 9044 6448
rect 8811 4892 8853 4901
rect 8811 4852 8812 4892
rect 8852 4852 8853 4892
rect 8811 4843 8853 4852
rect 9100 2540 9140 8128
rect 9196 8000 9236 8011
rect 9196 7925 9236 7960
rect 9195 7916 9237 7925
rect 9195 7876 9196 7916
rect 9236 7876 9237 7916
rect 9195 7867 9237 7876
rect 9195 7160 9237 7169
rect 9195 7120 9196 7160
rect 9236 7120 9237 7160
rect 9195 7111 9237 7120
rect 9196 7026 9236 7111
rect 9195 6572 9237 6581
rect 9195 6532 9196 6572
rect 9236 6532 9237 6572
rect 9195 6523 9237 6532
rect 9196 6438 9236 6523
rect 8620 2500 8756 2540
rect 8812 2500 9140 2540
rect 8620 1868 8660 2500
rect 8812 1877 8852 2500
rect 8620 1819 8660 1828
rect 8811 1868 8853 1877
rect 8811 1828 8812 1868
rect 8852 1828 8853 1868
rect 8811 1819 8853 1828
rect 9004 1868 9044 1877
rect 9004 1709 9044 1828
rect 8812 1700 8852 1709
rect 8524 1408 8660 1448
rect 8139 1280 8181 1289
rect 8139 1240 8140 1280
rect 8180 1240 8181 1280
rect 8139 1231 8181 1240
rect 8523 1196 8565 1205
rect 8523 1156 8524 1196
rect 8564 1156 8565 1196
rect 8523 1147 8565 1156
rect 8044 988 8372 1028
rect 7852 904 7988 944
rect 7948 80 7988 904
rect 8139 608 8181 617
rect 8139 568 8140 608
rect 8180 568 8181 608
rect 8139 559 8181 568
rect 8140 80 8180 559
rect 8332 80 8372 988
rect 8524 80 8564 1147
rect 8620 701 8660 1408
rect 8715 1280 8757 1289
rect 8715 1240 8716 1280
rect 8756 1240 8757 1280
rect 8715 1231 8757 1240
rect 8619 692 8661 701
rect 8619 652 8620 692
rect 8660 652 8661 692
rect 8619 643 8661 652
rect 8716 80 8756 1231
rect 8812 869 8852 1660
rect 9003 1700 9045 1709
rect 9196 1700 9236 1709
rect 9003 1660 9004 1700
rect 9044 1660 9045 1700
rect 9003 1651 9045 1660
rect 9100 1660 9196 1700
rect 9003 1196 9045 1205
rect 9003 1156 9004 1196
rect 9044 1156 9045 1196
rect 9003 1147 9045 1156
rect 9004 1062 9044 1147
rect 8811 860 8853 869
rect 8811 820 8812 860
rect 8852 820 8853 860
rect 8811 811 8853 820
rect 9100 785 9140 1660
rect 9196 1651 9236 1660
rect 9195 1532 9237 1541
rect 9195 1492 9196 1532
rect 9236 1492 9237 1532
rect 9195 1483 9237 1492
rect 9196 1112 9236 1483
rect 9292 1196 9332 12412
rect 9484 12293 9524 12496
rect 9483 12284 9525 12293
rect 9483 12244 9484 12284
rect 9524 12244 9525 12284
rect 9483 12235 9525 12244
rect 9388 11696 9428 11707
rect 9388 11621 9428 11656
rect 9387 11612 9429 11621
rect 9387 11572 9388 11612
rect 9428 11572 9429 11612
rect 9387 11563 9429 11572
rect 9580 11360 9620 13831
rect 9772 13208 9812 13219
rect 9772 13133 9812 13168
rect 9771 13124 9813 13133
rect 9771 13084 9772 13124
rect 9812 13084 9813 13124
rect 9771 13075 9813 13084
rect 9868 11873 9908 14008
rect 9964 14048 10004 15175
rect 10060 14981 10100 16183
rect 10156 15989 10196 17284
rect 10444 17240 10484 20308
rect 10540 20180 10580 20189
rect 10580 20140 10868 20180
rect 10540 20131 10580 20140
rect 10828 20096 10868 20140
rect 10828 20047 10868 20056
rect 10924 20096 10964 20105
rect 10635 19844 10677 19853
rect 10635 19804 10636 19844
rect 10676 19804 10677 19844
rect 10635 19795 10677 19804
rect 10636 18593 10676 19795
rect 10924 18845 10964 20056
rect 10923 18836 10965 18845
rect 10923 18796 10924 18836
rect 10964 18796 10965 18836
rect 10923 18787 10965 18796
rect 11020 18761 11060 20812
rect 11308 20012 11348 21055
rect 11403 20096 11445 20105
rect 11403 20056 11404 20096
rect 11444 20056 11445 20096
rect 11403 20047 11445 20056
rect 11211 19508 11253 19517
rect 11211 19468 11212 19508
rect 11252 19468 11253 19508
rect 11211 19459 11253 19468
rect 11212 19256 11252 19459
rect 11212 19181 11252 19216
rect 11211 19172 11253 19181
rect 11211 19132 11212 19172
rect 11252 19132 11253 19172
rect 11211 19123 11253 19132
rect 11212 19092 11252 19123
rect 11115 18836 11157 18845
rect 11115 18796 11116 18836
rect 11156 18796 11157 18836
rect 11115 18787 11157 18796
rect 11019 18752 11061 18761
rect 11019 18712 11020 18752
rect 11060 18712 11061 18752
rect 11019 18703 11061 18712
rect 10732 18668 10772 18677
rect 10772 18628 10964 18668
rect 10732 18619 10772 18628
rect 10540 18584 10580 18593
rect 10540 17837 10580 18544
rect 10635 18584 10677 18593
rect 10635 18544 10636 18584
rect 10676 18544 10677 18584
rect 10924 18584 10964 18628
rect 11020 18584 11060 18593
rect 10924 18544 11020 18584
rect 10635 18535 10677 18544
rect 11020 18535 11060 18544
rect 11116 18584 11156 18787
rect 11211 18668 11253 18677
rect 11211 18628 11212 18668
rect 11252 18628 11253 18668
rect 11211 18619 11253 18628
rect 10539 17828 10581 17837
rect 10539 17788 10540 17828
rect 10580 17788 10581 17828
rect 10539 17779 10581 17788
rect 10539 17408 10581 17417
rect 10539 17368 10540 17408
rect 10580 17368 10581 17408
rect 10539 17359 10581 17368
rect 10252 17200 10484 17240
rect 10155 15980 10197 15989
rect 10155 15940 10156 15980
rect 10196 15940 10197 15980
rect 10155 15931 10197 15940
rect 10059 14972 10101 14981
rect 10059 14932 10060 14972
rect 10100 14932 10101 14972
rect 10059 14923 10101 14932
rect 9964 13999 10004 14008
rect 10252 13805 10292 17200
rect 10444 17072 10484 17081
rect 10540 17072 10580 17359
rect 10484 17032 10580 17072
rect 10348 16241 10388 16326
rect 10347 16232 10389 16241
rect 10347 16192 10348 16232
rect 10388 16192 10389 16232
rect 10347 16183 10389 16192
rect 10444 15140 10484 17032
rect 10636 16988 10676 18535
rect 10731 18248 10773 18257
rect 10731 18208 10732 18248
rect 10772 18208 10773 18248
rect 10731 18199 10773 18208
rect 10348 15100 10484 15140
rect 10540 16948 10676 16988
rect 10251 13796 10293 13805
rect 10251 13756 10252 13796
rect 10292 13756 10293 13796
rect 10251 13747 10293 13756
rect 9963 12620 10005 12629
rect 9963 12580 9964 12620
rect 10004 12580 10005 12620
rect 9963 12571 10005 12580
rect 9867 11864 9909 11873
rect 9867 11824 9868 11864
rect 9908 11824 9909 11864
rect 9867 11815 9909 11824
rect 9868 11701 9908 11710
rect 9484 11320 9620 11360
rect 9675 11360 9717 11369
rect 9675 11320 9676 11360
rect 9716 11320 9717 11360
rect 9387 7076 9429 7085
rect 9387 7036 9388 7076
rect 9428 7036 9429 7076
rect 9387 7027 9429 7036
rect 9388 6488 9428 7027
rect 9388 6439 9428 6448
rect 9387 2792 9429 2801
rect 9387 2752 9388 2792
rect 9428 2752 9429 2792
rect 9387 2743 9429 2752
rect 9388 2624 9428 2743
rect 9388 2575 9428 2584
rect 9387 2372 9429 2381
rect 9387 2332 9388 2372
rect 9428 2332 9429 2372
rect 9387 2323 9429 2332
rect 9388 1952 9428 2323
rect 9484 2204 9524 11320
rect 9675 11311 9717 11320
rect 9579 8588 9621 8597
rect 9579 8548 9580 8588
rect 9620 8548 9621 8588
rect 9579 8539 9621 8548
rect 9580 8009 9620 8539
rect 9579 8000 9621 8009
rect 9579 7960 9580 8000
rect 9620 7960 9621 8000
rect 9579 7951 9621 7960
rect 9580 4136 9620 7951
rect 9676 7925 9716 11311
rect 9868 11201 9908 11661
rect 9867 11192 9909 11201
rect 9867 11152 9868 11192
rect 9908 11152 9909 11192
rect 9867 11143 9909 11152
rect 9964 11024 10004 12571
rect 9964 10193 10004 10984
rect 10060 11528 10100 11537
rect 10060 10949 10100 11488
rect 10348 11360 10388 15100
rect 10443 14972 10485 14981
rect 10443 14932 10444 14972
rect 10484 14932 10485 14972
rect 10443 14923 10485 14932
rect 10444 14048 10484 14923
rect 10444 13999 10484 14008
rect 10540 13880 10580 16948
rect 10732 16904 10772 18199
rect 11116 17660 11156 18544
rect 11020 17620 11156 17660
rect 10923 17156 10965 17165
rect 10923 17116 10924 17156
rect 10964 17116 10965 17156
rect 10923 17107 10965 17116
rect 10924 17067 10964 17107
rect 10924 17018 10964 17027
rect 11020 16913 11060 17620
rect 11212 17417 11252 18619
rect 11308 18584 11348 19972
rect 11404 19962 11444 20047
rect 11500 18584 11540 18593
rect 11308 18544 11500 18584
rect 11500 18535 11540 18544
rect 11595 18500 11637 18509
rect 11595 18460 11596 18500
rect 11636 18460 11637 18500
rect 11595 18451 11637 18460
rect 11596 18366 11636 18451
rect 11595 18164 11637 18173
rect 11595 18124 11596 18164
rect 11636 18124 11637 18164
rect 11595 18115 11637 18124
rect 11403 17828 11445 17837
rect 11403 17788 11404 17828
rect 11444 17788 11445 17828
rect 11403 17779 11445 17788
rect 11211 17408 11253 17417
rect 11211 17368 11212 17408
rect 11252 17368 11253 17408
rect 11211 17359 11253 17368
rect 11116 17156 11156 17165
rect 10444 13840 10580 13880
rect 10636 16864 10772 16904
rect 11019 16904 11061 16913
rect 11019 16864 11020 16904
rect 11060 16864 11061 16904
rect 10636 15560 10676 16864
rect 11019 16855 11061 16864
rect 11116 16316 11156 17116
rect 11307 17156 11349 17165
rect 11307 17116 11308 17156
rect 11348 17116 11349 17156
rect 11307 17107 11349 17116
rect 11308 17022 11348 17107
rect 11404 17072 11444 17779
rect 11596 17753 11636 18115
rect 11500 17744 11540 17753
rect 11500 17501 11540 17704
rect 11595 17744 11637 17753
rect 11595 17704 11596 17744
rect 11636 17704 11637 17744
rect 11595 17695 11637 17704
rect 11499 17492 11541 17501
rect 11499 17452 11500 17492
rect 11540 17452 11541 17492
rect 11499 17443 11541 17452
rect 11500 17249 11540 17443
rect 11499 17240 11541 17249
rect 11499 17200 11500 17240
rect 11540 17200 11541 17240
rect 11499 17191 11541 17200
rect 11500 17072 11540 17081
rect 11404 17032 11500 17072
rect 11500 17023 11540 17032
rect 11116 16276 11348 16316
rect 10876 16241 10916 16250
rect 10916 16201 11252 16232
rect 10876 16192 11252 16201
rect 11019 16064 11061 16073
rect 11019 16024 11020 16064
rect 11060 16024 11061 16064
rect 11019 16015 11061 16024
rect 11020 15930 11060 16015
rect 10444 11537 10484 13840
rect 10636 12788 10676 15520
rect 11212 14972 11252 16192
rect 11212 14923 11252 14932
rect 11019 14720 11061 14729
rect 11019 14680 11020 14720
rect 11060 14680 11061 14720
rect 11019 14671 11061 14680
rect 11020 14586 11060 14671
rect 11116 14132 11156 14141
rect 10540 12748 10676 12788
rect 10828 14092 11116 14132
rect 10540 11705 10580 12748
rect 10731 12620 10773 12629
rect 10731 12580 10732 12620
rect 10772 12580 10773 12620
rect 10731 12571 10773 12580
rect 10732 12536 10772 12571
rect 10732 12485 10772 12496
rect 10732 11780 10772 11789
rect 10828 11780 10868 14092
rect 11116 14083 11156 14092
rect 10972 14006 11012 14015
rect 10972 13964 11012 13966
rect 10972 13924 11252 13964
rect 11212 13460 11252 13924
rect 11212 13411 11252 13420
rect 11020 13229 11060 13312
rect 11019 13177 11020 13226
rect 11060 13177 11061 13226
rect 11019 13168 11061 13177
rect 11308 12704 11348 16276
rect 11596 14720 11636 17695
rect 11692 15485 11732 21904
rect 11691 15476 11733 15485
rect 11691 15436 11692 15476
rect 11732 15436 11733 15476
rect 11691 15427 11733 15436
rect 11788 15224 11828 22072
rect 12172 22062 12212 22147
rect 12075 21524 12117 21533
rect 12075 21484 12076 21524
rect 12116 21484 12117 21524
rect 12075 21475 12117 21484
rect 11884 20054 11924 20063
rect 11883 20014 11884 20021
rect 11924 20014 11925 20021
rect 11883 20012 11925 20014
rect 11883 19972 11884 20012
rect 11924 19972 12020 20012
rect 11883 19963 11925 19972
rect 11884 19919 11924 19963
rect 11980 18584 12020 19972
rect 12076 18752 12116 21475
rect 12268 20777 12308 23920
rect 12460 23920 12596 23960
rect 12747 23960 12789 23969
rect 12747 23920 12748 23960
rect 12788 23920 12789 23960
rect 12363 23876 12405 23885
rect 12363 23836 12364 23876
rect 12404 23836 12405 23876
rect 12363 23827 12405 23836
rect 12364 23792 12404 23827
rect 12364 23741 12404 23752
rect 12363 23120 12405 23129
rect 12363 23080 12364 23120
rect 12404 23080 12405 23120
rect 12363 23071 12405 23080
rect 12364 22986 12404 23071
rect 12460 22448 12500 23920
rect 12747 23911 12789 23920
rect 12652 23801 12692 23886
rect 12556 23792 12596 23801
rect 12556 23624 12596 23752
rect 12651 23792 12693 23801
rect 12651 23752 12652 23792
rect 12692 23752 12693 23792
rect 12651 23743 12693 23752
rect 12844 23624 12884 23633
rect 12556 23584 12844 23624
rect 12844 23575 12884 23584
rect 12555 23456 12597 23465
rect 12940 23456 12980 26776
rect 13228 26144 13268 27607
rect 13420 27497 13460 28960
rect 13516 28960 13604 29000
rect 13708 29000 13748 29884
rect 13900 29849 13940 30808
rect 13899 29840 13941 29849
rect 13899 29800 13900 29840
rect 13940 29800 13941 29840
rect 13899 29791 13941 29800
rect 13708 28960 13844 29000
rect 13516 28580 13556 28960
rect 13516 28531 13556 28540
rect 13419 27488 13461 27497
rect 13419 27448 13420 27488
rect 13460 27448 13461 27488
rect 13419 27439 13461 27448
rect 13420 26993 13460 27439
rect 13419 26984 13461 26993
rect 13419 26944 13420 26984
rect 13460 26944 13461 26984
rect 13419 26935 13461 26944
rect 13372 26825 13412 26834
rect 13412 26785 13460 26816
rect 13372 26776 13460 26785
rect 13420 26312 13460 26776
rect 13515 26648 13557 26657
rect 13515 26608 13516 26648
rect 13556 26608 13557 26648
rect 13515 26599 13557 26608
rect 13516 26514 13556 26599
rect 13420 26263 13460 26272
rect 13228 26095 13268 26104
rect 13131 25892 13173 25901
rect 13131 25852 13132 25892
rect 13172 25852 13173 25892
rect 13131 25843 13173 25852
rect 13132 25304 13172 25843
rect 13132 25255 13172 25264
rect 13132 24632 13172 24641
rect 13132 23969 13172 24592
rect 13707 24128 13749 24137
rect 13707 24088 13708 24128
rect 13748 24088 13749 24128
rect 13707 24079 13749 24088
rect 13131 23960 13173 23969
rect 13131 23920 13132 23960
rect 13172 23920 13173 23960
rect 13131 23911 13173 23920
rect 13515 23876 13557 23885
rect 13515 23836 13516 23876
rect 13556 23836 13557 23876
rect 13515 23827 13557 23836
rect 12555 23416 12556 23456
rect 12596 23416 12597 23456
rect 12555 23407 12597 23416
rect 12748 23416 12980 23456
rect 13036 23792 13076 23801
rect 12556 23297 12596 23407
rect 12555 23288 12597 23297
rect 12555 23248 12556 23288
rect 12596 23248 12597 23288
rect 12555 23239 12597 23248
rect 12364 22408 12500 22448
rect 12267 20768 12309 20777
rect 12267 20728 12268 20768
rect 12308 20728 12309 20768
rect 12267 20719 12309 20728
rect 12268 20634 12308 20719
rect 12364 20348 12404 22408
rect 12460 22280 12500 22289
rect 12460 21785 12500 22240
rect 12556 22196 12596 22207
rect 12556 22121 12596 22156
rect 12555 22112 12597 22121
rect 12555 22072 12556 22112
rect 12596 22072 12597 22112
rect 12555 22063 12597 22072
rect 12459 21776 12501 21785
rect 12459 21736 12460 21776
rect 12500 21736 12501 21776
rect 12459 21727 12501 21736
rect 12556 21449 12596 22063
rect 12652 21701 12692 21732
rect 12651 21692 12693 21701
rect 12651 21652 12652 21692
rect 12692 21652 12693 21692
rect 12651 21643 12693 21652
rect 12652 21608 12692 21643
rect 12748 21617 12788 23416
rect 12843 23288 12885 23297
rect 12843 23248 12844 23288
rect 12884 23248 12885 23288
rect 12843 23239 12885 23248
rect 12844 23120 12884 23239
rect 12844 23071 12884 23080
rect 12939 23036 12981 23045
rect 12939 22996 12940 23036
rect 12980 22996 12981 23036
rect 12939 22987 12981 22996
rect 12940 22902 12980 22987
rect 12844 22532 12884 22541
rect 13036 22532 13076 23752
rect 13132 23792 13172 23801
rect 13516 23792 13556 23827
rect 13172 23752 13460 23792
rect 13132 23743 13172 23752
rect 13131 23624 13173 23633
rect 13131 23584 13132 23624
rect 13172 23584 13173 23624
rect 13131 23575 13173 23584
rect 13132 22709 13172 23575
rect 13420 23213 13460 23752
rect 13516 23741 13556 23752
rect 13612 23792 13652 23801
rect 13515 23624 13557 23633
rect 13515 23584 13516 23624
rect 13556 23584 13557 23624
rect 13515 23575 13557 23584
rect 13419 23204 13461 23213
rect 13419 23164 13420 23204
rect 13460 23164 13461 23204
rect 13419 23155 13461 23164
rect 13324 23120 13364 23129
rect 13131 22700 13173 22709
rect 13131 22660 13132 22700
rect 13172 22660 13173 22700
rect 13131 22651 13173 22660
rect 12884 22492 13076 22532
rect 12844 22483 12884 22492
rect 13131 22448 13173 22457
rect 13131 22408 13132 22448
rect 13172 22408 13173 22448
rect 13324 22448 13364 23080
rect 13420 23120 13460 23155
rect 13420 23070 13460 23080
rect 13324 22408 13460 22448
rect 13131 22399 13173 22408
rect 13035 22280 13077 22289
rect 13035 22240 13036 22280
rect 13076 22240 13077 22280
rect 13035 22231 13077 22240
rect 12843 22196 12885 22205
rect 12843 22156 12844 22196
rect 12884 22156 12885 22196
rect 12843 22147 12885 22156
rect 12844 21776 12884 22147
rect 13036 22146 13076 22231
rect 13132 22196 13172 22399
rect 13228 22280 13268 22291
rect 13228 22205 13268 22240
rect 13323 22280 13365 22289
rect 13323 22240 13324 22280
rect 13364 22240 13365 22280
rect 13323 22231 13365 22240
rect 13132 22147 13172 22156
rect 13227 22196 13269 22205
rect 13227 22156 13228 22196
rect 13268 22156 13269 22196
rect 13227 22147 13269 22156
rect 13324 22146 13364 22231
rect 13131 21944 13173 21953
rect 13131 21904 13132 21944
rect 13172 21904 13173 21944
rect 13131 21895 13173 21904
rect 12844 21727 12884 21736
rect 12555 21440 12597 21449
rect 12555 21400 12556 21440
rect 12596 21400 12597 21440
rect 12555 21391 12597 21400
rect 12652 20777 12692 21568
rect 12747 21608 12789 21617
rect 12747 21568 12748 21608
rect 12788 21568 12789 21608
rect 12747 21559 12789 21568
rect 12843 21440 12885 21449
rect 12843 21400 12844 21440
rect 12884 21400 12885 21440
rect 12843 21391 12885 21400
rect 12651 20768 12693 20777
rect 12651 20728 12652 20768
rect 12692 20728 12693 20768
rect 12651 20719 12693 20728
rect 12172 20308 12404 20348
rect 12172 19937 12212 20308
rect 12267 20180 12309 20189
rect 12267 20140 12268 20180
rect 12308 20140 12309 20180
rect 12267 20138 12309 20140
rect 12556 20180 12596 20189
rect 12267 20131 12401 20138
rect 12268 20098 12401 20131
rect 12361 20095 12401 20098
rect 12361 20086 12404 20095
rect 12361 20046 12364 20086
rect 12364 20037 12404 20046
rect 12267 20012 12309 20021
rect 12267 19972 12268 20012
rect 12308 19972 12309 20012
rect 12267 19963 12309 19972
rect 12171 19928 12213 19937
rect 12171 19888 12172 19928
rect 12212 19888 12213 19928
rect 12171 19879 12213 19888
rect 12076 18712 12212 18752
rect 12076 18584 12116 18593
rect 11980 18544 12076 18584
rect 11883 15560 11925 15569
rect 11883 15520 11884 15560
rect 11924 15520 11925 15560
rect 11883 15511 11925 15520
rect 11884 15426 11924 15511
rect 11788 15184 11924 15224
rect 11788 14720 11828 14729
rect 11020 12664 11348 12704
rect 11500 14680 11788 14720
rect 10924 12284 10964 12293
rect 10924 12125 10964 12244
rect 10923 12116 10965 12125
rect 10923 12076 10924 12116
rect 10964 12076 10965 12116
rect 10923 12067 10965 12076
rect 10772 11740 10868 11780
rect 10732 11731 10772 11740
rect 10539 11696 10581 11705
rect 10539 11656 10540 11696
rect 10580 11656 10581 11696
rect 10539 11647 10581 11656
rect 10443 11528 10485 11537
rect 10443 11488 10444 11528
rect 10484 11488 10485 11528
rect 10443 11479 10485 11488
rect 10540 11528 10580 11537
rect 10540 11360 10580 11488
rect 10827 11444 10869 11453
rect 10827 11404 10828 11444
rect 10868 11404 10869 11444
rect 10827 11395 10869 11404
rect 10348 11320 10484 11360
rect 10540 11320 10772 11360
rect 10156 11201 10196 11286
rect 10155 11192 10197 11201
rect 10155 11152 10156 11192
rect 10196 11152 10197 11192
rect 10155 11143 10197 11152
rect 10251 11108 10293 11117
rect 10251 11068 10252 11108
rect 10292 11068 10293 11108
rect 10251 11059 10293 11068
rect 10155 11024 10197 11033
rect 10155 10984 10156 11024
rect 10196 10984 10197 11024
rect 10155 10975 10197 10984
rect 10059 10940 10101 10949
rect 10059 10900 10060 10940
rect 10100 10900 10101 10940
rect 10059 10891 10101 10900
rect 9963 10184 10005 10193
rect 9963 10144 9964 10184
rect 10004 10144 10005 10184
rect 9963 10135 10005 10144
rect 9771 9596 9813 9605
rect 9771 9556 9772 9596
rect 9812 9556 9813 9596
rect 9771 9547 9813 9556
rect 9772 8672 9812 9547
rect 9867 9512 9909 9521
rect 9867 9472 9868 9512
rect 9908 9472 9909 9512
rect 9867 9463 9909 9472
rect 9868 9378 9908 9463
rect 10059 8840 10101 8849
rect 10059 8800 10060 8840
rect 10100 8800 10101 8840
rect 10059 8791 10101 8800
rect 9772 8623 9812 8632
rect 9963 8672 10005 8681
rect 9963 8632 9964 8672
rect 10004 8632 10005 8672
rect 9963 8623 10005 8632
rect 10060 8672 10100 8791
rect 10156 8765 10196 10975
rect 10155 8756 10197 8765
rect 10155 8716 10156 8756
rect 10196 8716 10197 8756
rect 10155 8707 10197 8716
rect 10060 8623 10100 8632
rect 10252 8672 10292 11059
rect 10444 11033 10484 11320
rect 10636 11192 10676 11203
rect 10636 11117 10676 11152
rect 10635 11108 10677 11117
rect 10635 11068 10636 11108
rect 10676 11068 10677 11108
rect 10635 11059 10677 11068
rect 10348 11024 10388 11033
rect 10348 10352 10388 10984
rect 10443 11024 10485 11033
rect 10443 10984 10444 11024
rect 10484 10984 10485 11024
rect 10443 10975 10485 10984
rect 10444 10890 10484 10975
rect 10732 10865 10772 11320
rect 10731 10856 10773 10865
rect 10731 10816 10732 10856
rect 10772 10816 10773 10856
rect 10731 10807 10773 10816
rect 10828 10604 10868 11395
rect 10636 10564 10868 10604
rect 10540 10361 10580 10446
rect 10539 10352 10581 10361
rect 10348 10312 10484 10352
rect 10347 10184 10389 10193
rect 10347 10144 10348 10184
rect 10388 10144 10389 10184
rect 10347 10135 10389 10144
rect 10348 10050 10388 10135
rect 10347 9680 10389 9689
rect 10347 9640 10348 9680
rect 10388 9640 10389 9680
rect 10347 9631 10389 9640
rect 10348 9546 10388 9631
rect 10444 9428 10484 10312
rect 10539 10312 10540 10352
rect 10580 10312 10581 10352
rect 10539 10303 10581 10312
rect 10539 10184 10581 10193
rect 10539 10144 10540 10184
rect 10580 10144 10581 10184
rect 10539 10135 10581 10144
rect 10540 9512 10580 10135
rect 10540 9463 10580 9472
rect 10348 9388 10484 9428
rect 10348 9185 10388 9388
rect 10347 9176 10389 9185
rect 10347 9136 10348 9176
rect 10388 9136 10389 9176
rect 10347 9127 10389 9136
rect 10252 8623 10292 8632
rect 10348 8672 10388 9127
rect 10503 8765 10543 8780
rect 10502 8756 10544 8765
rect 10502 8716 10503 8756
rect 10543 8716 10545 8756
rect 10502 8707 10545 8716
rect 10505 8687 10545 8707
rect 10505 8638 10545 8647
rect 10348 8623 10388 8632
rect 9964 8538 10004 8623
rect 10059 8504 10101 8513
rect 10059 8464 10060 8504
rect 10100 8464 10101 8504
rect 10059 8455 10101 8464
rect 10156 8504 10196 8513
rect 10060 8261 10100 8455
rect 10059 8252 10101 8261
rect 10059 8212 10060 8252
rect 10100 8212 10101 8252
rect 10059 8203 10101 8212
rect 9675 7916 9717 7925
rect 9675 7876 9676 7916
rect 9716 7876 9717 7916
rect 9675 7867 9717 7876
rect 9771 7076 9813 7085
rect 9771 7036 9772 7076
rect 9812 7036 9813 7076
rect 9771 7027 9813 7036
rect 9772 5648 9812 7027
rect 10156 5909 10196 8464
rect 10347 8504 10389 8513
rect 10347 8464 10348 8504
rect 10388 8464 10389 8504
rect 10347 8455 10389 8464
rect 10251 7496 10293 7505
rect 10251 7456 10252 7496
rect 10292 7456 10293 7496
rect 10251 7447 10293 7456
rect 10252 6917 10292 7447
rect 10251 6908 10293 6917
rect 10251 6868 10252 6908
rect 10292 6868 10293 6908
rect 10251 6859 10293 6868
rect 10155 5900 10197 5909
rect 10155 5860 10156 5900
rect 10196 5860 10197 5900
rect 10155 5851 10197 5860
rect 9676 5608 9772 5648
rect 9676 4976 9716 5608
rect 9772 5599 9812 5608
rect 9867 5648 9909 5657
rect 9867 5608 9868 5648
rect 9908 5608 9909 5648
rect 9867 5599 9909 5608
rect 10156 5648 10196 5657
rect 9771 5144 9813 5153
rect 9771 5104 9772 5144
rect 9812 5104 9813 5144
rect 9771 5095 9813 5104
rect 9676 4649 9716 4936
rect 9675 4640 9717 4649
rect 9675 4600 9676 4640
rect 9716 4600 9717 4640
rect 9675 4591 9717 4600
rect 9580 4087 9620 4096
rect 9676 3893 9716 4591
rect 9772 4304 9812 5095
rect 9772 4255 9812 4264
rect 9868 5060 9908 5599
rect 9964 5573 10004 5604
rect 9963 5564 10005 5573
rect 9963 5524 9964 5564
rect 10004 5524 10005 5564
rect 9963 5515 10005 5524
rect 9771 4136 9813 4145
rect 9771 4096 9772 4136
rect 9812 4096 9813 4136
rect 9771 4087 9813 4096
rect 9868 4136 9908 5020
rect 9964 5480 10004 5515
rect 9964 4976 10004 5440
rect 10156 5153 10196 5608
rect 10251 5648 10293 5657
rect 10251 5608 10252 5648
rect 10292 5608 10293 5648
rect 10251 5599 10293 5608
rect 10252 5514 10292 5599
rect 10348 5312 10388 8455
rect 10636 8336 10676 10564
rect 10731 10436 10773 10445
rect 10731 10396 10732 10436
rect 10772 10396 10773 10436
rect 10731 10387 10773 10396
rect 10732 10016 10772 10387
rect 10876 10193 10916 10202
rect 10732 9967 10772 9976
rect 10828 10153 10876 10184
rect 10828 10144 10916 10153
rect 10828 9689 10868 10144
rect 10827 9680 10869 9689
rect 10827 9640 10828 9680
rect 10868 9640 10869 9680
rect 10827 9631 10869 9640
rect 10540 8296 10676 8336
rect 10828 8672 10868 8681
rect 10443 8252 10485 8261
rect 10443 8212 10444 8252
rect 10484 8212 10485 8252
rect 10443 8203 10485 8212
rect 10444 8000 10484 8203
rect 10444 7951 10484 7960
rect 10444 7160 10484 7171
rect 10444 7085 10484 7120
rect 10443 7076 10485 7085
rect 10443 7036 10444 7076
rect 10484 7036 10485 7076
rect 10443 7027 10485 7036
rect 10540 5993 10580 8296
rect 10636 8168 10676 8177
rect 10828 8168 10868 8632
rect 10924 8672 10964 8683
rect 10924 8597 10964 8632
rect 10923 8588 10965 8597
rect 10923 8548 10924 8588
rect 10964 8548 10965 8588
rect 10923 8539 10965 8548
rect 10923 8336 10965 8345
rect 10923 8296 10924 8336
rect 10964 8296 10965 8336
rect 10923 8287 10965 8296
rect 10676 8128 10868 8168
rect 10636 8119 10676 8128
rect 10924 7925 10964 8287
rect 11020 8177 11060 12664
rect 11212 12536 11252 12545
rect 11212 12125 11252 12496
rect 11308 12536 11348 12545
rect 11211 12116 11253 12125
rect 11211 12076 11212 12116
rect 11252 12076 11253 12116
rect 11211 12067 11253 12076
rect 11211 11864 11253 11873
rect 11211 11824 11212 11864
rect 11252 11824 11253 11864
rect 11211 11815 11253 11824
rect 11212 11696 11252 11815
rect 11212 11369 11252 11656
rect 11308 11453 11348 12496
rect 11307 11444 11349 11453
rect 11307 11404 11308 11444
rect 11348 11404 11349 11444
rect 11307 11395 11349 11404
rect 11211 11360 11253 11369
rect 11211 11320 11212 11360
rect 11252 11320 11253 11360
rect 11211 11311 11253 11320
rect 11115 10184 11157 10193
rect 11115 10144 11116 10184
rect 11156 10144 11157 10184
rect 11115 10135 11157 10144
rect 11019 8168 11061 8177
rect 11019 8128 11020 8168
rect 11060 8128 11061 8168
rect 11019 8119 11061 8128
rect 11020 8000 11060 8009
rect 10923 7916 10965 7925
rect 11020 7916 11060 7960
rect 10923 7876 10924 7916
rect 10964 7876 11060 7916
rect 10923 7867 10965 7876
rect 11116 7832 11156 10135
rect 11308 10109 11348 11395
rect 11500 11285 11540 14680
rect 11788 14671 11828 14680
rect 11691 14552 11733 14561
rect 11691 14512 11692 14552
rect 11732 14512 11733 14552
rect 11691 14503 11733 14512
rect 11692 12452 11732 14503
rect 11884 14048 11924 15184
rect 11692 11369 11732 12412
rect 11788 12452 11828 12461
rect 11691 11360 11733 11369
rect 11691 11320 11692 11360
rect 11732 11320 11733 11360
rect 11691 11311 11733 11320
rect 11499 11276 11541 11285
rect 11499 11236 11500 11276
rect 11540 11236 11541 11276
rect 11499 11227 11541 11236
rect 11691 11192 11733 11201
rect 11691 11152 11692 11192
rect 11732 11152 11733 11192
rect 11691 11143 11733 11152
rect 11499 11108 11541 11117
rect 11499 11068 11500 11108
rect 11540 11068 11541 11108
rect 11499 11059 11541 11068
rect 11403 11024 11445 11033
rect 11403 10984 11404 11024
rect 11444 10984 11445 11024
rect 11403 10975 11445 10984
rect 11404 10193 11444 10975
rect 11403 10184 11445 10193
rect 11403 10144 11404 10184
rect 11444 10144 11445 10184
rect 11403 10135 11445 10144
rect 11307 10100 11349 10109
rect 11307 10060 11308 10100
rect 11348 10060 11349 10100
rect 11307 10051 11349 10060
rect 11211 8756 11253 8765
rect 11211 8716 11212 8756
rect 11252 8716 11253 8756
rect 11211 8707 11253 8716
rect 11020 7792 11156 7832
rect 11020 7505 11060 7792
rect 11115 7580 11157 7589
rect 11115 7540 11116 7580
rect 11156 7540 11157 7580
rect 11115 7531 11157 7540
rect 11019 7496 11061 7505
rect 11019 7456 11020 7496
rect 11060 7456 11061 7496
rect 11019 7447 11061 7456
rect 11116 7412 11156 7531
rect 11116 7372 11163 7412
rect 10636 7328 10676 7337
rect 10676 7288 10875 7328
rect 10636 6908 10676 7288
rect 10835 7165 10875 7288
rect 11123 7165 11163 7372
rect 11212 7337 11252 8707
rect 11308 8672 11348 10051
rect 11404 10050 11444 10135
rect 11308 7505 11348 8632
rect 11404 8672 11444 8681
rect 11500 8672 11540 11059
rect 11444 8632 11540 8672
rect 11692 11024 11732 11143
rect 11404 8177 11444 8632
rect 11403 8168 11445 8177
rect 11403 8128 11404 8168
rect 11444 8128 11445 8168
rect 11403 8119 11445 8128
rect 11296 7496 11348 7505
rect 11296 7456 11297 7496
rect 11337 7456 11348 7496
rect 11296 7447 11338 7456
rect 11211 7328 11253 7337
rect 11211 7288 11212 7328
rect 11252 7288 11253 7328
rect 11211 7279 11253 7288
rect 11403 7328 11445 7337
rect 11403 7288 11404 7328
rect 11444 7288 11445 7328
rect 11403 7279 11445 7288
rect 10835 7116 10875 7125
rect 10931 7156 10971 7165
rect 11123 7116 11163 7125
rect 10931 7085 10971 7116
rect 10923 7076 10971 7085
rect 10923 7036 10924 7076
rect 10964 7036 10971 7076
rect 11211 7076 11253 7085
rect 11211 7036 11212 7076
rect 11252 7036 11253 7076
rect 10923 7027 10965 7036
rect 11211 7027 11253 7036
rect 11020 6992 11060 7001
rect 11020 6908 11060 6952
rect 10636 6868 10772 6908
rect 10635 6740 10677 6749
rect 10635 6700 10636 6740
rect 10676 6700 10677 6740
rect 10635 6691 10677 6700
rect 10636 6488 10676 6691
rect 10732 6497 10772 6868
rect 10924 6868 11060 6908
rect 10924 6740 10964 6868
rect 10828 6700 10964 6740
rect 10636 6439 10676 6448
rect 10731 6488 10773 6497
rect 10731 6448 10732 6488
rect 10772 6448 10773 6488
rect 10731 6439 10773 6448
rect 10828 6488 10868 6700
rect 11115 6656 11157 6665
rect 11115 6616 11116 6656
rect 11156 6616 11157 6656
rect 11115 6607 11157 6616
rect 10828 6439 10868 6448
rect 10923 6488 10965 6497
rect 10923 6448 10924 6488
rect 10964 6448 10965 6488
rect 10923 6439 10965 6448
rect 11116 6488 11156 6607
rect 11212 6581 11252 7027
rect 11211 6572 11253 6581
rect 11404 6572 11444 7279
rect 11499 7244 11541 7253
rect 11499 7204 11500 7244
rect 11540 7204 11541 7244
rect 11499 7195 11541 7204
rect 11500 7160 11540 7195
rect 11500 7109 11540 7120
rect 11692 7085 11732 10984
rect 11788 10436 11828 12412
rect 11884 10613 11924 14008
rect 11980 10697 12020 18544
rect 12076 18535 12116 18544
rect 12172 17753 12212 18712
rect 12171 17744 12213 17753
rect 12171 17704 12172 17744
rect 12212 17704 12213 17744
rect 12171 17695 12213 17704
rect 12268 15821 12308 19963
rect 12363 19928 12405 19937
rect 12363 19888 12364 19928
rect 12404 19888 12405 19928
rect 12363 19879 12405 19888
rect 12364 16829 12404 19879
rect 12556 19853 12596 20140
rect 12651 20180 12693 20189
rect 12651 20140 12652 20180
rect 12692 20140 12693 20180
rect 12651 20131 12693 20140
rect 12555 19844 12597 19853
rect 12555 19804 12556 19844
rect 12596 19804 12597 19844
rect 12555 19795 12597 19804
rect 12652 19508 12692 20131
rect 12652 19459 12692 19468
rect 12748 20096 12788 20105
rect 12460 19256 12500 19265
rect 12460 19013 12500 19216
rect 12555 19172 12597 19181
rect 12555 19132 12556 19172
rect 12596 19132 12597 19172
rect 12555 19123 12597 19132
rect 12459 19004 12501 19013
rect 12459 18964 12460 19004
rect 12500 18964 12501 19004
rect 12459 18955 12501 18964
rect 12556 18668 12596 19123
rect 12748 18929 12788 20056
rect 12747 18920 12789 18929
rect 12747 18880 12748 18920
rect 12788 18880 12789 18920
rect 12747 18871 12789 18880
rect 12651 18836 12693 18845
rect 12651 18796 12652 18836
rect 12692 18796 12693 18836
rect 12651 18787 12693 18796
rect 12460 18628 12596 18668
rect 12363 16820 12405 16829
rect 12363 16780 12364 16820
rect 12404 16780 12405 16820
rect 12363 16771 12405 16780
rect 12460 16232 12500 18628
rect 12556 18570 12596 18579
rect 12556 18005 12596 18530
rect 12652 18089 12692 18787
rect 12747 18668 12789 18677
rect 12747 18628 12748 18668
rect 12788 18628 12789 18668
rect 12747 18619 12789 18628
rect 12748 18534 12788 18619
rect 12747 18164 12789 18173
rect 12747 18124 12748 18164
rect 12788 18124 12789 18164
rect 12747 18115 12789 18124
rect 12651 18080 12693 18089
rect 12651 18040 12652 18080
rect 12692 18040 12693 18080
rect 12651 18031 12693 18040
rect 12555 17996 12597 18005
rect 12555 17956 12556 17996
rect 12596 17956 12597 17996
rect 12555 17947 12597 17956
rect 12500 16192 12596 16232
rect 12460 16183 12500 16192
rect 12267 15812 12309 15821
rect 12267 15772 12268 15812
rect 12308 15772 12309 15812
rect 12267 15763 12309 15772
rect 12076 15644 12116 15653
rect 12116 15604 12404 15644
rect 12076 15595 12116 15604
rect 12364 15560 12404 15604
rect 12364 15511 12404 15520
rect 12460 15560 12500 15569
rect 12075 15476 12117 15485
rect 12075 15436 12076 15476
rect 12116 15436 12117 15476
rect 12075 15427 12117 15436
rect 12076 10781 12116 15427
rect 12460 15392 12500 15520
rect 12172 15352 12500 15392
rect 12172 14813 12212 15352
rect 12171 14804 12213 14813
rect 12171 14764 12172 14804
rect 12212 14764 12213 14804
rect 12171 14755 12213 14764
rect 12075 10772 12117 10781
rect 12075 10732 12076 10772
rect 12116 10732 12117 10772
rect 12075 10723 12117 10732
rect 11979 10688 12021 10697
rect 11979 10648 11980 10688
rect 12020 10648 12021 10688
rect 11979 10639 12021 10648
rect 11883 10604 11925 10613
rect 11883 10564 11884 10604
rect 11924 10564 11925 10604
rect 11883 10555 11925 10564
rect 11980 10529 12020 10639
rect 12075 10604 12117 10613
rect 12075 10564 12076 10604
rect 12116 10564 12117 10604
rect 12075 10555 12117 10564
rect 11979 10520 12021 10529
rect 11979 10480 11980 10520
rect 12020 10480 12021 10520
rect 11979 10471 12021 10480
rect 11883 10436 11925 10445
rect 11788 10396 11884 10436
rect 11924 10396 11925 10436
rect 11883 10387 11925 10396
rect 11884 10268 11924 10387
rect 11884 10219 11924 10228
rect 11979 10184 12021 10193
rect 11979 10144 11980 10184
rect 12020 10144 12021 10184
rect 11979 10135 12021 10144
rect 11980 10050 12020 10135
rect 11787 9596 11829 9605
rect 11787 9556 11788 9596
rect 11828 9556 11829 9596
rect 11787 9547 11829 9556
rect 11788 9512 11828 9547
rect 11788 9428 11828 9472
rect 11980 9470 12020 9479
rect 11980 9428 12020 9430
rect 11788 9388 12020 9428
rect 11787 8840 11829 8849
rect 12076 8840 12116 10555
rect 11787 8800 11788 8840
rect 11828 8800 11829 8840
rect 11787 8791 11829 8800
rect 11980 8800 12116 8840
rect 11691 7076 11733 7085
rect 11691 7036 11692 7076
rect 11732 7036 11733 7076
rect 11691 7027 11733 7036
rect 11788 6665 11828 8791
rect 11884 8672 11924 8681
rect 11884 8513 11924 8632
rect 11883 8504 11925 8513
rect 11883 8464 11884 8504
rect 11924 8464 11925 8504
rect 11883 8455 11925 8464
rect 11884 8093 11924 8455
rect 11883 8084 11925 8093
rect 11883 8044 11884 8084
rect 11924 8044 11925 8084
rect 11883 8035 11925 8044
rect 11692 6656 11732 6665
rect 11211 6532 11212 6572
rect 11252 6532 11253 6572
rect 11211 6523 11253 6532
rect 11369 6532 11444 6572
rect 11500 6616 11692 6656
rect 11116 6439 11156 6448
rect 11212 6488 11252 6523
rect 10924 6354 10964 6439
rect 11212 6438 11252 6448
rect 11369 6481 11409 6532
rect 11369 6413 11409 6441
rect 11355 6404 11409 6413
rect 11355 6364 11356 6404
rect 11396 6364 11409 6404
rect 11355 6355 11409 6364
rect 11369 6346 11409 6355
rect 10731 6320 10773 6329
rect 10731 6280 10732 6320
rect 10772 6280 10773 6320
rect 10731 6271 10773 6280
rect 11019 6320 11061 6329
rect 11019 6280 11020 6320
rect 11060 6280 11061 6320
rect 11019 6271 11061 6280
rect 11211 6320 11253 6329
rect 11211 6280 11212 6320
rect 11252 6280 11253 6320
rect 11211 6271 11253 6280
rect 10539 5984 10581 5993
rect 10732 5984 10772 6271
rect 10828 6236 10868 6245
rect 10868 6196 10964 6236
rect 10828 6187 10868 6196
rect 10539 5944 10540 5984
rect 10580 5944 10581 5984
rect 10539 5935 10581 5944
rect 10697 5944 10772 5984
rect 10697 5663 10737 5944
rect 10252 5272 10388 5312
rect 10444 5648 10484 5657
rect 10155 5144 10197 5153
rect 10155 5104 10156 5144
rect 10196 5104 10197 5144
rect 10155 5095 10197 5104
rect 10060 4976 10100 4985
rect 9964 4936 10060 4976
rect 10060 4145 10100 4936
rect 10156 4976 10196 4985
rect 10156 4817 10196 4936
rect 10155 4808 10197 4817
rect 10155 4768 10156 4808
rect 10196 4768 10197 4808
rect 10155 4759 10197 4768
rect 9868 4087 9908 4096
rect 10059 4136 10101 4145
rect 10059 4096 10060 4136
rect 10100 4096 10101 4136
rect 10059 4087 10101 4096
rect 9772 4002 9812 4087
rect 10155 3968 10197 3977
rect 10155 3928 10156 3968
rect 10196 3928 10197 3968
rect 10155 3919 10197 3928
rect 9675 3884 9717 3893
rect 9675 3844 9676 3884
rect 9716 3844 9717 3884
rect 9675 3835 9717 3844
rect 10156 3834 10196 3919
rect 10252 3632 10292 5272
rect 10348 5144 10388 5153
rect 10444 5144 10484 5608
rect 10540 5648 10580 5659
rect 10697 5614 10737 5623
rect 10540 5573 10580 5608
rect 10539 5564 10581 5573
rect 10539 5524 10540 5564
rect 10580 5524 10581 5564
rect 10539 5515 10581 5524
rect 10636 5480 10676 5489
rect 10636 5144 10676 5440
rect 10827 5396 10869 5405
rect 10827 5356 10828 5396
rect 10868 5356 10869 5396
rect 10827 5347 10869 5356
rect 10388 5104 10484 5144
rect 10540 5104 10676 5144
rect 10348 5095 10388 5104
rect 10156 3592 10292 3632
rect 10348 4136 10388 4145
rect 9868 3464 9908 3473
rect 9908 3424 10004 3464
rect 9868 3415 9908 3424
rect 9867 3212 9909 3221
rect 9867 3172 9868 3212
rect 9908 3172 9909 3212
rect 9867 3163 9909 3172
rect 9580 2792 9620 2801
rect 9868 2792 9908 3163
rect 9964 2801 10004 3424
rect 10156 3305 10196 3592
rect 10252 3464 10292 3473
rect 10348 3464 10388 4096
rect 10443 4136 10485 4145
rect 10443 4096 10444 4136
rect 10484 4096 10485 4136
rect 10443 4087 10485 4096
rect 10444 4002 10484 4087
rect 10540 3632 10580 5104
rect 10636 4976 10676 4985
rect 10828 4976 10868 5347
rect 10676 4936 10868 4976
rect 10636 4927 10676 4936
rect 10635 4136 10677 4145
rect 10635 4096 10636 4136
rect 10676 4096 10677 4136
rect 10635 4087 10677 4096
rect 10732 4136 10772 4145
rect 10292 3424 10388 3464
rect 10252 3415 10292 3424
rect 10155 3296 10197 3305
rect 10155 3256 10156 3296
rect 10196 3256 10197 3296
rect 10155 3247 10197 3256
rect 10060 3212 10100 3221
rect 9620 2752 9908 2792
rect 9580 2381 9620 2752
rect 9868 2624 9908 2752
rect 9963 2792 10005 2801
rect 9963 2752 9964 2792
rect 10004 2752 10005 2792
rect 9963 2743 10005 2752
rect 10060 2633 10100 3172
rect 10155 3044 10197 3053
rect 10155 3004 10156 3044
rect 10196 3004 10197 3044
rect 10155 2995 10197 3004
rect 9868 2575 9908 2584
rect 10059 2624 10101 2633
rect 10059 2584 10060 2624
rect 10100 2584 10101 2624
rect 10059 2575 10101 2584
rect 10156 2624 10196 2995
rect 10156 2575 10196 2584
rect 10252 2540 10292 2580
rect 10252 2456 10292 2500
rect 10060 2416 10292 2456
rect 9579 2372 9621 2381
rect 9579 2332 9580 2372
rect 9620 2332 9621 2372
rect 9579 2323 9621 2332
rect 9484 2164 9620 2204
rect 9388 1903 9428 1912
rect 9484 1952 9524 1961
rect 9484 1709 9524 1912
rect 9483 1700 9525 1709
rect 9483 1660 9484 1700
rect 9524 1660 9525 1700
rect 9483 1651 9525 1660
rect 9483 1532 9525 1541
rect 9483 1492 9484 1532
rect 9524 1492 9525 1532
rect 9483 1483 9525 1492
rect 9388 1196 9428 1205
rect 9292 1156 9388 1196
rect 9388 1147 9428 1156
rect 9196 1072 9332 1112
rect 9195 944 9237 953
rect 9195 904 9196 944
rect 9236 904 9237 944
rect 9195 895 9237 904
rect 9196 810 9236 895
rect 9099 776 9141 785
rect 9099 736 9100 776
rect 9140 736 9141 776
rect 9099 727 9141 736
rect 9099 608 9141 617
rect 9099 568 9100 608
rect 9140 568 9141 608
rect 9099 559 9141 568
rect 8907 356 8949 365
rect 8907 316 8908 356
rect 8948 316 8949 356
rect 8907 307 8949 316
rect 8908 80 8948 307
rect 9100 80 9140 559
rect 9292 80 9332 1072
rect 9484 80 9524 1483
rect 9580 1196 9620 2164
rect 9676 2120 9716 2129
rect 9716 2080 10004 2120
rect 9676 2071 9716 2080
rect 9867 1952 9909 1961
rect 9867 1912 9868 1952
rect 9908 1912 9909 1952
rect 9867 1903 9909 1912
rect 9964 1952 10004 2080
rect 10060 2045 10100 2416
rect 10156 2120 10196 2129
rect 10348 2120 10388 3424
rect 10444 3592 10580 3632
rect 10444 2717 10484 3592
rect 10540 3464 10580 3473
rect 10636 3464 10676 4087
rect 10732 3641 10772 4096
rect 10731 3632 10773 3641
rect 10731 3592 10732 3632
rect 10772 3592 10773 3632
rect 10731 3583 10773 3592
rect 10828 3557 10868 4936
rect 10924 4397 10964 6196
rect 10923 4388 10965 4397
rect 10923 4348 10924 4388
rect 10964 4348 10965 4388
rect 10923 4339 10965 4348
rect 10827 3548 10869 3557
rect 10827 3508 10828 3548
rect 10868 3508 10869 3548
rect 10827 3499 10869 3508
rect 10580 3424 10676 3464
rect 10540 3415 10580 3424
rect 10539 3296 10581 3305
rect 10539 3256 10540 3296
rect 10580 3256 10581 3296
rect 10539 3247 10581 3256
rect 10540 3162 10580 3247
rect 10636 3044 10676 3424
rect 10732 3464 10772 3473
rect 10732 3221 10772 3424
rect 10923 3464 10965 3473
rect 10923 3424 10924 3464
rect 10964 3424 10965 3464
rect 10923 3415 10965 3424
rect 10924 3330 10964 3415
rect 10827 3296 10869 3305
rect 10827 3256 10828 3296
rect 10868 3256 10869 3296
rect 10827 3247 10869 3256
rect 10731 3212 10773 3221
rect 10731 3172 10732 3212
rect 10772 3172 10773 3212
rect 10731 3163 10773 3172
rect 10828 3162 10868 3247
rect 10636 3004 10868 3044
rect 10540 2792 10580 2801
rect 10580 2752 10772 2792
rect 10540 2743 10580 2752
rect 10443 2708 10485 2717
rect 10443 2668 10444 2708
rect 10484 2668 10485 2708
rect 10443 2659 10485 2668
rect 10732 2624 10772 2752
rect 10828 2708 10868 3004
rect 10924 2717 10964 2732
rect 10828 2659 10868 2668
rect 10923 2708 10965 2717
rect 10923 2668 10924 2708
rect 10964 2668 10965 2708
rect 10923 2659 10965 2668
rect 10924 2637 10964 2659
rect 10924 2588 10964 2597
rect 10732 2575 10772 2584
rect 10443 2540 10485 2549
rect 11020 2540 11060 6271
rect 11212 4817 11252 6271
rect 11307 5984 11349 5993
rect 11307 5944 11308 5984
rect 11348 5944 11349 5984
rect 11307 5935 11349 5944
rect 11308 5648 11348 5935
rect 11308 5599 11348 5608
rect 11211 4808 11253 4817
rect 11211 4768 11212 4808
rect 11252 4768 11253 4808
rect 11211 4759 11253 4768
rect 11500 4229 11540 6616
rect 11692 6607 11732 6616
rect 11787 6656 11829 6665
rect 11787 6616 11788 6656
rect 11828 6616 11829 6656
rect 11787 6607 11829 6616
rect 11630 6473 11670 6499
rect 11630 6413 11670 6433
rect 11788 6488 11828 6497
rect 11629 6404 11671 6413
rect 11629 6364 11630 6404
rect 11670 6364 11671 6404
rect 11629 6355 11671 6364
rect 11691 6236 11733 6245
rect 11691 6196 11692 6236
rect 11732 6196 11733 6236
rect 11691 6187 11733 6196
rect 11595 6152 11637 6161
rect 11595 6112 11596 6152
rect 11636 6112 11637 6152
rect 11595 6103 11637 6112
rect 11596 4313 11636 6103
rect 11595 4304 11637 4313
rect 11595 4264 11596 4304
rect 11636 4264 11637 4304
rect 11595 4255 11637 4264
rect 11499 4220 11541 4229
rect 11499 4180 11500 4220
rect 11540 4180 11541 4220
rect 11499 4171 11541 4180
rect 11211 3632 11253 3641
rect 11211 3592 11212 3632
rect 11252 3592 11348 3632
rect 11116 3557 11156 3588
rect 11211 3583 11253 3592
rect 11115 3548 11157 3557
rect 11115 3508 11116 3548
rect 11156 3508 11157 3548
rect 11115 3499 11157 3508
rect 11116 3464 11156 3499
rect 11116 3221 11156 3424
rect 11211 3296 11253 3305
rect 11211 3256 11212 3296
rect 11252 3256 11253 3296
rect 11211 3247 11253 3256
rect 11115 3212 11157 3221
rect 11115 3172 11116 3212
rect 11156 3172 11157 3212
rect 11115 3163 11157 3172
rect 10443 2500 10444 2540
rect 10484 2500 10485 2540
rect 10443 2491 10485 2500
rect 10828 2500 11060 2540
rect 10196 2080 10388 2120
rect 10156 2071 10196 2080
rect 10059 2036 10101 2045
rect 10059 1996 10060 2036
rect 10100 1996 10101 2036
rect 10059 1987 10101 1996
rect 9964 1903 10004 1912
rect 10156 1952 10196 1961
rect 10444 1952 10484 2491
rect 10539 2036 10581 2045
rect 10539 1996 10540 2036
rect 10580 1996 10581 2036
rect 10539 1987 10581 1996
rect 10196 1912 10484 1952
rect 10156 1903 10196 1912
rect 9868 1818 9908 1903
rect 10540 1868 10580 1987
rect 10540 1819 10580 1828
rect 10732 1700 10772 1709
rect 10539 1616 10581 1625
rect 10539 1576 10540 1616
rect 10580 1576 10581 1616
rect 10539 1567 10581 1576
rect 9867 1532 9909 1541
rect 9867 1492 9868 1532
rect 9908 1492 9909 1532
rect 9867 1483 9909 1492
rect 9772 1196 9812 1205
rect 9580 1156 9772 1196
rect 9772 1147 9812 1156
rect 9580 944 9620 953
rect 9620 904 9716 944
rect 9580 895 9620 904
rect 9676 80 9716 904
rect 9868 80 9908 1483
rect 10155 1196 10197 1205
rect 10155 1156 10156 1196
rect 10196 1156 10197 1196
rect 10155 1147 10197 1156
rect 10540 1196 10580 1567
rect 10732 1457 10772 1660
rect 10731 1448 10773 1457
rect 10731 1408 10732 1448
rect 10772 1408 10773 1448
rect 10731 1399 10773 1408
rect 10635 1364 10677 1373
rect 10635 1324 10636 1364
rect 10676 1324 10677 1364
rect 10635 1315 10677 1324
rect 10540 1147 10580 1156
rect 10156 1062 10196 1147
rect 9964 944 10004 953
rect 9964 449 10004 904
rect 10059 944 10101 953
rect 10059 904 10060 944
rect 10100 904 10101 944
rect 10059 895 10101 904
rect 10348 944 10388 953
rect 10388 904 10484 944
rect 10348 895 10388 904
rect 9963 440 10005 449
rect 9963 400 9964 440
rect 10004 400 10005 440
rect 9963 391 10005 400
rect 10060 80 10100 895
rect 10251 860 10293 869
rect 10251 820 10252 860
rect 10292 820 10293 860
rect 10251 811 10293 820
rect 10252 80 10292 811
rect 10444 80 10484 904
rect 10636 80 10676 1315
rect 10828 1205 10868 2500
rect 11116 2456 11156 2465
rect 11020 2416 11116 2456
rect 10923 2120 10965 2129
rect 10923 2080 10924 2120
rect 10964 2080 10965 2120
rect 10923 2071 10965 2080
rect 10924 1868 10964 2071
rect 10924 1819 10964 1828
rect 10923 1700 10965 1709
rect 10923 1660 10924 1700
rect 10964 1660 10965 1700
rect 10923 1651 10965 1660
rect 10827 1196 10869 1205
rect 10827 1156 10828 1196
rect 10868 1156 10869 1196
rect 10827 1147 10869 1156
rect 10924 1196 10964 1651
rect 10924 1147 10964 1156
rect 10732 944 10772 953
rect 10732 533 10772 904
rect 10731 524 10773 533
rect 10731 484 10732 524
rect 10772 484 10773 524
rect 10731 475 10773 484
rect 10827 440 10869 449
rect 10827 400 10828 440
rect 10868 400 10869 440
rect 10827 391 10869 400
rect 10828 80 10868 391
rect 11020 80 11060 2416
rect 11116 2407 11156 2416
rect 11212 1961 11252 3247
rect 11308 3137 11348 3592
rect 11307 3128 11349 3137
rect 11307 3088 11308 3128
rect 11348 3088 11349 3128
rect 11307 3079 11349 3088
rect 11307 2708 11349 2717
rect 11307 2668 11308 2708
rect 11348 2668 11349 2708
rect 11307 2659 11349 2668
rect 11308 2574 11348 2659
rect 11692 2540 11732 6187
rect 11788 5069 11828 6448
rect 11884 6488 11924 6497
rect 11884 5153 11924 6448
rect 11980 5405 12020 8800
rect 12172 6908 12212 14755
rect 12267 13376 12309 13385
rect 12267 13336 12268 13376
rect 12308 13336 12309 13376
rect 12267 13327 12309 13336
rect 12268 12536 12308 13327
rect 12268 12487 12308 12496
rect 12459 11696 12501 11705
rect 12459 11656 12460 11696
rect 12500 11656 12501 11696
rect 12459 11647 12501 11656
rect 12460 11562 12500 11647
rect 12556 11360 12596 16192
rect 12652 15317 12692 18031
rect 12748 17837 12788 18115
rect 12747 17828 12789 17837
rect 12747 17788 12748 17828
rect 12788 17788 12789 17828
rect 12747 17779 12789 17788
rect 12748 17744 12788 17779
rect 12748 17694 12788 17704
rect 12844 17660 12884 21391
rect 13035 18752 13077 18761
rect 13035 18712 13036 18752
rect 13076 18712 13077 18752
rect 13035 18703 13077 18712
rect 12939 17996 12981 18005
rect 12939 17956 12940 17996
rect 12980 17956 12981 17996
rect 12939 17947 12981 17956
rect 12940 17862 12980 17947
rect 12844 17620 12980 17660
rect 12748 17072 12788 17081
rect 12748 16745 12788 17032
rect 12747 16736 12789 16745
rect 12747 16696 12748 16736
rect 12788 16696 12789 16736
rect 12747 16687 12789 16696
rect 12747 15560 12789 15569
rect 12747 15520 12748 15560
rect 12788 15520 12789 15560
rect 12747 15511 12789 15520
rect 12651 15308 12693 15317
rect 12651 15268 12652 15308
rect 12692 15268 12693 15308
rect 12651 15259 12693 15268
rect 12652 12293 12692 15259
rect 12748 14729 12788 15511
rect 12844 15485 12884 15570
rect 12843 15476 12885 15485
rect 12843 15436 12844 15476
rect 12884 15436 12885 15476
rect 12843 15427 12885 15436
rect 12940 15476 12980 17620
rect 13036 16064 13076 18703
rect 13132 17585 13172 21895
rect 13420 21617 13460 22408
rect 13516 21953 13556 23575
rect 13612 23297 13652 23752
rect 13611 23288 13653 23297
rect 13611 23248 13612 23288
rect 13652 23248 13653 23288
rect 13611 23239 13653 23248
rect 13611 23120 13653 23129
rect 13611 23080 13612 23120
rect 13652 23080 13653 23120
rect 13611 23071 13653 23080
rect 13515 21944 13557 21953
rect 13515 21904 13516 21944
rect 13556 21904 13557 21944
rect 13515 21895 13557 21904
rect 13612 21776 13652 23071
rect 13708 22877 13748 24079
rect 13707 22868 13749 22877
rect 13707 22828 13708 22868
rect 13748 22828 13749 22868
rect 13707 22819 13749 22828
rect 13707 22280 13749 22289
rect 13707 22240 13708 22280
rect 13748 22240 13749 22280
rect 13707 22231 13749 22240
rect 13708 22146 13748 22231
rect 13612 21736 13748 21776
rect 13227 21608 13269 21617
rect 13419 21608 13461 21617
rect 13227 21568 13228 21608
rect 13268 21568 13269 21608
rect 13227 21559 13269 21568
rect 13324 21568 13420 21608
rect 13460 21568 13461 21608
rect 13228 17660 13268 21559
rect 13324 19349 13364 21568
rect 13419 21559 13461 21568
rect 13516 21608 13556 21617
rect 13419 21440 13461 21449
rect 13419 21400 13420 21440
rect 13460 21400 13461 21440
rect 13419 21391 13461 21400
rect 13323 19340 13365 19349
rect 13323 19300 13324 19340
rect 13364 19300 13365 19340
rect 13323 19291 13365 19300
rect 13228 17620 13364 17660
rect 13131 17576 13173 17585
rect 13131 17536 13132 17576
rect 13172 17536 13173 17576
rect 13131 17527 13173 17536
rect 13036 16024 13268 16064
rect 13131 15896 13173 15905
rect 13131 15856 13132 15896
rect 13172 15856 13173 15896
rect 13131 15847 13173 15856
rect 12843 14888 12885 14897
rect 12843 14848 12844 14888
rect 12884 14848 12885 14888
rect 12843 14839 12885 14848
rect 12747 14720 12789 14729
rect 12747 14680 12748 14720
rect 12788 14680 12789 14720
rect 12747 14671 12789 14680
rect 12748 12522 12788 12531
rect 12651 12284 12693 12293
rect 12651 12244 12652 12284
rect 12692 12244 12693 12284
rect 12651 12235 12693 12244
rect 12652 11948 12692 11957
rect 12748 11948 12788 12482
rect 12692 11908 12788 11948
rect 12652 11899 12692 11908
rect 12268 11320 12596 11360
rect 12268 8168 12308 11320
rect 12555 10772 12597 10781
rect 12555 10732 12556 10772
rect 12596 10732 12597 10772
rect 12555 10723 12597 10732
rect 12459 10352 12501 10361
rect 12459 10312 12460 10352
rect 12500 10312 12501 10352
rect 12459 10303 12501 10312
rect 12363 10184 12405 10193
rect 12363 10144 12364 10184
rect 12404 10144 12405 10184
rect 12363 10135 12405 10144
rect 12460 10184 12500 10303
rect 12460 10135 12500 10144
rect 12364 10050 12404 10135
rect 12556 10016 12596 10723
rect 12747 10604 12789 10613
rect 12747 10564 12748 10604
rect 12788 10564 12789 10604
rect 12747 10555 12789 10564
rect 12651 10184 12693 10193
rect 12651 10144 12652 10184
rect 12692 10144 12693 10184
rect 12651 10135 12693 10144
rect 12460 9976 12596 10016
rect 12460 8849 12500 9976
rect 12555 9008 12597 9017
rect 12555 8968 12556 9008
rect 12596 8968 12597 9008
rect 12555 8959 12597 8968
rect 12459 8840 12501 8849
rect 12459 8800 12460 8840
rect 12500 8800 12501 8840
rect 12459 8791 12501 8800
rect 12412 8681 12452 8690
rect 12452 8641 12500 8672
rect 12412 8632 12500 8641
rect 12460 8168 12500 8632
rect 12556 8588 12596 8959
rect 12556 8539 12596 8548
rect 12555 8252 12597 8261
rect 12555 8212 12556 8252
rect 12596 8212 12597 8252
rect 12555 8203 12597 8212
rect 12268 8128 12404 8168
rect 12268 8000 12308 8011
rect 12268 7925 12308 7960
rect 12267 7916 12309 7925
rect 12267 7876 12268 7916
rect 12308 7876 12309 7916
rect 12267 7867 12309 7876
rect 12364 7076 12404 8128
rect 12460 8119 12500 8128
rect 12556 7925 12596 8203
rect 12652 8009 12692 10135
rect 12748 8681 12788 10555
rect 12844 8765 12884 14839
rect 12940 14561 12980 15436
rect 13035 14720 13077 14729
rect 13035 14680 13036 14720
rect 13076 14680 13077 14720
rect 13035 14671 13077 14680
rect 12939 14552 12981 14561
rect 12939 14512 12940 14552
rect 12980 14512 12981 14552
rect 12939 14503 12981 14512
rect 13036 14048 13076 14671
rect 13132 14468 13172 15847
rect 13228 14897 13268 16024
rect 13227 14888 13269 14897
rect 13227 14848 13228 14888
rect 13268 14848 13269 14888
rect 13227 14839 13269 14848
rect 13324 14720 13364 17620
rect 13420 15905 13460 21391
rect 13516 21020 13556 21568
rect 13611 21608 13653 21617
rect 13611 21568 13612 21608
rect 13652 21568 13653 21608
rect 13611 21559 13653 21568
rect 13612 21474 13652 21559
rect 13708 21449 13748 21736
rect 13707 21440 13749 21449
rect 13707 21400 13708 21440
rect 13748 21400 13749 21440
rect 13707 21391 13749 21400
rect 13708 21020 13748 21029
rect 13516 20980 13708 21020
rect 13708 20971 13748 20980
rect 13515 20768 13557 20777
rect 13515 20728 13516 20768
rect 13556 20728 13748 20768
rect 13515 20719 13557 20728
rect 13516 20634 13556 20719
rect 13612 19349 13652 19380
rect 13611 19340 13653 19349
rect 13611 19300 13612 19340
rect 13652 19300 13653 19340
rect 13611 19291 13653 19300
rect 13515 19256 13557 19265
rect 13515 19216 13516 19256
rect 13556 19216 13557 19256
rect 13515 19207 13557 19216
rect 13612 19256 13652 19291
rect 13516 19122 13556 19207
rect 13516 17753 13556 17838
rect 13515 17744 13557 17753
rect 13515 17704 13516 17744
rect 13556 17704 13557 17744
rect 13515 17695 13557 17704
rect 13612 17576 13652 19216
rect 13708 19013 13748 20728
rect 13707 19004 13749 19013
rect 13707 18964 13708 19004
rect 13748 18964 13749 19004
rect 13707 18955 13749 18964
rect 13804 18761 13844 28960
rect 13900 23120 13940 29791
rect 14092 29000 14132 32824
rect 14379 32192 14421 32201
rect 14379 32152 14380 32192
rect 14420 32152 14421 32192
rect 14379 32143 14421 32152
rect 14476 32192 14516 32201
rect 14380 32058 14420 32143
rect 14187 31772 14229 31781
rect 14187 31732 14188 31772
rect 14228 31732 14229 31772
rect 14187 31723 14229 31732
rect 13996 28960 14132 29000
rect 14188 30680 14228 31723
rect 14379 31604 14421 31613
rect 14379 31564 14380 31604
rect 14420 31564 14421 31604
rect 14379 31555 14421 31564
rect 13996 23969 14036 28960
rect 14188 28337 14228 30640
rect 14284 30596 14324 30605
rect 14284 29000 14324 30556
rect 14380 29597 14420 31555
rect 14476 31529 14516 32152
rect 14572 31865 14612 34000
rect 14763 33991 14805 34000
rect 14668 33872 14708 33881
rect 14860 33872 14900 35839
rect 14955 34040 14997 34049
rect 14955 34000 14956 34040
rect 14996 34000 14997 34040
rect 14955 33991 14997 34000
rect 14708 33832 14900 33872
rect 14668 33713 14708 33832
rect 14667 33704 14709 33713
rect 14667 33664 14668 33704
rect 14708 33664 14709 33704
rect 14667 33655 14709 33664
rect 14860 33704 14900 33713
rect 14956 33704 14996 33991
rect 14900 33664 14996 33704
rect 14860 33655 14900 33664
rect 15244 32864 15284 39031
rect 15340 38492 15380 49288
rect 15532 49288 15668 49328
rect 15435 49160 15477 49169
rect 15435 49120 15436 49160
rect 15476 49120 15477 49160
rect 15435 49111 15477 49120
rect 15436 44969 15476 49111
rect 15532 47312 15572 49288
rect 15627 49160 15669 49169
rect 15627 49120 15628 49160
rect 15668 49120 15669 49160
rect 15627 49111 15669 49120
rect 15628 48824 15668 49111
rect 15628 48775 15668 48784
rect 15532 45716 15572 47272
rect 15628 47312 15668 47321
rect 15724 47312 15764 49447
rect 15820 49169 15860 49456
rect 15916 49446 15956 49531
rect 15819 49160 15861 49169
rect 15819 49120 15820 49160
rect 15860 49120 15861 49160
rect 15819 49111 15861 49120
rect 15820 48245 15860 49111
rect 15819 48236 15861 48245
rect 15819 48196 15820 48236
rect 15860 48196 15861 48236
rect 15819 48187 15861 48196
rect 15668 47272 15764 47312
rect 15628 47263 15668 47272
rect 15724 46145 15764 47272
rect 16012 46817 16052 49708
rect 16108 47312 16148 50716
rect 16204 50681 16244 50968
rect 16203 50672 16245 50681
rect 16203 50632 16204 50672
rect 16244 50632 16245 50672
rect 16203 50623 16245 50632
rect 16203 48908 16245 48917
rect 16203 48868 16204 48908
rect 16244 48868 16245 48908
rect 16203 48859 16245 48868
rect 16204 48236 16244 48859
rect 16204 48187 16244 48196
rect 16011 46808 16053 46817
rect 16011 46768 16012 46808
rect 16052 46768 16053 46808
rect 16011 46759 16053 46768
rect 16108 46229 16148 47272
rect 16107 46220 16149 46229
rect 16107 46180 16108 46220
rect 16148 46180 16149 46220
rect 16107 46171 16149 46180
rect 15723 46136 15765 46145
rect 15723 46096 15724 46136
rect 15764 46096 15765 46136
rect 15723 46087 15765 46096
rect 15724 45800 15764 46087
rect 16108 45800 16148 46171
rect 16204 45800 16244 45809
rect 16108 45760 16204 45800
rect 15724 45751 15764 45760
rect 16204 45751 16244 45760
rect 15628 45716 15668 45725
rect 15532 45676 15628 45716
rect 15531 45380 15573 45389
rect 15531 45340 15532 45380
rect 15572 45340 15573 45380
rect 15531 45331 15573 45340
rect 15435 44960 15477 44969
rect 15435 44920 15436 44960
rect 15476 44920 15477 44960
rect 15435 44911 15477 44920
rect 15435 44456 15477 44465
rect 15435 44416 15436 44456
rect 15476 44416 15477 44456
rect 15435 44407 15477 44416
rect 15436 44322 15476 44407
rect 15532 43205 15572 45331
rect 15531 43196 15573 43205
rect 15531 43156 15532 43196
rect 15572 43156 15573 43196
rect 15531 43147 15573 43156
rect 15330 38452 15380 38492
rect 15330 38408 15370 38452
rect 15330 38368 15380 38408
rect 15340 38240 15380 38368
rect 15340 38200 15476 38240
rect 15340 38145 15380 38154
rect 15340 36233 15380 38105
rect 15436 38072 15476 38200
rect 15532 38072 15572 38081
rect 15436 38032 15532 38072
rect 15532 38023 15572 38032
rect 15435 37904 15477 37913
rect 15435 37864 15436 37904
rect 15476 37864 15477 37904
rect 15435 37855 15477 37864
rect 15339 36224 15381 36233
rect 15339 36184 15340 36224
rect 15380 36184 15381 36224
rect 15339 36175 15381 36184
rect 15436 32864 15476 37855
rect 15531 35216 15573 35225
rect 15531 35176 15532 35216
rect 15572 35176 15573 35216
rect 15531 35167 15573 35176
rect 15532 34721 15572 35167
rect 15531 34712 15573 34721
rect 15531 34672 15532 34712
rect 15572 34672 15573 34712
rect 15531 34663 15573 34672
rect 15628 33368 15668 45676
rect 16011 45632 16053 45641
rect 16011 45592 16012 45632
rect 16052 45592 16053 45632
rect 16011 45583 16053 45592
rect 15723 44456 15765 44465
rect 15723 44416 15724 44456
rect 15764 44416 15765 44456
rect 15723 44407 15765 44416
rect 15724 44288 15764 44407
rect 15724 44239 15764 44248
rect 15820 44288 15860 44299
rect 15820 44213 15860 44248
rect 15819 44204 15861 44213
rect 15819 44164 15820 44204
rect 15860 44164 15861 44204
rect 15819 44155 15861 44164
rect 15819 43448 15861 43457
rect 15819 43408 15820 43448
rect 15860 43408 15861 43448
rect 15819 43399 15861 43408
rect 15820 43314 15860 43399
rect 15819 43196 15861 43205
rect 15819 43156 15820 43196
rect 15860 43156 15861 43196
rect 15819 43147 15861 43156
rect 15723 39752 15765 39761
rect 15723 39712 15724 39752
rect 15764 39712 15765 39752
rect 15723 39703 15765 39712
rect 15724 33713 15764 39703
rect 15820 37913 15860 43147
rect 16012 41525 16052 45583
rect 16107 44624 16149 44633
rect 16107 44584 16108 44624
rect 16148 44584 16149 44624
rect 16107 44575 16149 44584
rect 16108 43457 16148 44575
rect 16203 44372 16245 44381
rect 16203 44332 16204 44372
rect 16244 44332 16245 44372
rect 16203 44323 16245 44332
rect 16204 44288 16244 44323
rect 16204 44237 16244 44248
rect 16300 44288 16340 51556
rect 16396 49757 16436 55159
rect 16492 54867 16532 55336
rect 16588 55217 16628 55588
rect 16875 55588 16876 55628
rect 16916 55588 16917 55628
rect 16875 55579 16917 55588
rect 16876 55544 16916 55579
rect 16972 55553 17012 55915
rect 16876 55493 16916 55504
rect 16971 55544 17013 55553
rect 16971 55504 16972 55544
rect 17012 55504 17013 55544
rect 16971 55495 17013 55504
rect 16684 55376 16724 55385
rect 16587 55208 16629 55217
rect 16587 55168 16588 55208
rect 16628 55168 16629 55208
rect 16587 55159 16629 55168
rect 16684 54881 16724 55336
rect 16779 55376 16821 55385
rect 16779 55336 16780 55376
rect 16820 55336 16821 55376
rect 16779 55327 16821 55336
rect 16780 55040 16820 55327
rect 16780 54991 16820 55000
rect 16588 54867 16628 54876
rect 16492 54827 16588 54867
rect 16588 54818 16628 54827
rect 16683 54872 16725 54881
rect 16683 54832 16684 54872
rect 16724 54832 16725 54872
rect 16683 54823 16725 54832
rect 16972 54452 17012 55495
rect 16492 54412 17012 54452
rect 16492 50252 16532 54412
rect 16587 54284 16629 54293
rect 16587 54244 16588 54284
rect 16628 54244 16629 54284
rect 16587 54235 16629 54244
rect 16588 53117 16628 54235
rect 16779 54200 16821 54209
rect 16779 54160 16780 54200
rect 16820 54160 16821 54200
rect 16779 54151 16821 54160
rect 16780 54032 16820 54151
rect 16683 53864 16725 53873
rect 16683 53824 16684 53864
rect 16724 53824 16725 53864
rect 16683 53815 16725 53824
rect 16684 53355 16724 53815
rect 16684 53306 16724 53315
rect 16587 53108 16629 53117
rect 16587 53068 16588 53108
rect 16628 53068 16629 53108
rect 16587 53059 16629 53068
rect 16780 52940 16820 53992
rect 16972 53873 17012 53958
rect 16971 53864 17013 53873
rect 16971 53824 16972 53864
rect 17012 53824 17013 53864
rect 16971 53815 17013 53824
rect 16875 53528 16917 53537
rect 16875 53488 16876 53528
rect 16916 53488 16917 53528
rect 16875 53479 16917 53488
rect 16876 53394 16916 53479
rect 17068 53276 17108 56092
rect 17164 54368 17204 56260
rect 17260 54965 17300 56764
rect 17356 56309 17396 57016
rect 17452 56384 17492 57604
rect 17548 57065 17588 57688
rect 17547 57056 17589 57065
rect 17547 57016 17548 57056
rect 17588 57016 17589 57056
rect 17547 57007 17589 57016
rect 17452 56335 17492 56344
rect 17548 56384 17588 57007
rect 17355 56300 17397 56309
rect 17355 56260 17356 56300
rect 17396 56260 17397 56300
rect 17355 56251 17397 56260
rect 17451 55292 17493 55301
rect 17451 55252 17452 55292
rect 17492 55252 17493 55292
rect 17451 55243 17493 55252
rect 17259 54956 17301 54965
rect 17259 54916 17260 54956
rect 17300 54916 17301 54956
rect 17259 54907 17301 54916
rect 17355 54872 17397 54881
rect 17355 54832 17356 54872
rect 17396 54832 17397 54872
rect 17355 54823 17397 54832
rect 17452 54872 17492 55243
rect 17452 54823 17492 54832
rect 17356 54738 17396 54823
rect 17164 54328 17300 54368
rect 17164 54200 17204 54211
rect 17164 54125 17204 54160
rect 17163 54116 17205 54125
rect 17163 54076 17164 54116
rect 17204 54076 17205 54116
rect 17163 54067 17205 54076
rect 17260 53453 17300 54328
rect 17356 54116 17396 54125
rect 17356 53537 17396 54076
rect 17451 54116 17493 54125
rect 17451 54076 17452 54116
rect 17492 54076 17493 54116
rect 17451 54067 17493 54076
rect 17355 53528 17397 53537
rect 17355 53488 17356 53528
rect 17396 53488 17397 53528
rect 17355 53479 17397 53488
rect 17259 53444 17301 53453
rect 17259 53404 17260 53444
rect 17300 53404 17301 53444
rect 17259 53395 17301 53404
rect 17260 53276 17300 53285
rect 17068 53236 17204 53276
rect 17067 53108 17109 53117
rect 17067 53068 17068 53108
rect 17108 53068 17109 53108
rect 17067 53059 17109 53068
rect 17068 52974 17108 53059
rect 16780 52900 17012 52940
rect 16972 52184 17012 52900
rect 16972 52144 17108 52184
rect 16779 52100 16821 52109
rect 16779 52060 16780 52100
rect 16820 52060 16821 52100
rect 16779 52051 16821 52060
rect 16780 51848 16820 52051
rect 16971 52016 17013 52025
rect 16971 51976 16972 52016
rect 17012 51976 17013 52016
rect 16971 51967 17013 51976
rect 16820 51808 16916 51848
rect 16780 51799 16820 51808
rect 16779 51008 16821 51017
rect 16779 50968 16780 51008
rect 16820 50968 16821 51008
rect 16779 50959 16821 50968
rect 16683 50420 16725 50429
rect 16683 50380 16684 50420
rect 16724 50380 16725 50420
rect 16683 50371 16725 50380
rect 16492 50212 16628 50252
rect 16588 50093 16628 50212
rect 16492 50084 16532 50093
rect 16395 49748 16437 49757
rect 16395 49708 16396 49748
rect 16436 49708 16437 49748
rect 16395 49699 16437 49708
rect 16395 49496 16437 49505
rect 16395 49456 16396 49496
rect 16436 49456 16437 49496
rect 16395 49447 16437 49456
rect 16396 49362 16436 49447
rect 16396 48068 16436 48077
rect 16396 47489 16436 48028
rect 16395 47480 16437 47489
rect 16395 47440 16396 47480
rect 16436 47440 16437 47480
rect 16395 47431 16437 47440
rect 16492 46640 16532 50044
rect 16587 50084 16629 50093
rect 16587 50044 16588 50084
rect 16628 50044 16629 50084
rect 16587 50035 16629 50044
rect 16587 49748 16629 49757
rect 16587 49708 16588 49748
rect 16628 49708 16629 49748
rect 16587 49699 16629 49708
rect 16588 49505 16628 49699
rect 16587 49496 16629 49505
rect 16587 49456 16588 49496
rect 16628 49456 16629 49496
rect 16587 49447 16629 49456
rect 16588 47984 16628 47993
rect 16684 47984 16724 50371
rect 16780 48824 16820 50959
rect 16876 49757 16916 51808
rect 16972 50177 17012 51967
rect 17068 51101 17108 52144
rect 17067 51092 17109 51101
rect 17067 51052 17068 51092
rect 17108 51052 17109 51092
rect 17067 51043 17109 51052
rect 17068 50429 17108 51043
rect 17067 50420 17109 50429
rect 17067 50380 17068 50420
rect 17108 50380 17109 50420
rect 17067 50371 17109 50380
rect 17164 50336 17204 53236
rect 17260 52109 17300 53236
rect 17452 52949 17492 54067
rect 17451 52940 17493 52949
rect 17451 52900 17452 52940
rect 17492 52900 17493 52940
rect 17451 52891 17493 52900
rect 17452 52520 17492 52891
rect 17356 52480 17452 52520
rect 17259 52100 17301 52109
rect 17259 52060 17260 52100
rect 17300 52060 17301 52100
rect 17259 52051 17301 52060
rect 17260 51834 17300 51843
rect 17260 51269 17300 51794
rect 17259 51260 17301 51269
rect 17259 51220 17260 51260
rect 17300 51220 17301 51260
rect 17259 51211 17301 51220
rect 17259 50504 17301 50513
rect 17259 50464 17260 50504
rect 17300 50464 17301 50504
rect 17259 50455 17301 50464
rect 17164 50287 17204 50296
rect 17067 50252 17109 50261
rect 17067 50212 17068 50252
rect 17108 50212 17109 50252
rect 17067 50203 17109 50212
rect 16971 50168 17013 50177
rect 16971 50128 16972 50168
rect 17012 50128 17013 50168
rect 16971 50119 17013 50128
rect 16875 49748 16917 49757
rect 16875 49708 16876 49748
rect 16916 49708 16917 49748
rect 16875 49699 16917 49708
rect 16924 49505 16964 49514
rect 16964 49465 17012 49496
rect 16924 49456 17012 49465
rect 16972 48992 17012 49456
rect 17068 49412 17108 50203
rect 17163 50168 17205 50177
rect 17163 50128 17164 50168
rect 17204 50128 17205 50168
rect 17163 50119 17205 50128
rect 17068 49363 17108 49372
rect 17068 48992 17108 49001
rect 16972 48952 17068 48992
rect 17068 48943 17108 48952
rect 16876 48824 16916 48833
rect 16780 48784 16876 48824
rect 16876 47993 16916 48784
rect 16875 47984 16917 47993
rect 16628 47944 16820 47984
rect 16588 47935 16628 47944
rect 16780 47816 16820 47944
rect 16875 47944 16876 47984
rect 16916 47944 16917 47984
rect 16875 47935 16917 47944
rect 16780 47776 17108 47816
rect 16779 47480 16821 47489
rect 16779 47440 16780 47480
rect 16820 47440 16821 47480
rect 16779 47431 16821 47440
rect 16780 47346 16820 47431
rect 16971 47312 17013 47321
rect 16636 47270 16676 47279
rect 16971 47272 16972 47312
rect 17012 47272 17013 47312
rect 16971 47263 17013 47272
rect 16636 47228 16676 47230
rect 16636 47188 16724 47228
rect 16684 46724 16724 47188
rect 16972 47178 17012 47263
rect 16684 46675 16724 46684
rect 16300 44239 16340 44248
rect 16396 46600 16532 46640
rect 16107 43448 16149 43457
rect 16107 43408 16108 43448
rect 16148 43408 16149 43448
rect 16107 43399 16149 43408
rect 16011 41516 16053 41525
rect 16011 41476 16012 41516
rect 16052 41476 16053 41516
rect 16011 41467 16053 41476
rect 16299 39668 16341 39677
rect 16299 39628 16300 39668
rect 16340 39628 16341 39668
rect 16299 39619 16341 39628
rect 16300 39173 16340 39619
rect 16299 39164 16341 39173
rect 16299 39124 16300 39164
rect 16340 39124 16341 39164
rect 16299 39115 16341 39124
rect 15819 37904 15861 37913
rect 15819 37864 15820 37904
rect 15860 37864 15861 37904
rect 15819 37855 15861 37864
rect 16012 34376 16052 34385
rect 15723 33704 15765 33713
rect 15723 33664 15724 33704
rect 15764 33664 15765 33704
rect 15723 33655 15765 33664
rect 16012 33545 16052 34336
rect 16108 33704 16148 33713
rect 16011 33536 16053 33545
rect 16011 33496 16012 33536
rect 16052 33496 16053 33536
rect 16011 33487 16053 33496
rect 16108 33377 16148 33664
rect 16203 33704 16245 33713
rect 16203 33664 16204 33704
rect 16244 33664 16245 33704
rect 16203 33655 16245 33664
rect 16107 33368 16149 33377
rect 15628 33328 16052 33368
rect 15436 32824 15764 32864
rect 14763 32696 14805 32705
rect 14763 32656 14764 32696
rect 14804 32656 14805 32696
rect 14763 32647 14805 32656
rect 14668 32201 14708 32286
rect 14667 32192 14709 32201
rect 14667 32152 14668 32192
rect 14708 32152 14709 32192
rect 14667 32143 14709 32152
rect 14667 32024 14709 32033
rect 14667 31984 14668 32024
rect 14708 31984 14709 32024
rect 14667 31975 14709 31984
rect 14668 31890 14708 31975
rect 14571 31856 14613 31865
rect 14571 31816 14572 31856
rect 14612 31816 14613 31856
rect 14571 31807 14613 31816
rect 14475 31520 14517 31529
rect 14475 31480 14476 31520
rect 14516 31480 14517 31520
rect 14475 31471 14517 31480
rect 14764 31352 14804 32647
rect 14860 32192 14900 32201
rect 14860 32033 14900 32152
rect 15147 32192 15189 32201
rect 15147 32152 15148 32192
rect 15188 32152 15189 32192
rect 15147 32143 15189 32152
rect 14956 32108 14996 32117
rect 14996 32068 15092 32108
rect 14956 32059 14996 32068
rect 14859 32024 14901 32033
rect 14859 31984 14860 32024
rect 14900 31984 14901 32024
rect 14859 31975 14901 31984
rect 14859 31856 14901 31865
rect 14859 31816 14860 31856
rect 14900 31816 14901 31856
rect 14859 31807 14901 31816
rect 14668 31312 14764 31352
rect 14571 31100 14613 31109
rect 14571 31060 14572 31100
rect 14612 31060 14613 31100
rect 14571 31051 14613 31060
rect 14572 30689 14612 31051
rect 14571 30680 14613 30689
rect 14571 30640 14572 30680
rect 14612 30640 14613 30680
rect 14571 30631 14613 30640
rect 14475 29840 14517 29849
rect 14475 29800 14476 29840
rect 14516 29800 14517 29840
rect 14475 29791 14517 29800
rect 14476 29706 14516 29791
rect 14379 29588 14421 29597
rect 14379 29548 14380 29588
rect 14420 29548 14421 29588
rect 14379 29539 14421 29548
rect 14380 29168 14420 29539
rect 14476 29168 14516 29177
rect 14380 29128 14476 29168
rect 14476 29119 14516 29128
rect 14284 28960 14420 29000
rect 14187 28328 14229 28337
rect 14187 28288 14188 28328
rect 14228 28288 14229 28328
rect 14187 28279 14229 28288
rect 14283 27656 14325 27665
rect 14283 27616 14284 27656
rect 14324 27616 14325 27656
rect 14283 27607 14325 27616
rect 14284 27522 14324 27607
rect 14187 27068 14229 27077
rect 14187 27028 14188 27068
rect 14228 27028 14229 27068
rect 14187 27019 14229 27028
rect 14188 26816 14228 27019
rect 14188 26767 14228 26776
rect 14092 26144 14132 26153
rect 14092 25565 14132 26104
rect 14188 26144 14228 26153
rect 14380 26144 14420 28960
rect 14476 28328 14516 28337
rect 14476 27824 14516 28288
rect 14476 27775 14516 27784
rect 14572 28328 14612 30631
rect 14668 30428 14708 31312
rect 14764 31303 14804 31312
rect 14763 30680 14805 30689
rect 14763 30640 14764 30680
rect 14804 30640 14805 30680
rect 14763 30631 14805 30640
rect 14764 30546 14804 30631
rect 14668 30388 14804 30428
rect 14667 30260 14709 30269
rect 14667 30220 14668 30260
rect 14708 30220 14709 30260
rect 14667 30211 14709 30220
rect 14668 30101 14708 30211
rect 14667 30092 14709 30101
rect 14667 30052 14668 30092
rect 14708 30052 14709 30092
rect 14667 30043 14709 30052
rect 14668 29958 14708 30043
rect 14764 29849 14804 30388
rect 14763 29840 14805 29849
rect 14763 29800 14764 29840
rect 14804 29800 14805 29840
rect 14763 29791 14805 29800
rect 14475 27488 14517 27497
rect 14475 27448 14476 27488
rect 14516 27448 14517 27488
rect 14475 27439 14517 27448
rect 14228 26104 14420 26144
rect 14091 25556 14133 25565
rect 14091 25516 14092 25556
rect 14132 25516 14133 25556
rect 14091 25507 14133 25516
rect 14091 24884 14133 24893
rect 14091 24844 14092 24884
rect 14132 24844 14133 24884
rect 14091 24835 14133 24844
rect 13995 23960 14037 23969
rect 13995 23920 13996 23960
rect 14036 23920 14037 23960
rect 13995 23911 14037 23920
rect 13995 23792 14037 23801
rect 13995 23752 13996 23792
rect 14036 23752 14037 23792
rect 13995 23743 14037 23752
rect 14092 23792 14132 24835
rect 14188 24137 14228 26104
rect 14380 25304 14420 25315
rect 14380 25229 14420 25264
rect 14379 25220 14421 25229
rect 14379 25180 14380 25220
rect 14420 25180 14421 25220
rect 14379 25171 14421 25180
rect 14380 24641 14420 25171
rect 14379 24632 14421 24641
rect 14379 24592 14380 24632
rect 14420 24592 14421 24632
rect 14379 24583 14421 24592
rect 14380 24498 14420 24583
rect 14187 24128 14229 24137
rect 14187 24088 14188 24128
rect 14228 24088 14229 24128
rect 14187 24079 14229 24088
rect 14379 23960 14421 23969
rect 14379 23920 14380 23960
rect 14420 23920 14421 23960
rect 14379 23911 14421 23920
rect 13996 23658 14036 23743
rect 14092 23708 14132 23752
rect 14283 23792 14325 23801
rect 14283 23752 14284 23792
rect 14324 23752 14325 23792
rect 14283 23743 14325 23752
rect 14092 23668 14228 23708
rect 13996 23120 14036 23129
rect 13900 23080 13996 23120
rect 13900 19097 13940 23080
rect 13996 23071 14036 23080
rect 13995 22532 14037 22541
rect 13995 22492 13996 22532
rect 14036 22492 14037 22532
rect 13995 22483 14037 22492
rect 13996 21608 14036 22483
rect 14091 22364 14133 22373
rect 14091 22324 14092 22364
rect 14132 22324 14133 22364
rect 14091 22315 14133 22324
rect 14092 21869 14132 22315
rect 14091 21860 14133 21869
rect 14091 21820 14092 21860
rect 14132 21820 14133 21860
rect 14091 21811 14133 21820
rect 13996 21356 14036 21568
rect 14092 21608 14132 21811
rect 14092 21559 14132 21568
rect 13996 21316 14132 21356
rect 13995 20768 14037 20777
rect 13995 20728 13996 20768
rect 14036 20728 14037 20768
rect 13995 20719 14037 20728
rect 13996 20609 14036 20719
rect 13995 20600 14037 20609
rect 13995 20560 13996 20600
rect 14036 20560 14037 20600
rect 13995 20551 14037 20560
rect 13996 20096 14036 20551
rect 13996 20047 14036 20056
rect 14092 20021 14132 21316
rect 14188 20189 14228 23668
rect 14284 23045 14324 23743
rect 14283 23036 14325 23045
rect 14283 22996 14284 23036
rect 14324 22996 14325 23036
rect 14283 22987 14325 22996
rect 14187 20180 14229 20189
rect 14187 20140 14188 20180
rect 14228 20140 14229 20180
rect 14187 20131 14229 20140
rect 14091 20012 14133 20021
rect 14091 19972 14092 20012
rect 14132 19972 14133 20012
rect 14091 19963 14133 19972
rect 13995 19928 14037 19937
rect 13995 19888 13996 19928
rect 14036 19888 14037 19928
rect 13995 19879 14037 19888
rect 13996 19592 14036 19879
rect 14188 19844 14228 19853
rect 13996 19552 14132 19592
rect 13995 19340 14037 19349
rect 13995 19300 13996 19340
rect 14036 19300 14037 19340
rect 13995 19291 14037 19300
rect 13996 19206 14036 19291
rect 14092 19256 14132 19552
rect 14188 19265 14228 19804
rect 14284 19349 14324 22987
rect 14380 22625 14420 23911
rect 14379 22616 14421 22625
rect 14379 22576 14380 22616
rect 14420 22576 14421 22616
rect 14379 22567 14421 22576
rect 14379 21020 14421 21029
rect 14379 20980 14380 21020
rect 14420 20980 14421 21020
rect 14379 20971 14421 20980
rect 14380 20768 14420 20971
rect 14380 20719 14420 20728
rect 14476 20609 14516 27439
rect 14572 26573 14612 28288
rect 14763 27656 14805 27665
rect 14763 27616 14764 27656
rect 14804 27616 14805 27656
rect 14763 27607 14805 27616
rect 14667 27572 14709 27581
rect 14667 27532 14668 27572
rect 14708 27532 14709 27572
rect 14667 27523 14709 27532
rect 14571 26564 14613 26573
rect 14571 26524 14572 26564
rect 14612 26524 14613 26564
rect 14571 26515 14613 26524
rect 14668 26153 14708 27523
rect 14667 26144 14709 26153
rect 14667 26104 14668 26144
rect 14708 26104 14709 26144
rect 14667 26095 14709 26104
rect 14571 26060 14613 26069
rect 14571 26020 14572 26060
rect 14612 26020 14613 26060
rect 14571 26011 14613 26020
rect 14572 25926 14612 26011
rect 14668 26010 14708 26095
rect 14667 25640 14709 25649
rect 14667 25600 14668 25640
rect 14708 25600 14709 25640
rect 14667 25591 14709 25600
rect 14571 25556 14613 25565
rect 14571 25516 14572 25556
rect 14612 25516 14613 25556
rect 14571 25507 14613 25516
rect 14572 25422 14612 25507
rect 14572 24380 14612 24389
rect 14572 23969 14612 24340
rect 14571 23960 14613 23969
rect 14571 23920 14572 23960
rect 14612 23920 14613 23960
rect 14571 23911 14613 23920
rect 14571 23792 14613 23801
rect 14571 23752 14572 23792
rect 14612 23752 14613 23792
rect 14571 23743 14613 23752
rect 14572 23658 14612 23743
rect 14572 21608 14612 21617
rect 14475 20600 14517 20609
rect 14475 20560 14476 20600
rect 14516 20560 14517 20600
rect 14475 20551 14517 20560
rect 14379 20096 14421 20105
rect 14379 20056 14380 20096
rect 14420 20056 14421 20096
rect 14379 20047 14421 20056
rect 14380 19962 14420 20047
rect 14475 19844 14517 19853
rect 14475 19804 14476 19844
rect 14516 19804 14517 19844
rect 14475 19795 14517 19804
rect 14476 19710 14516 19795
rect 14379 19676 14421 19685
rect 14379 19636 14380 19676
rect 14420 19636 14421 19676
rect 14379 19627 14421 19636
rect 14283 19340 14325 19349
rect 14283 19300 14284 19340
rect 14324 19300 14325 19340
rect 14283 19291 14325 19300
rect 13899 19088 13941 19097
rect 13899 19048 13900 19088
rect 13940 19048 13941 19088
rect 13899 19039 13941 19048
rect 13803 18752 13845 18761
rect 13803 18712 13804 18752
rect 13844 18712 13845 18752
rect 13803 18703 13845 18712
rect 13803 18584 13845 18593
rect 13803 18544 13804 18584
rect 13844 18544 13845 18584
rect 13803 18535 13845 18544
rect 13804 18450 13844 18535
rect 14092 17660 14132 19216
rect 14187 19256 14229 19265
rect 14187 19216 14188 19256
rect 14228 19216 14229 19256
rect 14187 19207 14229 19216
rect 13516 17536 13652 17576
rect 13804 17620 14132 17660
rect 13516 17081 13556 17536
rect 13515 17072 13557 17081
rect 13515 17032 13516 17072
rect 13556 17032 13557 17072
rect 13515 17023 13557 17032
rect 13612 17072 13652 17081
rect 13419 15896 13461 15905
rect 13419 15856 13420 15896
rect 13460 15856 13461 15896
rect 13419 15847 13461 15856
rect 13420 15560 13460 15569
rect 13420 14972 13460 15520
rect 13612 15317 13652 17032
rect 13708 16232 13748 16241
rect 13708 15569 13748 16192
rect 13707 15560 13749 15569
rect 13707 15520 13708 15560
rect 13748 15520 13749 15560
rect 13707 15511 13749 15520
rect 13611 15308 13653 15317
rect 13611 15268 13612 15308
rect 13652 15268 13653 15308
rect 13611 15259 13653 15268
rect 13804 14972 13844 17620
rect 14187 16904 14229 16913
rect 14187 16864 14188 16904
rect 14228 16864 14229 16904
rect 14187 16855 14229 16864
rect 13900 16064 13940 16073
rect 13900 15555 13940 16024
rect 13995 15812 14037 15821
rect 13995 15772 13996 15812
rect 14036 15772 14037 15812
rect 13995 15763 14037 15772
rect 13900 15506 13940 15515
rect 13996 15224 14036 15763
rect 14091 15728 14133 15737
rect 14091 15688 14092 15728
rect 14132 15688 14133 15728
rect 14091 15679 14133 15688
rect 14092 15594 14132 15679
rect 13420 14932 13844 14972
rect 13516 14720 13556 14729
rect 13324 14680 13459 14720
rect 13228 14636 13268 14645
rect 13419 14636 13459 14680
rect 13268 14596 13364 14636
rect 13419 14596 13460 14636
rect 13228 14587 13268 14596
rect 13324 14477 13364 14596
rect 13323 14468 13365 14477
rect 13132 14428 13268 14468
rect 13132 14048 13172 14057
rect 13036 14008 13132 14048
rect 13132 13889 13172 14008
rect 13131 13880 13173 13889
rect 13131 13840 13132 13880
rect 13172 13840 13173 13880
rect 13131 13831 13173 13840
rect 13131 13208 13173 13217
rect 13131 13168 13132 13208
rect 13172 13168 13173 13208
rect 13131 13159 13173 13168
rect 12940 12620 12980 12629
rect 12940 11789 12980 12580
rect 13132 12536 13172 13159
rect 13228 13040 13268 14428
rect 13323 14428 13324 14468
rect 13364 14428 13365 14468
rect 13323 14419 13365 14428
rect 13324 13796 13364 13805
rect 13324 13208 13364 13756
rect 13420 13385 13460 14596
rect 13516 14477 13556 14680
rect 13612 14720 13652 14729
rect 13515 14468 13557 14477
rect 13515 14428 13516 14468
rect 13556 14428 13557 14468
rect 13515 14419 13557 14428
rect 13419 13376 13461 13385
rect 13419 13336 13420 13376
rect 13460 13336 13461 13376
rect 13419 13327 13461 13336
rect 13612 13301 13652 14680
rect 13804 14636 13844 14932
rect 13708 14596 13844 14636
rect 13900 15184 14036 15224
rect 13611 13292 13653 13301
rect 13611 13252 13612 13292
rect 13652 13252 13653 13292
rect 13611 13243 13653 13252
rect 13324 13159 13364 13168
rect 13419 13208 13461 13217
rect 13419 13168 13420 13208
rect 13460 13168 13461 13208
rect 13419 13159 13461 13168
rect 13420 13074 13460 13159
rect 13708 13040 13748 14596
rect 13900 14048 13940 15184
rect 14188 15140 14228 16855
rect 14284 15560 14324 15569
rect 14284 15317 14324 15520
rect 14283 15308 14325 15317
rect 14283 15268 14284 15308
rect 14324 15268 14325 15308
rect 14283 15259 14325 15268
rect 14188 15100 14324 15140
rect 13995 14888 14037 14897
rect 13995 14848 13996 14888
rect 14036 14848 14037 14888
rect 13995 14839 14037 14848
rect 13996 14804 14036 14839
rect 13996 14132 14036 14764
rect 14092 14720 14132 14729
rect 14132 14680 14228 14720
rect 14092 14671 14132 14680
rect 14188 14141 14228 14680
rect 14187 14132 14229 14141
rect 13996 14092 14132 14132
rect 13940 14008 14036 14048
rect 13900 13999 13940 14008
rect 13803 13712 13845 13721
rect 13803 13672 13804 13712
rect 13844 13672 13845 13712
rect 13803 13663 13845 13672
rect 13804 13292 13844 13663
rect 13804 13243 13844 13252
rect 13899 13292 13941 13301
rect 13899 13252 13900 13292
rect 13940 13252 13941 13292
rect 13899 13243 13941 13252
rect 13228 13000 13364 13040
rect 13132 12496 13268 12536
rect 13035 12284 13077 12293
rect 13035 12244 13036 12284
rect 13076 12244 13077 12284
rect 13035 12235 13077 12244
rect 12939 11780 12981 11789
rect 12939 11740 12940 11780
rect 12980 11740 12981 11780
rect 12939 11731 12981 11740
rect 13036 11033 13076 12235
rect 13132 11696 13172 11705
rect 13132 11192 13172 11656
rect 13228 11696 13268 12496
rect 13228 11647 13268 11656
rect 13324 11621 13364 13000
rect 13612 13000 13748 13040
rect 13612 12956 13652 13000
rect 13516 12916 13652 12956
rect 13419 12872 13461 12881
rect 13419 12832 13420 12872
rect 13460 12832 13461 12872
rect 13419 12823 13461 12832
rect 13323 11612 13365 11621
rect 13323 11572 13324 11612
rect 13364 11572 13365 11612
rect 13323 11563 13365 11572
rect 13420 11360 13460 12823
rect 13132 11143 13172 11152
rect 13324 11320 13460 11360
rect 12940 11024 12980 11033
rect 12940 10865 12980 10984
rect 13035 11024 13077 11033
rect 13035 10984 13036 11024
rect 13076 10984 13077 11024
rect 13035 10975 13077 10984
rect 12939 10856 12981 10865
rect 12939 10816 12940 10856
rect 12980 10816 12981 10856
rect 12939 10807 12981 10816
rect 12843 8756 12885 8765
rect 12843 8716 12844 8756
rect 12884 8716 12885 8756
rect 12843 8707 12885 8716
rect 12747 8672 12789 8681
rect 12747 8632 12748 8672
rect 12788 8632 12789 8672
rect 12747 8623 12789 8632
rect 12940 8261 12980 10807
rect 12939 8252 12981 8261
rect 12939 8212 12940 8252
rect 12980 8212 12981 8252
rect 12939 8203 12981 8212
rect 12651 8000 12693 8009
rect 12651 7960 12652 8000
rect 12692 7960 12693 8000
rect 12651 7951 12693 7960
rect 12844 8000 12884 8009
rect 12555 7916 12597 7925
rect 12555 7876 12556 7916
rect 12596 7876 12597 7916
rect 12555 7867 12597 7876
rect 12364 7036 12500 7076
rect 12167 6868 12212 6908
rect 12167 6824 12207 6868
rect 12167 6784 12404 6824
rect 12267 6656 12309 6665
rect 12267 6616 12268 6656
rect 12308 6616 12309 6656
rect 12267 6607 12309 6616
rect 12172 6497 12212 6582
rect 12076 6488 12116 6497
rect 11979 5396 12021 5405
rect 11979 5356 11980 5396
rect 12020 5356 12021 5396
rect 11979 5347 12021 5356
rect 11883 5144 11925 5153
rect 11883 5104 11884 5144
rect 11924 5104 11925 5144
rect 11883 5095 11925 5104
rect 11787 5060 11829 5069
rect 11787 5020 11788 5060
rect 11828 5020 11829 5060
rect 11787 5011 11829 5020
rect 12076 4985 12116 6448
rect 12171 6488 12213 6497
rect 12171 6448 12172 6488
rect 12212 6448 12213 6488
rect 12171 6439 12213 6448
rect 12268 5573 12308 6607
rect 12267 5564 12309 5573
rect 12267 5524 12268 5564
rect 12308 5524 12309 5564
rect 12267 5515 12309 5524
rect 12268 5153 12308 5238
rect 12267 5144 12309 5153
rect 12267 5104 12268 5144
rect 12308 5104 12309 5144
rect 12267 5095 12309 5104
rect 11884 4976 11924 4985
rect 11884 4892 11924 4936
rect 12075 4976 12117 4985
rect 12364 4976 12404 6784
rect 12460 5657 12500 7036
rect 12556 6665 12596 7867
rect 12555 6656 12597 6665
rect 12555 6616 12556 6656
rect 12596 6616 12597 6656
rect 12555 6607 12597 6616
rect 12556 6488 12596 6497
rect 12556 6320 12596 6448
rect 12652 6488 12692 7951
rect 12747 7496 12789 7505
rect 12747 7456 12748 7496
rect 12788 7456 12789 7496
rect 12747 7447 12789 7456
rect 12748 7160 12788 7447
rect 12844 7412 12884 7960
rect 12939 8000 12981 8009
rect 12939 7960 12940 8000
rect 12980 7960 12981 8000
rect 12939 7951 12981 7960
rect 12940 7866 12980 7951
rect 12940 7412 12980 7421
rect 12844 7372 12940 7412
rect 12940 7363 12980 7372
rect 12748 7111 12788 7120
rect 13036 6749 13076 10975
rect 13324 10352 13364 11320
rect 13419 11024 13461 11033
rect 13419 10984 13420 11024
rect 13460 10984 13461 11024
rect 13419 10975 13461 10984
rect 13420 10890 13460 10975
rect 13132 10312 13364 10352
rect 13132 7328 13172 10312
rect 13228 10184 13268 10193
rect 13228 9680 13268 10144
rect 13323 10184 13365 10193
rect 13323 10144 13324 10184
rect 13364 10144 13365 10184
rect 13323 10135 13365 10144
rect 13324 10050 13364 10135
rect 13420 9680 13460 9689
rect 13228 9640 13420 9680
rect 13420 9631 13460 9640
rect 13228 9512 13268 9521
rect 13228 9353 13268 9472
rect 13227 9344 13269 9353
rect 13227 9304 13228 9344
rect 13268 9304 13269 9344
rect 13227 9295 13269 9304
rect 13324 7916 13364 7925
rect 13132 7288 13268 7328
rect 13131 7160 13173 7169
rect 13131 7120 13132 7160
rect 13172 7120 13173 7160
rect 13131 7111 13173 7120
rect 13132 7026 13172 7111
rect 13035 6740 13077 6749
rect 13035 6700 13036 6740
rect 13076 6700 13077 6740
rect 13035 6691 13077 6700
rect 12652 6439 12692 6448
rect 12843 6488 12885 6497
rect 12843 6448 12844 6488
rect 12884 6448 12885 6488
rect 12843 6439 12885 6448
rect 13131 6488 13173 6497
rect 13131 6448 13132 6488
rect 13172 6448 13173 6488
rect 13131 6439 13173 6448
rect 12556 6280 12788 6320
rect 12748 5900 12788 6280
rect 12748 5851 12788 5860
rect 12459 5648 12501 5657
rect 12459 5608 12460 5648
rect 12500 5608 12501 5648
rect 12459 5599 12501 5608
rect 12556 5648 12596 5659
rect 12460 5237 12500 5599
rect 12556 5573 12596 5608
rect 12555 5564 12597 5573
rect 12555 5524 12556 5564
rect 12596 5524 12597 5564
rect 12555 5515 12597 5524
rect 12459 5228 12501 5237
rect 12459 5188 12460 5228
rect 12500 5188 12501 5228
rect 12556 5228 12596 5515
rect 12844 5480 12884 6439
rect 13035 6404 13077 6413
rect 13035 6364 13036 6404
rect 13076 6364 13077 6404
rect 13035 6355 13077 6364
rect 13036 6270 13076 6355
rect 13132 6354 13172 6439
rect 12940 5657 12980 5742
rect 12939 5648 12981 5657
rect 12939 5608 12940 5648
rect 12980 5608 12981 5648
rect 12939 5599 12981 5608
rect 12844 5440 12980 5480
rect 12556 5188 12692 5228
rect 12459 5179 12501 5188
rect 12555 5060 12597 5069
rect 12555 5020 12556 5060
rect 12596 5020 12597 5060
rect 12555 5011 12597 5020
rect 12075 4936 12076 4976
rect 12116 4936 12117 4976
rect 12075 4927 12117 4936
rect 12268 4936 12404 4976
rect 12460 4976 12500 4985
rect 11788 4852 11924 4892
rect 11788 4145 11828 4852
rect 12076 4808 12116 4927
rect 12171 4892 12213 4901
rect 12171 4852 12172 4892
rect 12212 4852 12213 4892
rect 12171 4843 12213 4852
rect 12076 4759 12116 4768
rect 12172 4388 12212 4843
rect 12172 4339 12212 4348
rect 11787 4136 11829 4145
rect 11787 4096 11788 4136
rect 11828 4096 11829 4136
rect 11787 4087 11829 4096
rect 11979 4136 12021 4145
rect 11979 4096 11980 4136
rect 12020 4096 12021 4136
rect 11979 4087 12021 4096
rect 11980 4002 12020 4087
rect 11692 2500 11828 2540
rect 11307 2204 11349 2213
rect 11307 2164 11308 2204
rect 11348 2164 11349 2204
rect 11307 2155 11349 2164
rect 11211 1952 11253 1961
rect 11211 1912 11212 1952
rect 11252 1912 11253 1952
rect 11211 1903 11253 1912
rect 11308 1868 11348 2155
rect 11788 1868 11828 2500
rect 12268 2036 12308 4936
rect 12460 4817 12500 4936
rect 12556 4976 12596 5011
rect 12556 4925 12596 4936
rect 12459 4808 12501 4817
rect 12652 4808 12692 5188
rect 12843 5060 12885 5069
rect 12843 5020 12844 5060
rect 12884 5020 12885 5060
rect 12843 5011 12885 5020
rect 12940 5060 12980 5440
rect 12940 5011 12980 5020
rect 12747 4976 12789 4985
rect 12747 4936 12748 4976
rect 12788 4936 12789 4976
rect 12747 4927 12789 4936
rect 12844 4976 12884 5011
rect 13036 4985 13076 5070
rect 12748 4842 12788 4927
rect 12844 4925 12884 4936
rect 13035 4976 13077 4985
rect 13035 4936 13036 4976
rect 13076 4936 13077 4976
rect 13035 4927 13077 4936
rect 13228 4808 13268 7288
rect 13324 7001 13364 7876
rect 13420 7916 13460 7927
rect 13420 7841 13460 7876
rect 13419 7832 13461 7841
rect 13419 7792 13420 7832
rect 13460 7792 13461 7832
rect 13419 7783 13461 7792
rect 13323 6992 13365 7001
rect 13323 6952 13324 6992
rect 13364 6952 13365 6992
rect 13323 6943 13365 6952
rect 13324 6413 13364 6943
rect 13516 6497 13556 12916
rect 13707 12872 13749 12881
rect 13707 12832 13708 12872
rect 13748 12832 13749 12872
rect 13707 12823 13749 12832
rect 13708 12536 13748 12823
rect 13900 12620 13940 13243
rect 13708 12487 13748 12496
rect 13804 12580 13940 12620
rect 13611 12284 13653 12293
rect 13611 12244 13612 12284
rect 13652 12244 13653 12284
rect 13611 12235 13653 12244
rect 13612 11780 13652 12235
rect 13612 11731 13652 11740
rect 13708 11780 13748 11789
rect 13804 11780 13844 12580
rect 13748 11740 13844 11780
rect 13708 10613 13748 11740
rect 13803 11612 13845 11621
rect 13803 11572 13804 11612
rect 13844 11572 13845 11612
rect 13803 11563 13845 11572
rect 13707 10604 13749 10613
rect 13707 10564 13708 10604
rect 13748 10564 13749 10604
rect 13707 10555 13749 10564
rect 13707 10352 13749 10361
rect 13707 10312 13708 10352
rect 13748 10312 13749 10352
rect 13707 10303 13749 10312
rect 13708 10268 13748 10303
rect 13708 10217 13748 10228
rect 13804 10184 13844 11563
rect 13611 9512 13653 9521
rect 13611 9472 13612 9512
rect 13652 9472 13653 9512
rect 13611 9463 13653 9472
rect 13612 9378 13652 9463
rect 13707 9260 13749 9269
rect 13707 9220 13708 9260
rect 13748 9220 13749 9260
rect 13707 9211 13749 9220
rect 13611 8252 13653 8261
rect 13611 8212 13612 8252
rect 13652 8212 13653 8252
rect 13611 8203 13653 8212
rect 13612 7169 13652 8203
rect 13611 7160 13653 7169
rect 13611 7120 13612 7160
rect 13652 7120 13653 7160
rect 13611 7111 13653 7120
rect 13611 6908 13653 6917
rect 13611 6868 13612 6908
rect 13652 6868 13653 6908
rect 13611 6859 13653 6868
rect 13515 6488 13557 6497
rect 13515 6448 13516 6488
rect 13556 6448 13557 6488
rect 13515 6439 13557 6448
rect 13612 6488 13652 6859
rect 13612 6439 13652 6448
rect 13323 6404 13365 6413
rect 13323 6364 13324 6404
rect 13364 6364 13365 6404
rect 13323 6355 13365 6364
rect 13708 6236 13748 9211
rect 13804 7841 13844 10144
rect 13996 10109 14036 14008
rect 14092 12293 14132 14092
rect 14187 14092 14188 14132
rect 14228 14092 14229 14132
rect 14187 14083 14229 14092
rect 14187 13376 14229 13385
rect 14187 13336 14188 13376
rect 14228 13336 14229 13376
rect 14187 13327 14229 13336
rect 14091 12284 14133 12293
rect 14091 12244 14092 12284
rect 14132 12244 14133 12284
rect 14091 12235 14133 12244
rect 14188 11696 14228 13327
rect 14284 13040 14324 15100
rect 14380 14804 14420 19627
rect 14572 19256 14612 21568
rect 14572 18929 14612 19216
rect 14571 18920 14613 18929
rect 14571 18880 14572 18920
rect 14612 18880 14613 18920
rect 14571 18871 14613 18880
rect 14668 17828 14708 25591
rect 14764 20777 14804 27607
rect 14763 20768 14805 20777
rect 14763 20728 14764 20768
rect 14804 20728 14805 20768
rect 14763 20719 14805 20728
rect 14763 20600 14805 20609
rect 14763 20560 14764 20600
rect 14804 20560 14805 20600
rect 14763 20551 14805 20560
rect 14572 17788 14708 17828
rect 14572 16997 14612 17788
rect 14764 17744 14804 20551
rect 14860 18341 14900 31807
rect 15052 31604 15092 32068
rect 15148 32058 15188 32143
rect 15052 31564 15188 31604
rect 14955 31520 14997 31529
rect 14955 31480 14956 31520
rect 14996 31480 15092 31520
rect 14955 31471 14997 31480
rect 14956 31386 14996 31471
rect 15052 30932 15092 31480
rect 15148 31352 15188 31564
rect 15244 31529 15284 32824
rect 15436 32696 15476 32705
rect 15339 32360 15381 32369
rect 15339 32320 15340 32360
rect 15380 32320 15381 32360
rect 15339 32311 15381 32320
rect 15340 32192 15380 32311
rect 15436 32201 15476 32656
rect 15340 32143 15380 32152
rect 15435 32192 15477 32201
rect 15435 32152 15436 32192
rect 15476 32152 15477 32192
rect 15435 32143 15477 32152
rect 15243 31520 15285 31529
rect 15628 31520 15668 31529
rect 15243 31480 15244 31520
rect 15284 31480 15285 31520
rect 15243 31471 15285 31480
rect 15436 31480 15628 31520
rect 15148 31303 15188 31312
rect 15244 31352 15284 31361
rect 15244 31193 15284 31312
rect 15436 31352 15476 31480
rect 15628 31471 15668 31480
rect 15628 31352 15668 31361
rect 15436 31303 15476 31312
rect 15532 31312 15628 31352
rect 15339 31268 15381 31277
rect 15339 31228 15340 31268
rect 15380 31228 15381 31268
rect 15339 31219 15381 31228
rect 15243 31184 15285 31193
rect 15243 31144 15244 31184
rect 15284 31144 15285 31184
rect 15243 31135 15285 31144
rect 15340 31134 15380 31219
rect 14956 30892 15284 30932
rect 14956 29840 14996 30892
rect 15147 30680 15189 30689
rect 15147 30640 15148 30680
rect 15188 30640 15189 30680
rect 15147 30631 15189 30640
rect 15244 30675 15284 30892
rect 15436 30848 15476 30857
rect 15532 30848 15572 31312
rect 15628 31303 15668 31312
rect 15724 30848 15764 32824
rect 15819 32192 15861 32201
rect 15819 32152 15820 32192
rect 15860 32152 15861 32192
rect 15819 32143 15861 32152
rect 15820 31352 15860 32143
rect 15915 32108 15957 32117
rect 15915 32068 15916 32108
rect 15956 32068 15957 32108
rect 15915 32059 15957 32068
rect 15820 31303 15860 31312
rect 15476 30808 15572 30848
rect 15628 30808 15764 30848
rect 15916 30848 15956 32059
rect 15436 30799 15476 30808
rect 15628 30764 15668 30808
rect 15916 30799 15956 30808
rect 15532 30724 15668 30764
rect 15532 30680 15572 30724
rect 15051 30512 15093 30521
rect 15051 30472 15052 30512
rect 15092 30472 15093 30512
rect 15051 30463 15093 30472
rect 14956 29791 14996 29800
rect 15052 28412 15092 30463
rect 15052 28363 15092 28372
rect 14955 28328 14997 28337
rect 14955 28288 14956 28328
rect 14996 28288 14997 28328
rect 14955 28279 14997 28288
rect 14956 26237 14996 28279
rect 15148 26312 15188 30631
rect 15244 30605 15284 30635
rect 15436 30640 15572 30680
rect 15724 30680 15764 30689
rect 15243 30596 15285 30605
rect 15243 30556 15244 30596
rect 15284 30556 15285 30596
rect 15243 30547 15285 30556
rect 15244 30511 15284 30547
rect 15243 30008 15285 30017
rect 15243 29968 15244 30008
rect 15284 29968 15285 30008
rect 15243 29959 15285 29968
rect 15244 29840 15284 29959
rect 15244 29791 15284 29800
rect 15339 29756 15381 29765
rect 15339 29716 15340 29756
rect 15380 29716 15381 29756
rect 15339 29707 15381 29716
rect 15340 29622 15380 29707
rect 15243 29588 15285 29597
rect 15243 29548 15244 29588
rect 15284 29548 15285 29588
rect 15243 29539 15285 29548
rect 15052 26272 15188 26312
rect 14955 26228 14997 26237
rect 14955 26188 14956 26228
rect 14996 26188 14997 26228
rect 14955 26179 14997 26188
rect 14955 25556 14997 25565
rect 14955 25516 14956 25556
rect 14996 25516 14997 25556
rect 14955 25507 14997 25516
rect 14956 25313 14996 25507
rect 14955 25304 14997 25313
rect 14955 25264 14956 25304
rect 14996 25264 14997 25304
rect 15052 25304 15092 26272
rect 15147 26144 15189 26153
rect 15147 26104 15148 26144
rect 15188 26104 15189 26144
rect 15147 26095 15189 26104
rect 15148 26010 15188 26095
rect 15244 25649 15284 29539
rect 15436 29000 15476 30640
rect 15628 30635 15668 30644
rect 15627 30556 15628 30605
rect 15668 30556 15669 30605
rect 15627 30547 15669 30556
rect 15628 30500 15668 30547
rect 15724 30521 15764 30640
rect 15820 30680 15860 30689
rect 15723 30512 15765 30521
rect 15723 30472 15724 30512
rect 15764 30472 15765 30512
rect 15723 30463 15765 30472
rect 15820 30269 15860 30640
rect 15819 30260 15861 30269
rect 15819 30220 15820 30260
rect 15860 30220 15861 30260
rect 15819 30211 15861 30220
rect 15723 30092 15765 30101
rect 15723 30052 15724 30092
rect 15764 30052 15765 30092
rect 15723 30043 15765 30052
rect 15628 30008 15668 30017
rect 15628 29849 15668 29968
rect 15627 29840 15669 29849
rect 15627 29800 15628 29840
rect 15668 29800 15669 29840
rect 15627 29791 15669 29800
rect 15724 29168 15764 30043
rect 15820 29840 15860 30211
rect 15820 29791 15860 29800
rect 15915 29840 15957 29849
rect 15915 29800 15916 29840
rect 15956 29800 15957 29840
rect 15915 29791 15957 29800
rect 15916 29706 15956 29791
rect 15819 29672 15861 29681
rect 15819 29632 15820 29672
rect 15860 29632 15861 29672
rect 15819 29623 15861 29632
rect 15724 29000 15764 29128
rect 15340 28960 15476 29000
rect 15628 28960 15764 29000
rect 15243 25640 15285 25649
rect 15243 25600 15244 25640
rect 15284 25600 15285 25640
rect 15243 25591 15285 25600
rect 15147 25556 15189 25565
rect 15147 25516 15148 25556
rect 15188 25516 15189 25556
rect 15147 25507 15189 25516
rect 15148 25422 15188 25507
rect 15340 25472 15380 28960
rect 15531 28916 15573 28925
rect 15531 28876 15532 28916
rect 15572 28876 15573 28916
rect 15531 28867 15573 28876
rect 15532 28328 15572 28867
rect 15532 28279 15572 28288
rect 15435 27992 15477 28001
rect 15435 27952 15436 27992
rect 15476 27952 15477 27992
rect 15435 27943 15477 27952
rect 15436 26816 15476 27943
rect 15628 27824 15668 28960
rect 15532 27784 15668 27824
rect 15532 27665 15572 27784
rect 15531 27656 15573 27665
rect 15531 27616 15532 27656
rect 15572 27616 15573 27656
rect 15531 27607 15573 27616
rect 15628 27656 15668 27667
rect 15628 27581 15668 27616
rect 15723 27656 15765 27665
rect 15723 27616 15724 27656
rect 15764 27616 15765 27656
rect 15723 27607 15765 27616
rect 15627 27572 15669 27581
rect 15627 27532 15628 27572
rect 15668 27532 15669 27572
rect 15627 27523 15669 27532
rect 15724 27522 15764 27607
rect 15820 26984 15860 29623
rect 16012 29000 16052 33328
rect 16107 33328 16108 33368
rect 16148 33328 16149 33368
rect 16107 33319 16149 33328
rect 16204 32957 16244 33655
rect 16203 32948 16245 32957
rect 16203 32908 16204 32948
rect 16244 32908 16245 32948
rect 16203 32899 16245 32908
rect 16204 32864 16244 32899
rect 16107 31940 16149 31949
rect 16107 31900 16108 31940
rect 16148 31900 16149 31940
rect 16107 31891 16149 31900
rect 16108 31352 16148 31891
rect 16204 31436 16244 32824
rect 16300 32369 16340 39115
rect 16396 35132 16436 46600
rect 16492 46472 16532 46481
rect 16492 44960 16532 46432
rect 16876 45884 16916 45893
rect 16916 45844 17012 45884
rect 16876 45835 16916 45844
rect 16779 45800 16821 45809
rect 16684 45786 16724 45795
rect 16779 45760 16780 45800
rect 16820 45760 16821 45800
rect 16779 45751 16821 45760
rect 16684 45212 16724 45746
rect 16684 45163 16724 45172
rect 16492 44885 16532 44920
rect 16491 44876 16533 44885
rect 16491 44836 16492 44876
rect 16532 44836 16533 44876
rect 16491 44827 16533 44836
rect 16780 44288 16820 45751
rect 16875 45212 16917 45221
rect 16875 45172 16876 45212
rect 16916 45172 16917 45212
rect 16875 45163 16917 45172
rect 16876 45078 16916 45163
rect 16972 45044 17012 45844
rect 17068 45800 17108 47776
rect 17068 45389 17108 45760
rect 17067 45380 17109 45389
rect 17067 45340 17068 45380
rect 17108 45340 17109 45380
rect 17067 45331 17109 45340
rect 17068 45044 17108 45053
rect 16972 45004 17068 45044
rect 17068 44995 17108 45004
rect 16780 37820 16820 44248
rect 17067 44288 17109 44297
rect 17067 44248 17068 44288
rect 17108 44248 17109 44288
rect 17067 44239 17109 44248
rect 17068 43448 17108 44239
rect 17164 44213 17204 50119
rect 17260 49748 17300 50455
rect 17356 50336 17396 52480
rect 17452 52471 17492 52480
rect 17451 52100 17493 52109
rect 17451 52060 17452 52100
rect 17492 52060 17493 52100
rect 17451 52051 17493 52060
rect 17452 52016 17492 52051
rect 17548 52025 17588 56344
rect 17740 56309 17780 59275
rect 17836 58157 17876 60460
rect 18028 60332 18068 63727
rect 18124 63272 18164 63904
rect 18220 63785 18260 63904
rect 18315 63944 18357 63953
rect 18315 63904 18316 63944
rect 18356 63904 18357 63944
rect 18315 63895 18357 63904
rect 18219 63776 18261 63785
rect 18219 63736 18220 63776
rect 18260 63736 18261 63776
rect 18219 63727 18261 63736
rect 18219 63356 18261 63365
rect 18219 63316 18220 63356
rect 18260 63316 18261 63356
rect 18219 63307 18261 63316
rect 18124 63223 18164 63232
rect 18124 63104 18164 63113
rect 18124 60509 18164 63064
rect 18220 63104 18260 63307
rect 18316 63113 18356 63895
rect 18412 63281 18452 64240
rect 18508 64240 18644 64280
rect 18411 63272 18453 63281
rect 18411 63232 18412 63272
rect 18452 63232 18453 63272
rect 18411 63223 18453 63232
rect 18220 63055 18260 63064
rect 18315 63104 18357 63113
rect 18412 63104 18452 63113
rect 18315 63064 18316 63104
rect 18356 63064 18412 63104
rect 18315 63055 18357 63064
rect 18412 63055 18452 63064
rect 18316 62970 18356 63055
rect 18220 60920 18260 60929
rect 18220 60761 18260 60880
rect 18219 60752 18261 60761
rect 18219 60712 18220 60752
rect 18260 60712 18261 60752
rect 18219 60703 18261 60712
rect 18123 60500 18165 60509
rect 18123 60460 18124 60500
rect 18164 60460 18165 60500
rect 18123 60451 18165 60460
rect 18028 60292 18164 60332
rect 18028 60080 18068 60089
rect 18028 59324 18068 60040
rect 18124 60080 18164 60292
rect 18124 59333 18164 60040
rect 17932 59284 18028 59324
rect 17835 58148 17877 58157
rect 17835 58108 17836 58148
rect 17876 58108 17877 58148
rect 17835 58099 17877 58108
rect 17835 57140 17877 57149
rect 17835 57100 17836 57140
rect 17876 57100 17877 57140
rect 17835 57091 17877 57100
rect 17836 57056 17876 57091
rect 17836 57005 17876 57016
rect 17932 56981 17972 59284
rect 18028 59275 18068 59284
rect 18123 59324 18165 59333
rect 18123 59284 18124 59324
rect 18164 59284 18165 59324
rect 18123 59275 18165 59284
rect 18124 59190 18164 59275
rect 18027 59156 18069 59165
rect 18027 59116 18028 59156
rect 18068 59116 18069 59156
rect 18027 59107 18069 59116
rect 18028 58568 18068 59107
rect 18220 58904 18260 60703
rect 18315 60416 18357 60425
rect 18315 60376 18316 60416
rect 18356 60376 18357 60416
rect 18315 60367 18357 60376
rect 18316 59249 18356 60367
rect 18315 59240 18357 59249
rect 18315 59200 18316 59240
rect 18356 59200 18357 59240
rect 18315 59191 18357 59200
rect 18028 58519 18068 58528
rect 18124 58864 18260 58904
rect 18124 58316 18164 58864
rect 18412 58568 18452 58577
rect 18220 58400 18260 58409
rect 18260 58360 18356 58400
rect 18220 58351 18260 58360
rect 18028 58276 18164 58316
rect 17931 56972 17973 56981
rect 17931 56932 17932 56972
rect 17972 56932 17973 56972
rect 17931 56923 17973 56932
rect 17835 56888 17877 56897
rect 17835 56848 17836 56888
rect 17876 56848 17877 56888
rect 17835 56839 17877 56848
rect 17739 56300 17781 56309
rect 17739 56260 17740 56300
rect 17780 56260 17781 56300
rect 17739 56251 17781 56260
rect 17836 55460 17876 56839
rect 17932 56384 17972 56923
rect 18028 56897 18068 58276
rect 18219 58232 18261 58241
rect 18219 58192 18220 58232
rect 18260 58192 18261 58232
rect 18219 58183 18261 58192
rect 18123 58148 18165 58157
rect 18123 58108 18124 58148
rect 18164 58108 18165 58148
rect 18123 58099 18165 58108
rect 18027 56888 18069 56897
rect 18027 56848 18028 56888
rect 18068 56848 18069 56888
rect 18027 56839 18069 56848
rect 17932 56335 17972 56344
rect 18027 56300 18069 56309
rect 18027 56260 18028 56300
rect 18068 56260 18069 56300
rect 18027 56251 18069 56260
rect 18028 56166 18068 56251
rect 18124 56225 18164 58099
rect 18123 56216 18165 56225
rect 18123 56176 18124 56216
rect 18164 56176 18165 56216
rect 18123 56167 18165 56176
rect 18124 55553 18164 55638
rect 18123 55544 18165 55553
rect 18123 55504 18124 55544
rect 18164 55504 18165 55544
rect 18123 55495 18165 55504
rect 17740 55420 17876 55460
rect 17643 55124 17685 55133
rect 17643 55084 17644 55124
rect 17684 55084 17685 55124
rect 17643 55075 17685 55084
rect 17644 54545 17684 55075
rect 17643 54536 17685 54545
rect 17643 54496 17644 54536
rect 17684 54496 17685 54536
rect 17643 54487 17685 54496
rect 17740 54032 17780 55420
rect 17931 54956 17973 54965
rect 17931 54916 17932 54956
rect 17972 54916 17973 54956
rect 17931 54907 17973 54916
rect 17932 54872 17972 54907
rect 17932 54821 17972 54832
rect 17836 54788 17876 54797
rect 17836 54200 17876 54748
rect 17836 54160 18068 54200
rect 17836 54032 17876 54041
rect 17740 53992 17836 54032
rect 17452 51965 17492 51976
rect 17547 52016 17589 52025
rect 17547 51976 17548 52016
rect 17588 51976 17589 52016
rect 17547 51967 17589 51976
rect 17739 51848 17781 51857
rect 17739 51808 17740 51848
rect 17780 51808 17781 51848
rect 17739 51799 17781 51808
rect 17643 51260 17685 51269
rect 17643 51220 17644 51260
rect 17684 51220 17685 51260
rect 17643 51211 17685 51220
rect 17644 51126 17684 51211
rect 17451 51008 17493 51017
rect 17451 50968 17452 51008
rect 17492 50968 17493 51008
rect 17451 50959 17493 50968
rect 17452 50874 17492 50959
rect 17547 50504 17589 50513
rect 17547 50464 17548 50504
rect 17588 50464 17589 50504
rect 17547 50455 17589 50464
rect 17451 50420 17493 50429
rect 17451 50380 17452 50420
rect 17492 50380 17493 50420
rect 17451 50371 17493 50380
rect 17355 50296 17396 50336
rect 17355 50252 17395 50296
rect 17355 50212 17396 50252
rect 17260 49699 17300 49708
rect 17356 49328 17396 50212
rect 17452 49496 17492 50371
rect 17548 50336 17588 50455
rect 17548 50287 17588 50296
rect 17644 50336 17684 50345
rect 17547 50084 17589 50093
rect 17547 50044 17548 50084
rect 17588 50044 17589 50084
rect 17547 50035 17589 50044
rect 17452 49447 17492 49456
rect 17260 49288 17396 49328
rect 17260 47321 17300 49288
rect 17355 49160 17397 49169
rect 17355 49120 17356 49160
rect 17396 49120 17397 49160
rect 17355 49111 17397 49120
rect 17259 47312 17301 47321
rect 17259 47272 17260 47312
rect 17300 47272 17301 47312
rect 17259 47263 17301 47272
rect 17260 44274 17300 44283
rect 17163 44204 17205 44213
rect 17163 44164 17164 44204
rect 17204 44164 17205 44204
rect 17163 44155 17205 44164
rect 17260 43700 17300 44234
rect 17260 43651 17300 43660
rect 17068 43399 17108 43408
rect 16971 42440 17013 42449
rect 16971 42400 16972 42440
rect 17012 42400 17013 42440
rect 16971 42391 17013 42400
rect 16972 42020 17012 42391
rect 17163 42188 17205 42197
rect 17163 42148 17164 42188
rect 17204 42148 17205 42188
rect 17163 42139 17205 42148
rect 17164 42054 17204 42139
rect 16972 41971 17012 41980
rect 16780 37780 16916 37820
rect 16396 35083 16436 35092
rect 16587 34964 16629 34973
rect 16587 34924 16588 34964
rect 16628 34924 16629 34964
rect 16587 34915 16629 34924
rect 16588 34830 16628 34915
rect 16491 33536 16533 33545
rect 16491 33496 16492 33536
rect 16532 33496 16533 33536
rect 16491 33487 16533 33496
rect 16299 32360 16341 32369
rect 16299 32320 16300 32360
rect 16340 32320 16341 32360
rect 16299 32311 16341 32320
rect 16204 31396 16340 31436
rect 16108 31303 16148 31312
rect 16204 31332 16244 31341
rect 16107 31184 16149 31193
rect 16107 31144 16108 31184
rect 16148 31144 16149 31184
rect 16107 31135 16149 31144
rect 16108 29672 16148 31135
rect 16204 31109 16244 31292
rect 16203 31100 16245 31109
rect 16203 31060 16204 31100
rect 16244 31060 16245 31100
rect 16203 31051 16245 31060
rect 16204 30269 16244 31051
rect 16203 30260 16245 30269
rect 16203 30220 16204 30260
rect 16244 30220 16245 30260
rect 16203 30211 16245 30220
rect 16108 29623 16148 29632
rect 16300 29597 16340 31396
rect 16492 30680 16532 33487
rect 16587 32696 16629 32705
rect 16587 32656 16588 32696
rect 16628 32656 16629 32696
rect 16587 32647 16629 32656
rect 16588 32192 16628 32647
rect 16588 32143 16628 32152
rect 16779 31940 16821 31949
rect 16779 31900 16780 31940
rect 16820 31900 16821 31940
rect 16779 31891 16821 31900
rect 16780 31806 16820 31891
rect 16588 31352 16628 31361
rect 16588 31025 16628 31312
rect 16684 31352 16724 31361
rect 16587 31016 16629 31025
rect 16587 30976 16588 31016
rect 16628 30976 16629 31016
rect 16587 30967 16629 30976
rect 16299 29588 16341 29597
rect 16299 29548 16300 29588
rect 16340 29548 16341 29588
rect 16299 29539 16341 29548
rect 16492 29429 16532 30640
rect 16588 30521 16628 30967
rect 16587 30512 16629 30521
rect 16587 30472 16588 30512
rect 16628 30472 16629 30512
rect 16587 30463 16629 30472
rect 16684 29933 16724 31312
rect 16683 29924 16725 29933
rect 16683 29884 16684 29924
rect 16724 29884 16725 29924
rect 16683 29875 16725 29884
rect 16491 29420 16533 29429
rect 16491 29380 16492 29420
rect 16532 29380 16533 29420
rect 16491 29371 16533 29380
rect 16299 29336 16341 29345
rect 16299 29296 16300 29336
rect 16340 29296 16341 29336
rect 16299 29287 16341 29296
rect 16683 29336 16725 29345
rect 16683 29296 16684 29336
rect 16724 29296 16725 29336
rect 16300 29202 16340 29287
rect 16492 29261 16532 29292
rect 16683 29287 16725 29296
rect 16491 29252 16533 29261
rect 16491 29212 16492 29252
rect 16532 29212 16533 29252
rect 16491 29203 16533 29212
rect 16204 29168 16244 29177
rect 16204 29000 16244 29128
rect 16396 29168 16436 29179
rect 16396 29093 16436 29128
rect 16492 29168 16532 29203
rect 16395 29084 16437 29093
rect 16395 29044 16396 29084
rect 16436 29044 16437 29084
rect 16395 29035 16437 29044
rect 16012 28960 16148 29000
rect 16204 28960 16340 29000
rect 15916 28916 15956 28925
rect 15956 28876 16052 28916
rect 15916 28867 15956 28876
rect 16012 28342 16052 28876
rect 16012 28293 16052 28302
rect 15916 27656 15956 27667
rect 15916 27581 15956 27616
rect 15915 27572 15957 27581
rect 15915 27532 15916 27572
rect 15956 27532 15957 27572
rect 15915 27523 15957 27532
rect 16108 26993 16148 28960
rect 16204 28160 16244 28169
rect 16204 27749 16244 28120
rect 16203 27740 16245 27749
rect 16203 27700 16204 27740
rect 16244 27700 16245 27740
rect 16203 27691 16245 27700
rect 15436 26153 15476 26776
rect 15532 26944 15860 26984
rect 16107 26984 16149 26993
rect 16107 26944 16108 26984
rect 16148 26944 16149 26984
rect 15435 26144 15477 26153
rect 15435 26104 15436 26144
rect 15476 26104 15477 26144
rect 15435 26095 15477 26104
rect 15244 25432 15380 25472
rect 15148 25304 15188 25313
rect 15052 25264 15148 25304
rect 14955 25255 14997 25264
rect 14956 25170 14996 25255
rect 14955 24632 14997 24641
rect 14955 24592 14956 24632
rect 14996 24592 14997 24632
rect 14955 24583 14997 24592
rect 14956 23465 14996 24583
rect 15148 24305 15188 25264
rect 15147 24296 15189 24305
rect 15147 24256 15148 24296
rect 15188 24256 15189 24296
rect 15147 24247 15189 24256
rect 15052 23801 15092 23887
rect 15244 23876 15284 25432
rect 15339 25304 15381 25313
rect 15339 25264 15340 25304
rect 15380 25264 15381 25304
rect 15339 25255 15381 25264
rect 15340 25170 15380 25255
rect 15436 25229 15476 26095
rect 15532 25304 15572 26944
rect 16107 26935 16149 26944
rect 15820 26816 15860 26825
rect 15628 26732 15668 26741
rect 15820 26732 15860 26776
rect 15668 26692 15860 26732
rect 16012 26816 16052 26825
rect 15628 26139 15668 26692
rect 15915 26648 15957 26657
rect 15915 26608 15916 26648
rect 15956 26608 15957 26648
rect 15915 26599 15957 26608
rect 15916 26514 15956 26599
rect 15819 26228 15861 26237
rect 15819 26188 15820 26228
rect 15860 26188 15861 26228
rect 15819 26179 15861 26188
rect 15628 26090 15668 26099
rect 15820 26094 15860 26179
rect 16012 26060 16052 26776
rect 15916 26020 16052 26060
rect 16108 26816 16148 26825
rect 15628 25556 15668 25565
rect 15916 25556 15956 26020
rect 16011 25892 16053 25901
rect 16011 25852 16012 25892
rect 16052 25852 16053 25892
rect 16011 25843 16053 25852
rect 16012 25758 16052 25843
rect 16108 25565 16148 26776
rect 16204 26153 16244 26238
rect 16203 26144 16245 26153
rect 16203 26104 16204 26144
rect 16244 26104 16245 26144
rect 16203 26095 16245 26104
rect 16300 25976 16340 28960
rect 16396 28580 16436 28589
rect 16492 28580 16532 29128
rect 16684 29168 16724 29287
rect 16684 29119 16724 29128
rect 16779 29168 16821 29177
rect 16779 29128 16780 29168
rect 16820 29128 16821 29168
rect 16779 29119 16821 29128
rect 16780 29034 16820 29119
rect 16683 28916 16725 28925
rect 16683 28876 16684 28916
rect 16724 28876 16725 28916
rect 16683 28867 16725 28876
rect 16684 28782 16724 28867
rect 16436 28540 16532 28580
rect 16396 28531 16436 28540
rect 16588 28328 16628 28337
rect 16588 27497 16628 28288
rect 16587 27488 16629 27497
rect 16587 27448 16588 27488
rect 16628 27448 16629 27488
rect 16587 27439 16629 27448
rect 16587 26984 16629 26993
rect 16587 26944 16588 26984
rect 16628 26944 16629 26984
rect 16587 26935 16629 26944
rect 16204 25936 16340 25976
rect 15668 25516 15956 25556
rect 16107 25556 16149 25565
rect 16107 25516 16108 25556
rect 16148 25516 16149 25556
rect 15628 25507 15668 25516
rect 16107 25507 16149 25516
rect 15628 25304 15668 25313
rect 15916 25304 15956 25313
rect 15532 25264 15628 25304
rect 15435 25220 15477 25229
rect 15435 25180 15436 25220
rect 15476 25180 15477 25220
rect 15435 25171 15477 25180
rect 15628 24800 15668 25264
rect 15436 24760 15668 24800
rect 15820 25264 15916 25304
rect 15340 24641 15380 24726
rect 15339 24632 15381 24641
rect 15339 24592 15340 24632
rect 15380 24592 15381 24632
rect 15339 24583 15381 24592
rect 15148 23836 15284 23876
rect 15051 23797 15093 23801
rect 15051 23752 15052 23797
rect 15092 23752 15093 23797
rect 15051 23743 15093 23752
rect 14955 23456 14997 23465
rect 14955 23416 14956 23456
rect 14996 23416 14997 23456
rect 14955 23407 14997 23416
rect 15148 22952 15188 23836
rect 15243 23708 15285 23717
rect 15243 23668 15244 23708
rect 15284 23668 15285 23708
rect 15243 23659 15285 23668
rect 15244 23574 15284 23659
rect 15436 23624 15476 24760
rect 15531 24296 15573 24305
rect 15531 24256 15532 24296
rect 15572 24256 15573 24296
rect 15531 24247 15573 24256
rect 15532 23876 15572 24247
rect 15628 24053 15668 24138
rect 15627 24044 15669 24053
rect 15627 24004 15628 24044
rect 15668 24004 15669 24044
rect 15627 23995 15669 24004
rect 15723 23876 15765 23885
rect 15532 23836 15668 23876
rect 15532 23781 15572 23790
rect 15532 23717 15572 23741
rect 15531 23708 15573 23717
rect 15531 23668 15532 23708
rect 15572 23668 15573 23708
rect 15531 23659 15573 23668
rect 15532 23646 15572 23659
rect 15340 23584 15476 23624
rect 15243 23456 15285 23465
rect 15243 23416 15244 23456
rect 15284 23416 15285 23456
rect 15243 23407 15285 23416
rect 15244 23213 15284 23407
rect 15243 23204 15285 23213
rect 15243 23164 15244 23204
rect 15284 23164 15285 23204
rect 15243 23155 15285 23164
rect 15244 23120 15284 23155
rect 15244 23070 15284 23080
rect 15148 22912 15284 22952
rect 14956 22280 14996 22289
rect 14956 21701 14996 22240
rect 15148 22112 15188 22121
rect 14955 21692 14997 21701
rect 14955 21652 14956 21692
rect 14996 21652 14997 21692
rect 14955 21643 14997 21652
rect 15148 21608 15188 22072
rect 15244 21776 15284 22912
rect 15244 21727 15284 21736
rect 15100 21598 15188 21608
rect 15140 21568 15188 21598
rect 15100 21549 15140 21558
rect 14955 20768 14997 20777
rect 14955 20728 14956 20768
rect 14996 20728 14997 20768
rect 14955 20719 14997 20728
rect 14956 18584 14996 20719
rect 15340 20180 15380 23584
rect 15531 23456 15573 23465
rect 15531 23416 15532 23456
rect 15572 23416 15573 23456
rect 15531 23407 15573 23416
rect 15435 23288 15477 23297
rect 15435 23248 15436 23288
rect 15476 23248 15477 23288
rect 15435 23239 15477 23248
rect 15436 23154 15476 23239
rect 15532 23129 15572 23407
rect 15531 23120 15573 23129
rect 15531 23080 15532 23120
rect 15572 23080 15573 23120
rect 15531 23071 15573 23080
rect 15435 23036 15477 23045
rect 15435 22996 15436 23036
rect 15476 22996 15477 23036
rect 15435 22987 15477 22996
rect 15436 21365 15476 22987
rect 15531 22952 15573 22961
rect 15531 22912 15532 22952
rect 15572 22912 15573 22952
rect 15531 22903 15573 22912
rect 15435 21356 15477 21365
rect 15435 21316 15436 21356
rect 15476 21316 15477 21356
rect 15435 21307 15477 21316
rect 15532 20936 15572 22903
rect 15628 22793 15668 23836
rect 15723 23836 15724 23876
rect 15764 23836 15765 23876
rect 15723 23827 15765 23836
rect 15724 23120 15764 23827
rect 15820 23801 15860 25264
rect 15916 25255 15956 25264
rect 16012 25304 16052 25313
rect 16012 24044 16052 25264
rect 16108 25304 16148 25313
rect 16108 24809 16148 25264
rect 16107 24800 16149 24809
rect 16107 24760 16108 24800
rect 16148 24760 16149 24800
rect 16107 24751 16149 24760
rect 16012 24004 16148 24044
rect 15915 23876 15957 23885
rect 15915 23836 15916 23876
rect 15956 23836 15957 23876
rect 15915 23827 15957 23836
rect 15819 23792 15861 23801
rect 15819 23752 15820 23792
rect 15860 23752 15861 23792
rect 15819 23743 15861 23752
rect 15916 23792 15956 23827
rect 15820 23297 15860 23743
rect 15916 23741 15956 23752
rect 16012 23792 16052 23801
rect 15819 23288 15861 23297
rect 16012 23288 16052 23752
rect 16108 23633 16148 24004
rect 16107 23624 16149 23633
rect 16107 23584 16108 23624
rect 16148 23584 16149 23624
rect 16107 23575 16149 23584
rect 16107 23456 16149 23465
rect 16107 23416 16108 23456
rect 16148 23416 16149 23456
rect 16107 23407 16149 23416
rect 15819 23248 15820 23288
rect 15860 23248 15861 23288
rect 15819 23239 15861 23248
rect 15916 23248 16052 23288
rect 15724 23071 15764 23080
rect 15916 22952 15956 23248
rect 16108 23204 16148 23407
rect 16012 23164 16148 23204
rect 16012 23147 16052 23164
rect 16012 23098 16052 23107
rect 16108 23078 16148 23087
rect 16108 23036 16148 23038
rect 15724 22912 15956 22952
rect 16012 22996 16148 23036
rect 15627 22784 15669 22793
rect 15627 22744 15628 22784
rect 15668 22744 15669 22784
rect 15627 22735 15669 22744
rect 15724 21617 15764 22912
rect 15915 22784 15957 22793
rect 15915 22744 15916 22784
rect 15956 22744 15957 22784
rect 15915 22735 15957 22744
rect 15628 21608 15668 21617
rect 15628 21020 15668 21568
rect 15723 21608 15765 21617
rect 15723 21568 15724 21608
rect 15764 21568 15765 21608
rect 15723 21559 15765 21568
rect 15724 21474 15764 21559
rect 15820 21020 15860 21029
rect 15628 20980 15820 21020
rect 15532 20896 15764 20936
rect 15627 20768 15669 20777
rect 15627 20728 15628 20768
rect 15668 20728 15669 20768
rect 15627 20719 15669 20728
rect 15628 20634 15668 20719
rect 15340 20140 15476 20180
rect 15100 19265 15140 19274
rect 15140 19225 15188 19256
rect 15100 19216 15188 19225
rect 15148 18752 15188 19216
rect 15244 19088 15284 19097
rect 15284 19048 15380 19088
rect 15244 19039 15284 19048
rect 15244 18752 15284 18761
rect 15148 18712 15244 18752
rect 15244 18703 15284 18712
rect 15052 18584 15092 18593
rect 14956 18544 15052 18584
rect 14859 18332 14901 18341
rect 14859 18292 14860 18332
rect 14900 18292 14901 18332
rect 14859 18283 14901 18292
rect 14956 18173 14996 18544
rect 15052 18535 15092 18544
rect 15243 18332 15285 18341
rect 15243 18292 15244 18332
rect 15284 18292 15285 18332
rect 15243 18283 15285 18292
rect 14955 18164 14997 18173
rect 14955 18124 14956 18164
rect 14996 18124 14997 18164
rect 14955 18115 14997 18124
rect 14955 17996 14997 18005
rect 14955 17956 14956 17996
rect 14996 17956 14997 17996
rect 14955 17947 14997 17956
rect 14956 17862 14996 17947
rect 15244 17921 15284 18283
rect 15243 17912 15285 17921
rect 15243 17872 15244 17912
rect 15284 17872 15285 17912
rect 15243 17863 15285 17872
rect 15148 17744 15188 17753
rect 14804 17704 15092 17744
rect 14764 17695 14804 17704
rect 14667 17660 14709 17669
rect 14667 17620 14668 17660
rect 14708 17620 14709 17660
rect 14667 17611 14709 17620
rect 14571 16988 14613 16997
rect 14571 16948 14572 16988
rect 14612 16948 14613 16988
rect 14571 16939 14613 16948
rect 14571 16820 14613 16829
rect 14571 16780 14572 16820
rect 14612 16780 14613 16820
rect 14571 16771 14613 16780
rect 14476 16232 14516 16241
rect 14572 16232 14612 16771
rect 14668 16400 14708 17611
rect 14956 17576 14996 17585
rect 14956 17492 14996 17536
rect 14668 16351 14708 16360
rect 14764 17452 14996 17492
rect 14668 16232 14708 16241
rect 14572 16192 14668 16232
rect 14476 14888 14516 16192
rect 14668 16183 14708 16192
rect 14764 16232 14804 17452
rect 15052 17408 15092 17704
rect 15148 17585 15188 17704
rect 15244 17744 15284 17863
rect 15244 17695 15284 17704
rect 15147 17576 15189 17585
rect 15147 17536 15148 17576
rect 15188 17536 15189 17576
rect 15147 17527 15189 17536
rect 14860 17368 15092 17408
rect 14860 17072 14900 17368
rect 15052 17240 15092 17249
rect 15148 17240 15188 17527
rect 15092 17200 15188 17240
rect 15052 17191 15092 17200
rect 14860 16913 14900 17032
rect 15243 17072 15285 17081
rect 15243 17032 15244 17072
rect 15284 17032 15285 17072
rect 15243 17023 15285 17032
rect 14955 16988 14997 16997
rect 14955 16948 14956 16988
rect 14996 16948 14997 16988
rect 14955 16939 14997 16948
rect 14859 16904 14901 16913
rect 14859 16864 14860 16904
rect 14900 16864 14901 16904
rect 14859 16855 14901 16864
rect 14764 16183 14804 16192
rect 14956 16232 14996 16939
rect 15244 16938 15284 17023
rect 15051 16820 15093 16829
rect 15051 16780 15052 16820
rect 15092 16780 15093 16820
rect 15051 16771 15093 16780
rect 15052 16686 15092 16771
rect 15147 16484 15189 16493
rect 15147 16444 15148 16484
rect 15188 16444 15189 16484
rect 15147 16435 15189 16444
rect 14476 14848 14708 14888
rect 14380 14764 14612 14804
rect 14380 14636 14420 14764
rect 14572 14720 14612 14764
rect 14572 14671 14612 14680
rect 14380 14596 14516 14636
rect 14379 13376 14421 13385
rect 14379 13336 14380 13376
rect 14420 13336 14421 13376
rect 14379 13327 14421 13336
rect 14380 13208 14420 13327
rect 14380 13159 14420 13168
rect 14284 13000 14420 13040
rect 14188 11647 14228 11656
rect 14091 11528 14133 11537
rect 14091 11488 14092 11528
rect 14132 11488 14133 11528
rect 14091 11479 14133 11488
rect 13995 10100 14037 10109
rect 13995 10060 13996 10100
rect 14036 10060 14037 10100
rect 13995 10051 14037 10060
rect 13899 8084 13941 8093
rect 13899 8044 13900 8084
rect 13940 8044 13941 8084
rect 13899 8035 13941 8044
rect 13900 8000 13940 8035
rect 13900 7949 13940 7960
rect 13803 7832 13845 7841
rect 13803 7792 13804 7832
rect 13844 7792 13845 7832
rect 13803 7783 13845 7792
rect 13803 7160 13845 7169
rect 13803 7120 13804 7160
rect 13844 7120 13845 7160
rect 13803 7111 13845 7120
rect 12459 4768 12460 4808
rect 12500 4768 12501 4808
rect 12459 4759 12501 4768
rect 12556 4768 12692 4808
rect 12940 4768 13268 4808
rect 12363 4640 12405 4649
rect 12363 4600 12364 4640
rect 12404 4600 12405 4640
rect 12363 4591 12405 4600
rect 12364 3464 12404 4591
rect 12556 4145 12596 4768
rect 12555 4136 12597 4145
rect 12555 4096 12556 4136
rect 12596 4096 12597 4136
rect 12555 4087 12597 4096
rect 12940 4136 12980 4768
rect 13035 4556 13077 4565
rect 13035 4516 13036 4556
rect 13076 4516 13077 4556
rect 13035 4507 13077 4516
rect 12940 4087 12980 4096
rect 12556 3548 12596 3557
rect 12596 3508 12884 3548
rect 12556 3499 12596 3508
rect 12364 3389 12404 3424
rect 12844 3464 12884 3508
rect 12844 3415 12884 3424
rect 12940 3464 12980 3473
rect 12363 3380 12405 3389
rect 12363 3340 12364 3380
rect 12404 3340 12405 3380
rect 12363 3331 12405 3340
rect 12940 2960 12980 3424
rect 12844 2920 12980 2960
rect 12844 2381 12884 2920
rect 12939 2708 12981 2717
rect 12939 2668 12940 2708
rect 12980 2668 12981 2708
rect 12939 2659 12981 2668
rect 12940 2624 12980 2659
rect 12940 2573 12980 2584
rect 12843 2372 12885 2381
rect 12843 2332 12844 2372
rect 12884 2332 12885 2372
rect 12843 2323 12885 2332
rect 12172 1996 12308 2036
rect 11884 1868 11924 1877
rect 11788 1828 11884 1868
rect 11308 1819 11348 1828
rect 11884 1819 11924 1828
rect 11116 1700 11156 1709
rect 11116 1289 11156 1660
rect 11499 1700 11541 1709
rect 11499 1660 11500 1700
rect 11540 1660 11541 1700
rect 11499 1651 11541 1660
rect 11692 1700 11732 1709
rect 12076 1700 12116 1709
rect 11500 1566 11540 1651
rect 11692 1373 11732 1660
rect 11884 1660 12076 1700
rect 11691 1364 11733 1373
rect 11691 1324 11692 1364
rect 11732 1324 11733 1364
rect 11691 1315 11733 1324
rect 11115 1280 11157 1289
rect 11115 1240 11116 1280
rect 11156 1240 11157 1280
rect 11115 1231 11157 1240
rect 11884 1112 11924 1660
rect 12076 1651 12116 1660
rect 11979 1448 12021 1457
rect 12172 1448 12212 1996
rect 12267 1868 12309 1877
rect 12267 1828 12268 1868
rect 12308 1828 12309 1868
rect 12267 1819 12309 1828
rect 12268 1734 12308 1819
rect 12844 1793 12884 2323
rect 12939 1868 12981 1877
rect 12939 1828 12940 1868
rect 12980 1828 12981 1868
rect 12939 1819 12981 1828
rect 12843 1784 12885 1793
rect 12843 1744 12844 1784
rect 12884 1744 12885 1784
rect 12843 1735 12885 1744
rect 12940 1734 12980 1819
rect 12363 1700 12405 1709
rect 12363 1660 12364 1700
rect 12404 1660 12405 1700
rect 12363 1651 12405 1660
rect 12748 1700 12788 1709
rect 11979 1408 11980 1448
rect 12020 1408 12021 1448
rect 11979 1399 12021 1408
rect 12076 1408 12212 1448
rect 11404 1072 11924 1112
rect 11115 944 11157 953
rect 11115 904 11116 944
rect 11156 904 11157 944
rect 11115 895 11157 904
rect 11116 810 11156 895
rect 11211 776 11253 785
rect 11211 736 11212 776
rect 11252 736 11253 776
rect 11211 727 11253 736
rect 11212 80 11252 727
rect 11404 80 11444 1072
rect 11787 944 11829 953
rect 11787 904 11788 944
rect 11828 904 11829 944
rect 11787 895 11829 904
rect 11595 524 11637 533
rect 11595 484 11596 524
rect 11636 484 11637 524
rect 11595 475 11637 484
rect 11596 80 11636 475
rect 11788 80 11828 895
rect 11980 80 12020 1399
rect 12076 281 12116 1408
rect 12171 1280 12213 1289
rect 12171 1240 12172 1280
rect 12212 1240 12213 1280
rect 12171 1231 12213 1240
rect 12075 272 12117 281
rect 12075 232 12076 272
rect 12116 232 12117 272
rect 12075 223 12117 232
rect 12172 80 12212 1231
rect 12364 80 12404 1651
rect 12748 1541 12788 1660
rect 13036 1616 13076 4507
rect 13131 4472 13173 4481
rect 13131 4432 13132 4472
rect 13172 4432 13173 4472
rect 13131 4423 13173 4432
rect 12940 1576 13076 1616
rect 12747 1532 12789 1541
rect 12747 1492 12748 1532
rect 12788 1492 12789 1532
rect 12747 1483 12789 1492
rect 12747 1280 12789 1289
rect 12747 1240 12748 1280
rect 12788 1240 12789 1280
rect 12747 1231 12789 1240
rect 12555 1112 12597 1121
rect 12555 1072 12556 1112
rect 12596 1072 12597 1112
rect 12555 1063 12597 1072
rect 12556 80 12596 1063
rect 12748 80 12788 1231
rect 12940 80 12980 1576
rect 13132 80 13172 4423
rect 13228 3137 13268 4768
rect 13324 6196 13748 6236
rect 13324 3464 13364 6196
rect 13804 5153 13844 7111
rect 13899 6404 13941 6413
rect 13899 6364 13900 6404
rect 13940 6364 13941 6404
rect 13899 6355 13941 6364
rect 13803 5144 13845 5153
rect 13708 5104 13804 5144
rect 13844 5104 13845 5144
rect 13708 4733 13748 5104
rect 13803 5095 13845 5104
rect 13803 4976 13845 4985
rect 13803 4936 13804 4976
rect 13844 4936 13845 4976
rect 13803 4927 13845 4936
rect 13707 4724 13749 4733
rect 13707 4684 13708 4724
rect 13748 4684 13749 4724
rect 13707 4675 13749 4684
rect 13707 4136 13749 4145
rect 13707 4096 13708 4136
rect 13748 4096 13749 4136
rect 13707 4087 13749 4096
rect 13324 3415 13364 3424
rect 13419 3464 13461 3473
rect 13419 3424 13420 3464
rect 13460 3424 13461 3464
rect 13419 3415 13461 3424
rect 13420 3330 13460 3415
rect 13227 3128 13269 3137
rect 13227 3088 13228 3128
rect 13268 3088 13269 3128
rect 13227 3079 13269 3088
rect 13228 2717 13268 3079
rect 13227 2708 13269 2717
rect 13227 2668 13228 2708
rect 13268 2668 13269 2708
rect 13227 2659 13269 2668
rect 13227 2540 13269 2549
rect 13227 2500 13228 2540
rect 13268 2500 13269 2540
rect 13227 2491 13269 2500
rect 13228 1868 13268 2491
rect 13708 2381 13748 4087
rect 13804 3641 13844 4927
rect 13803 3632 13845 3641
rect 13803 3592 13804 3632
rect 13844 3592 13845 3632
rect 13803 3583 13845 3592
rect 13900 3464 13940 6355
rect 13900 3415 13940 3424
rect 13996 2969 14036 10051
rect 14092 7757 14132 11479
rect 14380 11201 14420 13000
rect 14379 11192 14421 11201
rect 14379 11152 14380 11192
rect 14420 11152 14421 11192
rect 14379 11143 14421 11152
rect 14379 11024 14421 11033
rect 14379 10984 14380 11024
rect 14420 10984 14421 11024
rect 14379 10975 14421 10984
rect 14187 10940 14229 10949
rect 14187 10900 14188 10940
rect 14228 10900 14229 10940
rect 14187 10891 14229 10900
rect 14188 9689 14228 10891
rect 14283 10520 14325 10529
rect 14283 10480 14284 10520
rect 14324 10480 14325 10520
rect 14283 10471 14325 10480
rect 14284 10193 14324 10471
rect 14283 10184 14325 10193
rect 14283 10144 14284 10184
rect 14324 10144 14325 10184
rect 14283 10135 14325 10144
rect 14284 10050 14324 10135
rect 14187 9680 14229 9689
rect 14187 9640 14188 9680
rect 14228 9640 14229 9680
rect 14187 9631 14229 9640
rect 14188 8849 14228 9631
rect 14187 8840 14229 8849
rect 14380 8840 14420 10975
rect 14187 8800 14188 8840
rect 14228 8800 14229 8840
rect 14187 8791 14229 8800
rect 14284 8800 14420 8840
rect 14188 8672 14228 8791
rect 14188 8623 14228 8632
rect 14284 7832 14324 8800
rect 14476 8093 14516 14596
rect 14571 14552 14613 14561
rect 14571 14512 14572 14552
rect 14612 14512 14613 14552
rect 14571 14503 14613 14512
rect 14572 9521 14612 14503
rect 14668 13805 14708 14848
rect 14956 14561 14996 16192
rect 15051 15308 15093 15317
rect 15051 15268 15052 15308
rect 15092 15268 15093 15308
rect 15051 15259 15093 15268
rect 15052 14734 15092 15259
rect 15052 14685 15092 14694
rect 14955 14552 14997 14561
rect 14955 14512 14956 14552
rect 14996 14512 14997 14552
rect 14955 14503 14997 14512
rect 15148 14048 15188 16435
rect 15243 15392 15285 15401
rect 15243 15352 15244 15392
rect 15284 15352 15285 15392
rect 15243 15343 15285 15352
rect 15244 14636 15284 15343
rect 15244 14587 15284 14596
rect 15340 14384 15380 19048
rect 15436 18845 15476 20140
rect 15628 20096 15668 20105
rect 15628 19601 15668 20056
rect 15627 19592 15669 19601
rect 15627 19552 15628 19592
rect 15668 19552 15669 19592
rect 15627 19543 15669 19552
rect 15724 19013 15764 20896
rect 15820 20777 15860 20980
rect 15819 20768 15861 20777
rect 15819 20728 15820 20768
rect 15860 20728 15861 20768
rect 15819 20719 15861 20728
rect 15819 19844 15861 19853
rect 15819 19804 15820 19844
rect 15860 19804 15861 19844
rect 15819 19795 15861 19804
rect 15723 19004 15765 19013
rect 15723 18964 15724 19004
rect 15764 18964 15765 19004
rect 15723 18955 15765 18964
rect 15627 18920 15669 18929
rect 15627 18880 15628 18920
rect 15668 18880 15669 18920
rect 15627 18871 15669 18880
rect 15435 18836 15477 18845
rect 15435 18796 15436 18836
rect 15476 18796 15477 18836
rect 15435 18787 15477 18796
rect 15628 18752 15668 18871
rect 15724 18752 15764 18761
rect 15628 18712 15724 18752
rect 15724 18703 15764 18712
rect 15436 18584 15476 18593
rect 15724 18584 15764 18593
rect 15436 17837 15476 18544
rect 15532 18569 15572 18578
rect 15435 17828 15477 17837
rect 15435 17788 15436 17828
rect 15476 17788 15477 17828
rect 15435 17779 15477 17788
rect 15532 17660 15572 18529
rect 15627 18248 15669 18257
rect 15627 18208 15628 18248
rect 15668 18208 15669 18248
rect 15627 18199 15669 18208
rect 15628 17744 15668 18199
rect 15724 18005 15764 18544
rect 15820 18584 15860 19795
rect 15916 18761 15956 22735
rect 16012 22121 16052 22996
rect 16107 22868 16149 22877
rect 16107 22828 16108 22868
rect 16148 22828 16149 22868
rect 16204 22868 16244 25936
rect 16299 25472 16341 25481
rect 16299 25432 16300 25472
rect 16340 25432 16341 25472
rect 16299 25423 16341 25432
rect 16300 25338 16340 25423
rect 16491 25220 16533 25229
rect 16491 25180 16492 25220
rect 16532 25180 16533 25220
rect 16491 25171 16533 25180
rect 16492 24632 16532 25171
rect 16588 25136 16628 26935
rect 16683 25892 16725 25901
rect 16683 25852 16684 25892
rect 16724 25852 16725 25892
rect 16683 25843 16725 25852
rect 16684 25304 16724 25843
rect 16684 25255 16724 25264
rect 16588 25096 16724 25136
rect 16588 24632 16628 24641
rect 16492 24592 16588 24632
rect 16588 24583 16628 24592
rect 16491 24464 16533 24473
rect 16684 24464 16724 25096
rect 16779 24800 16821 24809
rect 16779 24760 16780 24800
rect 16820 24760 16821 24800
rect 16779 24751 16821 24760
rect 16780 24666 16820 24751
rect 16876 24641 16916 37780
rect 17164 31352 17204 31361
rect 17164 29345 17204 31312
rect 17356 30101 17396 49111
rect 17548 44633 17588 50035
rect 17644 49421 17684 50296
rect 17643 49412 17685 49421
rect 17643 49372 17644 49412
rect 17684 49372 17685 49412
rect 17643 49363 17685 49372
rect 17643 48824 17685 48833
rect 17643 48784 17644 48824
rect 17684 48784 17685 48824
rect 17643 48775 17685 48784
rect 17547 44624 17589 44633
rect 17547 44584 17548 44624
rect 17588 44584 17589 44624
rect 17547 44575 17589 44584
rect 17644 44549 17684 48775
rect 17740 47825 17780 51799
rect 17836 50177 17876 53992
rect 17932 51008 17972 51017
rect 17932 50597 17972 50968
rect 17931 50588 17973 50597
rect 17931 50548 17932 50588
rect 17972 50548 17973 50588
rect 17931 50539 17973 50548
rect 18028 50420 18068 54160
rect 18220 53285 18260 58183
rect 18316 57070 18356 58360
rect 18412 58325 18452 58528
rect 18411 58316 18453 58325
rect 18411 58276 18412 58316
rect 18452 58276 18453 58316
rect 18411 58267 18453 58276
rect 18316 57021 18356 57030
rect 18508 56972 18548 64240
rect 18700 64196 18740 68188
rect 18891 68179 18933 68188
rect 18808 68060 19176 68069
rect 18848 68020 18890 68060
rect 18930 68020 18972 68060
rect 19012 68020 19054 68060
rect 19094 68020 19136 68060
rect 18808 68011 19176 68020
rect 18987 67892 19029 67901
rect 19276 67892 19316 68188
rect 18987 67852 18988 67892
rect 19028 67852 19029 67892
rect 18987 67843 19029 67852
rect 19084 67852 19316 67892
rect 18988 66968 19028 67843
rect 19084 67645 19124 67852
rect 19084 67136 19124 67605
rect 19275 67556 19317 67565
rect 19275 67516 19276 67556
rect 19316 67516 19317 67556
rect 19275 67507 19317 67516
rect 19276 67422 19316 67507
rect 19372 67304 19412 68272
rect 19563 68144 19605 68153
rect 19563 68104 19564 68144
rect 19604 68104 19605 68144
rect 19563 68095 19605 68104
rect 19467 67640 19509 67649
rect 19467 67600 19468 67640
rect 19508 67600 19509 67640
rect 19467 67591 19509 67600
rect 19564 67640 19604 68095
rect 19756 67724 19796 68440
rect 19753 67684 19796 67724
rect 19564 67591 19604 67600
rect 19659 67640 19701 67649
rect 19659 67600 19660 67640
rect 19700 67600 19701 67640
rect 19753 67640 19793 67684
rect 19851 67640 19893 67649
rect 19948 67640 19988 67649
rect 19753 67600 19796 67640
rect 19659 67591 19701 67600
rect 19468 67506 19508 67591
rect 19660 67506 19700 67591
rect 19756 67556 19796 67600
rect 19851 67600 19852 67640
rect 19892 67600 19948 67640
rect 19851 67591 19893 67600
rect 19948 67591 19988 67600
rect 20236 67640 20276 67651
rect 19756 67507 19796 67516
rect 19755 67388 19797 67397
rect 19755 67348 19756 67388
rect 19796 67348 19797 67388
rect 19755 67339 19797 67348
rect 19372 67264 19604 67304
rect 19468 67136 19508 67145
rect 19084 67096 19468 67136
rect 19468 67087 19508 67096
rect 19276 66968 19316 66977
rect 18988 66928 19276 66968
rect 19316 66928 19508 66968
rect 19276 66919 19316 66928
rect 19371 66800 19413 66809
rect 19371 66760 19372 66800
rect 19412 66760 19413 66800
rect 19371 66751 19413 66760
rect 18808 66548 19176 66557
rect 18848 66508 18890 66548
rect 18930 66508 18972 66548
rect 19012 66508 19054 66548
rect 19094 66508 19136 66548
rect 18808 66499 19176 66508
rect 18808 65036 19176 65045
rect 18848 64996 18890 65036
rect 18930 64996 18972 65036
rect 19012 64996 19054 65036
rect 19094 64996 19136 65036
rect 18808 64987 19176 64996
rect 18604 64156 18740 64196
rect 18604 60341 18644 64156
rect 18808 63524 19176 63533
rect 18848 63484 18890 63524
rect 18930 63484 18972 63524
rect 19012 63484 19054 63524
rect 19094 63484 19136 63524
rect 18808 63475 19176 63484
rect 18699 63272 18741 63281
rect 18699 63232 18700 63272
rect 18740 63232 18741 63272
rect 18699 63223 18741 63232
rect 18603 60332 18645 60341
rect 18603 60292 18604 60332
rect 18644 60292 18645 60332
rect 18603 60283 18645 60292
rect 18604 60080 18644 60089
rect 18604 59408 18644 60040
rect 18700 59921 18740 63223
rect 18808 62012 19176 62021
rect 18848 61972 18890 62012
rect 18930 61972 18972 62012
rect 19012 61972 19054 62012
rect 19094 61972 19136 62012
rect 18808 61963 19176 61972
rect 19372 60584 19412 66751
rect 19468 66128 19508 66928
rect 19564 66800 19604 67264
rect 19756 66968 19796 67339
rect 19756 66919 19796 66928
rect 19756 66800 19796 66809
rect 19564 66760 19756 66800
rect 19756 66751 19796 66760
rect 19852 66380 19892 67591
rect 20044 67481 20084 67566
rect 20236 67565 20276 67600
rect 20235 67556 20277 67565
rect 20235 67516 20236 67556
rect 20276 67516 20277 67556
rect 20235 67507 20277 67516
rect 20043 67472 20085 67481
rect 20043 67432 20044 67472
rect 20084 67432 20085 67472
rect 20043 67423 20085 67432
rect 20048 67304 20416 67313
rect 20088 67264 20130 67304
rect 20170 67264 20212 67304
rect 20252 67264 20294 67304
rect 20334 67264 20376 67304
rect 20048 67255 20416 67264
rect 19947 66800 19989 66809
rect 19947 66760 19948 66800
rect 19988 66760 19989 66800
rect 19947 66751 19989 66760
rect 19948 66666 19988 66751
rect 19852 66331 19892 66340
rect 19660 66128 19700 66137
rect 19468 66088 19660 66128
rect 19660 64709 19700 66088
rect 20048 65792 20416 65801
rect 20088 65752 20130 65792
rect 20170 65752 20212 65792
rect 20252 65752 20294 65792
rect 20334 65752 20376 65792
rect 20048 65743 20416 65752
rect 19659 64700 19701 64709
rect 19659 64660 19660 64700
rect 19700 64660 19701 64700
rect 19659 64651 19701 64660
rect 19660 64280 19700 64651
rect 19468 64240 19700 64280
rect 20048 64280 20416 64289
rect 20088 64240 20130 64280
rect 20170 64240 20212 64280
rect 20252 64240 20294 64280
rect 20334 64240 20376 64280
rect 19468 60929 19508 64240
rect 20048 64231 20416 64240
rect 19947 63020 19989 63029
rect 19947 62980 19948 63020
rect 19988 62980 19989 63020
rect 19947 62971 19989 62980
rect 19467 60920 19509 60929
rect 19467 60880 19468 60920
rect 19508 60880 19604 60920
rect 19467 60871 19509 60880
rect 19468 60786 19508 60871
rect 19372 60544 19508 60584
rect 18808 60500 19176 60509
rect 18848 60460 18890 60500
rect 18930 60460 18972 60500
rect 19012 60460 19054 60500
rect 19094 60460 19136 60500
rect 18808 60451 19176 60460
rect 19083 60164 19125 60173
rect 19083 60124 19084 60164
rect 19124 60124 19125 60164
rect 19083 60115 19125 60124
rect 19084 60094 19124 60115
rect 19084 60029 19124 60054
rect 18699 59912 18741 59921
rect 18699 59872 18700 59912
rect 18740 59872 18741 59912
rect 18699 59863 18741 59872
rect 19275 59912 19317 59921
rect 19275 59872 19276 59912
rect 19316 59872 19317 59912
rect 19275 59863 19317 59872
rect 18604 57149 18644 59368
rect 18700 58241 18740 59863
rect 19276 59778 19316 59863
rect 19275 59492 19317 59501
rect 19275 59452 19276 59492
rect 19316 59452 19317 59492
rect 19275 59443 19317 59452
rect 19084 59394 19124 59403
rect 19276 59358 19316 59443
rect 19084 59165 19124 59354
rect 19083 59156 19125 59165
rect 19083 59116 19084 59156
rect 19124 59116 19125 59156
rect 19083 59107 19125 59116
rect 18808 58988 19176 58997
rect 18848 58948 18890 58988
rect 18930 58948 18972 58988
rect 19012 58948 19054 58988
rect 19094 58948 19136 58988
rect 18808 58939 19176 58948
rect 18699 58232 18741 58241
rect 18699 58192 18700 58232
rect 18740 58192 18741 58232
rect 18699 58183 18741 58192
rect 19275 57980 19317 57989
rect 19275 57940 19276 57980
rect 19316 57940 19317 57980
rect 19275 57931 19317 57940
rect 18808 57476 19176 57485
rect 18848 57436 18890 57476
rect 18930 57436 18972 57476
rect 19012 57436 19054 57476
rect 19094 57436 19136 57476
rect 18808 57427 19176 57436
rect 18891 57224 18933 57233
rect 18891 57184 18892 57224
rect 18932 57184 18933 57224
rect 18891 57175 18933 57184
rect 18603 57140 18645 57149
rect 18603 57100 18604 57140
rect 18644 57100 18645 57140
rect 18603 57091 18645 57100
rect 18316 56932 18508 56972
rect 18316 54797 18356 56932
rect 18508 56923 18548 56932
rect 18508 56384 18548 56393
rect 18604 56384 18644 57091
rect 18892 57056 18932 57175
rect 18892 57007 18932 57016
rect 18700 56888 18740 56897
rect 18740 56848 18836 56888
rect 18700 56839 18740 56848
rect 18796 56636 18836 56848
rect 18796 56596 19028 56636
rect 18548 56344 18644 56384
rect 18988 56379 19028 56596
rect 19179 56468 19221 56477
rect 19179 56428 19180 56468
rect 19220 56428 19221 56468
rect 19179 56419 19221 56428
rect 18508 56335 18548 56344
rect 18988 56330 19028 56339
rect 19180 56334 19220 56419
rect 18603 56216 18645 56225
rect 18603 56176 18604 56216
rect 18644 56176 18645 56216
rect 18603 56167 18645 56176
rect 18412 54872 18452 54881
rect 18315 54788 18357 54797
rect 18315 54748 18316 54788
rect 18356 54748 18357 54788
rect 18315 54739 18357 54748
rect 18316 54293 18356 54739
rect 18412 54704 18452 54832
rect 18604 54704 18644 56167
rect 18808 55964 19176 55973
rect 18848 55924 18890 55964
rect 18930 55924 18972 55964
rect 19012 55924 19054 55964
rect 19094 55924 19136 55964
rect 18808 55915 19176 55924
rect 19276 55628 19316 57931
rect 19372 56300 19412 56309
rect 19372 55805 19412 56260
rect 19371 55796 19413 55805
rect 19371 55756 19372 55796
rect 19412 55756 19413 55796
rect 19371 55747 19413 55756
rect 19372 55628 19412 55637
rect 19276 55588 19372 55628
rect 19372 55579 19412 55588
rect 19468 55460 19508 60544
rect 19564 58568 19604 60880
rect 19660 60668 19700 60677
rect 19660 60173 19700 60628
rect 19659 60164 19701 60173
rect 19659 60124 19660 60164
rect 19700 60124 19701 60164
rect 19659 60115 19701 60124
rect 19851 59156 19893 59165
rect 19851 59116 19852 59156
rect 19892 59116 19893 59156
rect 19851 59107 19893 59116
rect 19852 58820 19892 59107
rect 19852 58771 19892 58780
rect 19660 58568 19700 58577
rect 19564 58528 19660 58568
rect 19564 57233 19604 58528
rect 19660 58519 19700 58528
rect 19851 57560 19893 57569
rect 19851 57520 19852 57560
rect 19892 57520 19893 57560
rect 19851 57511 19893 57520
rect 19563 57224 19605 57233
rect 19563 57184 19564 57224
rect 19604 57184 19605 57224
rect 19563 57175 19605 57184
rect 19563 57056 19605 57065
rect 19563 57016 19564 57056
rect 19604 57016 19605 57056
rect 19563 57007 19605 57016
rect 19564 56552 19604 57007
rect 19564 56503 19604 56512
rect 19563 55712 19605 55721
rect 19563 55672 19564 55712
rect 19604 55672 19605 55712
rect 19563 55663 19605 55672
rect 19564 55578 19604 55663
rect 19468 55420 19604 55460
rect 19084 54956 19124 54965
rect 19124 54916 19508 54956
rect 19084 54907 19124 54916
rect 18940 54830 18980 54839
rect 18940 54788 18980 54790
rect 19468 54788 19508 54916
rect 18940 54748 19412 54788
rect 18412 54664 18644 54704
rect 18507 54536 18549 54545
rect 18507 54496 18508 54536
rect 18548 54496 18549 54536
rect 18507 54487 18549 54496
rect 18315 54284 18357 54293
rect 18315 54244 18316 54284
rect 18356 54244 18357 54284
rect 18315 54235 18357 54244
rect 18508 53360 18548 54487
rect 18219 53276 18261 53285
rect 18219 53236 18220 53276
rect 18260 53236 18261 53276
rect 18219 53227 18261 53236
rect 17932 50380 18068 50420
rect 17835 50168 17877 50177
rect 17835 50128 17836 50168
rect 17876 50128 17877 50168
rect 17835 50119 17877 50128
rect 17932 49841 17972 50380
rect 18124 50336 18164 50345
rect 18220 50336 18260 53227
rect 18315 51932 18357 51941
rect 18315 51892 18316 51932
rect 18356 51892 18357 51932
rect 18315 51883 18357 51892
rect 18316 51848 18356 51883
rect 18412 51857 18452 51942
rect 18316 51797 18356 51808
rect 18411 51848 18453 51857
rect 18411 51808 18412 51848
rect 18452 51808 18453 51848
rect 18411 51799 18453 51808
rect 18164 50296 18260 50336
rect 18028 50252 18068 50261
rect 17931 49832 17973 49841
rect 17931 49792 17932 49832
rect 17972 49792 17973 49832
rect 17931 49783 17973 49792
rect 18028 49589 18068 50212
rect 18124 49841 18164 50296
rect 18219 50168 18261 50177
rect 18508 50168 18548 53320
rect 18604 50513 18644 54664
rect 19275 54620 19317 54629
rect 19275 54580 19276 54620
rect 19316 54580 19317 54620
rect 19275 54571 19317 54580
rect 19276 54486 19316 54571
rect 18808 54452 19176 54461
rect 18848 54412 18890 54452
rect 18930 54412 18972 54452
rect 19012 54412 19054 54452
rect 19094 54412 19136 54452
rect 18808 54403 19176 54412
rect 19179 54284 19221 54293
rect 19179 54244 19180 54284
rect 19220 54244 19221 54284
rect 19179 54235 19221 54244
rect 19276 54284 19316 54293
rect 19372 54284 19412 54748
rect 19468 54739 19508 54748
rect 19316 54244 19412 54284
rect 19276 54235 19316 54244
rect 19180 54116 19220 54235
rect 19468 54116 19508 54125
rect 19180 54076 19316 54116
rect 19083 54032 19125 54041
rect 19083 53992 19084 54032
rect 19124 53992 19125 54032
rect 19083 53983 19125 53992
rect 19084 53898 19124 53983
rect 18699 53360 18741 53369
rect 18699 53320 18700 53360
rect 18740 53320 18741 53360
rect 18699 53311 18741 53320
rect 18700 52520 18740 53311
rect 18808 52940 19176 52949
rect 18848 52900 18890 52940
rect 18930 52900 18972 52940
rect 19012 52900 19054 52940
rect 19094 52900 19136 52940
rect 18808 52891 19176 52900
rect 19276 52772 19316 54076
rect 19468 53621 19508 54076
rect 19467 53612 19509 53621
rect 19467 53572 19468 53612
rect 19508 53572 19509 53612
rect 19467 53563 19509 53572
rect 19564 52772 19604 55420
rect 19852 54797 19892 57511
rect 19660 54788 19700 54797
rect 19660 54545 19700 54748
rect 19851 54788 19893 54797
rect 19851 54748 19852 54788
rect 19892 54748 19893 54788
rect 19851 54739 19893 54748
rect 19852 54620 19892 54629
rect 19659 54536 19701 54545
rect 19659 54496 19660 54536
rect 19700 54496 19701 54536
rect 19659 54487 19701 54496
rect 19852 54377 19892 54580
rect 19851 54368 19893 54377
rect 19851 54328 19852 54368
rect 19892 54328 19893 54368
rect 19851 54319 19893 54328
rect 19851 54116 19893 54125
rect 19851 54076 19852 54116
rect 19892 54076 19893 54116
rect 19851 54067 19893 54076
rect 19852 53982 19892 54067
rect 18603 50504 18645 50513
rect 18603 50464 18604 50504
rect 18644 50464 18645 50504
rect 18603 50455 18645 50464
rect 18604 50336 18644 50455
rect 18604 50287 18644 50296
rect 18700 50168 18740 52480
rect 18988 52732 19316 52772
rect 19468 52732 19604 52772
rect 19660 53864 19700 53873
rect 18892 52352 18932 52361
rect 18796 52312 18892 52352
rect 18796 51941 18836 52312
rect 18892 52303 18932 52312
rect 18795 51932 18837 51941
rect 18795 51892 18796 51932
rect 18836 51892 18837 51932
rect 18795 51883 18837 51892
rect 18892 51848 18932 51857
rect 18988 51848 19028 52732
rect 19372 52352 19412 52361
rect 19275 52184 19317 52193
rect 19275 52144 19276 52184
rect 19316 52144 19317 52184
rect 19275 52135 19317 52144
rect 18932 51808 19028 51848
rect 19276 51848 19316 52135
rect 19372 52109 19412 52312
rect 19371 52100 19413 52109
rect 19371 52060 19372 52100
rect 19412 52060 19413 52100
rect 19371 52051 19413 52060
rect 19372 51848 19412 51857
rect 19276 51808 19372 51848
rect 18892 51799 18932 51808
rect 18795 51764 18837 51773
rect 18795 51724 18796 51764
rect 18836 51724 18837 51764
rect 18795 51715 18837 51724
rect 18796 51630 18836 51715
rect 18808 51428 19176 51437
rect 18848 51388 18890 51428
rect 18930 51388 18972 51428
rect 19012 51388 19054 51428
rect 19094 51388 19136 51428
rect 18808 51379 19176 51388
rect 19179 51092 19221 51101
rect 19179 51052 19180 51092
rect 19220 51052 19221 51092
rect 19179 51043 19221 51052
rect 19180 51008 19220 51043
rect 19180 50957 19220 50968
rect 19179 50840 19221 50849
rect 19179 50800 19180 50840
rect 19220 50800 19221 50840
rect 19179 50791 19221 50800
rect 19180 50336 19220 50791
rect 19276 50672 19316 51808
rect 19372 51799 19412 51808
rect 19372 50849 19412 50934
rect 19371 50840 19413 50849
rect 19371 50800 19372 50840
rect 19412 50800 19413 50840
rect 19371 50791 19413 50800
rect 19276 50632 19412 50672
rect 19275 50504 19317 50513
rect 19275 50464 19276 50504
rect 19316 50464 19317 50504
rect 19275 50455 19317 50464
rect 19276 50370 19316 50455
rect 19132 50326 19220 50336
rect 19172 50296 19220 50326
rect 19132 50277 19172 50286
rect 18219 50128 18220 50168
rect 18260 50128 18261 50168
rect 18219 50119 18261 50128
rect 18412 50128 18548 50168
rect 18604 50128 18740 50168
rect 18123 49832 18165 49841
rect 18123 49792 18124 49832
rect 18164 49792 18165 49832
rect 18123 49783 18165 49792
rect 18027 49580 18069 49589
rect 18027 49540 18028 49580
rect 18068 49540 18069 49580
rect 18027 49531 18069 49540
rect 18123 49412 18165 49421
rect 18123 49372 18124 49412
rect 18164 49372 18165 49412
rect 18123 49363 18165 49372
rect 18028 48824 18068 48833
rect 18028 48236 18068 48784
rect 18124 48824 18164 49363
rect 18124 48775 18164 48784
rect 18220 48656 18260 50119
rect 18412 48917 18452 50128
rect 18507 49832 18549 49841
rect 18507 49792 18508 49832
rect 18548 49792 18549 49832
rect 18507 49783 18549 49792
rect 18508 48992 18548 49783
rect 18604 49328 18644 50128
rect 18808 49916 19176 49925
rect 18848 49876 18890 49916
rect 18930 49876 18972 49916
rect 19012 49876 19054 49916
rect 19094 49876 19136 49916
rect 18808 49867 19176 49876
rect 19372 49832 19412 50632
rect 19468 50420 19508 52732
rect 19564 52604 19604 52613
rect 19564 52025 19604 52564
rect 19660 52361 19700 53824
rect 19755 53360 19797 53369
rect 19755 53320 19756 53360
rect 19796 53320 19797 53360
rect 19755 53311 19797 53320
rect 19756 53226 19796 53311
rect 19948 53276 19988 62971
rect 20048 62768 20416 62777
rect 20088 62728 20130 62768
rect 20170 62728 20212 62768
rect 20252 62728 20294 62768
rect 20334 62728 20376 62768
rect 20048 62719 20416 62728
rect 20524 62525 20564 76495
rect 20715 74528 20757 74537
rect 20715 74488 20716 74528
rect 20756 74488 20757 74528
rect 20715 74479 20757 74488
rect 20716 63449 20756 74479
rect 20715 63440 20757 63449
rect 20715 63400 20716 63440
rect 20756 63400 20757 63440
rect 20715 63391 20757 63400
rect 20523 62516 20565 62525
rect 20523 62476 20524 62516
rect 20564 62476 20565 62516
rect 20523 62467 20565 62476
rect 20715 61760 20757 61769
rect 20715 61720 20716 61760
rect 20756 61720 20757 61760
rect 20715 61711 20757 61720
rect 20048 61256 20416 61265
rect 20088 61216 20130 61256
rect 20170 61216 20212 61256
rect 20252 61216 20294 61256
rect 20334 61216 20376 61256
rect 20048 61207 20416 61216
rect 20048 59744 20416 59753
rect 20088 59704 20130 59744
rect 20170 59704 20212 59744
rect 20252 59704 20294 59744
rect 20334 59704 20376 59744
rect 20048 59695 20416 59704
rect 20619 59744 20661 59753
rect 20619 59704 20620 59744
rect 20660 59704 20661 59744
rect 20619 59695 20661 59704
rect 20048 58232 20416 58241
rect 20088 58192 20130 58232
rect 20170 58192 20212 58232
rect 20252 58192 20294 58232
rect 20334 58192 20376 58232
rect 20048 58183 20416 58192
rect 20043 57980 20085 57989
rect 20043 57940 20044 57980
rect 20084 57940 20085 57980
rect 20043 57931 20085 57940
rect 20044 57476 20084 57931
rect 20044 57436 20180 57476
rect 20140 57098 20180 57436
rect 20140 57049 20180 57058
rect 20048 56720 20416 56729
rect 20088 56680 20130 56720
rect 20170 56680 20212 56720
rect 20252 56680 20294 56720
rect 20334 56680 20376 56720
rect 20048 56671 20416 56680
rect 20048 55208 20416 55217
rect 20088 55168 20130 55208
rect 20170 55168 20212 55208
rect 20252 55168 20294 55208
rect 20334 55168 20376 55208
rect 20048 55159 20416 55168
rect 20235 55040 20277 55049
rect 20235 55000 20236 55040
rect 20276 55000 20277 55040
rect 20235 54991 20277 55000
rect 20236 54906 20276 54991
rect 20043 54788 20085 54797
rect 20043 54748 20044 54788
rect 20084 54748 20085 54788
rect 20043 54739 20085 54748
rect 20044 54654 20084 54739
rect 20044 53873 20084 53958
rect 20043 53864 20085 53873
rect 20043 53824 20044 53864
rect 20084 53824 20085 53864
rect 20043 53815 20085 53824
rect 20048 53696 20416 53705
rect 20088 53656 20130 53696
rect 20170 53656 20212 53696
rect 20252 53656 20294 53696
rect 20334 53656 20376 53696
rect 20048 53647 20416 53656
rect 19948 53236 20084 53276
rect 19948 53108 19988 53117
rect 19852 53068 19948 53108
rect 19755 52772 19797 52781
rect 19755 52732 19756 52772
rect 19796 52732 19797 52772
rect 19755 52723 19797 52732
rect 19756 52604 19796 52723
rect 19756 52555 19796 52564
rect 19755 52436 19797 52445
rect 19755 52396 19756 52436
rect 19796 52396 19797 52436
rect 19755 52387 19797 52396
rect 19659 52352 19701 52361
rect 19659 52312 19660 52352
rect 19700 52312 19701 52352
rect 19659 52303 19701 52312
rect 19659 52100 19701 52109
rect 19659 52060 19660 52100
rect 19700 52060 19701 52100
rect 19659 52051 19701 52060
rect 19563 52016 19605 52025
rect 19563 51976 19564 52016
rect 19604 51976 19605 52016
rect 19563 51967 19605 51976
rect 19563 50840 19605 50849
rect 19563 50800 19564 50840
rect 19604 50800 19605 50840
rect 19563 50791 19605 50800
rect 19564 50706 19604 50791
rect 19468 50380 19604 50420
rect 19468 50252 19508 50261
rect 19468 50093 19508 50212
rect 19467 50084 19509 50093
rect 19467 50044 19468 50084
rect 19508 50044 19509 50084
rect 19467 50035 19509 50044
rect 19276 49792 19412 49832
rect 18987 49748 19029 49757
rect 18987 49708 18988 49748
rect 19028 49708 19029 49748
rect 18987 49699 19029 49708
rect 18988 49614 19028 49699
rect 18700 49505 18740 49590
rect 19180 49580 19220 49589
rect 18699 49496 18741 49505
rect 18699 49456 18700 49496
rect 18740 49456 18741 49496
rect 18699 49447 18741 49456
rect 18604 49288 18740 49328
rect 18508 48952 18647 48992
rect 18411 48908 18453 48917
rect 18607 48908 18647 48952
rect 18411 48868 18412 48908
rect 18452 48868 18453 48908
rect 18411 48859 18453 48868
rect 18604 48868 18647 48908
rect 18315 48824 18357 48833
rect 18315 48784 18316 48824
rect 18356 48784 18357 48824
rect 18315 48775 18357 48784
rect 18604 48824 18644 48868
rect 18604 48775 18644 48784
rect 18028 48187 18068 48196
rect 18124 48616 18260 48656
rect 17835 47984 17877 47993
rect 17835 47944 17836 47984
rect 17876 47944 17877 47984
rect 17835 47935 17877 47944
rect 17836 47850 17876 47935
rect 17739 47816 17781 47825
rect 17739 47776 17740 47816
rect 17780 47776 17781 47816
rect 17739 47767 17781 47776
rect 18027 47816 18069 47825
rect 18027 47776 18028 47816
rect 18068 47776 18069 47816
rect 18027 47767 18069 47776
rect 17931 47060 17973 47069
rect 17931 47020 17932 47060
rect 17972 47020 17973 47060
rect 17931 47011 17973 47020
rect 17932 46472 17972 47011
rect 17932 46423 17972 46432
rect 18028 46472 18068 47767
rect 17835 45380 17877 45389
rect 17835 45340 17836 45380
rect 17876 45340 17877 45380
rect 17835 45331 17877 45340
rect 17739 44960 17781 44969
rect 17739 44920 17740 44960
rect 17780 44920 17781 44960
rect 17739 44911 17781 44920
rect 17643 44540 17685 44549
rect 17643 44500 17644 44540
rect 17684 44500 17685 44540
rect 17643 44491 17685 44500
rect 17452 44372 17492 44381
rect 17492 44332 17684 44372
rect 17452 44323 17492 44332
rect 17451 43784 17493 43793
rect 17451 43744 17452 43784
rect 17492 43744 17493 43784
rect 17451 43735 17493 43744
rect 17452 43700 17492 43735
rect 17452 43649 17492 43660
rect 17644 43532 17684 44332
rect 17740 44129 17780 44911
rect 17739 44120 17781 44129
rect 17739 44080 17740 44120
rect 17780 44080 17781 44120
rect 17739 44071 17781 44080
rect 17644 43483 17684 43492
rect 17739 43532 17781 43541
rect 17739 43492 17740 43532
rect 17780 43492 17781 43532
rect 17739 43483 17781 43492
rect 17836 43532 17876 45331
rect 17931 45212 17973 45221
rect 17931 45172 17932 45212
rect 17972 45172 17973 45212
rect 17931 45163 17973 45172
rect 17932 44960 17972 45163
rect 17932 44911 17972 44920
rect 18028 44960 18068 46432
rect 18124 45137 18164 48616
rect 18220 47984 18260 47993
rect 18316 47984 18356 48775
rect 18260 47944 18356 47984
rect 18508 48740 18548 48749
rect 18220 47935 18260 47944
rect 18315 47816 18357 47825
rect 18315 47776 18316 47816
rect 18356 47776 18357 47816
rect 18315 47767 18357 47776
rect 18220 47312 18260 47323
rect 18220 47237 18260 47272
rect 18219 47228 18261 47237
rect 18219 47188 18220 47228
rect 18260 47188 18261 47228
rect 18219 47179 18261 47188
rect 18316 47060 18356 47767
rect 18220 47020 18356 47060
rect 18411 47060 18453 47069
rect 18411 47020 18412 47060
rect 18452 47020 18453 47060
rect 18220 45725 18260 47020
rect 18411 47011 18453 47020
rect 18412 46926 18452 47011
rect 18315 46892 18357 46901
rect 18315 46852 18316 46892
rect 18356 46852 18357 46892
rect 18315 46843 18357 46852
rect 18316 45800 18356 46843
rect 18508 46640 18548 48700
rect 18603 48656 18645 48665
rect 18603 48616 18604 48656
rect 18644 48616 18645 48656
rect 18603 48607 18645 48616
rect 18604 47312 18644 48607
rect 18604 47263 18644 47272
rect 18700 46901 18740 49288
rect 19180 49001 19220 49540
rect 19179 48992 19221 49001
rect 19179 48952 19180 48992
rect 19220 48952 19221 48992
rect 19179 48943 19221 48952
rect 19084 48824 19124 48833
rect 19276 48824 19316 49792
rect 19371 49664 19413 49673
rect 19371 49624 19372 49664
rect 19412 49624 19413 49664
rect 19371 49615 19413 49624
rect 19372 49580 19412 49615
rect 19372 49529 19412 49540
rect 19564 49496 19604 50380
rect 19660 50345 19700 52051
rect 19756 51260 19796 52387
rect 19852 51843 19892 53068
rect 19948 53059 19988 53068
rect 20044 52445 20084 53236
rect 20043 52436 20085 52445
rect 20043 52396 20044 52436
rect 20084 52396 20085 52436
rect 20043 52387 20085 52396
rect 19852 51794 19892 51803
rect 19948 52352 19988 52361
rect 19948 51689 19988 52312
rect 20048 52184 20416 52193
rect 20088 52144 20130 52184
rect 20170 52144 20212 52184
rect 20252 52144 20294 52184
rect 20334 52144 20376 52184
rect 20048 52135 20416 52144
rect 20043 52016 20085 52025
rect 20043 51976 20044 52016
rect 20084 51976 20085 52016
rect 20043 51967 20085 51976
rect 20044 51882 20084 51967
rect 19947 51680 19989 51689
rect 19947 51640 19948 51680
rect 19988 51640 19989 51680
rect 19947 51631 19989 51640
rect 19947 51344 19989 51353
rect 19947 51304 19948 51344
rect 19988 51304 19989 51344
rect 19947 51295 19989 51304
rect 19756 51220 19892 51260
rect 19756 51092 19796 51101
rect 19756 50513 19796 51052
rect 19755 50504 19797 50513
rect 19755 50464 19756 50504
rect 19796 50464 19797 50504
rect 19755 50455 19797 50464
rect 19852 50429 19892 51220
rect 19948 51092 19988 51295
rect 19948 51043 19988 51052
rect 20139 51008 20181 51017
rect 20139 50968 20140 51008
rect 20180 50968 20181 51008
rect 20139 50959 20181 50968
rect 20140 50840 20180 50959
rect 20140 50791 20180 50800
rect 19947 50672 19989 50681
rect 19947 50632 19948 50672
rect 19988 50632 19989 50672
rect 19947 50623 19989 50632
rect 20048 50672 20416 50681
rect 20088 50632 20130 50672
rect 20170 50632 20212 50672
rect 20252 50632 20294 50672
rect 20334 50632 20376 50672
rect 20048 50623 20416 50632
rect 19851 50420 19893 50429
rect 19851 50380 19852 50420
rect 19892 50380 19893 50420
rect 19851 50371 19893 50380
rect 19659 50336 19701 50345
rect 19659 50296 19660 50336
rect 19700 50296 19701 50336
rect 19659 50287 19701 50296
rect 19852 50252 19892 50263
rect 19852 50177 19892 50212
rect 19851 50168 19893 50177
rect 19851 50128 19852 50168
rect 19892 50128 19893 50168
rect 19851 50119 19893 50128
rect 19660 50084 19700 50093
rect 19660 49673 19700 50044
rect 19659 49664 19701 49673
rect 19659 49624 19660 49664
rect 19700 49624 19701 49664
rect 19659 49615 19701 49624
rect 19756 49580 19796 49589
rect 19948 49580 19988 50623
rect 20043 50336 20085 50345
rect 20043 50296 20044 50336
rect 20084 50296 20085 50336
rect 20043 50287 20085 50296
rect 20044 50168 20084 50287
rect 20044 50119 20084 50128
rect 19796 49540 19988 49580
rect 19756 49531 19796 49540
rect 19468 49456 19604 49496
rect 19468 49076 19508 49456
rect 19564 49328 19604 49337
rect 19948 49328 19988 49337
rect 19604 49288 19892 49328
rect 19564 49279 19604 49288
rect 19124 48784 19316 48824
rect 19084 48775 19124 48784
rect 18808 48404 19176 48413
rect 18848 48364 18890 48404
rect 18930 48364 18972 48404
rect 19012 48364 19054 48404
rect 19094 48364 19136 48404
rect 18808 48355 19176 48364
rect 19276 47573 19316 48784
rect 19372 49036 19508 49076
rect 19275 47564 19317 47573
rect 19275 47524 19276 47564
rect 19316 47524 19317 47564
rect 19275 47515 19317 47524
rect 19275 47396 19317 47405
rect 19275 47356 19276 47396
rect 19316 47356 19317 47396
rect 19275 47347 19317 47356
rect 18699 46892 18741 46901
rect 18699 46852 18700 46892
rect 18740 46852 18741 46892
rect 18699 46843 18741 46852
rect 18808 46892 19176 46901
rect 18848 46852 18890 46892
rect 18930 46852 18972 46892
rect 19012 46852 19054 46892
rect 19094 46852 19136 46892
rect 18808 46843 19176 46852
rect 18987 46724 19029 46733
rect 18987 46684 18988 46724
rect 19028 46684 19029 46724
rect 18987 46675 19029 46684
rect 18219 45716 18261 45725
rect 18219 45676 18220 45716
rect 18260 45676 18261 45716
rect 18219 45667 18261 45676
rect 18123 45128 18165 45137
rect 18123 45088 18124 45128
rect 18164 45088 18165 45128
rect 18123 45079 18165 45088
rect 18028 43952 18068 44920
rect 18316 44885 18356 45760
rect 18412 46600 18548 46640
rect 18412 46556 18452 46600
rect 18412 45044 18452 46516
rect 18507 46472 18549 46481
rect 18988 46472 19028 46675
rect 18507 46432 18508 46472
rect 18548 46432 18644 46472
rect 18507 46423 18549 46432
rect 18508 46338 18548 46423
rect 18508 45548 18548 45557
rect 18508 45221 18548 45508
rect 18507 45212 18549 45221
rect 18507 45172 18508 45212
rect 18548 45172 18549 45212
rect 18507 45163 18549 45172
rect 18315 44876 18357 44885
rect 18315 44836 18316 44876
rect 18356 44836 18357 44876
rect 18315 44827 18357 44836
rect 18123 44540 18165 44549
rect 18123 44500 18124 44540
rect 18164 44500 18165 44540
rect 18123 44491 18165 44500
rect 18124 44288 18164 44491
rect 18316 44297 18356 44827
rect 18124 44239 18164 44248
rect 18315 44288 18357 44297
rect 18315 44248 18316 44288
rect 18356 44248 18357 44288
rect 18315 44239 18357 44248
rect 18219 44204 18261 44213
rect 18219 44164 18220 44204
rect 18260 44164 18261 44204
rect 18219 44155 18261 44164
rect 18028 43912 18164 43952
rect 17836 43483 17876 43492
rect 17547 42860 17589 42869
rect 17547 42820 17548 42860
rect 17588 42820 17589 42860
rect 17547 42811 17589 42820
rect 17452 32864 17492 32873
rect 17452 32705 17492 32824
rect 17451 32696 17493 32705
rect 17451 32656 17452 32696
rect 17492 32656 17493 32696
rect 17451 32647 17493 32656
rect 17355 30092 17397 30101
rect 17548 30092 17588 42811
rect 17740 40433 17780 43483
rect 18028 43280 18068 43289
rect 18028 42953 18068 43240
rect 18027 42944 18069 42953
rect 18027 42904 18028 42944
rect 18068 42904 18069 42944
rect 18027 42895 18069 42904
rect 17931 42272 17973 42281
rect 17931 42232 17932 42272
rect 17972 42232 17973 42272
rect 17931 42223 17973 42232
rect 17739 40424 17781 40433
rect 17739 40384 17740 40424
rect 17780 40384 17781 40424
rect 17739 40375 17781 40384
rect 17644 32696 17684 32705
rect 17644 31366 17684 32656
rect 17644 31317 17684 31326
rect 17739 31352 17781 31361
rect 17739 31312 17740 31352
rect 17780 31312 17781 31352
rect 17739 31303 17781 31312
rect 17740 30773 17780 31303
rect 17835 31268 17877 31277
rect 17835 31228 17836 31268
rect 17876 31228 17877 31268
rect 17835 31219 17877 31228
rect 17836 31134 17876 31219
rect 17932 31016 17972 42223
rect 18027 42020 18069 42029
rect 18027 41980 18028 42020
rect 18068 41980 18069 42020
rect 18027 41971 18069 41980
rect 17836 30976 17972 31016
rect 17739 30764 17781 30773
rect 17739 30724 17740 30764
rect 17780 30724 17781 30764
rect 17739 30715 17781 30724
rect 17740 30680 17780 30715
rect 17643 30260 17685 30269
rect 17643 30220 17644 30260
rect 17684 30220 17685 30260
rect 17643 30211 17685 30220
rect 17355 30052 17356 30092
rect 17396 30052 17397 30092
rect 17355 30043 17397 30052
rect 17452 30052 17588 30092
rect 17452 29672 17492 30052
rect 17548 29849 17588 29934
rect 17547 29840 17589 29849
rect 17547 29800 17548 29840
rect 17588 29800 17589 29840
rect 17547 29791 17589 29800
rect 17644 29840 17684 30211
rect 17644 29791 17684 29800
rect 17452 29632 17588 29672
rect 17163 29336 17205 29345
rect 17163 29296 17164 29336
rect 17204 29296 17205 29336
rect 17163 29287 17205 29296
rect 16971 29252 17013 29261
rect 16971 29212 16972 29252
rect 17012 29212 17013 29252
rect 16971 29203 17013 29212
rect 16972 29168 17012 29203
rect 16972 29117 17012 29128
rect 17068 29168 17108 29177
rect 17068 27665 17108 29128
rect 17220 29168 17396 29188
rect 17452 29168 17492 29177
rect 17260 29148 17452 29168
rect 17356 29128 17452 29148
rect 17220 29093 17260 29128
rect 17219 29084 17261 29093
rect 17219 29044 17220 29084
rect 17260 29044 17261 29084
rect 17219 29035 17261 29044
rect 17220 29004 17260 29035
rect 17356 27824 17396 27833
rect 17452 27824 17492 29128
rect 17548 29168 17588 29632
rect 17740 29513 17780 30640
rect 17739 29504 17781 29513
rect 17739 29464 17740 29504
rect 17780 29464 17781 29504
rect 17739 29455 17781 29464
rect 17643 29420 17685 29429
rect 17643 29380 17644 29420
rect 17684 29380 17685 29420
rect 17643 29371 17685 29380
rect 17548 29093 17588 29128
rect 17547 29084 17589 29093
rect 17547 29044 17548 29084
rect 17588 29044 17589 29084
rect 17547 29035 17589 29044
rect 17548 29004 17588 29035
rect 17644 28916 17684 29371
rect 17740 29336 17780 29345
rect 17740 29177 17780 29296
rect 17739 29168 17781 29177
rect 17739 29128 17740 29168
rect 17780 29128 17781 29168
rect 17739 29119 17781 29128
rect 17396 27784 17492 27824
rect 17548 28876 17684 28916
rect 17356 27775 17396 27784
rect 17067 27656 17109 27665
rect 17067 27616 17068 27656
rect 17108 27616 17109 27656
rect 17067 27607 17109 27616
rect 17164 27656 17204 27665
rect 17164 27497 17204 27616
rect 17163 27488 17205 27497
rect 17163 27448 17164 27488
rect 17204 27448 17205 27488
rect 17163 27439 17205 27448
rect 17259 27320 17301 27329
rect 17259 27280 17260 27320
rect 17300 27280 17301 27320
rect 17259 27271 17301 27280
rect 17067 26648 17109 26657
rect 17067 26608 17068 26648
rect 17108 26608 17109 26648
rect 17067 26599 17109 26608
rect 16971 26228 17013 26237
rect 16971 26188 16972 26228
rect 17012 26188 17013 26228
rect 16971 26179 17013 26188
rect 16972 25304 17012 26179
rect 16972 25255 17012 25264
rect 17068 25304 17108 26599
rect 17260 26144 17300 27271
rect 17356 26816 17396 26827
rect 17356 26741 17396 26776
rect 17452 26816 17492 26825
rect 17355 26732 17397 26741
rect 17355 26692 17356 26732
rect 17396 26692 17397 26732
rect 17355 26683 17397 26692
rect 17452 26573 17492 26776
rect 17451 26564 17493 26573
rect 17451 26524 17452 26564
rect 17492 26524 17493 26564
rect 17451 26515 17493 26524
rect 17452 26144 17492 26153
rect 17260 26104 17452 26144
rect 17452 26095 17492 26104
rect 17163 25472 17205 25481
rect 17163 25432 17164 25472
rect 17204 25432 17205 25472
rect 17163 25423 17205 25432
rect 17356 25472 17396 25481
rect 17068 25255 17108 25264
rect 16971 24800 17013 24809
rect 16971 24760 16972 24800
rect 17012 24760 17013 24800
rect 16971 24751 17013 24760
rect 16875 24632 16917 24641
rect 16875 24592 16876 24632
rect 16916 24592 16917 24632
rect 16875 24583 16917 24592
rect 16972 24632 17012 24751
rect 16972 24583 17012 24592
rect 17068 24632 17108 24641
rect 16491 24424 16492 24464
rect 16532 24424 16533 24464
rect 16491 24415 16533 24424
rect 16588 24424 16724 24464
rect 16492 23876 16532 24415
rect 16492 23827 16532 23836
rect 16396 23792 16436 23801
rect 16299 23624 16341 23633
rect 16299 23584 16300 23624
rect 16340 23584 16341 23624
rect 16299 23575 16341 23584
rect 16300 22952 16340 23575
rect 16396 23381 16436 23752
rect 16395 23372 16437 23381
rect 16395 23332 16396 23372
rect 16436 23332 16437 23372
rect 16395 23323 16437 23332
rect 16396 22952 16436 22961
rect 16300 22912 16396 22952
rect 16396 22903 16436 22912
rect 16204 22828 16340 22868
rect 16107 22819 16149 22828
rect 16011 22112 16053 22121
rect 16011 22072 16012 22112
rect 16052 22072 16053 22112
rect 16011 22063 16053 22072
rect 16012 21533 16052 22063
rect 16108 21608 16148 22819
rect 16203 22700 16245 22709
rect 16203 22660 16204 22700
rect 16244 22660 16245 22700
rect 16203 22651 16245 22660
rect 16204 21869 16244 22651
rect 16203 21860 16245 21869
rect 16203 21820 16204 21860
rect 16244 21820 16245 21860
rect 16203 21811 16245 21820
rect 16108 21559 16148 21568
rect 16204 21608 16244 21811
rect 16204 21559 16244 21568
rect 16011 21524 16053 21533
rect 16011 21484 16012 21524
rect 16052 21484 16053 21524
rect 16011 21475 16053 21484
rect 16107 21440 16149 21449
rect 16107 21400 16108 21440
rect 16148 21400 16149 21440
rect 16107 21391 16149 21400
rect 16011 21356 16053 21365
rect 16011 21316 16012 21356
rect 16052 21316 16053 21356
rect 16011 21307 16053 21316
rect 15915 18752 15957 18761
rect 15915 18712 15916 18752
rect 15956 18712 15957 18752
rect 15915 18703 15957 18712
rect 15921 18584 15961 18593
rect 15820 18535 15860 18544
rect 15916 18544 15921 18584
rect 15916 18535 15961 18544
rect 15723 17996 15765 18005
rect 15723 17956 15724 17996
rect 15764 17956 15765 17996
rect 15723 17947 15765 17956
rect 15819 17912 15861 17921
rect 15819 17872 15820 17912
rect 15860 17872 15861 17912
rect 15819 17863 15861 17872
rect 15628 17695 15668 17704
rect 15436 17620 15572 17660
rect 15436 17576 15476 17620
rect 15436 17527 15476 17536
rect 15435 17240 15477 17249
rect 15435 17200 15436 17240
rect 15476 17200 15477 17240
rect 15435 17191 15477 17200
rect 15436 14897 15476 17191
rect 15532 15560 15572 15569
rect 15435 14888 15477 14897
rect 15435 14848 15436 14888
rect 15476 14848 15477 14888
rect 15435 14839 15477 14848
rect 15532 14729 15572 15520
rect 15723 15308 15765 15317
rect 15723 15268 15724 15308
rect 15764 15268 15765 15308
rect 15723 15259 15765 15268
rect 15724 15174 15764 15259
rect 15531 14720 15573 14729
rect 15531 14680 15532 14720
rect 15572 14680 15573 14720
rect 15531 14671 15573 14680
rect 14667 13796 14709 13805
rect 14667 13756 14668 13796
rect 14708 13756 14709 13796
rect 14667 13747 14709 13756
rect 15148 13385 15188 14008
rect 15244 14344 15380 14384
rect 15147 13376 15189 13385
rect 15147 13336 15148 13376
rect 15188 13336 15189 13376
rect 15147 13327 15189 13336
rect 14908 13217 14948 13226
rect 14948 13177 15188 13208
rect 14908 13168 15188 13177
rect 15051 13040 15093 13049
rect 15051 13000 15052 13040
rect 15092 13000 15093 13040
rect 15051 12991 15093 13000
rect 15052 12906 15092 12991
rect 15148 12620 15188 13168
rect 15244 12629 15284 14344
rect 15340 14132 15380 14141
rect 15380 14092 15668 14132
rect 15340 14083 15380 14092
rect 15628 14048 15668 14092
rect 15628 13999 15668 14008
rect 15724 14048 15764 14057
rect 15339 13880 15381 13889
rect 15339 13840 15340 13880
rect 15380 13840 15381 13880
rect 15339 13831 15381 13840
rect 15148 12571 15188 12580
rect 15243 12620 15285 12629
rect 15243 12580 15244 12620
rect 15284 12580 15285 12620
rect 15243 12571 15285 12580
rect 14956 12536 14996 12545
rect 14716 11705 14756 11714
rect 14956 11705 14996 12496
rect 14955 11696 14997 11705
rect 14756 11665 14804 11696
rect 14716 11656 14804 11665
rect 14764 11192 14804 11656
rect 14955 11656 14956 11696
rect 14996 11656 14997 11696
rect 14955 11647 14997 11656
rect 14859 11528 14901 11537
rect 14859 11488 14860 11528
rect 14900 11488 14901 11528
rect 14859 11479 14901 11488
rect 14860 11394 14900 11479
rect 14860 11192 14900 11201
rect 14764 11152 14860 11192
rect 14860 11143 14900 11152
rect 14956 11033 14996 11647
rect 15340 11360 15380 13831
rect 15435 13796 15477 13805
rect 15435 13756 15436 13796
rect 15476 13756 15477 13796
rect 15435 13747 15477 13756
rect 15148 11320 15380 11360
rect 14668 11024 14708 11033
rect 14668 10865 14708 10984
rect 14955 11024 14997 11033
rect 14955 10984 14956 11024
rect 14996 10984 14997 11024
rect 14955 10975 14997 10984
rect 15052 11024 15092 11035
rect 15052 10949 15092 10984
rect 15051 10940 15093 10949
rect 15051 10900 15052 10940
rect 15092 10900 15093 10940
rect 15051 10891 15093 10900
rect 14667 10856 14709 10865
rect 14667 10816 14668 10856
rect 14708 10816 14709 10856
rect 14667 10807 14709 10816
rect 14667 10268 14709 10277
rect 14667 10228 14668 10268
rect 14708 10228 14709 10268
rect 14667 10219 14709 10228
rect 14668 10100 14708 10219
rect 14812 10193 14852 10202
rect 14852 10153 15092 10184
rect 14812 10144 15092 10153
rect 14668 10060 14996 10100
rect 14956 10016 14996 10060
rect 14956 9967 14996 9976
rect 14667 9932 14709 9941
rect 14667 9892 14668 9932
rect 14708 9892 14709 9932
rect 14667 9883 14709 9892
rect 14571 9512 14613 9521
rect 14571 9472 14572 9512
rect 14612 9472 14613 9512
rect 14571 9463 14613 9472
rect 14571 8420 14613 8429
rect 14571 8380 14572 8420
rect 14612 8380 14613 8420
rect 14571 8371 14613 8380
rect 14572 8168 14612 8371
rect 14572 8119 14612 8128
rect 14475 8084 14517 8093
rect 14475 8044 14476 8084
rect 14516 8044 14517 8084
rect 14475 8035 14517 8044
rect 14428 7958 14468 7967
rect 14428 7916 14468 7918
rect 14428 7876 14612 7916
rect 14284 7792 14420 7832
rect 14091 7748 14133 7757
rect 14091 7708 14092 7748
rect 14132 7708 14133 7748
rect 14091 7699 14133 7708
rect 14380 7505 14420 7792
rect 14379 7496 14421 7505
rect 14379 7456 14380 7496
rect 14420 7456 14421 7496
rect 14379 7447 14421 7456
rect 14283 7412 14325 7421
rect 14283 7372 14284 7412
rect 14324 7372 14325 7412
rect 14283 7363 14325 7372
rect 14284 6656 14324 7363
rect 14380 7160 14420 7447
rect 14572 7412 14612 7876
rect 14572 7363 14612 7372
rect 14668 7244 14708 9883
rect 15052 9680 15092 10144
rect 15052 9631 15092 9640
rect 14859 9512 14901 9521
rect 14859 9472 14860 9512
rect 14900 9472 14901 9512
rect 14859 9463 14901 9472
rect 14860 9353 14900 9463
rect 14859 9344 14901 9353
rect 14859 9304 14860 9344
rect 14900 9304 14901 9344
rect 14859 9295 14901 9304
rect 15148 8261 15188 11320
rect 15436 10352 15476 13747
rect 15627 13376 15669 13385
rect 15627 13336 15628 13376
rect 15668 13336 15669 13376
rect 15627 13327 15669 13336
rect 15531 13208 15573 13217
rect 15531 13168 15532 13208
rect 15572 13168 15573 13208
rect 15531 13159 15573 13168
rect 15244 10312 15476 10352
rect 15147 8252 15189 8261
rect 15147 8212 15148 8252
rect 15188 8212 15189 8252
rect 15147 8203 15189 8212
rect 15052 8000 15092 8009
rect 14764 7960 15052 8000
rect 14764 7412 14804 7960
rect 15052 7951 15092 7960
rect 15148 8000 15188 8009
rect 15244 8000 15284 10312
rect 15340 10184 15380 10193
rect 15340 8933 15380 10144
rect 15436 10184 15476 10312
rect 15436 10135 15476 10144
rect 15339 8924 15381 8933
rect 15339 8884 15340 8924
rect 15380 8884 15381 8924
rect 15339 8875 15381 8884
rect 15435 8756 15477 8765
rect 15435 8716 15436 8756
rect 15476 8716 15477 8756
rect 15435 8707 15477 8716
rect 15188 7960 15284 8000
rect 15148 7951 15188 7960
rect 14764 7363 14804 7372
rect 14860 7288 15092 7328
rect 14860 7244 14900 7288
rect 14668 7204 14900 7244
rect 14380 6917 14420 7120
rect 14955 7160 14997 7169
rect 14955 7120 14956 7160
rect 14996 7120 14997 7160
rect 14955 7111 14997 7120
rect 14379 6908 14421 6917
rect 14379 6868 14380 6908
rect 14420 6868 14421 6908
rect 14379 6859 14421 6868
rect 14284 6607 14324 6616
rect 14140 6478 14420 6488
rect 14180 6448 14420 6478
rect 14140 6429 14180 6438
rect 14380 5900 14420 6448
rect 14380 5851 14420 5860
rect 14188 5648 14228 5657
rect 14188 5573 14228 5608
rect 14187 5564 14229 5573
rect 14187 5524 14188 5564
rect 14228 5524 14229 5564
rect 14187 5515 14229 5524
rect 14188 5237 14228 5515
rect 14763 5396 14805 5405
rect 14763 5356 14764 5396
rect 14804 5356 14805 5396
rect 14763 5347 14805 5356
rect 14187 5228 14229 5237
rect 14187 5188 14188 5228
rect 14228 5188 14229 5228
rect 14187 5179 14229 5188
rect 14187 4220 14229 4229
rect 14187 4180 14188 4220
rect 14228 4180 14229 4220
rect 14187 4171 14229 4180
rect 14188 4136 14228 4171
rect 14764 4145 14804 5347
rect 14956 4229 14996 7111
rect 15052 4976 15092 7288
rect 15148 5648 15188 5657
rect 15148 5144 15188 5608
rect 15244 5648 15284 7960
rect 15436 8672 15476 8707
rect 15532 8681 15572 13159
rect 15628 12629 15668 13327
rect 15724 13217 15764 14008
rect 15723 13208 15765 13217
rect 15723 13168 15724 13208
rect 15764 13168 15765 13208
rect 15723 13159 15765 13168
rect 15627 12620 15669 12629
rect 15627 12580 15628 12620
rect 15668 12580 15669 12620
rect 15627 12571 15669 12580
rect 15723 10436 15765 10445
rect 15723 10396 15724 10436
rect 15764 10396 15765 10436
rect 15820 10436 15860 17863
rect 15916 17585 15956 18535
rect 16012 17753 16052 21307
rect 16011 17744 16053 17753
rect 16011 17704 16012 17744
rect 16052 17704 16053 17744
rect 16011 17695 16053 17704
rect 15915 17576 15957 17585
rect 15915 17536 15916 17576
rect 15956 17536 15957 17576
rect 15915 17527 15957 17536
rect 15915 17156 15957 17165
rect 15915 17116 15916 17156
rect 15956 17116 15957 17156
rect 15915 17107 15957 17116
rect 15916 13721 15956 17107
rect 16012 13889 16052 17695
rect 16108 14552 16148 21391
rect 16203 20768 16245 20777
rect 16203 20728 16204 20768
rect 16244 20728 16245 20768
rect 16203 20719 16245 20728
rect 16204 20634 16244 20719
rect 16300 20525 16340 22828
rect 16395 22616 16437 22625
rect 16395 22576 16396 22616
rect 16436 22576 16437 22616
rect 16395 22567 16437 22576
rect 16396 22289 16436 22567
rect 16395 22280 16437 22289
rect 16395 22240 16396 22280
rect 16436 22240 16437 22280
rect 16395 22231 16437 22240
rect 16396 21449 16436 22231
rect 16588 21869 16628 24424
rect 17068 23969 17108 24592
rect 17164 24632 17204 25423
rect 17356 24809 17396 25432
rect 17355 24800 17397 24809
rect 17355 24760 17356 24800
rect 17396 24760 17397 24800
rect 17355 24751 17397 24760
rect 17164 24583 17204 24592
rect 17260 24632 17300 24641
rect 17260 24137 17300 24592
rect 17259 24128 17301 24137
rect 17259 24088 17260 24128
rect 17300 24088 17301 24128
rect 17259 24079 17301 24088
rect 17067 23960 17109 23969
rect 17548 23960 17588 28876
rect 17836 28421 17876 30976
rect 18028 30521 18068 41971
rect 18027 30512 18069 30521
rect 18027 30472 18028 30512
rect 18068 30472 18069 30512
rect 18027 30463 18069 30472
rect 17932 30428 17972 30439
rect 17932 30353 17972 30388
rect 17931 30344 17973 30353
rect 17931 30304 17932 30344
rect 17972 30304 17973 30344
rect 17931 30295 17973 30304
rect 18124 30176 18164 43912
rect 18220 37820 18260 44155
rect 18316 42020 18356 42029
rect 18316 41021 18356 41980
rect 18412 41600 18452 45004
rect 18508 45044 18548 45053
rect 18604 45044 18644 46432
rect 19028 46432 19124 46472
rect 18988 46423 19028 46432
rect 18891 45968 18933 45977
rect 18891 45928 18892 45968
rect 18932 45928 18933 45968
rect 18891 45919 18933 45928
rect 18892 45809 18932 45919
rect 18891 45800 18933 45809
rect 18891 45760 18892 45800
rect 18932 45760 18933 45800
rect 18891 45751 18933 45760
rect 18988 45725 19028 45810
rect 18699 45716 18741 45725
rect 18699 45676 18700 45716
rect 18740 45676 18741 45716
rect 18699 45667 18741 45676
rect 18987 45716 19029 45725
rect 18987 45676 18988 45716
rect 19028 45676 19029 45716
rect 18987 45667 19029 45676
rect 18548 45004 18644 45044
rect 18508 44995 18548 45004
rect 18604 42692 18644 42701
rect 18508 42652 18604 42692
rect 18508 42029 18548 42652
rect 18604 42643 18644 42652
rect 18700 42524 18740 45667
rect 18796 45557 18836 45642
rect 19084 45557 19124 46432
rect 19180 45968 19220 45977
rect 19276 45968 19316 47347
rect 19372 46388 19412 49036
rect 19755 48992 19797 49001
rect 19755 48952 19756 48992
rect 19796 48952 19797 48992
rect 19755 48943 19797 48952
rect 19756 48858 19796 48943
rect 19612 48782 19652 48791
rect 19612 48740 19652 48742
rect 19612 48700 19700 48740
rect 19660 48236 19700 48700
rect 19852 48329 19892 49288
rect 19948 49001 19988 49288
rect 20048 49160 20416 49169
rect 20088 49120 20130 49160
rect 20170 49120 20212 49160
rect 20252 49120 20294 49160
rect 20334 49120 20376 49160
rect 20048 49111 20416 49120
rect 19947 48992 19989 49001
rect 19947 48952 19948 48992
rect 19988 48952 19989 48992
rect 19947 48943 19989 48952
rect 19948 48740 19988 48749
rect 19948 48497 19988 48700
rect 20140 48572 20180 48581
rect 19947 48488 19989 48497
rect 19947 48448 19948 48488
rect 19988 48448 19989 48488
rect 19947 48439 19989 48448
rect 19851 48320 19893 48329
rect 19851 48280 19852 48320
rect 19892 48280 19893 48320
rect 19851 48271 19893 48280
rect 19660 48187 19700 48196
rect 19851 48068 19893 48077
rect 19851 48028 19852 48068
rect 19892 48028 19893 48068
rect 19851 48019 19893 48028
rect 19467 47984 19509 47993
rect 19467 47944 19468 47984
rect 19508 47944 19509 47984
rect 19467 47935 19509 47944
rect 19468 47850 19508 47935
rect 19852 47934 19892 48019
rect 20140 47825 20180 48532
rect 20044 47816 20084 47825
rect 19948 47776 20044 47816
rect 19467 47564 19509 47573
rect 19467 47524 19468 47564
rect 19508 47524 19509 47564
rect 19467 47515 19509 47524
rect 19468 46733 19508 47515
rect 19852 47312 19892 47323
rect 19852 47237 19892 47272
rect 19851 47228 19893 47237
rect 19851 47188 19852 47228
rect 19892 47188 19893 47228
rect 19851 47179 19893 47188
rect 19948 46985 19988 47776
rect 20044 47767 20084 47776
rect 20139 47816 20181 47825
rect 20139 47776 20140 47816
rect 20180 47776 20181 47816
rect 20139 47767 20181 47776
rect 20048 47648 20416 47657
rect 20088 47608 20130 47648
rect 20170 47608 20212 47648
rect 20252 47608 20294 47648
rect 20334 47608 20376 47648
rect 20048 47599 20416 47608
rect 20044 47060 20084 47069
rect 19947 46976 19989 46985
rect 19947 46936 19948 46976
rect 19988 46936 19989 46976
rect 19947 46927 19989 46936
rect 20044 46808 20084 47020
rect 19564 46768 20084 46808
rect 19467 46724 19509 46733
rect 19467 46684 19468 46724
rect 19508 46684 19509 46724
rect 19467 46675 19509 46684
rect 19564 46556 19604 46768
rect 19516 46516 19604 46556
rect 19851 46556 19893 46565
rect 19851 46516 19852 46556
rect 19892 46516 19893 46556
rect 19516 46514 19556 46516
rect 19851 46507 19893 46516
rect 19516 46465 19556 46474
rect 19852 46422 19892 46507
rect 19372 46348 19508 46388
rect 19220 45928 19316 45968
rect 19180 45919 19220 45928
rect 19275 45800 19317 45809
rect 19275 45760 19276 45800
rect 19316 45760 19317 45800
rect 19275 45751 19317 45760
rect 18795 45548 18837 45557
rect 18795 45508 18796 45548
rect 18836 45508 18837 45548
rect 18795 45499 18837 45508
rect 19083 45548 19125 45557
rect 19083 45508 19084 45548
rect 19124 45508 19125 45548
rect 19083 45499 19125 45508
rect 18808 45380 19176 45389
rect 18848 45340 18890 45380
rect 18930 45340 18972 45380
rect 19012 45340 19054 45380
rect 19094 45340 19136 45380
rect 18808 45331 19176 45340
rect 18891 45212 18933 45221
rect 18891 45172 18892 45212
rect 18932 45172 18933 45212
rect 18891 45163 18933 45172
rect 18892 44801 18932 45163
rect 18987 45128 19029 45137
rect 18987 45088 18988 45128
rect 19028 45088 19029 45128
rect 18987 45079 19029 45088
rect 18988 44969 19028 45079
rect 18987 44960 19029 44969
rect 18987 44920 18988 44960
rect 19028 44920 19029 44960
rect 18987 44911 19029 44920
rect 18988 44826 19028 44911
rect 18891 44792 18933 44801
rect 18891 44752 18892 44792
rect 18932 44752 18933 44792
rect 18891 44743 18933 44752
rect 18808 43868 19176 43877
rect 18848 43828 18890 43868
rect 18930 43828 18972 43868
rect 19012 43828 19054 43868
rect 19094 43828 19136 43868
rect 18808 43819 19176 43828
rect 19179 43700 19221 43709
rect 19179 43660 19180 43700
rect 19220 43660 19221 43700
rect 19179 43651 19221 43660
rect 19180 43566 19220 43651
rect 18987 43532 19029 43541
rect 18987 43492 18988 43532
rect 19028 43492 19029 43532
rect 19276 43532 19316 45751
rect 19372 45716 19412 45725
rect 19372 45557 19412 45676
rect 19371 45548 19413 45557
rect 19371 45508 19372 45548
rect 19412 45508 19413 45548
rect 19371 45499 19413 45508
rect 19468 45128 19508 46348
rect 20044 46313 20084 46398
rect 19660 46304 19700 46313
rect 19563 45884 19605 45893
rect 19563 45844 19564 45884
rect 19604 45844 19605 45884
rect 19563 45835 19605 45844
rect 19564 45716 19604 45835
rect 19660 45725 19700 46264
rect 20043 46304 20085 46313
rect 20043 46264 20044 46304
rect 20084 46264 20085 46304
rect 20043 46255 20085 46264
rect 20048 46136 20416 46145
rect 20088 46096 20130 46136
rect 20170 46096 20212 46136
rect 20252 46096 20294 46136
rect 20334 46096 20376 46136
rect 20048 46087 20416 46096
rect 19564 45667 19604 45676
rect 19659 45716 19701 45725
rect 19659 45676 19660 45716
rect 19700 45676 19701 45716
rect 19659 45667 19701 45676
rect 19659 45548 19701 45557
rect 19659 45508 19660 45548
rect 19700 45508 19701 45548
rect 19659 45499 19701 45508
rect 19756 45548 19796 45557
rect 19372 45088 19508 45128
rect 19372 44456 19412 45088
rect 19516 44969 19556 44978
rect 19556 44929 19604 44960
rect 19516 44920 19604 44929
rect 19564 44456 19604 44920
rect 19660 44876 19700 45499
rect 19756 44969 19796 45508
rect 19851 45044 19893 45053
rect 19851 45004 19852 45044
rect 19892 45004 19893 45044
rect 19851 44995 19893 45004
rect 19755 44960 19797 44969
rect 19755 44920 19756 44960
rect 19796 44920 19797 44960
rect 19755 44911 19797 44920
rect 19852 44910 19892 44995
rect 19660 44827 19700 44836
rect 19851 44792 19893 44801
rect 20044 44792 20084 44801
rect 19851 44752 19852 44792
rect 19892 44752 19893 44792
rect 19851 44743 19893 44752
rect 19948 44752 20044 44792
rect 19755 44540 19797 44549
rect 19755 44500 19756 44540
rect 19796 44500 19797 44540
rect 19755 44491 19797 44500
rect 19372 44416 19508 44456
rect 19371 44288 19413 44297
rect 19371 44248 19372 44288
rect 19412 44248 19413 44288
rect 19371 44239 19413 44248
rect 19372 44154 19412 44239
rect 19372 43532 19412 43541
rect 19276 43492 19372 43532
rect 18987 43483 19029 43492
rect 19372 43483 19412 43492
rect 18988 43398 19028 43483
rect 18988 42692 19028 42701
rect 18796 42533 18836 42618
rect 18988 42533 19028 42652
rect 19180 42617 19220 42702
rect 19372 42692 19412 42701
rect 19179 42608 19221 42617
rect 19179 42568 19180 42608
rect 19220 42568 19221 42608
rect 19179 42559 19221 42568
rect 18604 42484 18740 42524
rect 18795 42524 18837 42533
rect 18795 42484 18796 42524
rect 18836 42484 18837 42524
rect 18507 42020 18549 42029
rect 18507 41980 18508 42020
rect 18548 41980 18549 42020
rect 18507 41971 18549 41980
rect 18508 41777 18548 41862
rect 18507 41768 18549 41777
rect 18507 41728 18508 41768
rect 18548 41728 18549 41768
rect 18507 41719 18549 41728
rect 18412 41560 18548 41600
rect 18315 41012 18357 41021
rect 18315 40972 18316 41012
rect 18356 40972 18357 41012
rect 18315 40963 18357 40972
rect 18220 37780 18452 37820
rect 18315 35048 18357 35057
rect 18315 35008 18316 35048
rect 18356 35008 18357 35048
rect 18315 34999 18357 35008
rect 18316 33545 18356 34999
rect 18315 33536 18357 33545
rect 18315 33496 18316 33536
rect 18356 33496 18357 33536
rect 18315 33487 18357 33496
rect 18219 33368 18261 33377
rect 18219 33328 18220 33368
rect 18260 33328 18261 33368
rect 18219 33319 18261 33328
rect 18220 31352 18260 33319
rect 18220 31303 18260 31312
rect 18412 31277 18452 37780
rect 18411 31268 18453 31277
rect 18411 31228 18412 31268
rect 18452 31228 18453 31268
rect 18411 31219 18453 31228
rect 18412 30680 18452 30689
rect 18412 30269 18452 30640
rect 18411 30260 18453 30269
rect 18411 30220 18412 30260
rect 18452 30220 18453 30260
rect 18411 30211 18453 30220
rect 17932 30136 18164 30176
rect 17835 28412 17877 28421
rect 17835 28372 17836 28412
rect 17876 28372 17877 28412
rect 17835 28363 17877 28372
rect 17836 28328 17876 28363
rect 17836 28278 17876 28288
rect 17835 27824 17877 27833
rect 17835 27784 17836 27824
rect 17876 27784 17877 27824
rect 17835 27775 17877 27784
rect 17739 27740 17781 27749
rect 17739 27700 17740 27740
rect 17780 27700 17781 27740
rect 17739 27691 17781 27700
rect 17643 26732 17685 26741
rect 17643 26692 17644 26732
rect 17684 26692 17685 26732
rect 17643 26683 17685 26692
rect 17644 26312 17684 26683
rect 17644 26263 17684 26272
rect 17740 26144 17780 27691
rect 17836 26900 17876 27775
rect 17932 26984 17972 30136
rect 18123 29924 18165 29933
rect 18123 29884 18124 29924
rect 18164 29884 18165 29924
rect 18123 29875 18165 29884
rect 18315 29924 18357 29933
rect 18315 29884 18316 29924
rect 18356 29884 18357 29924
rect 18315 29875 18357 29884
rect 18028 29840 18068 29849
rect 18028 29420 18068 29800
rect 18124 29790 18164 29875
rect 18123 29672 18165 29681
rect 18123 29632 18124 29672
rect 18164 29632 18165 29672
rect 18316 29672 18356 29875
rect 18412 29849 18452 30211
rect 18411 29840 18453 29849
rect 18411 29800 18412 29840
rect 18452 29800 18453 29840
rect 18411 29791 18453 29800
rect 18316 29632 18452 29672
rect 18123 29623 18165 29632
rect 18124 29504 18164 29623
rect 18124 29464 18356 29504
rect 18028 29380 18260 29420
rect 18123 29252 18165 29261
rect 18123 29212 18124 29252
rect 18164 29212 18165 29252
rect 18123 29203 18165 29212
rect 18027 29168 18069 29177
rect 18027 29128 18028 29168
rect 18068 29128 18069 29168
rect 18027 29119 18069 29128
rect 18124 29168 18164 29203
rect 18028 29034 18068 29119
rect 18124 29117 18164 29128
rect 18220 29000 18260 29380
rect 18316 29168 18356 29464
rect 18316 29119 18356 29128
rect 18124 28960 18260 29000
rect 18124 27833 18164 28960
rect 18220 28328 18260 28337
rect 18123 27824 18165 27833
rect 18123 27784 18124 27824
rect 18164 27784 18165 27824
rect 18123 27775 18165 27784
rect 18124 27656 18164 27665
rect 18028 27616 18124 27656
rect 18028 27245 18068 27616
rect 18124 27607 18164 27616
rect 18220 27581 18260 28288
rect 18315 27992 18357 28001
rect 18315 27952 18316 27992
rect 18356 27952 18357 27992
rect 18315 27943 18357 27952
rect 18219 27572 18261 27581
rect 18219 27532 18220 27572
rect 18260 27532 18261 27572
rect 18219 27523 18261 27532
rect 18027 27236 18069 27245
rect 18027 27196 18028 27236
rect 18068 27196 18069 27236
rect 18027 27187 18069 27196
rect 17932 26944 18068 26984
rect 17836 26851 17876 26860
rect 17931 26816 17973 26825
rect 17931 26776 17932 26816
rect 17972 26776 17973 26816
rect 17931 26767 17973 26776
rect 17932 26682 17972 26767
rect 18028 26564 18068 26944
rect 17932 26524 18068 26564
rect 17836 26144 17876 26153
rect 17740 26104 17836 26144
rect 17836 25229 17876 26104
rect 17835 25220 17877 25229
rect 17835 25180 17836 25220
rect 17876 25180 17877 25220
rect 17835 25171 17877 25180
rect 17836 23969 17876 25171
rect 17067 23920 17068 23960
rect 17108 23920 17109 23960
rect 17067 23911 17109 23920
rect 17356 23920 17588 23960
rect 17835 23960 17877 23969
rect 17835 23920 17836 23960
rect 17876 23920 17877 23960
rect 16972 23792 17012 23801
rect 16779 23540 16821 23549
rect 16779 23500 16780 23540
rect 16820 23500 16821 23540
rect 16779 23491 16821 23500
rect 16683 23456 16725 23465
rect 16683 23416 16684 23456
rect 16724 23416 16725 23456
rect 16683 23407 16725 23416
rect 16587 21860 16629 21869
rect 16587 21820 16588 21860
rect 16628 21820 16629 21860
rect 16587 21811 16629 21820
rect 16491 21776 16533 21785
rect 16491 21736 16492 21776
rect 16532 21736 16533 21776
rect 16491 21727 16533 21736
rect 16395 21440 16437 21449
rect 16395 21400 16396 21440
rect 16436 21400 16437 21440
rect 16395 21391 16437 21400
rect 16492 20768 16532 21727
rect 16684 21608 16724 23407
rect 16780 23120 16820 23491
rect 16780 23071 16820 23080
rect 16972 22709 17012 23752
rect 16971 22700 17013 22709
rect 16971 22660 16972 22700
rect 17012 22660 17013 22700
rect 16971 22651 17013 22660
rect 17356 22625 17396 23920
rect 17835 23911 17877 23920
rect 17452 23797 17492 23806
rect 17452 23297 17492 23757
rect 17643 23708 17685 23717
rect 17643 23668 17644 23708
rect 17684 23668 17685 23708
rect 17643 23659 17685 23668
rect 17644 23574 17684 23659
rect 17836 23549 17876 23911
rect 17835 23540 17877 23549
rect 17835 23500 17836 23540
rect 17876 23500 17877 23540
rect 17835 23491 17877 23500
rect 17835 23372 17877 23381
rect 17835 23332 17836 23372
rect 17876 23332 17877 23372
rect 17835 23323 17877 23332
rect 17451 23288 17493 23297
rect 17451 23248 17452 23288
rect 17492 23248 17588 23288
rect 17451 23239 17493 23248
rect 17355 22616 17397 22625
rect 17355 22576 17356 22616
rect 17396 22576 17397 22616
rect 17355 22567 17397 22576
rect 17451 22532 17493 22541
rect 17451 22492 17452 22532
rect 17492 22492 17493 22532
rect 17451 22483 17493 22492
rect 16684 21559 16724 21568
rect 16972 22280 17012 22289
rect 16587 21524 16629 21533
rect 16587 21484 16588 21524
rect 16628 21484 16629 21524
rect 16587 21475 16629 21484
rect 16299 20516 16341 20525
rect 16299 20476 16300 20516
rect 16340 20476 16341 20516
rect 16299 20467 16341 20476
rect 16492 20180 16532 20728
rect 16588 20768 16628 21475
rect 16876 20936 16916 20945
rect 16876 20777 16916 20896
rect 16588 20719 16628 20728
rect 16875 20768 16917 20777
rect 16875 20728 16876 20768
rect 16916 20728 16917 20768
rect 16875 20719 16917 20728
rect 16779 20684 16821 20693
rect 16779 20644 16780 20684
rect 16820 20644 16821 20684
rect 16779 20635 16821 20644
rect 16396 20140 16532 20180
rect 16299 19004 16341 19013
rect 16299 18964 16300 19004
rect 16340 18964 16341 19004
rect 16299 18955 16341 18964
rect 16203 18752 16245 18761
rect 16203 18712 16204 18752
rect 16244 18712 16245 18752
rect 16203 18703 16245 18712
rect 16204 17165 16244 18703
rect 16203 17156 16245 17165
rect 16203 17116 16204 17156
rect 16244 17116 16245 17156
rect 16203 17107 16245 17116
rect 16203 16904 16245 16913
rect 16203 16864 16204 16904
rect 16244 16864 16245 16904
rect 16203 16855 16245 16864
rect 16204 16409 16244 16855
rect 16300 16493 16340 18955
rect 16299 16484 16341 16493
rect 16299 16444 16300 16484
rect 16340 16444 16341 16484
rect 16396 16484 16436 20140
rect 16780 17660 16820 20635
rect 16972 20609 17012 22240
rect 17452 22280 17492 22483
rect 17068 22112 17108 22121
rect 16971 20600 17013 20609
rect 16971 20560 16972 20600
rect 17012 20560 17013 20600
rect 16971 20551 17013 20560
rect 16876 20096 16916 20107
rect 16876 20021 16916 20056
rect 16875 20012 16917 20021
rect 16875 19972 16876 20012
rect 16916 19972 16917 20012
rect 16875 19963 16917 19972
rect 16972 19928 17012 20551
rect 17068 20105 17108 22072
rect 17356 21692 17396 21701
rect 17164 21594 17204 21603
rect 17164 21449 17204 21554
rect 17163 21440 17205 21449
rect 17163 21400 17164 21440
rect 17204 21400 17205 21440
rect 17163 21391 17205 21400
rect 17356 20861 17396 21652
rect 17163 20852 17205 20861
rect 17163 20812 17164 20852
rect 17204 20812 17205 20852
rect 17163 20803 17205 20812
rect 17355 20852 17397 20861
rect 17355 20812 17356 20852
rect 17396 20812 17397 20852
rect 17355 20803 17397 20812
rect 17164 20768 17204 20803
rect 17164 20717 17204 20728
rect 17452 20768 17492 22240
rect 17548 22280 17588 23248
rect 17548 22231 17588 22240
rect 17739 22112 17781 22121
rect 17739 22072 17740 22112
rect 17780 22072 17781 22112
rect 17739 22063 17781 22072
rect 17740 21978 17780 22063
rect 17740 21608 17780 21617
rect 17836 21608 17876 23323
rect 17780 21568 17876 21608
rect 17740 21524 17780 21568
rect 17644 21484 17780 21524
rect 17547 21440 17589 21449
rect 17547 21400 17548 21440
rect 17588 21400 17589 21440
rect 17547 21391 17589 21400
rect 17548 21306 17588 21391
rect 17452 20719 17492 20728
rect 17547 20684 17589 20693
rect 17547 20644 17548 20684
rect 17588 20644 17589 20684
rect 17547 20635 17589 20644
rect 17548 20550 17588 20635
rect 17163 20516 17205 20525
rect 17163 20476 17164 20516
rect 17204 20476 17205 20516
rect 17163 20467 17205 20476
rect 17067 20096 17109 20105
rect 17067 20056 17068 20096
rect 17108 20056 17109 20096
rect 17067 20047 17109 20056
rect 17068 19928 17108 19937
rect 16972 19888 17068 19928
rect 17068 19879 17108 19888
rect 16875 19760 16917 19769
rect 16875 19720 16876 19760
rect 16916 19720 16917 19760
rect 16875 19711 16917 19720
rect 16876 19349 16916 19711
rect 16875 19340 16917 19349
rect 16875 19300 16876 19340
rect 16916 19300 16917 19340
rect 16875 19291 16917 19300
rect 16684 17620 16820 17660
rect 16876 17744 16916 19291
rect 16972 18584 17012 18593
rect 16972 17996 17012 18544
rect 17068 18584 17108 18593
rect 17164 18584 17204 20467
rect 17355 20348 17397 20357
rect 17355 20308 17356 20348
rect 17396 20308 17397 20348
rect 17644 20348 17684 21484
rect 17836 20936 17876 20945
rect 17740 20896 17836 20936
rect 17740 20525 17780 20896
rect 17836 20887 17876 20896
rect 17835 20684 17877 20693
rect 17835 20644 17836 20684
rect 17876 20644 17877 20684
rect 17835 20635 17877 20644
rect 17739 20516 17781 20525
rect 17739 20476 17740 20516
rect 17780 20476 17781 20516
rect 17739 20467 17781 20476
rect 17836 20432 17876 20635
rect 17932 20516 17972 26524
rect 18316 26480 18356 27943
rect 18412 27161 18452 29632
rect 18411 27152 18453 27161
rect 18411 27112 18412 27152
rect 18452 27112 18453 27152
rect 18411 27103 18453 27112
rect 18412 26816 18452 27103
rect 18412 26767 18452 26776
rect 18124 26440 18356 26480
rect 18124 24464 18164 26440
rect 18219 25220 18261 25229
rect 18219 25180 18220 25220
rect 18260 25180 18261 25220
rect 18219 25171 18261 25180
rect 18220 24632 18260 25171
rect 18508 24632 18548 41560
rect 18604 38156 18644 42484
rect 18795 42475 18837 42484
rect 18987 42524 19029 42533
rect 18987 42484 18988 42524
rect 19028 42484 19029 42524
rect 18987 42475 19029 42484
rect 18808 42356 19176 42365
rect 18848 42316 18890 42356
rect 18930 42316 18972 42356
rect 19012 42316 19054 42356
rect 19094 42316 19136 42356
rect 18808 42307 19176 42316
rect 19275 42188 19317 42197
rect 19275 42148 19276 42188
rect 19316 42148 19317 42188
rect 19275 42139 19317 42148
rect 18891 42104 18933 42113
rect 18891 42064 18892 42104
rect 18932 42064 18933 42104
rect 18891 42055 18933 42064
rect 18700 42020 18740 42029
rect 18700 41861 18740 41980
rect 18892 41970 18932 42055
rect 19276 42054 19316 42139
rect 19084 42020 19124 42029
rect 18988 41980 19084 42020
rect 18699 41852 18741 41861
rect 18699 41812 18700 41852
rect 18740 41812 18741 41852
rect 18699 41803 18741 41812
rect 18891 41432 18933 41441
rect 18988 41432 19028 41980
rect 19084 41971 19124 41980
rect 19372 41609 19412 42652
rect 19468 42608 19508 44416
rect 19564 44407 19604 44416
rect 19756 44204 19796 44491
rect 19756 44155 19796 44164
rect 19564 43280 19604 43289
rect 19604 43240 19700 43280
rect 19564 43231 19604 43240
rect 19564 42608 19604 42617
rect 19468 42568 19564 42608
rect 19564 42559 19604 42568
rect 19660 42281 19700 43240
rect 19755 42692 19797 42701
rect 19755 42652 19756 42692
rect 19796 42652 19797 42692
rect 19755 42643 19797 42652
rect 19756 42558 19796 42643
rect 19659 42272 19701 42281
rect 19659 42232 19660 42272
rect 19700 42232 19701 42272
rect 19659 42223 19701 42232
rect 19852 42197 19892 44743
rect 19948 44297 19988 44752
rect 20044 44743 20084 44752
rect 20048 44624 20416 44633
rect 20088 44584 20130 44624
rect 20170 44584 20212 44624
rect 20252 44584 20294 44624
rect 20334 44584 20376 44624
rect 20048 44575 20416 44584
rect 19947 44288 19989 44297
rect 19947 44248 19948 44288
rect 19988 44248 19989 44288
rect 19947 44239 19989 44248
rect 19948 44036 19988 44045
rect 19948 43625 19988 43996
rect 19947 43616 19989 43625
rect 19947 43576 19948 43616
rect 19988 43576 19989 43616
rect 19947 43567 19989 43576
rect 19947 43280 19989 43289
rect 19947 43240 19948 43280
rect 19988 43240 19989 43280
rect 19947 43231 19989 43240
rect 19948 42692 19988 43231
rect 20048 43112 20416 43121
rect 20088 43072 20130 43112
rect 20170 43072 20212 43112
rect 20252 43072 20294 43112
rect 20334 43072 20376 43112
rect 20048 43063 20416 43072
rect 19948 42652 20084 42692
rect 19948 42524 19988 42533
rect 19851 42188 19893 42197
rect 19851 42148 19852 42188
rect 19892 42148 19893 42188
rect 19851 42139 19893 42148
rect 19468 42020 19508 42029
rect 19852 42020 19892 42029
rect 19508 41980 19604 42020
rect 19468 41971 19508 41980
rect 19371 41600 19413 41609
rect 19371 41560 19372 41600
rect 19412 41560 19413 41600
rect 19371 41551 19413 41560
rect 18891 41392 18892 41432
rect 18932 41392 19028 41432
rect 18891 41383 18933 41392
rect 18892 41180 18932 41189
rect 18892 41021 18932 41140
rect 18988 41105 19028 41392
rect 19083 41432 19125 41441
rect 19083 41392 19084 41432
rect 19124 41392 19125 41432
rect 19083 41383 19125 41392
rect 19084 41298 19124 41383
rect 19371 41348 19413 41357
rect 19371 41308 19372 41348
rect 19412 41308 19413 41348
rect 19371 41299 19413 41308
rect 19275 41180 19317 41189
rect 19275 41140 19276 41180
rect 19316 41140 19317 41180
rect 19275 41131 19317 41140
rect 18987 41096 19029 41105
rect 18987 41056 18988 41096
rect 19028 41056 19029 41096
rect 18987 41047 19029 41056
rect 19276 41046 19316 41131
rect 18891 41012 18933 41021
rect 18891 40972 18892 41012
rect 18932 40972 18933 41012
rect 18891 40963 18933 40972
rect 18808 40844 19176 40853
rect 18848 40804 18890 40844
rect 18930 40804 18972 40844
rect 19012 40804 19054 40844
rect 19094 40804 19136 40844
rect 18808 40795 19176 40804
rect 19083 40676 19125 40685
rect 19083 40636 19084 40676
rect 19124 40636 19125 40676
rect 19083 40627 19125 40636
rect 19084 40542 19124 40627
rect 18892 40508 18932 40517
rect 18892 39500 18932 40468
rect 19276 40508 19316 40517
rect 19372 40508 19412 41299
rect 19467 41012 19509 41021
rect 19467 40972 19468 41012
rect 19508 40972 19509 41012
rect 19467 40963 19509 40972
rect 19468 40878 19508 40963
rect 19467 40676 19509 40685
rect 19467 40636 19468 40676
rect 19508 40636 19509 40676
rect 19467 40627 19509 40636
rect 19468 40542 19508 40627
rect 19564 40601 19604 41980
rect 19756 41980 19852 42020
rect 19659 41768 19701 41777
rect 19659 41728 19660 41768
rect 19700 41728 19701 41768
rect 19659 41719 19701 41728
rect 19660 41634 19700 41719
rect 19659 41516 19701 41525
rect 19659 41476 19660 41516
rect 19700 41476 19701 41516
rect 19659 41467 19701 41476
rect 19660 41180 19700 41467
rect 19660 41131 19700 41140
rect 19563 40592 19605 40601
rect 19563 40552 19564 40592
rect 19604 40552 19605 40592
rect 19563 40543 19605 40552
rect 19316 40468 19412 40508
rect 19659 40508 19701 40517
rect 19659 40468 19660 40508
rect 19700 40468 19701 40508
rect 19276 40459 19316 40468
rect 19659 40459 19701 40468
rect 19660 40374 19700 40459
rect 18987 40172 19029 40181
rect 18987 40132 18988 40172
rect 19028 40132 19029 40172
rect 18987 40123 19029 40132
rect 18988 39668 19028 40123
rect 19563 40004 19605 40013
rect 19563 39964 19564 40004
rect 19604 39964 19605 40004
rect 19563 39955 19605 39964
rect 19564 39920 19604 39955
rect 19564 39869 19604 39880
rect 19756 39836 19796 41980
rect 19852 41971 19892 41980
rect 19851 41852 19893 41861
rect 19851 41812 19852 41852
rect 19892 41812 19893 41852
rect 19851 41803 19893 41812
rect 19852 41516 19892 41803
rect 19948 41693 19988 42484
rect 20044 42188 20084 42652
rect 20044 42139 20084 42148
rect 19947 41684 19989 41693
rect 19947 41644 19948 41684
rect 19988 41644 19989 41684
rect 19947 41635 19989 41644
rect 20048 41600 20416 41609
rect 20088 41560 20130 41600
rect 20170 41560 20212 41600
rect 20252 41560 20294 41600
rect 20334 41560 20376 41600
rect 20048 41551 20416 41560
rect 19852 41476 19988 41516
rect 19851 41012 19893 41021
rect 19851 40972 19852 41012
rect 19892 40972 19893 41012
rect 19851 40963 19893 40972
rect 19852 40878 19892 40963
rect 19948 40517 19988 41476
rect 20043 41264 20085 41273
rect 20043 41224 20044 41264
rect 20084 41224 20085 41264
rect 20043 41215 20085 41224
rect 19947 40508 19989 40517
rect 19947 40468 19948 40508
rect 19988 40468 19989 40508
rect 19947 40459 19989 40468
rect 20044 40508 20084 41215
rect 20044 40459 20084 40468
rect 19851 40256 19893 40265
rect 19851 40216 19852 40256
rect 19892 40216 19893 40256
rect 19851 40207 19893 40216
rect 20236 40256 20276 40265
rect 20276 40216 20564 40256
rect 20236 40207 20276 40216
rect 19852 40122 19892 40207
rect 20048 40088 20416 40097
rect 20088 40048 20130 40088
rect 20170 40048 20212 40088
rect 20252 40048 20294 40088
rect 20334 40048 20376 40088
rect 20048 40039 20416 40048
rect 19947 39920 19989 39929
rect 19947 39880 19948 39920
rect 19988 39880 19989 39920
rect 19947 39871 19989 39880
rect 19660 39796 19796 39836
rect 19371 39752 19413 39761
rect 19371 39712 19372 39752
rect 19412 39712 19413 39752
rect 19371 39703 19413 39712
rect 19563 39752 19605 39761
rect 19563 39712 19564 39752
rect 19604 39712 19605 39752
rect 19563 39703 19605 39712
rect 18988 39619 19028 39628
rect 19372 39668 19412 39703
rect 19372 39617 19412 39628
rect 18700 39460 18932 39500
rect 19180 39500 19220 39509
rect 19371 39500 19413 39509
rect 19220 39460 19316 39500
rect 18700 38501 18740 39460
rect 19180 39451 19220 39460
rect 18808 39332 19176 39341
rect 18848 39292 18890 39332
rect 18930 39292 18972 39332
rect 19012 39292 19054 39332
rect 19094 39292 19136 39332
rect 18808 39283 19176 39292
rect 19276 38921 19316 39460
rect 19371 39460 19372 39500
rect 19412 39460 19413 39500
rect 19371 39451 19413 39460
rect 19372 38996 19412 39451
rect 19564 39248 19604 39703
rect 19660 39425 19700 39796
rect 19948 39786 19988 39871
rect 19755 39668 19797 39677
rect 19755 39628 19756 39668
rect 19796 39628 19797 39668
rect 19755 39619 19797 39628
rect 19756 39534 19796 39619
rect 20524 39593 20564 40216
rect 20523 39584 20565 39593
rect 20523 39544 20524 39584
rect 20564 39544 20565 39584
rect 20523 39535 20565 39544
rect 19659 39416 19701 39425
rect 19659 39376 19660 39416
rect 19700 39376 19701 39416
rect 19659 39367 19701 39376
rect 19564 39208 19700 39248
rect 19372 38947 19412 38956
rect 19275 38912 19317 38921
rect 19275 38872 19276 38912
rect 19316 38872 19317 38912
rect 19275 38863 19317 38872
rect 19564 38744 19604 38753
rect 18699 38492 18741 38501
rect 18699 38452 18700 38492
rect 18740 38452 18741 38492
rect 18699 38443 18741 38452
rect 19275 38408 19317 38417
rect 19275 38368 19276 38408
rect 19316 38368 19317 38408
rect 19275 38359 19317 38368
rect 18604 38107 18644 38116
rect 18796 37988 18836 37997
rect 18700 37948 18796 37988
rect 18700 37577 18740 37948
rect 18796 37939 18836 37948
rect 18808 37820 19176 37829
rect 18848 37780 18890 37820
rect 18930 37780 18972 37820
rect 19012 37780 19054 37820
rect 19094 37780 19136 37820
rect 18808 37771 19176 37780
rect 18699 37568 18741 37577
rect 18699 37528 18700 37568
rect 18740 37528 18741 37568
rect 18699 37519 18741 37528
rect 18988 37484 19028 37493
rect 19276 37484 19316 38359
rect 19564 38249 19604 38704
rect 19563 38240 19605 38249
rect 19563 38200 19564 38240
rect 19604 38200 19605 38240
rect 19563 38191 19605 38200
rect 19372 38156 19412 38165
rect 19372 37820 19412 38116
rect 19563 38072 19605 38081
rect 19563 38032 19564 38072
rect 19604 38032 19605 38072
rect 19563 38023 19605 38032
rect 19564 37938 19604 38023
rect 19372 37780 19508 37820
rect 19028 37444 19316 37484
rect 19372 37484 19412 37493
rect 18988 37435 19028 37444
rect 18987 37316 19029 37325
rect 18987 37276 18988 37316
rect 19028 37276 19029 37316
rect 18987 37267 19029 37276
rect 18891 37232 18933 37241
rect 18891 37192 18892 37232
rect 18932 37192 18933 37232
rect 18891 37183 18933 37192
rect 18892 36485 18932 37183
rect 18988 36644 19028 37267
rect 19180 37232 19220 37241
rect 19180 36905 19220 37192
rect 19179 36896 19221 36905
rect 19179 36856 19180 36896
rect 19220 36856 19221 36896
rect 19179 36847 19221 36856
rect 19372 36812 19412 37444
rect 19468 37241 19508 37780
rect 19564 37568 19604 37579
rect 19564 37493 19604 37528
rect 19563 37484 19605 37493
rect 19563 37444 19564 37484
rect 19604 37444 19605 37484
rect 19563 37435 19605 37444
rect 19660 37325 19700 39208
rect 20048 38576 20416 38585
rect 20088 38536 20130 38576
rect 20170 38536 20212 38576
rect 20252 38536 20294 38576
rect 20334 38536 20376 38576
rect 20048 38527 20416 38536
rect 19947 37652 19989 37661
rect 19947 37612 19948 37652
rect 19988 37612 19989 37652
rect 19947 37603 19989 37612
rect 19948 37518 19988 37603
rect 19756 37484 19796 37493
rect 19659 37316 19701 37325
rect 19659 37276 19660 37316
rect 19700 37276 19701 37316
rect 19659 37267 19701 37276
rect 19467 37232 19509 37241
rect 19467 37192 19468 37232
rect 19508 37192 19509 37232
rect 19467 37183 19509 37192
rect 19756 37157 19796 37444
rect 19755 37148 19797 37157
rect 19755 37108 19756 37148
rect 19796 37108 19797 37148
rect 19755 37099 19797 37108
rect 20048 37064 20416 37073
rect 20088 37024 20130 37064
rect 20170 37024 20212 37064
rect 20252 37024 20294 37064
rect 20334 37024 20376 37064
rect 20048 37015 20416 37024
rect 19564 36896 19604 36907
rect 19564 36821 19604 36856
rect 19563 36812 19605 36821
rect 19372 36772 19508 36812
rect 18988 36595 19028 36604
rect 19371 36644 19413 36653
rect 19371 36604 19372 36644
rect 19412 36604 19413 36644
rect 19371 36595 19413 36604
rect 19372 36510 19412 36595
rect 18891 36476 18933 36485
rect 18891 36436 18892 36476
rect 18932 36436 18933 36476
rect 18891 36427 18933 36436
rect 19180 36476 19220 36485
rect 19220 36436 19316 36476
rect 19180 36427 19220 36436
rect 18808 36308 19176 36317
rect 18848 36268 18890 36308
rect 18930 36268 18972 36308
rect 19012 36268 19054 36308
rect 19094 36268 19136 36308
rect 18808 36259 19176 36268
rect 19276 36233 19316 36436
rect 19275 36224 19317 36233
rect 19275 36184 19276 36224
rect 19316 36184 19317 36224
rect 19275 36175 19317 36184
rect 19179 36056 19221 36065
rect 19179 36016 19180 36056
rect 19220 36016 19221 36056
rect 19179 36007 19221 36016
rect 18988 35972 19028 35981
rect 18892 35932 18988 35972
rect 18892 34964 18932 35932
rect 18988 35923 19028 35932
rect 19180 35922 19220 36007
rect 19372 35972 19412 35981
rect 19276 35932 19372 35972
rect 19179 35300 19221 35309
rect 19179 35260 19180 35300
rect 19220 35260 19221 35300
rect 19179 35251 19221 35260
rect 18988 35132 19028 35141
rect 18988 35057 19028 35092
rect 18977 35048 19028 35057
rect 18977 35008 18978 35048
rect 19018 35008 19028 35048
rect 19180 35048 19220 35251
rect 18977 34999 19019 35008
rect 19180 34999 19220 35008
rect 18700 34924 18932 34964
rect 18700 33377 18740 34924
rect 18808 34796 19176 34805
rect 18848 34756 18890 34796
rect 18930 34756 18972 34796
rect 19012 34756 19054 34796
rect 19094 34756 19136 34796
rect 18808 34747 19176 34756
rect 18699 33368 18741 33377
rect 18699 33328 18700 33368
rect 18740 33328 18741 33368
rect 18699 33319 18741 33328
rect 18808 33284 19176 33293
rect 18848 33244 18890 33284
rect 18930 33244 18972 33284
rect 19012 33244 19054 33284
rect 19094 33244 19136 33284
rect 18808 33235 19176 33244
rect 18808 31772 19176 31781
rect 18848 31732 18890 31772
rect 18930 31732 18972 31772
rect 19012 31732 19054 31772
rect 19094 31732 19136 31772
rect 18808 31723 19176 31732
rect 19276 31613 19316 35932
rect 19372 35923 19412 35932
rect 19371 35132 19413 35141
rect 19371 35092 19372 35132
rect 19412 35092 19413 35132
rect 19371 35083 19413 35092
rect 19372 34998 19412 35083
rect 19468 34889 19508 36772
rect 19563 36772 19564 36812
rect 19604 36772 19605 36812
rect 19563 36763 19605 36772
rect 19659 36644 19701 36653
rect 19659 36604 19660 36644
rect 19700 36604 19701 36644
rect 19659 36595 19701 36604
rect 19563 36308 19605 36317
rect 19563 36268 19564 36308
rect 19604 36268 19605 36308
rect 19563 36259 19605 36268
rect 19564 36140 19604 36259
rect 19564 36091 19604 36100
rect 19563 35048 19605 35057
rect 19563 35008 19564 35048
rect 19604 35008 19605 35048
rect 19563 34999 19605 35008
rect 19564 34914 19604 34999
rect 19467 34880 19509 34889
rect 19467 34840 19468 34880
rect 19508 34840 19509 34880
rect 19467 34831 19509 34840
rect 19563 34628 19605 34637
rect 19563 34588 19564 34628
rect 19604 34588 19605 34628
rect 19563 34579 19605 34588
rect 19564 34494 19604 34579
rect 19372 34460 19412 34469
rect 19372 34049 19412 34420
rect 19371 34040 19413 34049
rect 19371 34000 19372 34040
rect 19412 34000 19413 34040
rect 19371 33991 19413 34000
rect 19660 32285 19700 36595
rect 20620 36065 20660 59695
rect 20716 48581 20756 61711
rect 20812 59837 20852 78511
rect 20907 75872 20949 75881
rect 20907 75832 20908 75872
rect 20948 75832 20949 75872
rect 20907 75823 20949 75832
rect 20811 59828 20853 59837
rect 20811 59788 20812 59828
rect 20852 59788 20853 59828
rect 20811 59779 20853 59788
rect 20908 56813 20948 75823
rect 21387 75200 21429 75209
rect 21387 75160 21388 75200
rect 21428 75160 21429 75200
rect 21387 75151 21429 75160
rect 21003 73184 21045 73193
rect 21003 73144 21004 73184
rect 21044 73144 21045 73184
rect 21003 73135 21045 73144
rect 21004 62693 21044 73135
rect 21099 63776 21141 63785
rect 21099 63736 21100 63776
rect 21140 63736 21141 63776
rect 21099 63727 21141 63736
rect 21003 62684 21045 62693
rect 21003 62644 21004 62684
rect 21044 62644 21045 62684
rect 21003 62635 21045 62644
rect 21003 59072 21045 59081
rect 21003 59032 21004 59072
rect 21044 59032 21045 59072
rect 21003 59023 21045 59032
rect 20907 56804 20949 56813
rect 20907 56764 20908 56804
rect 20948 56764 20949 56804
rect 20907 56755 20949 56764
rect 20715 48572 20757 48581
rect 20715 48532 20716 48572
rect 20756 48532 20757 48572
rect 20715 48523 20757 48532
rect 20619 36056 20661 36065
rect 20619 36016 20620 36056
rect 20660 36016 20661 36056
rect 20619 36007 20661 36016
rect 19756 35972 19796 35981
rect 19756 35225 19796 35932
rect 19948 35720 19988 35731
rect 19948 35645 19988 35680
rect 19947 35636 19989 35645
rect 19947 35596 19948 35636
rect 19988 35596 19989 35636
rect 19947 35587 19989 35596
rect 20048 35552 20416 35561
rect 20088 35512 20130 35552
rect 20170 35512 20212 35552
rect 20252 35512 20294 35552
rect 20334 35512 20376 35552
rect 20048 35503 20416 35512
rect 21004 35309 21044 59023
rect 21100 36317 21140 63727
rect 21291 62432 21333 62441
rect 21291 62392 21292 62432
rect 21332 62392 21333 62432
rect 21291 62383 21333 62392
rect 21195 61088 21237 61097
rect 21195 61048 21196 61088
rect 21236 61048 21237 61088
rect 21195 61039 21237 61048
rect 21196 39929 21236 61039
rect 21195 39920 21237 39929
rect 21195 39880 21196 39920
rect 21236 39880 21237 39920
rect 21195 39871 21237 39880
rect 21292 38837 21332 62383
rect 21388 61601 21428 75151
rect 21387 61592 21429 61601
rect 21387 61552 21388 61592
rect 21428 61552 21429 61592
rect 21387 61543 21429 61552
rect 21291 38828 21333 38837
rect 21291 38788 21292 38828
rect 21332 38788 21333 38828
rect 21291 38779 21333 38788
rect 21099 36308 21141 36317
rect 21099 36268 21100 36308
rect 21140 36268 21141 36308
rect 21099 36259 21141 36268
rect 21387 35804 21429 35813
rect 21387 35764 21388 35804
rect 21428 35764 21429 35804
rect 21387 35755 21429 35764
rect 21388 35561 21428 35755
rect 21387 35552 21429 35561
rect 21387 35512 21388 35552
rect 21428 35512 21429 35552
rect 21387 35503 21429 35512
rect 21003 35300 21045 35309
rect 21003 35260 21004 35300
rect 21044 35260 21045 35300
rect 21003 35251 21045 35260
rect 19755 35216 19797 35225
rect 19755 35176 19756 35216
rect 19796 35176 19797 35216
rect 19755 35167 19797 35176
rect 19755 34544 19797 34553
rect 19755 34504 19756 34544
rect 19796 34504 19797 34544
rect 19755 34495 19797 34504
rect 19756 34376 19796 34495
rect 19756 34327 19796 34336
rect 19851 34208 19893 34217
rect 19851 34168 19852 34208
rect 19892 34168 19893 34208
rect 19851 34159 19893 34168
rect 19852 34074 19892 34159
rect 20048 34040 20416 34049
rect 20088 34000 20130 34040
rect 20170 34000 20212 34040
rect 20252 34000 20294 34040
rect 20334 34000 20376 34040
rect 20048 33991 20416 34000
rect 20048 32528 20416 32537
rect 20088 32488 20130 32528
rect 20170 32488 20212 32528
rect 20252 32488 20294 32528
rect 20334 32488 20376 32528
rect 20048 32479 20416 32488
rect 19659 32276 19701 32285
rect 19659 32236 19660 32276
rect 19700 32236 19701 32276
rect 19659 32227 19701 32236
rect 19275 31604 19317 31613
rect 19275 31564 19276 31604
rect 19316 31564 19317 31604
rect 19275 31555 19317 31564
rect 19468 31361 19508 31446
rect 19467 31352 19509 31361
rect 19852 31352 19892 31361
rect 19467 31312 19468 31352
rect 19508 31312 19509 31352
rect 19467 31303 19509 31312
rect 19564 31312 19852 31352
rect 19564 31184 19604 31312
rect 19852 31303 19892 31312
rect 20044 31352 20084 31361
rect 20044 31193 20084 31312
rect 19372 31144 19604 31184
rect 19660 31184 19700 31193
rect 19948 31184 19988 31193
rect 19700 31144 19892 31184
rect 18699 31016 18741 31025
rect 18699 30976 18700 31016
rect 18740 30976 18741 31016
rect 18699 30967 18741 30976
rect 19275 31016 19317 31025
rect 19275 30976 19276 31016
rect 19316 30976 19317 31016
rect 19275 30967 19317 30976
rect 18603 30680 18645 30689
rect 18603 30640 18604 30680
rect 18644 30640 18645 30680
rect 18603 30631 18645 30640
rect 18700 30680 18740 30967
rect 18795 30932 18837 30941
rect 18795 30892 18796 30932
rect 18836 30892 18837 30932
rect 18795 30883 18837 30892
rect 18796 30764 18836 30883
rect 18796 30715 18836 30724
rect 18700 30631 18740 30640
rect 19276 30680 19316 30967
rect 19276 30631 19316 30640
rect 18604 29840 18644 30631
rect 18699 30512 18741 30521
rect 18699 30472 18700 30512
rect 18740 30472 18741 30512
rect 18699 30463 18741 30472
rect 18604 29791 18644 29800
rect 18603 29504 18645 29513
rect 18603 29464 18604 29504
rect 18644 29464 18645 29504
rect 18603 29455 18645 29464
rect 18220 24583 18260 24592
rect 18316 24592 18548 24632
rect 18124 24424 18260 24464
rect 18028 24380 18068 24389
rect 18028 23885 18068 24340
rect 18027 23876 18069 23885
rect 18027 23836 18028 23876
rect 18068 23836 18069 23876
rect 18027 23827 18069 23836
rect 18124 23801 18164 23886
rect 18123 23792 18165 23801
rect 18123 23752 18124 23792
rect 18164 23752 18165 23792
rect 18123 23743 18165 23752
rect 18220 23624 18260 24424
rect 18124 23584 18260 23624
rect 18027 23540 18069 23549
rect 18027 23500 18028 23540
rect 18068 23500 18069 23540
rect 18027 23491 18069 23500
rect 18028 23120 18068 23491
rect 18028 23071 18068 23080
rect 18027 21440 18069 21449
rect 18027 21400 18028 21440
rect 18068 21400 18069 21440
rect 18027 21391 18069 21400
rect 18028 20768 18068 21391
rect 18124 21113 18164 23584
rect 18219 23288 18261 23297
rect 18219 23248 18220 23288
rect 18260 23248 18261 23288
rect 18219 23239 18261 23248
rect 18220 23154 18260 23239
rect 18123 21104 18165 21113
rect 18123 21064 18124 21104
rect 18164 21064 18165 21104
rect 18123 21055 18165 21064
rect 18028 20693 18068 20728
rect 18123 20768 18165 20777
rect 18123 20728 18124 20768
rect 18164 20728 18165 20768
rect 18316 20768 18356 24592
rect 18604 23381 18644 29455
rect 18700 27581 18740 30463
rect 19084 30437 19124 30522
rect 19275 30512 19317 30521
rect 19275 30472 19276 30512
rect 19316 30472 19317 30512
rect 19275 30463 19317 30472
rect 19083 30428 19125 30437
rect 19083 30388 19084 30428
rect 19124 30388 19125 30428
rect 19083 30379 19125 30388
rect 19276 30378 19316 30463
rect 18808 30260 19176 30269
rect 18848 30220 18890 30260
rect 18930 30220 18972 30260
rect 19012 30220 19054 30260
rect 19094 30220 19136 30260
rect 18808 30211 19176 30220
rect 19084 29845 19124 29854
rect 19084 29681 19124 29805
rect 19276 29756 19316 29765
rect 19372 29756 19412 31144
rect 19660 31135 19700 31144
rect 19756 30848 19796 30857
rect 19468 30808 19756 30848
rect 19852 30848 19892 31144
rect 19948 31025 19988 31144
rect 20043 31184 20085 31193
rect 20043 31144 20044 31184
rect 20084 31144 20085 31184
rect 20043 31135 20085 31144
rect 19947 31016 19989 31025
rect 19947 30976 19948 31016
rect 19988 30976 19989 31016
rect 19947 30967 19989 30976
rect 20048 31016 20416 31025
rect 20088 30976 20130 31016
rect 20170 30976 20212 31016
rect 20252 30976 20294 31016
rect 20334 30976 20376 31016
rect 20048 30967 20416 30976
rect 19852 30808 20084 30848
rect 19468 30680 19508 30808
rect 19756 30799 19796 30808
rect 19468 30631 19508 30640
rect 19564 30680 19604 30689
rect 19947 30680 19989 30689
rect 19604 30640 19796 30680
rect 19564 30631 19604 30640
rect 19659 30260 19701 30269
rect 19659 30220 19660 30260
rect 19700 30220 19701 30260
rect 19659 30211 19701 30220
rect 19467 30008 19509 30017
rect 19467 29968 19468 30008
rect 19508 29968 19509 30008
rect 19467 29959 19509 29968
rect 19316 29716 19412 29756
rect 19276 29707 19316 29716
rect 19083 29672 19125 29681
rect 19083 29632 19084 29672
rect 19124 29632 19125 29672
rect 19083 29623 19125 29632
rect 19468 29000 19508 29959
rect 19563 29840 19605 29849
rect 19563 29800 19564 29840
rect 19604 29800 19605 29840
rect 19563 29791 19605 29800
rect 19564 29706 19604 29791
rect 19563 29504 19605 29513
rect 19563 29464 19564 29504
rect 19604 29464 19605 29504
rect 19563 29455 19605 29464
rect 19564 29168 19604 29455
rect 19660 29261 19700 30211
rect 19756 29336 19796 30640
rect 19947 30640 19948 30680
rect 19988 30640 19989 30680
rect 19947 30631 19989 30640
rect 20044 30680 20084 30808
rect 19948 30546 19988 30631
rect 19851 30008 19893 30017
rect 19851 29968 19852 30008
rect 19892 29968 19893 30008
rect 19851 29959 19893 29968
rect 19852 29840 19892 29959
rect 19852 29791 19892 29800
rect 19947 29756 19989 29765
rect 19947 29716 19948 29756
rect 19988 29716 19989 29756
rect 19947 29707 19989 29716
rect 19948 29622 19988 29707
rect 20044 29681 20084 30640
rect 20235 30680 20277 30689
rect 20235 30640 20236 30680
rect 20276 30640 20277 30680
rect 20235 30631 20277 30640
rect 20236 30092 20276 30631
rect 20619 30512 20661 30521
rect 20619 30472 20620 30512
rect 20660 30472 20661 30512
rect 20619 30463 20661 30472
rect 20523 30428 20565 30437
rect 20523 30388 20524 30428
rect 20564 30388 20565 30428
rect 20523 30379 20565 30388
rect 20236 30043 20276 30052
rect 20043 29672 20085 29681
rect 20043 29632 20044 29672
rect 20084 29632 20085 29672
rect 20043 29623 20085 29632
rect 20048 29504 20416 29513
rect 20088 29464 20130 29504
rect 20170 29464 20212 29504
rect 20252 29464 20294 29504
rect 20334 29464 20376 29504
rect 20048 29455 20416 29464
rect 20044 29336 20084 29345
rect 19756 29296 20044 29336
rect 20044 29287 20084 29296
rect 20139 29336 20181 29345
rect 20139 29296 20140 29336
rect 20180 29296 20181 29336
rect 20139 29287 20181 29296
rect 19659 29252 19701 29261
rect 19659 29212 19660 29252
rect 19700 29212 19701 29252
rect 19659 29203 19701 29212
rect 19564 29119 19604 29128
rect 19276 28960 19508 29000
rect 19660 29000 19700 29203
rect 19947 29168 19989 29177
rect 19947 29128 19948 29168
rect 19988 29128 19989 29168
rect 19947 29119 19989 29128
rect 20140 29168 20180 29287
rect 20140 29119 20180 29128
rect 20236 29168 20276 29177
rect 20524 29168 20564 30379
rect 20276 29128 20564 29168
rect 20236 29119 20276 29128
rect 19948 29034 19988 29119
rect 19756 29000 19796 29009
rect 19660 28960 19756 29000
rect 18808 28748 19176 28757
rect 18848 28708 18890 28748
rect 18930 28708 18972 28748
rect 19012 28708 19054 28748
rect 19094 28708 19136 28748
rect 18808 28699 19176 28708
rect 18699 27572 18741 27581
rect 18699 27532 18700 27572
rect 18740 27532 18741 27572
rect 18699 27523 18741 27532
rect 19276 27488 19316 28960
rect 19756 28951 19796 28960
rect 20043 28496 20085 28505
rect 20043 28456 20044 28496
rect 20084 28456 20085 28496
rect 20043 28447 20085 28456
rect 19948 28337 19988 28422
rect 19468 28328 19508 28337
rect 19468 27917 19508 28288
rect 19852 28328 19892 28337
rect 19660 28160 19700 28169
rect 19467 27908 19509 27917
rect 19467 27868 19468 27908
rect 19508 27868 19509 27908
rect 19467 27859 19509 27868
rect 19468 27740 19508 27859
rect 19440 27700 19508 27740
rect 19440 27656 19480 27700
rect 19372 27635 19480 27656
rect 19412 27616 19480 27635
rect 19372 27586 19412 27595
rect 19660 27488 19700 28120
rect 19755 27992 19797 28001
rect 19755 27952 19756 27992
rect 19796 27952 19797 27992
rect 19755 27943 19797 27952
rect 19756 27657 19796 27943
rect 19852 27833 19892 28288
rect 19947 28328 19989 28337
rect 19947 28288 19948 28328
rect 19988 28288 19989 28328
rect 19947 28279 19989 28288
rect 20044 28328 20084 28447
rect 20044 28279 20084 28288
rect 20140 28160 20180 28169
rect 19948 28120 20140 28160
rect 19851 27824 19893 27833
rect 19851 27784 19852 27824
rect 19892 27784 19893 27824
rect 19851 27775 19893 27784
rect 19756 27608 19796 27617
rect 19852 27656 19892 27665
rect 19276 27448 19412 27488
rect 19660 27448 19796 27488
rect 18808 27236 19176 27245
rect 18848 27196 18890 27236
rect 18930 27196 18972 27236
rect 19012 27196 19054 27236
rect 19094 27196 19136 27236
rect 18808 27187 19176 27196
rect 19275 27236 19317 27245
rect 19275 27196 19276 27236
rect 19316 27196 19317 27236
rect 19275 27187 19317 27196
rect 18940 26825 18980 26834
rect 19276 26825 19316 27187
rect 19372 26825 19412 27448
rect 19564 27404 19604 27413
rect 19604 27364 19700 27404
rect 19564 27355 19604 27364
rect 19467 27320 19509 27329
rect 19467 27280 19468 27320
rect 19508 27280 19509 27320
rect 19467 27271 19509 27280
rect 18699 26816 18741 26825
rect 18699 26776 18700 26816
rect 18740 26776 18741 26816
rect 18980 26816 19316 26825
rect 18980 26785 19276 26816
rect 18940 26776 18980 26785
rect 18699 26767 18741 26776
rect 19276 26767 19316 26776
rect 19371 26816 19413 26825
rect 19371 26776 19372 26816
rect 19412 26776 19413 26816
rect 19371 26767 19413 26776
rect 19468 26816 19508 27271
rect 19660 27245 19700 27364
rect 19659 27236 19701 27245
rect 19659 27196 19660 27236
rect 19700 27196 19701 27236
rect 19659 27187 19701 27196
rect 19756 27068 19796 27448
rect 19852 27245 19892 27616
rect 19948 27497 19988 28120
rect 20140 28111 20180 28120
rect 20048 27992 20416 28001
rect 20088 27952 20130 27992
rect 20170 27952 20212 27992
rect 20252 27952 20294 27992
rect 20334 27952 20376 27992
rect 20048 27943 20416 27952
rect 20044 27824 20084 27833
rect 19947 27488 19989 27497
rect 19947 27448 19948 27488
rect 19988 27448 19989 27488
rect 19947 27439 19989 27448
rect 20044 27413 20084 27784
rect 20139 27740 20181 27749
rect 20139 27700 20140 27740
rect 20180 27700 20181 27740
rect 20139 27691 20181 27700
rect 20043 27404 20085 27413
rect 20043 27364 20044 27404
rect 20084 27364 20085 27404
rect 20043 27355 20085 27364
rect 19851 27236 19893 27245
rect 20140 27236 20180 27691
rect 19851 27196 19852 27236
rect 19892 27196 19893 27236
rect 19851 27187 19893 27196
rect 20044 27196 20180 27236
rect 19468 26767 19508 26776
rect 19660 27028 19892 27068
rect 18700 24044 18740 26767
rect 19084 26648 19124 26657
rect 19563 26648 19605 26657
rect 19124 26608 19508 26648
rect 19084 26599 19124 26608
rect 19083 26480 19125 26489
rect 19083 26440 19084 26480
rect 19124 26440 19125 26480
rect 19083 26431 19125 26440
rect 19275 26480 19317 26489
rect 19275 26440 19276 26480
rect 19316 26440 19317 26480
rect 19275 26431 19317 26440
rect 19084 26144 19124 26431
rect 19276 26312 19316 26431
rect 19276 26263 19316 26272
rect 19468 26144 19508 26608
rect 19563 26608 19564 26648
rect 19604 26608 19605 26648
rect 19563 26599 19605 26608
rect 19564 26514 19604 26599
rect 19124 26104 19316 26144
rect 19084 26095 19124 26104
rect 18808 25724 19176 25733
rect 18848 25684 18890 25724
rect 18930 25684 18972 25724
rect 19012 25684 19054 25724
rect 19094 25684 19136 25724
rect 18808 25675 19176 25684
rect 18808 24212 19176 24221
rect 18848 24172 18890 24212
rect 18930 24172 18972 24212
rect 19012 24172 19054 24212
rect 19094 24172 19136 24212
rect 18808 24163 19176 24172
rect 19276 24044 19316 26104
rect 19468 26095 19508 26104
rect 19564 26144 19604 26153
rect 19660 26144 19700 27028
rect 19755 26816 19797 26825
rect 19755 26776 19756 26816
rect 19796 26776 19797 26816
rect 19755 26767 19797 26776
rect 19852 26816 19892 27028
rect 19852 26767 19892 26776
rect 19756 26682 19796 26767
rect 19947 26732 19989 26741
rect 19947 26692 19948 26732
rect 19988 26692 19989 26732
rect 19947 26683 19989 26692
rect 19604 26104 19700 26144
rect 19564 26095 19604 26104
rect 18700 24004 18836 24044
rect 18603 23372 18645 23381
rect 18603 23332 18604 23372
rect 18644 23332 18645 23372
rect 18603 23323 18645 23332
rect 18411 23288 18453 23297
rect 18411 23248 18412 23288
rect 18452 23248 18453 23288
rect 18411 23239 18453 23248
rect 18412 23120 18452 23239
rect 18412 23071 18452 23080
rect 18508 23120 18548 23129
rect 18508 21785 18548 23080
rect 18604 23120 18644 23129
rect 18604 22121 18644 23080
rect 18699 23120 18741 23129
rect 18699 23080 18700 23120
rect 18740 23080 18741 23120
rect 18699 23071 18741 23080
rect 18700 22986 18740 23071
rect 18796 22868 18836 24004
rect 18700 22828 18836 22868
rect 19084 24004 19316 24044
rect 19468 24632 19508 24641
rect 19084 22868 19124 24004
rect 19371 23960 19413 23969
rect 19371 23920 19372 23960
rect 19412 23920 19413 23960
rect 19371 23911 19413 23920
rect 19179 23876 19221 23885
rect 19179 23836 19180 23876
rect 19220 23836 19221 23876
rect 19179 23827 19221 23836
rect 19180 23120 19220 23827
rect 19372 23792 19412 23911
rect 19372 23743 19412 23752
rect 19275 23624 19317 23633
rect 19275 23584 19276 23624
rect 19316 23584 19317 23624
rect 19275 23575 19317 23584
rect 19180 23071 19220 23080
rect 19276 23120 19316 23575
rect 19468 23456 19508 24592
rect 19756 23792 19796 23801
rect 19563 23624 19605 23633
rect 19756 23624 19796 23752
rect 19852 23792 19892 23803
rect 19852 23717 19892 23752
rect 19851 23708 19893 23717
rect 19851 23668 19852 23708
rect 19892 23668 19893 23708
rect 19851 23659 19893 23668
rect 19563 23584 19564 23624
rect 19604 23584 19796 23624
rect 19563 23575 19605 23584
rect 19564 23490 19604 23575
rect 19851 23540 19893 23549
rect 19851 23500 19852 23540
rect 19892 23500 19893 23540
rect 19851 23491 19893 23500
rect 19276 23071 19316 23080
rect 19372 23416 19508 23456
rect 19084 22828 19316 22868
rect 18603 22112 18645 22121
rect 18603 22072 18604 22112
rect 18644 22072 18645 22112
rect 18603 22063 18645 22072
rect 18507 21776 18549 21785
rect 18507 21736 18508 21776
rect 18548 21736 18549 21776
rect 18507 21727 18549 21736
rect 18700 21020 18740 22828
rect 18808 22700 19176 22709
rect 18848 22660 18890 22700
rect 18930 22660 18972 22700
rect 19012 22660 19054 22700
rect 19094 22660 19136 22700
rect 18808 22651 19176 22660
rect 19276 21701 19316 22828
rect 19275 21692 19317 21701
rect 19275 21652 19276 21692
rect 19316 21652 19317 21692
rect 19275 21643 19317 21652
rect 18987 21608 19029 21617
rect 18987 21568 18988 21608
rect 19028 21568 19029 21608
rect 18987 21559 19029 21568
rect 18988 21474 19028 21559
rect 18808 21188 19176 21197
rect 18848 21148 18890 21188
rect 18930 21148 18972 21188
rect 19012 21148 19054 21188
rect 19094 21148 19136 21188
rect 18808 21139 19176 21148
rect 18700 20980 18836 21020
rect 18507 20852 18549 20861
rect 18507 20812 18508 20852
rect 18548 20812 18549 20852
rect 18507 20803 18549 20812
rect 18508 20768 18548 20803
rect 18316 20728 18452 20768
rect 18123 20719 18165 20728
rect 18027 20684 18069 20693
rect 18027 20644 18028 20684
rect 18068 20644 18069 20684
rect 18027 20635 18069 20644
rect 18124 20634 18164 20719
rect 18316 20600 18356 20609
rect 18412 20600 18452 20728
rect 18508 20717 18548 20728
rect 18700 20768 18740 20777
rect 18700 20609 18740 20728
rect 18604 20600 18644 20609
rect 18412 20560 18548 20600
rect 18123 20516 18165 20525
rect 17932 20476 18068 20516
rect 17836 20392 17972 20432
rect 17644 20308 17876 20348
rect 17355 20299 17397 20308
rect 17260 20096 17300 20105
rect 17356 20096 17396 20299
rect 17739 20096 17781 20105
rect 17356 20091 17475 20096
rect 17356 20082 17492 20091
rect 17356 20056 17452 20082
rect 17260 20012 17300 20056
rect 17435 20046 17452 20056
rect 17545 20077 17684 20096
rect 17545 20042 17552 20077
rect 17452 20033 17492 20042
rect 17592 20056 17684 20077
rect 17552 20028 17592 20037
rect 17260 19972 17396 20012
rect 17356 19853 17396 19972
rect 17108 18544 17204 18584
rect 17068 18535 17108 18544
rect 17068 17996 17108 18005
rect 16972 17956 17068 17996
rect 17068 17947 17108 17956
rect 16491 17576 16533 17585
rect 16491 17536 16492 17576
rect 16532 17536 16533 17576
rect 16491 17527 16533 17536
rect 16492 17072 16532 17527
rect 16684 17417 16724 17620
rect 16876 17585 16916 17704
rect 17164 17660 17204 18544
rect 17068 17620 17204 17660
rect 17260 19844 17300 19853
rect 16875 17576 16917 17585
rect 16875 17536 16876 17576
rect 16916 17536 16917 17576
rect 16875 17527 16917 17536
rect 16683 17408 16725 17417
rect 16683 17368 16684 17408
rect 16724 17368 16725 17408
rect 16683 17359 16725 17368
rect 16492 17023 16532 17032
rect 16684 17116 17012 17156
rect 16684 16904 16724 17116
rect 16972 17072 17012 17116
rect 17068 17081 17108 17620
rect 16972 17023 17012 17032
rect 17067 17072 17109 17081
rect 17067 17032 17068 17072
rect 17108 17032 17109 17072
rect 17067 17023 17109 17032
rect 16779 16988 16821 16997
rect 16779 16948 16780 16988
rect 16820 16948 16821 16988
rect 16779 16939 16821 16948
rect 16684 16855 16724 16864
rect 16396 16444 16532 16484
rect 16299 16435 16341 16444
rect 16203 16400 16245 16409
rect 16203 16360 16204 16400
rect 16244 16360 16245 16400
rect 16203 16351 16245 16360
rect 16204 16232 16244 16351
rect 16395 16316 16437 16325
rect 16395 16276 16396 16316
rect 16436 16276 16437 16316
rect 16395 16267 16437 16276
rect 16204 16183 16244 16192
rect 16396 16148 16436 16267
rect 16396 16099 16436 16108
rect 16492 15980 16532 16444
rect 16683 16316 16725 16325
rect 16683 16276 16684 16316
rect 16724 16276 16725 16316
rect 16683 16267 16725 16276
rect 16684 16232 16724 16267
rect 16684 16181 16724 16192
rect 16780 16232 16820 16939
rect 16875 16904 16917 16913
rect 16875 16864 16876 16904
rect 16916 16864 16917 16904
rect 16875 16855 16917 16864
rect 16396 15940 16532 15980
rect 16108 14512 16340 14552
rect 16107 14132 16149 14141
rect 16107 14092 16108 14132
rect 16148 14092 16149 14132
rect 16107 14083 16149 14092
rect 16108 14048 16148 14083
rect 16108 13997 16148 14008
rect 16204 13964 16244 13973
rect 16011 13880 16053 13889
rect 16011 13840 16012 13880
rect 16052 13840 16053 13880
rect 16011 13831 16053 13840
rect 16204 13721 16244 13924
rect 15915 13712 15957 13721
rect 15915 13672 15916 13712
rect 15956 13672 15957 13712
rect 15915 13663 15957 13672
rect 16203 13712 16245 13721
rect 16203 13672 16204 13712
rect 16244 13672 16245 13712
rect 16203 13663 16245 13672
rect 15915 13292 15957 13301
rect 15915 13252 15916 13292
rect 15956 13252 15957 13292
rect 15915 13243 15957 13252
rect 15916 13208 15956 13243
rect 15916 13157 15956 13168
rect 16300 12545 16340 14512
rect 16396 13301 16436 15940
rect 16588 15569 16628 15654
rect 16587 15560 16629 15569
rect 16587 15520 16588 15560
rect 16628 15520 16629 15560
rect 16587 15511 16629 15520
rect 16587 15308 16629 15317
rect 16587 15268 16588 15308
rect 16628 15268 16629 15308
rect 16587 15259 16629 15268
rect 16491 14888 16533 14897
rect 16491 14848 16492 14888
rect 16532 14848 16533 14888
rect 16491 14839 16533 14848
rect 16492 14561 16532 14839
rect 16491 14552 16533 14561
rect 16491 14512 16492 14552
rect 16532 14512 16533 14552
rect 16491 14503 16533 14512
rect 16395 13292 16437 13301
rect 16395 13252 16396 13292
rect 16436 13252 16437 13292
rect 16395 13243 16437 13252
rect 15915 12536 15957 12545
rect 15915 12496 15916 12536
rect 15956 12496 15957 12536
rect 15915 12487 15957 12496
rect 16012 12536 16052 12545
rect 16299 12536 16341 12545
rect 16052 12496 16300 12536
rect 16340 12496 16341 12536
rect 16012 12487 16052 12496
rect 15916 12368 15956 12487
rect 15916 12328 16148 12368
rect 16108 11957 16148 12328
rect 16107 11948 16149 11957
rect 16107 11908 16108 11948
rect 16148 11908 16149 11948
rect 16107 11899 16149 11908
rect 15916 11696 15956 11705
rect 15916 11201 15956 11656
rect 16012 11696 16052 11705
rect 15915 11192 15957 11201
rect 15915 11152 15916 11192
rect 15956 11152 15957 11192
rect 15915 11143 15957 11152
rect 16012 10445 16052 11656
rect 16011 10436 16053 10445
rect 15820 10396 15956 10436
rect 15723 10387 15765 10396
rect 15724 10268 15764 10387
rect 15820 10268 15860 10277
rect 15724 10228 15820 10268
rect 15627 8924 15669 8933
rect 15627 8884 15628 8924
rect 15668 8884 15669 8924
rect 15627 8875 15669 8884
rect 15628 8840 15668 8875
rect 15628 8789 15668 8800
rect 15436 7169 15476 8632
rect 15531 8672 15573 8681
rect 15531 8632 15532 8672
rect 15572 8632 15573 8672
rect 15531 8623 15573 8632
rect 15724 8084 15764 10228
rect 15820 10219 15860 10228
rect 15916 10184 15956 10396
rect 16011 10396 16012 10436
rect 16052 10396 16053 10436
rect 16011 10387 16053 10396
rect 15820 9512 15860 9521
rect 15820 9101 15860 9472
rect 15819 9092 15861 9101
rect 15819 9052 15820 9092
rect 15860 9052 15861 9092
rect 15819 9043 15861 9052
rect 15532 8044 15764 8084
rect 15532 7916 15572 8044
rect 15435 7160 15477 7169
rect 15435 7120 15436 7160
rect 15476 7120 15477 7160
rect 15435 7111 15477 7120
rect 15435 6992 15477 7001
rect 15435 6952 15436 6992
rect 15476 6952 15477 6992
rect 15435 6943 15477 6952
rect 15436 6488 15476 6943
rect 15436 6439 15476 6448
rect 15532 5648 15572 7876
rect 15628 7916 15668 7925
rect 15916 7916 15956 10144
rect 16011 9512 16053 9521
rect 16108 9512 16148 11899
rect 16011 9472 16012 9512
rect 16052 9472 16148 9512
rect 16011 9463 16053 9472
rect 15668 7876 15956 7916
rect 15628 7867 15668 7876
rect 15628 5648 15668 5657
rect 15244 5405 15284 5608
rect 15436 5608 15628 5648
rect 15243 5396 15285 5405
rect 15243 5356 15244 5396
rect 15284 5356 15285 5396
rect 15243 5347 15285 5356
rect 15244 5144 15284 5153
rect 15148 5104 15244 5144
rect 15244 5095 15284 5104
rect 15436 4976 15476 5608
rect 15628 5599 15668 5608
rect 15724 5648 15764 7876
rect 15764 5608 15860 5648
rect 15724 5599 15764 5608
rect 15723 5480 15765 5489
rect 15723 5440 15724 5480
rect 15764 5440 15765 5480
rect 15723 5431 15765 5440
rect 15531 5060 15573 5069
rect 15531 5020 15532 5060
rect 15572 5020 15573 5060
rect 15531 5011 15573 5020
rect 14955 4220 14997 4229
rect 14955 4180 14956 4220
rect 14996 4180 14997 4220
rect 14955 4171 14997 4180
rect 14188 4085 14228 4096
rect 14668 4136 14708 4145
rect 14380 4052 14420 4061
rect 14668 4052 14708 4096
rect 14763 4136 14805 4145
rect 14763 4096 14764 4136
rect 14804 4096 14805 4136
rect 14763 4087 14805 4096
rect 14420 4012 14708 4052
rect 14380 4003 14420 4012
rect 14764 4002 14804 4087
rect 14572 3548 14612 3557
rect 14380 3450 14420 3459
rect 14187 3380 14229 3389
rect 14187 3340 14188 3380
rect 14228 3340 14229 3380
rect 14187 3331 14229 3340
rect 13995 2960 14037 2969
rect 13995 2920 13996 2960
rect 14036 2920 14037 2960
rect 13995 2911 14037 2920
rect 14188 2633 14228 3331
rect 14380 2876 14420 3410
rect 14572 3305 14612 3508
rect 14571 3296 14613 3305
rect 14571 3256 14572 3296
rect 14612 3256 14613 3296
rect 14571 3247 14613 3256
rect 14859 3212 14901 3221
rect 14859 3172 14860 3212
rect 14900 3172 14901 3212
rect 14859 3163 14901 3172
rect 14380 2827 14420 2836
rect 14187 2624 14229 2633
rect 14187 2584 14188 2624
rect 14228 2584 14229 2624
rect 14187 2575 14229 2584
rect 14860 2624 14900 3163
rect 15052 2801 15092 4936
rect 15148 4936 15476 4976
rect 15532 4976 15572 5011
rect 15148 4136 15188 4936
rect 15532 4925 15572 4936
rect 15051 2792 15093 2801
rect 15051 2752 15052 2792
rect 15092 2752 15093 2792
rect 15051 2743 15093 2752
rect 15148 2637 15188 4096
rect 15243 4136 15285 4145
rect 15243 4096 15244 4136
rect 15284 4096 15285 4136
rect 15243 4087 15285 4096
rect 15724 4136 15764 5431
rect 15820 4145 15860 5608
rect 15915 5060 15957 5069
rect 15915 5020 15916 5060
rect 15956 5020 15957 5060
rect 15915 5011 15957 5020
rect 15724 4087 15764 4096
rect 15819 4136 15861 4145
rect 15819 4096 15820 4136
rect 15860 4096 15861 4136
rect 15819 4087 15861 4096
rect 15244 3473 15284 4087
rect 15243 3464 15285 3473
rect 15243 3424 15244 3464
rect 15284 3424 15285 3464
rect 15243 3415 15285 3424
rect 15436 3464 15476 3473
rect 15436 2969 15476 3424
rect 15435 2960 15477 2969
rect 15435 2920 15436 2960
rect 15476 2920 15477 2960
rect 15435 2911 15477 2920
rect 15531 2792 15573 2801
rect 15531 2752 15532 2792
rect 15572 2752 15573 2792
rect 15531 2743 15573 2752
rect 14860 2575 14900 2584
rect 14956 2597 15188 2637
rect 14667 2456 14709 2465
rect 14667 2416 14668 2456
rect 14708 2416 14709 2456
rect 14667 2407 14709 2416
rect 13707 2372 13749 2381
rect 13707 2332 13708 2372
rect 13748 2332 13749 2372
rect 13707 2323 13749 2332
rect 14284 1877 14324 1962
rect 13228 1819 13268 1828
rect 13899 1868 13941 1877
rect 13899 1828 13900 1868
rect 13940 1828 13941 1868
rect 13899 1819 13941 1828
rect 14283 1868 14325 1877
rect 14283 1828 14284 1868
rect 14324 1828 14325 1868
rect 14283 1819 14325 1828
rect 14668 1868 14708 2407
rect 14668 1819 14708 1828
rect 13900 1734 13940 1819
rect 13420 1700 13460 1709
rect 13323 1616 13365 1625
rect 13323 1576 13324 1616
rect 13364 1576 13365 1616
rect 13323 1567 13365 1576
rect 13324 80 13364 1567
rect 13420 785 13460 1660
rect 14092 1700 14132 1709
rect 14476 1700 14516 1709
rect 14860 1700 14900 1709
rect 14132 1660 14420 1700
rect 14092 1651 14132 1660
rect 14283 1448 14325 1457
rect 14283 1408 14284 1448
rect 14324 1408 14325 1448
rect 14283 1399 14325 1408
rect 13899 1280 13941 1289
rect 13899 1240 13900 1280
rect 13940 1240 13941 1280
rect 13899 1231 13941 1240
rect 13707 860 13749 869
rect 13707 820 13708 860
rect 13748 820 13749 860
rect 13707 811 13749 820
rect 13419 776 13461 785
rect 13419 736 13420 776
rect 13460 736 13461 776
rect 13419 727 13461 736
rect 13515 692 13557 701
rect 13515 652 13516 692
rect 13556 652 13557 692
rect 13515 643 13557 652
rect 13516 80 13556 643
rect 13708 80 13748 811
rect 13900 80 13940 1231
rect 14091 776 14133 785
rect 14091 736 14092 776
rect 14132 736 14133 776
rect 14091 727 14133 736
rect 14092 80 14132 727
rect 14284 80 14324 1399
rect 14380 1112 14420 1660
rect 14516 1660 14804 1700
rect 14476 1651 14516 1660
rect 14380 1072 14708 1112
rect 14475 944 14517 953
rect 14475 904 14476 944
rect 14516 904 14517 944
rect 14475 895 14517 904
rect 14476 80 14516 895
rect 14668 80 14708 1072
rect 14764 860 14804 1660
rect 14860 1037 14900 1660
rect 14956 1121 14996 2597
rect 15243 1868 15285 1877
rect 15243 1828 15244 1868
rect 15284 1828 15285 1868
rect 15243 1819 15285 1828
rect 15244 1734 15284 1819
rect 15052 1700 15092 1709
rect 14955 1112 14997 1121
rect 14955 1072 14956 1112
rect 14996 1072 14997 1112
rect 14955 1063 14997 1072
rect 14859 1028 14901 1037
rect 14859 988 14860 1028
rect 14900 988 14901 1028
rect 14859 979 14901 988
rect 14955 944 14997 953
rect 14955 904 14956 944
rect 14996 904 14997 944
rect 14955 895 14997 904
rect 14764 820 14900 860
rect 14860 80 14900 820
rect 14956 810 14996 895
rect 15052 692 15092 1660
rect 15436 1700 15476 1709
rect 15436 1457 15476 1660
rect 15435 1448 15477 1457
rect 15435 1408 15436 1448
rect 15476 1408 15477 1448
rect 15435 1399 15477 1408
rect 15147 1196 15189 1205
rect 15147 1156 15148 1196
rect 15188 1156 15189 1196
rect 15147 1147 15189 1156
rect 15148 1062 15188 1147
rect 15435 1028 15477 1037
rect 15435 988 15436 1028
rect 15476 988 15477 1028
rect 15435 979 15477 988
rect 15243 860 15285 869
rect 15243 820 15244 860
rect 15284 820 15285 860
rect 15243 811 15285 820
rect 14956 652 15092 692
rect 14956 365 14996 652
rect 15051 524 15093 533
rect 15051 484 15052 524
rect 15092 484 15093 524
rect 15051 475 15093 484
rect 14955 356 14997 365
rect 14955 316 14956 356
rect 14996 316 14997 356
rect 14955 307 14997 316
rect 15052 80 15092 475
rect 15244 80 15284 811
rect 15436 80 15476 979
rect 15532 365 15572 2743
rect 15627 1868 15669 1877
rect 15627 1828 15628 1868
rect 15668 1828 15669 1868
rect 15627 1819 15669 1828
rect 15628 1734 15668 1819
rect 15820 1700 15860 1709
rect 15724 1660 15820 1700
rect 15627 1280 15669 1289
rect 15627 1240 15628 1280
rect 15668 1240 15669 1280
rect 15627 1231 15669 1240
rect 15531 356 15573 365
rect 15531 316 15532 356
rect 15572 316 15573 356
rect 15531 307 15573 316
rect 15628 80 15668 1231
rect 15724 785 15764 1660
rect 15820 1651 15860 1660
rect 15916 1196 15956 5011
rect 16012 2036 16052 9463
rect 16107 8000 16149 8009
rect 16107 7960 16108 8000
rect 16148 7960 16149 8000
rect 16107 7951 16149 7960
rect 16108 7866 16148 7951
rect 16204 7328 16244 12496
rect 16299 12487 16341 12496
rect 16300 12402 16340 12487
rect 16395 11780 16437 11789
rect 16395 11740 16396 11780
rect 16436 11740 16437 11780
rect 16395 11731 16437 11740
rect 16492 11780 16532 14503
rect 16492 11731 16532 11740
rect 16299 11024 16341 11033
rect 16299 10984 16300 11024
rect 16340 10984 16341 11024
rect 16299 10975 16341 10984
rect 16300 10890 16340 10975
rect 16396 10184 16436 11731
rect 16491 11192 16533 11201
rect 16491 11152 16492 11192
rect 16532 11152 16533 11192
rect 16491 11143 16533 11152
rect 16492 11058 16532 11143
rect 16299 8672 16341 8681
rect 16299 8632 16300 8672
rect 16340 8632 16341 8672
rect 16299 8623 16341 8632
rect 16108 7288 16244 7328
rect 16108 4985 16148 7288
rect 16204 7160 16244 7169
rect 16204 6749 16244 7120
rect 16203 6740 16245 6749
rect 16203 6700 16204 6740
rect 16244 6700 16245 6740
rect 16203 6691 16245 6700
rect 16300 5909 16340 8623
rect 16396 8009 16436 10144
rect 16588 8084 16628 15259
rect 16780 14729 16820 16192
rect 16779 14720 16821 14729
rect 16779 14680 16780 14720
rect 16820 14680 16821 14720
rect 16779 14671 16821 14680
rect 16683 14216 16725 14225
rect 16683 14176 16684 14216
rect 16724 14176 16725 14216
rect 16683 14167 16725 14176
rect 16684 14048 16724 14167
rect 16684 13999 16724 14008
rect 16780 13880 16820 14671
rect 16684 13840 16820 13880
rect 16684 8261 16724 13840
rect 16876 10352 16916 16855
rect 17260 16484 17300 19804
rect 17355 19844 17397 19853
rect 17355 19804 17356 19844
rect 17396 19804 17397 19844
rect 17644 19844 17684 20056
rect 17739 20056 17740 20096
rect 17780 20056 17781 20096
rect 17739 20047 17781 20056
rect 17740 19962 17780 20047
rect 17836 20021 17876 20308
rect 17932 20096 17972 20392
rect 18028 20273 18068 20476
rect 18123 20476 18124 20516
rect 18164 20476 18165 20516
rect 18123 20467 18165 20476
rect 18027 20264 18069 20273
rect 18027 20224 18028 20264
rect 18068 20224 18069 20264
rect 18027 20215 18069 20224
rect 18124 20180 18164 20467
rect 18316 20357 18356 20560
rect 18411 20432 18453 20441
rect 18411 20392 18412 20432
rect 18452 20392 18453 20432
rect 18411 20383 18453 20392
rect 18315 20348 18357 20357
rect 18315 20308 18316 20348
rect 18356 20308 18357 20348
rect 18315 20299 18357 20308
rect 18121 20140 18164 20180
rect 18315 20180 18357 20189
rect 18315 20140 18316 20180
rect 18356 20140 18357 20180
rect 18121 20138 18161 20140
rect 17932 20047 17972 20056
rect 18028 20098 18161 20138
rect 18315 20131 18357 20140
rect 18028 20096 18068 20098
rect 18028 20047 18068 20056
rect 17835 20012 17877 20021
rect 17835 19972 17836 20012
rect 17876 19972 17877 20012
rect 17835 19963 17877 19972
rect 17740 19844 17780 19853
rect 17644 19804 17740 19844
rect 17355 19795 17397 19804
rect 17740 19795 17780 19804
rect 17451 19256 17493 19265
rect 17451 19216 17452 19256
rect 17492 19216 17493 19256
rect 17451 19207 17493 19216
rect 17452 19122 17492 19207
rect 17355 19088 17397 19097
rect 17355 19048 17356 19088
rect 17396 19048 17397 19088
rect 17355 19039 17397 19048
rect 17164 16444 17300 16484
rect 17164 16400 17204 16444
rect 17068 16360 17204 16400
rect 17068 15317 17108 16360
rect 17164 16232 17204 16241
rect 17164 15560 17204 16192
rect 17260 16232 17300 16243
rect 17260 16157 17300 16192
rect 17259 16148 17301 16157
rect 17259 16108 17260 16148
rect 17300 16108 17301 16148
rect 17259 16099 17301 16108
rect 17164 15520 17300 15560
rect 17067 15308 17109 15317
rect 17067 15268 17068 15308
rect 17108 15268 17109 15308
rect 17067 15259 17109 15268
rect 17260 14813 17300 15520
rect 17259 14804 17301 14813
rect 17259 14764 17260 14804
rect 17300 14764 17301 14804
rect 17259 14755 17301 14764
rect 17068 14720 17108 14729
rect 17068 13469 17108 14680
rect 17163 14720 17205 14729
rect 17163 14680 17164 14720
rect 17204 14680 17205 14720
rect 17163 14671 17205 14680
rect 17164 14586 17204 14671
rect 17356 14552 17396 19039
rect 17547 18668 17589 18677
rect 17547 18628 17548 18668
rect 17588 18628 17589 18668
rect 17547 18619 17589 18628
rect 17548 18584 17588 18619
rect 17452 18500 17492 18509
rect 17452 16988 17492 18460
rect 17452 14804 17492 16948
rect 17548 16988 17588 18544
rect 17643 17744 17685 17753
rect 17643 17704 17644 17744
rect 17684 17704 17685 17744
rect 17643 17695 17685 17704
rect 17644 17610 17684 17695
rect 17548 16157 17588 16948
rect 17836 16913 17876 19963
rect 18028 18584 18068 18593
rect 18028 17072 18068 18544
rect 17835 16904 17877 16913
rect 17835 16864 17836 16904
rect 17876 16864 17877 16904
rect 17835 16855 17877 16864
rect 17835 16400 17877 16409
rect 17835 16360 17836 16400
rect 17876 16360 17877 16400
rect 17835 16351 17877 16360
rect 17739 16232 17781 16241
rect 17739 16192 17740 16232
rect 17780 16192 17781 16232
rect 17739 16183 17781 16192
rect 17547 16148 17589 16157
rect 17547 16108 17548 16148
rect 17588 16108 17589 16148
rect 17547 16099 17589 16108
rect 17548 15140 17588 16099
rect 17740 16098 17780 16183
rect 17836 15560 17876 16351
rect 18028 16241 18068 17032
rect 18027 16232 18069 16241
rect 17932 16192 18028 16232
rect 18068 16192 18069 16232
rect 17932 15560 17972 16192
rect 18027 16183 18069 16192
rect 18220 16237 18260 16246
rect 18028 15728 18068 15737
rect 18220 15728 18260 16197
rect 18068 15688 18260 15728
rect 18028 15679 18068 15688
rect 17932 15520 18164 15560
rect 17836 15511 17876 15520
rect 17548 15100 17684 15140
rect 17547 14804 17589 14813
rect 17452 14764 17548 14804
rect 17588 14764 17589 14804
rect 17547 14755 17589 14764
rect 17548 14670 17588 14755
rect 17644 14729 17684 15100
rect 17643 14720 17685 14729
rect 17643 14680 17644 14720
rect 17684 14680 17685 14720
rect 17643 14671 17685 14680
rect 18124 14720 18164 15520
rect 18124 14671 18164 14680
rect 18219 14720 18261 14729
rect 18219 14680 18220 14720
rect 18260 14680 18261 14720
rect 18219 14671 18261 14680
rect 17644 14586 17684 14671
rect 17356 14512 17588 14552
rect 17355 14300 17397 14309
rect 17355 14260 17356 14300
rect 17396 14260 17397 14300
rect 17355 14251 17397 14260
rect 17356 14216 17396 14251
rect 17356 14165 17396 14176
rect 17212 14038 17252 14047
rect 17252 13998 17492 14034
rect 17212 13994 17492 13998
rect 17212 13989 17252 13994
rect 17163 13880 17205 13889
rect 17163 13840 17164 13880
rect 17204 13840 17205 13880
rect 17163 13831 17205 13840
rect 17067 13460 17109 13469
rect 17067 13420 17068 13460
rect 17108 13420 17109 13460
rect 17067 13411 17109 13420
rect 17067 13292 17109 13301
rect 17067 13252 17068 13292
rect 17108 13252 17109 13292
rect 17067 13243 17109 13252
rect 16972 11696 17012 11705
rect 16972 11537 17012 11656
rect 16971 11528 17013 11537
rect 16971 11488 16972 11528
rect 17012 11488 17013 11528
rect 16971 11479 17013 11488
rect 17068 10361 17108 13243
rect 17164 13208 17204 13831
rect 17355 13460 17397 13469
rect 17355 13420 17356 13460
rect 17396 13420 17397 13460
rect 17355 13411 17397 13420
rect 17356 13326 17396 13411
rect 16780 10312 16916 10352
rect 17067 10352 17109 10361
rect 17067 10312 17068 10352
rect 17108 10312 17109 10352
rect 16780 10100 16820 10312
rect 17067 10303 17109 10312
rect 16924 10193 16964 10202
rect 16964 10153 17012 10184
rect 16924 10144 17012 10153
rect 16780 10060 16916 10100
rect 16683 8252 16725 8261
rect 16683 8212 16684 8252
rect 16724 8212 16725 8252
rect 16683 8203 16725 8212
rect 16779 8168 16821 8177
rect 16779 8128 16780 8168
rect 16820 8128 16821 8168
rect 16779 8119 16821 8128
rect 16492 8044 16628 8084
rect 16395 8000 16437 8009
rect 16395 7960 16396 8000
rect 16436 7960 16437 8000
rect 16395 7951 16437 7960
rect 16395 7832 16437 7841
rect 16395 7792 16396 7832
rect 16436 7792 16437 7832
rect 16395 7783 16437 7792
rect 16299 5900 16341 5909
rect 16299 5860 16300 5900
rect 16340 5860 16341 5900
rect 16299 5851 16341 5860
rect 16204 5648 16244 5657
rect 16204 5489 16244 5608
rect 16203 5480 16245 5489
rect 16203 5440 16204 5480
rect 16244 5440 16245 5480
rect 16203 5431 16245 5440
rect 16107 4976 16149 4985
rect 16107 4936 16108 4976
rect 16148 4936 16149 4976
rect 16107 4927 16149 4936
rect 16107 4220 16149 4229
rect 16107 4180 16108 4220
rect 16148 4180 16149 4220
rect 16107 4171 16149 4180
rect 16108 2624 16148 4171
rect 16252 4145 16292 4154
rect 16292 4105 16340 4136
rect 16252 4096 16340 4105
rect 16300 2876 16340 4096
rect 16396 4052 16436 7783
rect 16492 5069 16532 8044
rect 16780 8034 16820 8119
rect 16876 8000 16916 10060
rect 16972 9773 17012 10144
rect 17068 10058 17108 10303
rect 17068 10009 17108 10018
rect 16971 9764 17013 9773
rect 16971 9724 16972 9764
rect 17012 9724 17013 9764
rect 16971 9715 17013 9724
rect 17068 9512 17108 9521
rect 17164 9512 17204 13168
rect 17259 12620 17301 12629
rect 17259 12580 17260 12620
rect 17300 12580 17301 12620
rect 17259 12571 17301 12580
rect 17452 12620 17492 13994
rect 17452 12571 17492 12580
rect 17260 12536 17300 12571
rect 17260 12485 17300 12496
rect 17548 12452 17588 14512
rect 17740 14048 17780 14057
rect 17643 13964 17685 13973
rect 17740 13964 17780 14008
rect 17643 13924 17644 13964
rect 17684 13924 17780 13964
rect 17643 13915 17685 13924
rect 17356 12412 17588 12452
rect 17836 12452 17876 12461
rect 17260 10184 17300 10195
rect 17260 10109 17300 10144
rect 17259 10100 17301 10109
rect 17259 10060 17260 10100
rect 17300 10060 17301 10100
rect 17259 10051 17301 10060
rect 17259 9764 17301 9773
rect 17259 9724 17260 9764
rect 17300 9724 17301 9764
rect 17259 9715 17301 9724
rect 17260 9680 17300 9715
rect 17260 9629 17300 9640
rect 17108 9472 17204 9512
rect 17068 8765 17108 9472
rect 17163 8840 17205 8849
rect 17163 8800 17164 8840
rect 17204 8800 17205 8840
rect 17163 8791 17205 8800
rect 17067 8756 17109 8765
rect 17067 8716 17068 8756
rect 17108 8716 17109 8756
rect 17067 8707 17109 8716
rect 16972 8177 17012 8262
rect 16971 8168 17013 8177
rect 16971 8128 16972 8168
rect 17012 8128 17013 8168
rect 16971 8119 17013 8128
rect 17164 8000 17204 8791
rect 17259 8252 17301 8261
rect 17259 8212 17260 8252
rect 17300 8212 17301 8252
rect 17259 8203 17301 8212
rect 16636 7958 16676 7967
rect 16876 7960 17012 8000
rect 16636 7916 16676 7918
rect 16636 7876 16916 7916
rect 16683 7160 16725 7169
rect 16683 7120 16684 7160
rect 16724 7120 16725 7160
rect 16683 7111 16725 7120
rect 16587 6908 16629 6917
rect 16587 6868 16588 6908
rect 16628 6868 16629 6908
rect 16587 6859 16629 6868
rect 16491 5060 16533 5069
rect 16491 5020 16492 5060
rect 16532 5020 16533 5060
rect 16491 5011 16533 5020
rect 16396 4003 16436 4012
rect 16300 2827 16340 2836
rect 16108 2540 16148 2584
rect 16108 2500 16340 2540
rect 16012 1996 16148 2036
rect 16011 1868 16053 1877
rect 16011 1828 16012 1868
rect 16052 1828 16053 1868
rect 16011 1819 16053 1828
rect 16012 1734 16052 1819
rect 16012 1196 16052 1205
rect 15916 1156 16012 1196
rect 16012 1147 16052 1156
rect 16011 1028 16053 1037
rect 16011 988 16012 1028
rect 16052 988 16053 1028
rect 16011 979 16053 988
rect 15820 944 15860 953
rect 15723 776 15765 785
rect 15723 736 15724 776
rect 15764 736 15765 776
rect 15723 727 15765 736
rect 15820 533 15860 904
rect 15819 524 15861 533
rect 15819 484 15820 524
rect 15860 484 15861 524
rect 15819 475 15861 484
rect 15819 356 15861 365
rect 15819 316 15820 356
rect 15860 316 15861 356
rect 15819 307 15861 316
rect 15820 80 15860 307
rect 16012 80 16052 979
rect 16108 692 16148 1996
rect 16204 1700 16244 1709
rect 16204 869 16244 1660
rect 16300 1037 16340 2500
rect 16396 1877 16436 1962
rect 16395 1868 16437 1877
rect 16395 1828 16396 1868
rect 16436 1828 16437 1868
rect 16395 1819 16437 1828
rect 16588 1700 16628 6859
rect 16684 6488 16724 7111
rect 16876 6656 16916 7876
rect 16876 6607 16916 6616
rect 16684 6439 16724 6448
rect 16875 6488 16917 6497
rect 16875 6448 16876 6488
rect 16916 6448 16917 6488
rect 16875 6439 16917 6448
rect 16732 5657 16772 5666
rect 16772 5617 16820 5648
rect 16732 5608 16820 5617
rect 16683 5228 16725 5237
rect 16683 5188 16684 5228
rect 16724 5188 16725 5228
rect 16780 5228 16820 5608
rect 16876 5564 16916 6439
rect 16876 5515 16916 5524
rect 16972 5405 17012 7960
rect 17164 7925 17204 7960
rect 17163 7916 17205 7925
rect 17163 7876 17164 7916
rect 17204 7876 17205 7916
rect 17163 7867 17205 7876
rect 17163 7328 17205 7337
rect 17163 7288 17164 7328
rect 17204 7288 17205 7328
rect 17163 7279 17205 7288
rect 17164 6488 17204 7279
rect 17164 6439 17204 6448
rect 17164 5648 17204 5657
rect 17068 5608 17164 5648
rect 16971 5396 17013 5405
rect 16971 5356 16972 5396
rect 17012 5356 17013 5396
rect 16971 5347 17013 5356
rect 17068 5228 17108 5608
rect 17164 5599 17204 5608
rect 17260 5648 17300 8203
rect 17260 5573 17300 5608
rect 17259 5564 17301 5573
rect 17259 5524 17260 5564
rect 17300 5524 17301 5564
rect 17259 5515 17301 5524
rect 17259 5396 17301 5405
rect 17259 5356 17260 5396
rect 17300 5356 17301 5396
rect 17259 5347 17301 5356
rect 16780 5188 16916 5228
rect 16683 5179 16725 5188
rect 16684 4808 16724 5179
rect 16780 4985 16820 5070
rect 16779 4976 16821 4985
rect 16779 4936 16780 4976
rect 16820 4936 16821 4976
rect 16779 4927 16821 4936
rect 16684 4768 16820 4808
rect 16684 3464 16724 3473
rect 16684 2801 16724 3424
rect 16683 2792 16725 2801
rect 16683 2752 16684 2792
rect 16724 2752 16725 2792
rect 16683 2743 16725 2752
rect 16396 1660 16628 1700
rect 16299 1028 16341 1037
rect 16299 988 16300 1028
rect 16340 988 16341 1028
rect 16299 979 16341 988
rect 16203 860 16245 869
rect 16203 820 16204 860
rect 16244 820 16245 860
rect 16203 811 16245 820
rect 16108 652 16244 692
rect 16204 80 16244 652
rect 16396 80 16436 1660
rect 16780 1616 16820 4768
rect 16876 3632 16916 5188
rect 16972 5188 17108 5228
rect 16972 5144 17012 5188
rect 16972 5095 17012 5104
rect 17260 5060 17300 5347
rect 17068 5020 17300 5060
rect 16971 4976 17013 4985
rect 16971 4936 16972 4976
rect 17012 4936 17013 4976
rect 16971 4927 17013 4936
rect 16876 3583 16916 3592
rect 16972 3464 17012 4927
rect 16876 3424 17012 3464
rect 16876 2633 16916 3424
rect 16875 2624 16917 2633
rect 16875 2584 16876 2624
rect 16916 2584 16917 2624
rect 16875 2575 16917 2584
rect 16588 1576 16820 1616
rect 16588 80 16628 1576
rect 16876 1532 16916 2575
rect 17068 2540 17108 5020
rect 17356 2540 17396 12412
rect 17643 12368 17685 12377
rect 17643 12328 17644 12368
rect 17684 12328 17685 12368
rect 17643 12319 17685 12328
rect 17644 12234 17684 12319
rect 17836 12032 17876 12412
rect 18124 12284 18164 12293
rect 17644 11992 17876 12032
rect 17932 12244 18124 12284
rect 17452 11701 17492 11710
rect 17452 11621 17492 11661
rect 17451 11612 17493 11621
rect 17451 11572 17452 11612
rect 17492 11572 17493 11612
rect 17451 11563 17493 11572
rect 17547 11528 17589 11537
rect 17547 11488 17548 11528
rect 17588 11488 17589 11528
rect 17547 11479 17589 11488
rect 17644 11528 17684 11992
rect 17835 11612 17877 11621
rect 17835 11572 17836 11612
rect 17876 11572 17877 11612
rect 17835 11563 17877 11572
rect 17644 11479 17684 11488
rect 17548 11360 17588 11479
rect 17836 11478 17876 11563
rect 17548 11320 17876 11360
rect 17740 11108 17780 11117
rect 17644 11068 17740 11108
rect 17644 9437 17684 11068
rect 17740 11059 17780 11068
rect 17739 9680 17781 9689
rect 17739 9640 17740 9680
rect 17780 9640 17781 9680
rect 17739 9631 17781 9640
rect 17740 9512 17780 9631
rect 17740 9463 17780 9472
rect 17643 9428 17685 9437
rect 17643 9388 17644 9428
rect 17684 9388 17685 9428
rect 17643 9379 17685 9388
rect 17739 8924 17781 8933
rect 17739 8884 17740 8924
rect 17780 8884 17781 8924
rect 17739 8875 17781 8884
rect 17452 8672 17492 8681
rect 17452 8177 17492 8632
rect 17547 8672 17589 8681
rect 17547 8632 17548 8672
rect 17588 8632 17589 8672
rect 17547 8623 17589 8632
rect 17451 8168 17493 8177
rect 17451 8128 17452 8168
rect 17492 8128 17493 8168
rect 17451 8119 17493 8128
rect 17548 8009 17588 8623
rect 17547 8000 17589 8009
rect 17547 7960 17548 8000
rect 17588 7960 17589 8000
rect 17547 7951 17589 7960
rect 17643 7328 17685 7337
rect 17643 7288 17644 7328
rect 17684 7288 17685 7328
rect 17643 7279 17685 7288
rect 17644 6833 17684 7279
rect 17643 6824 17685 6833
rect 17643 6784 17644 6824
rect 17684 6784 17685 6824
rect 17643 6775 17685 6784
rect 17644 5732 17684 6775
rect 17644 5683 17684 5692
rect 17740 5732 17780 8875
rect 17836 8756 17876 11320
rect 17932 11019 17972 12244
rect 18124 12235 18164 12244
rect 18220 12116 18260 14671
rect 18316 13385 18356 20131
rect 18412 16148 18452 20383
rect 18508 18761 18548 20560
rect 18604 19853 18644 20560
rect 18699 20600 18741 20609
rect 18699 20560 18700 20600
rect 18740 20560 18741 20600
rect 18699 20551 18741 20560
rect 18796 20180 18836 20980
rect 18700 20140 18836 20180
rect 18603 19844 18645 19853
rect 18603 19804 18604 19844
rect 18644 19804 18645 19844
rect 18603 19795 18645 19804
rect 18700 19508 18740 20140
rect 18808 19676 19176 19685
rect 18848 19636 18890 19676
rect 18930 19636 18972 19676
rect 19012 19636 19054 19676
rect 19094 19636 19136 19676
rect 18808 19627 19176 19636
rect 18700 19468 18836 19508
rect 18699 19340 18741 19349
rect 18699 19300 18700 19340
rect 18740 19300 18741 19340
rect 18699 19291 18741 19300
rect 18700 19256 18740 19291
rect 18700 19205 18740 19216
rect 18603 19088 18645 19097
rect 18603 19048 18604 19088
rect 18644 19048 18645 19088
rect 18603 19039 18645 19048
rect 18507 18752 18549 18761
rect 18507 18712 18508 18752
rect 18548 18712 18549 18752
rect 18507 18703 18549 18712
rect 18604 18584 18644 19039
rect 18556 18574 18644 18584
rect 18596 18544 18644 18574
rect 18700 18668 18740 18677
rect 18796 18668 18836 19468
rect 18891 19088 18933 19097
rect 18891 19048 18892 19088
rect 18932 19048 18933 19088
rect 18891 19039 18933 19048
rect 18892 18954 18932 19039
rect 18740 18628 18836 18668
rect 18556 18525 18596 18534
rect 18507 17660 18549 17669
rect 18507 17620 18508 17660
rect 18548 17620 18549 17660
rect 18507 17611 18549 17620
rect 18508 17067 18548 17611
rect 18700 17324 18740 18628
rect 18808 18164 19176 18173
rect 18848 18124 18890 18164
rect 18930 18124 18972 18164
rect 19012 18124 19054 18164
rect 19094 18124 19136 18164
rect 18808 18115 19176 18124
rect 18892 17744 18932 17753
rect 18892 17585 18932 17704
rect 19083 17660 19125 17669
rect 19083 17620 19084 17660
rect 19124 17620 19125 17660
rect 19083 17611 19125 17620
rect 18891 17576 18933 17585
rect 18891 17536 18892 17576
rect 18932 17536 18933 17576
rect 18891 17527 18933 17536
rect 19084 17526 19124 17611
rect 19275 17576 19317 17585
rect 19275 17536 19276 17576
rect 19316 17536 19317 17576
rect 19275 17527 19317 17536
rect 18508 17018 18548 17027
rect 18604 17284 18740 17324
rect 18507 16904 18549 16913
rect 18507 16864 18508 16904
rect 18548 16864 18549 16904
rect 18507 16855 18549 16864
rect 18315 13376 18357 13385
rect 18315 13336 18316 13376
rect 18356 13336 18357 13376
rect 18315 13327 18357 13336
rect 18124 12076 18260 12116
rect 18316 12536 18356 12545
rect 18028 11696 18068 11705
rect 18028 11444 18068 11656
rect 18027 11404 18068 11444
rect 18027 11360 18067 11404
rect 18027 11320 18068 11360
rect 18028 11033 18068 11320
rect 17932 10970 17972 10979
rect 18027 11024 18069 11033
rect 18027 10984 18028 11024
rect 18068 10984 18069 11024
rect 18027 10975 18069 10984
rect 18027 10604 18069 10613
rect 18027 10564 18028 10604
rect 18068 10564 18069 10604
rect 18027 10555 18069 10564
rect 17932 8756 17972 8765
rect 17836 8716 17932 8756
rect 17932 8707 17972 8716
rect 18028 8756 18068 10555
rect 18124 8933 18164 12076
rect 18316 11033 18356 12496
rect 18412 11537 18452 16108
rect 18411 11528 18453 11537
rect 18411 11488 18412 11528
rect 18452 11488 18453 11528
rect 18411 11479 18453 11488
rect 18508 11360 18548 16855
rect 18604 16652 18644 17284
rect 18699 17156 18741 17165
rect 18699 17116 18700 17156
rect 18740 17116 18741 17156
rect 18699 17107 18741 17116
rect 18700 17022 18740 17107
rect 18808 16652 19176 16661
rect 18604 16612 18740 16652
rect 18604 14725 18644 14734
rect 18604 14225 18644 14685
rect 18603 14216 18645 14225
rect 18603 14176 18604 14216
rect 18644 14176 18645 14216
rect 18603 14167 18645 14176
rect 18700 14141 18740 16612
rect 18848 16612 18890 16652
rect 18930 16612 18972 16652
rect 19012 16612 19054 16652
rect 19094 16612 19136 16652
rect 18808 16603 19176 16612
rect 18808 15140 19176 15149
rect 18848 15100 18890 15140
rect 18930 15100 18972 15140
rect 19012 15100 19054 15140
rect 19094 15100 19136 15140
rect 18808 15091 19176 15100
rect 19276 14972 19316 17527
rect 19372 17501 19412 23416
rect 19468 23288 19508 23297
rect 19508 23248 19700 23288
rect 19468 23239 19508 23248
rect 19660 23120 19700 23248
rect 19660 23071 19700 23080
rect 19755 23120 19797 23129
rect 19755 23080 19756 23120
rect 19796 23080 19797 23120
rect 19755 23071 19797 23080
rect 19852 23120 19892 23491
rect 19948 23288 19988 26683
rect 20044 26648 20084 27196
rect 20620 27152 20660 30463
rect 21387 30008 21429 30017
rect 21387 29968 21388 30008
rect 21428 29968 21429 30008
rect 21387 29959 21429 29968
rect 20044 26599 20084 26608
rect 20524 27112 20660 27152
rect 20048 26480 20416 26489
rect 20088 26440 20130 26480
rect 20170 26440 20212 26480
rect 20252 26440 20294 26480
rect 20334 26440 20376 26480
rect 20048 26431 20416 26440
rect 20048 24968 20416 24977
rect 20088 24928 20130 24968
rect 20170 24928 20212 24968
rect 20252 24928 20294 24968
rect 20334 24928 20376 24968
rect 20048 24919 20416 24928
rect 20044 23633 20084 23718
rect 20043 23624 20085 23633
rect 20043 23584 20044 23624
rect 20084 23584 20085 23624
rect 20043 23575 20085 23584
rect 20048 23456 20416 23465
rect 20088 23416 20130 23456
rect 20170 23416 20212 23456
rect 20252 23416 20294 23456
rect 20334 23416 20376 23456
rect 20048 23407 20416 23416
rect 19948 23239 19988 23248
rect 19852 23071 19892 23080
rect 19756 22986 19796 23071
rect 20048 21944 20416 21953
rect 20088 21904 20130 21944
rect 20170 21904 20212 21944
rect 20252 21904 20294 21944
rect 20334 21904 20376 21944
rect 20048 21895 20416 21904
rect 20048 20432 20416 20441
rect 20088 20392 20130 20432
rect 20170 20392 20212 20432
rect 20252 20392 20294 20432
rect 20334 20392 20376 20432
rect 20048 20383 20416 20392
rect 20048 18920 20416 18929
rect 20088 18880 20130 18920
rect 20170 18880 20212 18920
rect 20252 18880 20294 18920
rect 20334 18880 20376 18920
rect 20048 18871 20416 18880
rect 19371 17492 19413 17501
rect 19371 17452 19372 17492
rect 19412 17452 19413 17492
rect 19371 17443 19413 17452
rect 20048 17408 20416 17417
rect 20088 17368 20130 17408
rect 20170 17368 20212 17408
rect 20252 17368 20294 17408
rect 20334 17368 20376 17408
rect 20048 17359 20416 17368
rect 20048 15896 20416 15905
rect 20088 15856 20130 15896
rect 20170 15856 20212 15896
rect 20252 15856 20294 15896
rect 20334 15856 20376 15896
rect 20048 15847 20416 15856
rect 18988 14932 19316 14972
rect 18795 14552 18837 14561
rect 18795 14512 18796 14552
rect 18836 14512 18837 14552
rect 18795 14503 18837 14512
rect 18796 14418 18836 14503
rect 18699 14132 18741 14141
rect 18699 14092 18700 14132
rect 18740 14092 18741 14132
rect 18699 14083 18741 14092
rect 18988 14048 19028 14932
rect 20048 14384 20416 14393
rect 20088 14344 20130 14384
rect 20170 14344 20212 14384
rect 20252 14344 20294 14384
rect 20334 14344 20376 14384
rect 20048 14335 20416 14344
rect 19179 14216 19221 14225
rect 19179 14176 19180 14216
rect 19220 14176 19221 14216
rect 19179 14167 19221 14176
rect 19180 14082 19220 14167
rect 19275 14132 19317 14141
rect 19275 14092 19276 14132
rect 19316 14092 19317 14132
rect 19275 14083 19317 14092
rect 18988 13889 19028 14008
rect 18987 13880 19029 13889
rect 18987 13840 18988 13880
rect 19028 13840 19029 13880
rect 18987 13831 19029 13840
rect 18808 13628 19176 13637
rect 18848 13588 18890 13628
rect 18930 13588 18972 13628
rect 19012 13588 19054 13628
rect 19094 13588 19136 13628
rect 18808 13579 19176 13588
rect 18808 12116 19176 12125
rect 18848 12076 18890 12116
rect 18930 12076 18972 12116
rect 19012 12076 19054 12116
rect 19094 12076 19136 12116
rect 18808 12067 19176 12076
rect 19276 11948 19316 14083
rect 20048 12872 20416 12881
rect 20088 12832 20130 12872
rect 20170 12832 20212 12872
rect 20252 12832 20294 12872
rect 20334 12832 20376 12872
rect 20048 12823 20416 12832
rect 19563 12536 19605 12545
rect 19563 12496 19564 12536
rect 19604 12496 19605 12536
rect 19563 12487 19605 12496
rect 19564 12402 19604 12487
rect 18988 11908 19316 11948
rect 18508 11320 18644 11360
rect 18315 11024 18357 11033
rect 18315 10984 18316 11024
rect 18356 10984 18357 11024
rect 18315 10975 18357 10984
rect 18412 11024 18452 11033
rect 18412 10193 18452 10984
rect 18507 11024 18549 11033
rect 18507 10984 18508 11024
rect 18548 10984 18549 11024
rect 18507 10975 18549 10984
rect 18411 10184 18453 10193
rect 18411 10144 18412 10184
rect 18452 10144 18453 10184
rect 18411 10135 18453 10144
rect 18508 10184 18548 10975
rect 18508 10135 18548 10144
rect 18315 9512 18357 9521
rect 18315 9472 18316 9512
rect 18356 9472 18357 9512
rect 18315 9463 18357 9472
rect 18316 9101 18356 9463
rect 18315 9092 18357 9101
rect 18315 9052 18316 9092
rect 18356 9052 18357 9092
rect 18315 9043 18357 9052
rect 18123 8924 18165 8933
rect 18123 8884 18124 8924
rect 18164 8884 18165 8924
rect 18123 8875 18165 8884
rect 18068 8716 18260 8756
rect 18028 8707 18068 8716
rect 17740 5683 17780 5692
rect 18220 5648 18260 8716
rect 18316 8000 18356 9043
rect 18412 8672 18452 10135
rect 18508 8672 18548 8681
rect 18412 8632 18508 8672
rect 18508 8623 18548 8632
rect 18412 8000 18452 8009
rect 18316 7960 18412 8000
rect 18412 7951 18452 7960
rect 18604 7916 18644 11320
rect 18988 11024 19028 11908
rect 18988 10975 19028 10984
rect 19276 11696 19316 11705
rect 18892 10940 18932 10949
rect 18700 10900 18892 10940
rect 18700 10613 18740 10900
rect 18892 10891 18932 10900
rect 18699 10604 18741 10613
rect 18699 10564 18700 10604
rect 18740 10564 18741 10604
rect 18699 10555 18741 10564
rect 18808 10604 19176 10613
rect 18848 10564 18890 10604
rect 18930 10564 18972 10604
rect 19012 10564 19054 10604
rect 19094 10564 19136 10604
rect 18808 10555 19176 10564
rect 18699 10436 18741 10445
rect 18699 10396 18700 10436
rect 18740 10396 18741 10436
rect 18699 10387 18741 10396
rect 18700 10302 18740 10387
rect 19276 9521 19316 11656
rect 20048 11360 20416 11369
rect 20088 11320 20130 11360
rect 20170 11320 20212 11360
rect 20252 11320 20294 11360
rect 20334 11320 20376 11360
rect 20048 11311 20416 11320
rect 19372 11024 19412 11033
rect 18988 9512 19028 9521
rect 18988 9260 19028 9472
rect 19275 9512 19317 9521
rect 19275 9472 19276 9512
rect 19316 9472 19317 9512
rect 19275 9463 19317 9472
rect 18700 9220 19028 9260
rect 19180 9260 19220 9269
rect 19220 9220 19316 9260
rect 18700 8849 18740 9220
rect 19180 9211 19220 9220
rect 18808 9092 19176 9101
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 18808 9043 19176 9052
rect 18699 8840 18741 8849
rect 18699 8800 18700 8840
rect 18740 8800 18741 8840
rect 18699 8791 18741 8800
rect 19036 8681 19076 8690
rect 19276 8672 19316 9220
rect 19076 8641 19316 8672
rect 19036 8632 19316 8641
rect 19180 8504 19220 8513
rect 19180 7925 19220 8464
rect 19372 8009 19412 10984
rect 19468 11024 19508 11033
rect 19468 10445 19508 10984
rect 19467 10436 19509 10445
rect 19467 10396 19468 10436
rect 19508 10396 19509 10436
rect 19467 10387 19509 10396
rect 20048 9848 20416 9857
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20048 9799 20416 9808
rect 20048 8336 20416 8345
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20048 8287 20416 8296
rect 19371 8000 19413 8009
rect 19371 7960 19372 8000
rect 19412 7960 19413 8000
rect 19371 7951 19413 7960
rect 18508 7876 18644 7916
rect 18795 7916 18837 7925
rect 18795 7876 18796 7916
rect 18836 7876 18837 7916
rect 18508 7832 18548 7876
rect 18795 7867 18837 7876
rect 19179 7916 19221 7925
rect 19179 7876 19180 7916
rect 19220 7876 19221 7916
rect 19179 7867 19221 7876
rect 18220 5599 18260 5608
rect 18412 7792 18548 7832
rect 18412 6488 18452 7792
rect 18796 7782 18836 7867
rect 18604 7748 18644 7757
rect 18412 4985 18452 6448
rect 18508 7708 18604 7748
rect 18508 6329 18548 7708
rect 18604 7699 18644 7708
rect 18808 7580 19176 7589
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 18808 7531 19176 7540
rect 20048 6824 20416 6833
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20048 6775 20416 6784
rect 18507 6320 18549 6329
rect 18507 6280 18508 6320
rect 18548 6280 18549 6320
rect 18507 6271 18549 6280
rect 18604 6236 18644 6245
rect 18644 6196 18740 6236
rect 18604 6187 18644 6196
rect 18700 5662 18740 6196
rect 18808 6068 19176 6077
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 18808 6019 19176 6028
rect 18700 5613 18740 5622
rect 18892 5480 18932 5489
rect 18892 5321 18932 5440
rect 18891 5312 18933 5321
rect 18891 5272 18892 5312
rect 18932 5272 18933 5312
rect 18891 5263 18933 5272
rect 20048 5312 20416 5321
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20048 5263 20416 5272
rect 18411 4976 18453 4985
rect 18411 4936 18412 4976
rect 18452 4936 18453 4976
rect 18411 4927 18453 4936
rect 18808 4556 19176 4565
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 18808 4507 19176 4516
rect 20048 3800 20416 3809
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20048 3751 20416 3760
rect 18808 3044 19176 3053
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 18808 2995 19176 3004
rect 16780 1492 16916 1532
rect 16972 2500 17108 2540
rect 17164 2500 17396 2540
rect 16780 80 16820 1492
rect 16972 80 17012 2500
rect 17164 80 17204 2500
rect 20048 2288 20416 2297
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20048 2239 20416 2248
rect 20524 1877 20564 27112
rect 21291 24548 21333 24557
rect 21291 24508 21292 24548
rect 21332 24508 21333 24548
rect 21291 24499 21333 24508
rect 20619 24044 20661 24053
rect 20619 24004 20620 24044
rect 20660 24004 20661 24044
rect 20619 23995 20661 24004
rect 20620 23465 20660 23995
rect 20619 23456 20661 23465
rect 20619 23416 20620 23456
rect 20660 23416 20661 23456
rect 20619 23407 20661 23416
rect 20619 18584 20661 18593
rect 20619 18544 20620 18584
rect 20660 18544 20661 18584
rect 20619 18535 20661 18544
rect 20620 16073 20660 18535
rect 20619 16064 20661 16073
rect 20619 16024 20620 16064
rect 20660 16024 20661 16064
rect 20619 16015 20661 16024
rect 21292 15401 21332 24499
rect 21388 18089 21428 29959
rect 21387 18080 21429 18089
rect 21387 18040 21388 18080
rect 21428 18040 21429 18080
rect 21387 18031 21429 18040
rect 21291 15392 21333 15401
rect 21291 15352 21292 15392
rect 21332 15352 21333 15392
rect 21291 15343 21333 15352
rect 21387 8672 21429 8681
rect 21387 8632 21388 8672
rect 21428 8632 21429 8672
rect 21387 8623 21429 8632
rect 21388 8177 21428 8623
rect 21387 8168 21429 8177
rect 21387 8128 21388 8168
rect 21428 8128 21429 8168
rect 21387 8119 21429 8128
rect 20523 1868 20565 1877
rect 20523 1828 20524 1868
rect 20564 1828 20565 1868
rect 20523 1819 20565 1828
rect 18808 1532 19176 1541
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 18808 1483 19176 1492
rect 17355 1280 17397 1289
rect 17355 1240 17356 1280
rect 17396 1240 17397 1280
rect 17355 1231 17397 1240
rect 17547 1280 17589 1289
rect 17547 1240 17548 1280
rect 17588 1240 17589 1280
rect 17547 1231 17589 1240
rect 18123 1280 18165 1289
rect 18123 1240 18124 1280
rect 18164 1240 18165 1280
rect 18123 1231 18165 1240
rect 18507 1280 18549 1289
rect 18507 1240 18508 1280
rect 18548 1240 18549 1280
rect 18507 1231 18549 1240
rect 19275 1280 19317 1289
rect 19275 1240 19276 1280
rect 19316 1240 19317 1280
rect 19275 1231 19317 1240
rect 19467 1280 19509 1289
rect 19467 1240 19468 1280
rect 19508 1240 19509 1280
rect 19467 1231 19509 1240
rect 17356 80 17396 1231
rect 17548 80 17588 1231
rect 17931 1028 17973 1037
rect 17931 988 17932 1028
rect 17972 988 17973 1028
rect 17931 979 17973 988
rect 17739 860 17781 869
rect 17739 820 17740 860
rect 17780 820 17781 860
rect 17739 811 17781 820
rect 17740 80 17780 811
rect 17932 80 17972 979
rect 18124 80 18164 1231
rect 18315 944 18357 953
rect 18315 904 18316 944
rect 18356 904 18357 944
rect 18315 895 18357 904
rect 18316 80 18356 895
rect 18508 80 18548 1231
rect 19083 1196 19125 1205
rect 19083 1156 19084 1196
rect 19124 1156 19125 1196
rect 19083 1147 19125 1156
rect 18891 1112 18933 1121
rect 18891 1072 18892 1112
rect 18932 1072 18933 1112
rect 18891 1063 18933 1072
rect 18699 608 18741 617
rect 18699 568 18700 608
rect 18740 568 18741 608
rect 18699 559 18741 568
rect 18700 80 18740 559
rect 18892 80 18932 1063
rect 19084 80 19124 1147
rect 19276 80 19316 1231
rect 19468 80 19508 1231
rect 20048 776 20416 785
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20048 727 20416 736
rect 4532 64 4552 80
rect 4472 0 4552 64
rect 4664 0 4744 80
rect 4856 0 4936 80
rect 5048 0 5128 80
rect 5240 0 5320 80
rect 5432 0 5512 80
rect 5624 0 5704 80
rect 5816 0 5896 80
rect 6008 0 6088 80
rect 6200 0 6280 80
rect 6392 0 6472 80
rect 6584 0 6664 80
rect 6776 0 6856 80
rect 6968 0 7048 80
rect 7160 0 7240 80
rect 7352 0 7432 80
rect 7544 0 7624 80
rect 7736 0 7816 80
rect 7928 0 8008 80
rect 8120 0 8200 80
rect 8312 0 8392 80
rect 8504 0 8584 80
rect 8696 0 8776 80
rect 8888 0 8968 80
rect 9080 0 9160 80
rect 9272 0 9352 80
rect 9464 0 9544 80
rect 9656 0 9736 80
rect 9848 0 9928 80
rect 10040 0 10120 80
rect 10232 0 10312 80
rect 10424 0 10504 80
rect 10616 0 10696 80
rect 10808 0 10888 80
rect 11000 0 11080 80
rect 11192 0 11272 80
rect 11384 0 11464 80
rect 11576 0 11656 80
rect 11768 0 11848 80
rect 11960 0 12040 80
rect 12152 0 12232 80
rect 12344 0 12424 80
rect 12536 0 12616 80
rect 12728 0 12808 80
rect 12920 0 13000 80
rect 13112 0 13192 80
rect 13304 0 13384 80
rect 13496 0 13576 80
rect 13688 0 13768 80
rect 13880 0 13960 80
rect 14072 0 14152 80
rect 14264 0 14344 80
rect 14456 0 14536 80
rect 14648 0 14728 80
rect 14840 0 14920 80
rect 15032 0 15112 80
rect 15224 0 15304 80
rect 15416 0 15496 80
rect 15608 0 15688 80
rect 15800 0 15880 80
rect 15992 0 16072 80
rect 16184 0 16264 80
rect 16376 0 16456 80
rect 16568 0 16648 80
rect 16760 0 16840 80
rect 16952 0 17032 80
rect 17144 0 17224 80
rect 17336 0 17416 80
rect 17528 0 17608 80
rect 17720 0 17800 80
rect 17912 0 17992 80
rect 18104 0 18184 80
rect 18296 0 18376 80
rect 18488 0 18568 80
rect 18680 0 18760 80
rect 18872 0 18952 80
rect 19064 0 19144 80
rect 19256 0 19336 80
rect 19448 0 19528 80
<< via2 >>
rect 268 85744 308 85784
rect 76 83728 116 83768
rect 1324 84064 1364 84104
rect 1132 82048 1172 82088
rect 364 79696 404 79736
rect 172 76336 212 76376
rect 268 72892 308 72932
rect 460 75076 500 75116
rect 940 75076 980 75116
rect 556 74320 596 74360
rect 364 72724 404 72764
rect 556 67348 596 67388
rect 1228 81964 1268 82004
rect 1228 81124 1268 81164
rect 1228 79360 1268 79400
rect 1804 83980 1844 84020
rect 2188 85912 2228 85952
rect 2092 84400 2132 84440
rect 2668 85240 2708 85280
rect 2188 83812 2228 83852
rect 3148 85240 3188 85280
rect 2956 84568 2996 84608
rect 3244 84316 3284 84356
rect 3052 83728 3092 83768
rect 1708 83476 1748 83516
rect 1708 82216 1748 82256
rect 1516 81124 1556 81164
rect 1420 80620 1460 80660
rect 1420 79360 1460 79400
rect 1612 80536 1652 80576
rect 1612 76000 1652 76040
rect 1804 81964 1844 82004
rect 1900 80452 1940 80492
rect 1804 80368 1844 80408
rect 1900 78940 1940 78980
rect 1804 78100 1844 78140
rect 1804 75916 1844 75956
rect 1420 74824 1460 74864
rect 1420 74488 1460 74528
rect 1228 74236 1268 74276
rect 1132 73312 1172 73352
rect 1036 72892 1076 72932
rect 1324 73984 1364 74024
rect 1324 73480 1364 73520
rect 2860 83476 2900 83516
rect 2572 82552 2612 82592
rect 3148 82552 3188 82592
rect 2476 82216 2516 82256
rect 2668 80704 2708 80744
rect 2572 80368 2612 80408
rect 2380 79108 2420 79148
rect 2284 76756 2324 76796
rect 2188 76252 2228 76292
rect 1900 75412 1940 75452
rect 1804 74824 1844 74864
rect 1708 74740 1748 74780
rect 1612 74320 1652 74360
rect 1708 74236 1748 74276
rect 1612 73648 1652 73688
rect 1516 73396 1556 73436
rect 1228 72976 1268 73016
rect 1132 72304 1172 72344
rect 1612 72640 1652 72680
rect 1420 72136 1460 72176
rect 1228 70540 1268 70580
rect 1324 69952 1364 69992
rect 1132 69196 1172 69236
rect 1036 68440 1076 68480
rect 1132 67600 1172 67640
rect 940 66928 980 66968
rect 172 65164 212 65204
rect 1228 66844 1268 66884
rect 1324 64996 1364 65036
rect 1516 72052 1556 72092
rect 2188 75916 2228 75956
rect 2092 75412 2132 75452
rect 1996 73900 2036 73940
rect 1900 73816 1940 73856
rect 1804 73480 1844 73520
rect 2188 73900 2228 73940
rect 1900 72136 1940 72176
rect 2092 72136 2132 72176
rect 2668 79696 2708 79736
rect 2668 79024 2708 79064
rect 2668 78856 2708 78896
rect 2572 78352 2612 78392
rect 2668 78100 2708 78140
rect 3148 81376 3188 81416
rect 2860 80620 2900 80660
rect 2860 79108 2900 79148
rect 2956 78016 2996 78056
rect 2956 77512 2996 77552
rect 2476 76756 2516 76796
rect 2572 75916 2612 75956
rect 2380 75160 2420 75200
rect 2764 75160 2804 75200
rect 2284 73816 2324 73856
rect 2380 73648 2420 73688
rect 2572 74824 2612 74864
rect 2668 74572 2708 74612
rect 2860 74740 2900 74780
rect 2860 74488 2900 74528
rect 2764 74404 2804 74444
rect 2764 74236 2804 74276
rect 2572 73732 2612 73772
rect 2284 72052 2324 72092
rect 1804 67768 1844 67808
rect 1708 66928 1748 66968
rect 1612 65416 1652 65456
rect 1708 65332 1748 65372
rect 1804 65248 1844 65288
rect 1516 64996 1556 65036
rect 1804 64996 1844 65036
rect 1132 63736 1172 63776
rect 1324 64576 1364 64616
rect 1420 62980 1460 63020
rect 1708 62392 1748 62432
rect 1612 61888 1652 61928
rect 1612 59956 1652 59996
rect 1516 59704 1556 59744
rect 1996 67600 2036 67640
rect 1900 64156 1940 64196
rect 2188 71380 2228 71420
rect 2188 68188 2228 68228
rect 2476 72976 2516 73016
rect 2476 72052 2516 72092
rect 2476 71884 2516 71924
rect 2668 71380 2708 71420
rect 2668 71212 2708 71252
rect 2572 70624 2612 70664
rect 2380 70540 2420 70580
rect 2476 69952 2516 69992
rect 2668 69952 2708 69992
rect 2668 69700 2708 69740
rect 2860 74152 2900 74192
rect 3148 79360 3188 79400
rect 3148 79024 3188 79064
rect 3436 84568 3476 84608
rect 3724 85828 3764 85868
rect 4300 85744 4340 85784
rect 3688 84652 3728 84692
rect 3770 84652 3810 84692
rect 3852 84652 3892 84692
rect 3934 84652 3974 84692
rect 4016 84652 4056 84692
rect 3628 84148 3668 84188
rect 4204 84820 4244 84860
rect 4300 83728 4340 83768
rect 3628 83308 3668 83348
rect 3688 83140 3728 83180
rect 3770 83140 3810 83180
rect 3852 83140 3892 83180
rect 3934 83140 3974 83180
rect 4016 83140 4056 83180
rect 3436 82048 3476 82088
rect 3436 81712 3476 81752
rect 3340 80032 3380 80072
rect 3724 82048 3764 82088
rect 4108 82720 4148 82760
rect 4108 82552 4148 82592
rect 3820 81880 3860 81920
rect 4108 81796 4148 81836
rect 3688 81628 3728 81668
rect 3770 81628 3810 81668
rect 3852 81628 3892 81668
rect 3934 81628 3974 81668
rect 4016 81628 4056 81668
rect 4012 81460 4052 81500
rect 3724 80368 3764 80408
rect 4396 83476 4436 83516
rect 4684 84820 4724 84860
rect 5260 84400 5300 84440
rect 5068 84064 5108 84104
rect 4928 83896 4968 83936
rect 5010 83896 5050 83936
rect 5092 83896 5132 83936
rect 5174 83896 5214 83936
rect 5256 83896 5296 83936
rect 6028 84484 6068 84524
rect 6604 84484 6644 84524
rect 5644 84400 5684 84440
rect 5836 84400 5876 84440
rect 6220 84400 6260 84440
rect 6412 84400 6452 84440
rect 6796 84400 6836 84440
rect 6988 84400 7028 84440
rect 5548 84232 5588 84272
rect 5548 83812 5588 83852
rect 6412 83980 6452 84020
rect 6220 83812 6260 83852
rect 7180 83812 7220 83852
rect 6988 83728 7028 83768
rect 5644 83644 5684 83684
rect 4972 83308 5012 83348
rect 4684 82468 4724 82508
rect 3688 80116 3728 80156
rect 3770 80116 3810 80156
rect 3852 80116 3892 80156
rect 3934 80116 3974 80156
rect 4016 80116 4056 80156
rect 3724 79612 3764 79652
rect 3148 78016 3188 78056
rect 3052 75244 3092 75284
rect 3052 74572 3092 74612
rect 3052 74404 3092 74444
rect 2956 73396 2996 73436
rect 3340 78184 3380 78224
rect 3340 77932 3380 77972
rect 3436 77596 3476 77636
rect 3436 77428 3476 77468
rect 3340 76756 3380 76796
rect 4108 79780 4148 79820
rect 4204 79696 4244 79736
rect 4300 79612 4340 79652
rect 4204 78940 4244 78980
rect 3688 78604 3728 78644
rect 3770 78604 3810 78644
rect 3852 78604 3892 78644
rect 3934 78604 3974 78644
rect 4016 78604 4056 78644
rect 3916 78436 3956 78476
rect 3688 77092 3728 77132
rect 3770 77092 3810 77132
rect 3852 77092 3892 77132
rect 3934 77092 3974 77132
rect 4016 77092 4056 77132
rect 4300 78016 4340 78056
rect 4204 77596 4244 77636
rect 4108 76672 4148 76712
rect 3244 76252 3284 76292
rect 3244 74488 3284 74528
rect 3148 73564 3188 73604
rect 3148 73396 3188 73436
rect 3052 73144 3092 73184
rect 2860 72724 2900 72764
rect 2956 72388 2996 72428
rect 3532 76504 3572 76544
rect 3688 75580 3728 75620
rect 3770 75580 3810 75620
rect 3852 75580 3892 75620
rect 3934 75580 3974 75620
rect 4016 75580 4056 75620
rect 3724 75412 3764 75452
rect 4108 74992 4148 75032
rect 4108 74488 4148 74528
rect 3532 74320 3572 74360
rect 3724 74320 3764 74360
rect 3436 74236 3476 74276
rect 3688 74068 3728 74108
rect 3770 74068 3810 74108
rect 3852 74068 3892 74108
rect 3934 74068 3974 74108
rect 4016 74068 4056 74108
rect 3340 73480 3380 73520
rect 3532 73060 3572 73100
rect 3436 72724 3476 72764
rect 3340 72556 3380 72596
rect 3244 72388 3284 72428
rect 2956 72052 2996 72092
rect 2860 71464 2900 71504
rect 3052 71212 3092 71252
rect 2860 71128 2900 71168
rect 2956 70708 2996 70748
rect 2860 70624 2900 70664
rect 2860 70036 2900 70076
rect 3052 69952 3092 69992
rect 3244 72052 3284 72092
rect 2860 69700 2900 69740
rect 2476 69196 2516 69236
rect 2572 68860 2612 68900
rect 2380 68440 2420 68480
rect 2380 68188 2420 68228
rect 2092 66508 2132 66548
rect 2476 67768 2516 67808
rect 2476 67600 2516 67640
rect 2572 67516 2612 67556
rect 2572 67096 2612 67136
rect 2284 66508 2324 66548
rect 2572 66172 2612 66212
rect 2188 65752 2228 65792
rect 2092 65584 2132 65624
rect 2956 68944 2996 68984
rect 2860 67768 2900 67808
rect 2860 67516 2900 67556
rect 2668 65920 2708 65960
rect 2572 65248 2612 65288
rect 2092 65080 2132 65120
rect 2476 65080 2516 65120
rect 1996 62560 2036 62600
rect 2572 64996 2612 65036
rect 2668 64660 2708 64700
rect 2284 64492 2324 64532
rect 2380 63148 2420 63188
rect 556 57856 596 57896
rect 748 56848 788 56888
rect 556 53740 596 53780
rect 1516 58276 1556 58316
rect 1900 58864 1940 58904
rect 2764 64576 2804 64616
rect 2476 62644 2516 62684
rect 2380 61636 2420 61676
rect 2188 61552 2228 61592
rect 2284 60544 2324 60584
rect 2764 64324 2804 64364
rect 2668 64240 2708 64280
rect 2956 67348 2996 67388
rect 2956 67012 2996 67052
rect 2956 66676 2996 66716
rect 2956 65332 2996 65372
rect 2956 64660 2996 64700
rect 2956 63232 2996 63272
rect 2956 63064 2996 63104
rect 2668 62896 2708 62936
rect 3148 68524 3188 68564
rect 3244 67516 3284 67556
rect 3148 67012 3188 67052
rect 3148 65584 3188 65624
rect 3688 72556 3728 72596
rect 3770 72556 3810 72596
rect 3852 72556 3892 72596
rect 3934 72556 3974 72596
rect 4016 72556 4056 72596
rect 3724 71968 3764 72008
rect 3916 71884 3956 71924
rect 3628 71800 3668 71840
rect 3532 71464 3572 71504
rect 3916 71464 3956 71504
rect 4108 71464 4148 71504
rect 3628 71212 3668 71252
rect 3688 71044 3728 71084
rect 3770 71044 3810 71084
rect 3852 71044 3892 71084
rect 3934 71044 3974 71084
rect 4016 71044 4056 71084
rect 3532 70624 3572 70664
rect 3724 70792 3764 70832
rect 3436 68944 3476 68984
rect 4012 70708 4052 70748
rect 4588 80452 4628 80492
rect 4492 78856 4532 78896
rect 4928 82384 4968 82424
rect 5010 82384 5050 82424
rect 5092 82384 5132 82424
rect 5174 82384 5214 82424
rect 5256 82384 5296 82424
rect 4972 81796 5012 81836
rect 4928 80872 4968 80912
rect 5010 80872 5050 80912
rect 5092 80872 5132 80912
rect 5174 80872 5214 80912
rect 5256 80872 5296 80912
rect 4972 80620 5012 80660
rect 4972 80452 5012 80492
rect 5164 80284 5204 80324
rect 5740 83476 5780 83516
rect 5740 80620 5780 80660
rect 5452 80284 5492 80324
rect 4928 79360 4968 79400
rect 5010 79360 5050 79400
rect 5092 79360 5132 79400
rect 5174 79360 5214 79400
rect 5256 79360 5296 79400
rect 5260 79108 5300 79148
rect 4876 78856 4916 78896
rect 5260 78520 5300 78560
rect 5548 79948 5588 79988
rect 5548 79360 5588 79400
rect 5452 79276 5492 79316
rect 6508 83056 6548 83096
rect 6316 81712 6356 81752
rect 6028 80452 6068 80492
rect 5932 80368 5972 80408
rect 5548 79108 5588 79148
rect 5452 79024 5492 79064
rect 5356 78352 5396 78392
rect 5932 79192 5972 79232
rect 5836 79024 5876 79064
rect 4876 78100 4916 78140
rect 4588 76840 4628 76880
rect 4492 76756 4532 76796
rect 4396 76672 4436 76712
rect 4396 76000 4436 76040
rect 4396 74992 4436 75032
rect 4300 74236 4340 74276
rect 4972 78016 5012 78056
rect 4928 77848 4968 77888
rect 5010 77848 5050 77888
rect 5092 77848 5132 77888
rect 5174 77848 5214 77888
rect 5256 77848 5296 77888
rect 5836 78856 5876 78896
rect 5644 78352 5684 78392
rect 5260 77512 5300 77552
rect 5356 76672 5396 76712
rect 4928 76336 4968 76376
rect 5010 76336 5050 76376
rect 5092 76336 5132 76376
rect 5174 76336 5214 76376
rect 5256 76336 5296 76376
rect 5452 76252 5492 76292
rect 5068 76000 5108 76040
rect 4972 75832 5012 75872
rect 4876 75580 4916 75620
rect 4780 75496 4820 75536
rect 5644 76756 5684 76796
rect 5644 76504 5684 76544
rect 5452 75916 5492 75956
rect 5548 75748 5588 75788
rect 6028 77680 6068 77720
rect 6028 77512 6068 77552
rect 6220 80536 6260 80576
rect 5836 76504 5876 76544
rect 5740 76168 5780 76208
rect 5644 75580 5684 75620
rect 5452 75496 5492 75536
rect 5356 75412 5396 75452
rect 5260 75160 5300 75200
rect 4780 74908 4820 74948
rect 4928 74824 4968 74864
rect 5010 74824 5050 74864
rect 5092 74824 5132 74864
rect 5174 74824 5214 74864
rect 5256 74824 5296 74864
rect 5452 74740 5492 74780
rect 5644 75328 5684 75368
rect 5548 74572 5588 74612
rect 5452 74488 5492 74528
rect 5548 74320 5588 74360
rect 5452 74236 5492 74276
rect 5356 73900 5396 73940
rect 5260 73732 5300 73772
rect 5836 74824 5876 74864
rect 5740 74740 5780 74780
rect 4684 73312 4724 73352
rect 4492 72976 4532 73016
rect 4588 72388 4628 72428
rect 4588 71968 4628 72008
rect 4928 73312 4968 73352
rect 5010 73312 5050 73352
rect 5092 73312 5132 73352
rect 5174 73312 5214 73352
rect 5256 73312 5296 73352
rect 4780 71884 4820 71924
rect 4684 71548 4724 71588
rect 4108 69952 4148 69992
rect 4300 69952 4340 69992
rect 3724 69700 3764 69740
rect 3688 69532 3728 69572
rect 3770 69532 3810 69572
rect 3852 69532 3892 69572
rect 3934 69532 3974 69572
rect 4016 69532 4056 69572
rect 3628 69364 3668 69404
rect 3820 68692 3860 68732
rect 3628 68524 3668 68564
rect 3820 68440 3860 68480
rect 3820 68188 3860 68228
rect 4684 70036 4724 70076
rect 4588 69952 4628 69992
rect 4108 68524 4148 68564
rect 4204 68440 4244 68480
rect 3688 68020 3728 68060
rect 3770 68020 3810 68060
rect 3852 68020 3892 68060
rect 3934 68020 3974 68060
rect 4016 68020 4056 68060
rect 4204 68020 4244 68060
rect 3628 67600 3668 67640
rect 3532 67516 3572 67556
rect 3436 67432 3476 67472
rect 3532 67012 3572 67052
rect 3436 66760 3476 66800
rect 4492 68440 4532 68480
rect 4684 69280 4724 69320
rect 4928 71800 4968 71840
rect 5010 71800 5050 71840
rect 5092 71800 5132 71840
rect 5174 71800 5214 71840
rect 5256 71800 5296 71840
rect 5068 71464 5108 71504
rect 5260 71380 5300 71420
rect 5836 73900 5876 73940
rect 6796 83224 6836 83264
rect 6892 82804 6932 82844
rect 6604 81880 6644 81920
rect 6796 80620 6836 80660
rect 6412 80032 6452 80072
rect 6412 77512 6452 77552
rect 6316 76840 6356 76880
rect 6220 76756 6260 76796
rect 6124 76672 6164 76712
rect 6028 76588 6068 76628
rect 6220 76504 6260 76544
rect 6028 75076 6068 75116
rect 5740 72556 5780 72596
rect 5932 72724 5972 72764
rect 6220 75160 6260 75200
rect 5836 72472 5876 72512
rect 6124 72472 6164 72512
rect 5932 72388 5972 72428
rect 5644 72136 5684 72176
rect 5452 72052 5492 72092
rect 6604 77680 6644 77720
rect 6508 76924 6548 76964
rect 6508 76672 6548 76712
rect 7372 83392 7412 83432
rect 7756 83728 7796 83768
rect 7756 83476 7796 83516
rect 8332 84316 8372 84356
rect 8332 84148 8372 84188
rect 8140 83728 8180 83768
rect 8140 83224 8180 83264
rect 7468 83140 7508 83180
rect 8044 83140 8084 83180
rect 7276 82804 7316 82844
rect 7948 82720 7988 82760
rect 6988 81040 7028 81080
rect 6988 79024 7028 79064
rect 6988 78772 7028 78812
rect 6892 77512 6932 77552
rect 6700 77176 6740 77216
rect 7372 81712 7412 81752
rect 7372 81292 7412 81332
rect 7564 81040 7604 81080
rect 7276 79276 7316 79316
rect 7180 79192 7220 79232
rect 7180 78184 7220 78224
rect 8044 79276 8084 79316
rect 7372 79192 7412 79232
rect 7948 79192 7988 79232
rect 7468 79024 7508 79064
rect 7468 78184 7508 78224
rect 7276 77176 7316 77216
rect 6604 76504 6644 76544
rect 7276 77008 7316 77048
rect 6700 76420 6740 76460
rect 6700 76168 6740 76208
rect 6604 76084 6644 76124
rect 6508 76035 6548 76040
rect 6508 76000 6548 76035
rect 6508 75580 6548 75620
rect 6412 74404 6452 74444
rect 6412 74236 6452 74276
rect 6412 73732 6452 73772
rect 6316 73396 6356 73436
rect 6316 72724 6356 72764
rect 5447 71464 5452 71504
rect 5452 71464 5487 71504
rect 5548 71464 5588 71504
rect 5740 71380 5780 71420
rect 5260 70792 5300 70832
rect 5164 70624 5204 70664
rect 5356 70624 5396 70664
rect 4928 70288 4968 70328
rect 5010 70288 5050 70328
rect 5092 70288 5132 70328
rect 5174 70288 5214 70328
rect 5256 70288 5296 70328
rect 5260 69028 5300 69068
rect 4928 68776 4968 68816
rect 5010 68776 5050 68816
rect 5092 68776 5132 68816
rect 5174 68776 5214 68816
rect 5256 68776 5296 68816
rect 4684 68524 4724 68564
rect 4492 68020 4532 68060
rect 4588 67852 4628 67892
rect 4492 67600 4532 67640
rect 4108 67432 4148 67472
rect 3688 66508 3728 66548
rect 3770 66508 3810 66548
rect 3852 66508 3892 66548
rect 3934 66508 3974 66548
rect 4016 66508 4056 66548
rect 5164 68608 5204 68648
rect 4876 67852 4916 67892
rect 5260 67852 5300 67892
rect 4928 67264 4968 67304
rect 5010 67264 5050 67304
rect 5092 67264 5132 67304
rect 5174 67264 5214 67304
rect 5256 67264 5296 67304
rect 5932 71548 5972 71588
rect 6028 71380 6068 71420
rect 5740 70792 5780 70832
rect 5644 70036 5684 70076
rect 5548 69616 5588 69656
rect 5452 69280 5492 69320
rect 5452 69028 5492 69068
rect 5356 67180 5396 67220
rect 4492 66760 4532 66800
rect 4396 66676 4436 66716
rect 4300 66340 4340 66380
rect 3724 66172 3764 66212
rect 3628 66088 3668 66128
rect 3532 66004 3572 66044
rect 3916 66088 3956 66128
rect 3340 65668 3380 65708
rect 3340 65500 3380 65540
rect 4108 66088 4148 66128
rect 4204 65752 4244 65792
rect 3532 65668 3572 65708
rect 4012 65668 4052 65708
rect 3436 65416 3476 65456
rect 3532 65332 3572 65372
rect 4300 65332 4340 65372
rect 3532 65164 3572 65204
rect 3688 64996 3728 65036
rect 3770 64996 3810 65036
rect 3852 64996 3892 65036
rect 3934 64996 3974 65036
rect 4016 64996 4056 65036
rect 4012 64660 4052 64700
rect 3532 64576 3572 64616
rect 3244 64324 3284 64364
rect 3148 63904 3188 63944
rect 3052 62980 3092 63020
rect 2764 62728 2804 62768
rect 2764 60964 2804 61004
rect 2668 60880 2708 60920
rect 3052 62728 3092 62768
rect 2956 61048 2996 61088
rect 2956 60376 2996 60416
rect 3340 63316 3380 63356
rect 3340 63148 3380 63188
rect 3148 62140 3188 62180
rect 3244 61636 3284 61676
rect 3148 61216 3188 61256
rect 2668 59788 2708 59828
rect 2956 59956 2996 59996
rect 3820 64072 3860 64112
rect 4492 66172 4532 66212
rect 4492 65332 4532 65372
rect 3688 63484 3728 63524
rect 3770 63484 3810 63524
rect 3852 63484 3892 63524
rect 3934 63484 3974 63524
rect 4016 63484 4056 63524
rect 3724 63316 3764 63356
rect 3532 63232 3572 63272
rect 3436 61804 3476 61844
rect 2860 59872 2900 59912
rect 2956 59788 2996 59828
rect 2668 59452 2708 59492
rect 2092 59284 2132 59324
rect 2572 58696 2612 58736
rect 1804 57520 1844 57560
rect 1612 56512 1652 56552
rect 1324 53908 1364 53948
rect 748 52900 788 52940
rect 1324 52648 1364 52688
rect 1228 51304 1268 51344
rect 1228 48616 1268 48656
rect 1228 46264 1268 46304
rect 1228 45760 1268 45800
rect 1516 53320 1556 53360
rect 1708 53824 1748 53864
rect 1420 52564 1460 52604
rect 1804 53488 1844 53528
rect 2092 55672 2132 55712
rect 1996 55084 2036 55124
rect 1996 54748 2036 54788
rect 1900 52732 1940 52772
rect 1804 52396 1844 52436
rect 1420 52144 1460 52184
rect 1420 51892 1460 51932
rect 1516 50800 1556 50840
rect 1516 50380 1556 50420
rect 1516 49456 1556 49496
rect 1516 48448 1556 48488
rect 1420 47944 1460 47984
rect 1708 52312 1748 52352
rect 1996 52564 2036 52604
rect 3436 60880 3476 60920
rect 3340 60544 3380 60584
rect 3340 59956 3380 59996
rect 3340 58612 3380 58652
rect 3724 62728 3764 62768
rect 3688 61972 3728 62012
rect 3770 61972 3810 62012
rect 3852 61972 3892 62012
rect 3934 61972 3974 62012
rect 4016 61972 4056 62012
rect 3724 61804 3764 61844
rect 3916 61720 3956 61760
rect 3820 61636 3860 61676
rect 4588 63904 4628 63944
rect 4492 62980 4532 63020
rect 4300 62644 4340 62684
rect 4204 62392 4244 62432
rect 4108 60712 4148 60752
rect 3688 60460 3728 60500
rect 3770 60460 3810 60500
rect 3852 60460 3892 60500
rect 3934 60460 3974 60500
rect 4016 60460 4056 60500
rect 3628 60292 3668 60332
rect 4492 62560 4532 62600
rect 4588 60964 4628 61004
rect 4780 66760 4820 66800
rect 5356 66760 5396 66800
rect 5740 68776 5780 68816
rect 5740 68608 5780 68648
rect 5548 68020 5588 68060
rect 4972 66676 5012 66716
rect 5068 66172 5108 66212
rect 4780 66004 4820 66044
rect 5452 66676 5492 66716
rect 5740 67600 5780 67640
rect 5740 66844 5780 66884
rect 5548 66256 5588 66296
rect 5164 66004 5204 66044
rect 5452 66004 5492 66044
rect 4972 65920 5012 65960
rect 5356 65836 5396 65876
rect 4928 65752 4968 65792
rect 5010 65752 5050 65792
rect 5092 65752 5132 65792
rect 5174 65752 5214 65792
rect 5256 65752 5296 65792
rect 4780 65248 4820 65288
rect 5164 65248 5204 65288
rect 4780 65080 4820 65120
rect 4780 64660 4820 64700
rect 5260 64912 5300 64952
rect 6508 73648 6548 73688
rect 6508 73480 6548 73520
rect 7084 76840 7124 76880
rect 6988 76000 7028 76040
rect 7180 76000 7220 76040
rect 7468 77260 7508 77300
rect 8140 78856 8180 78896
rect 7852 78772 7892 78812
rect 8428 83728 8468 83768
rect 8716 84904 8756 84944
rect 8812 84316 8852 84356
rect 9100 84904 9140 84944
rect 8524 83392 8564 83432
rect 8332 78520 8372 78560
rect 9004 83308 9044 83348
rect 8908 82216 8948 82256
rect 9004 80536 9044 80576
rect 8908 78940 8948 78980
rect 7948 78184 7988 78224
rect 7852 77512 7892 77552
rect 7756 76756 7796 76796
rect 7756 76168 7796 76208
rect 7468 76000 7508 76040
rect 7948 76756 7988 76796
rect 8524 77512 8564 77552
rect 8332 77428 8372 77468
rect 8428 77260 8468 77300
rect 8332 77176 8372 77216
rect 8236 76672 8276 76712
rect 7372 75832 7412 75872
rect 7564 75832 7604 75872
rect 6988 75580 7028 75620
rect 6892 74236 6932 74276
rect 6796 74152 6836 74192
rect 7361 75664 7401 75704
rect 6892 74068 6932 74108
rect 6796 73900 6836 73940
rect 6604 73312 6644 73352
rect 6508 73228 6548 73268
rect 6604 73144 6644 73184
rect 6412 72136 6452 72176
rect 6892 72640 6932 72680
rect 6316 72052 6356 72092
rect 6220 71968 6260 72008
rect 6412 71800 6452 71840
rect 6220 71296 6260 71336
rect 6028 70540 6068 70580
rect 6508 71380 6548 71420
rect 7564 75664 7604 75704
rect 7468 75580 7508 75620
rect 7564 74656 7604 74696
rect 7468 74152 7508 74192
rect 7372 74068 7412 74108
rect 7180 73648 7220 73688
rect 7281 73396 7321 73436
rect 7180 73312 7220 73352
rect 7084 73228 7124 73268
rect 6988 72052 7028 72092
rect 6796 71968 6836 72008
rect 7180 72388 7220 72428
rect 7084 71548 7124 71588
rect 6700 71464 6740 71504
rect 6604 71296 6644 71336
rect 6988 71296 7028 71336
rect 6892 71128 6932 71168
rect 6700 70792 6740 70832
rect 5932 70120 5972 70160
rect 6124 69868 6164 69908
rect 5932 69364 5972 69404
rect 6316 69952 6356 69992
rect 6316 69616 6356 69656
rect 6220 69280 6260 69320
rect 6124 68692 6164 68732
rect 5932 67768 5972 67808
rect 6028 67516 6068 67556
rect 6028 67264 6068 67304
rect 6220 68475 6260 68480
rect 6220 68440 6260 68475
rect 6124 67180 6164 67220
rect 5932 66592 5972 66632
rect 6028 66093 6068 66128
rect 6028 66088 6068 66093
rect 6508 69952 6548 69992
rect 6412 69112 6452 69152
rect 6796 70540 6836 70580
rect 7180 71128 7220 71168
rect 7372 71296 7412 71336
rect 7852 74236 7892 74276
rect 7756 74152 7796 74192
rect 7660 73396 7700 73436
rect 7756 71716 7796 71756
rect 7660 71296 7700 71336
rect 7084 70792 7124 70832
rect 7276 70792 7316 70832
rect 7180 70708 7220 70748
rect 7084 70624 7124 70664
rect 6892 70036 6932 70076
rect 6796 69952 6836 69992
rect 6892 69868 6932 69908
rect 6604 69616 6644 69656
rect 6700 69280 6740 69320
rect 6316 66592 6356 66632
rect 6700 68188 6740 68228
rect 6700 67852 6740 67892
rect 6604 67096 6644 67136
rect 6604 66760 6644 66800
rect 6508 66340 6548 66380
rect 6316 66088 6356 66128
rect 6220 65920 6260 65960
rect 5932 65752 5972 65792
rect 5740 65164 5780 65204
rect 5548 65080 5588 65120
rect 5356 64408 5396 64448
rect 4928 64240 4968 64280
rect 5010 64240 5050 64280
rect 5092 64240 5132 64280
rect 5174 64240 5214 64280
rect 5256 64240 5296 64280
rect 4928 62728 4968 62768
rect 5010 62728 5050 62768
rect 5092 62728 5132 62768
rect 5174 62728 5214 62768
rect 5256 62728 5296 62768
rect 4780 62560 4820 62600
rect 4780 61636 4820 61676
rect 4684 60376 4724 60416
rect 4928 61216 4968 61256
rect 5010 61216 5050 61256
rect 5092 61216 5132 61256
rect 5174 61216 5214 61256
rect 5256 61216 5296 61256
rect 5068 60880 5108 60920
rect 5452 64072 5492 64112
rect 5548 63904 5588 63944
rect 6508 66088 6548 66128
rect 6220 65500 6260 65540
rect 6028 64408 6068 64448
rect 5932 64324 5972 64364
rect 5836 64072 5876 64112
rect 5740 63904 5780 63944
rect 5452 62644 5492 62684
rect 5164 60628 5204 60668
rect 5356 60544 5396 60584
rect 5260 60460 5300 60500
rect 5164 60376 5204 60416
rect 4396 59704 4436 59744
rect 4396 59536 4436 59576
rect 3688 58948 3728 58988
rect 3770 58948 3810 58988
rect 3852 58948 3892 58988
rect 3934 58948 3974 58988
rect 4016 58948 4056 58988
rect 3724 58780 3764 58820
rect 3724 58276 3764 58316
rect 4300 58024 4340 58064
rect 3628 57856 3668 57896
rect 4108 57772 4148 57812
rect 2956 57016 2996 57056
rect 3436 57016 3476 57056
rect 3688 57436 3728 57476
rect 3770 57436 3810 57476
rect 3852 57436 3892 57476
rect 3934 57436 3974 57476
rect 4016 57436 4056 57476
rect 2860 56512 2900 56552
rect 2764 56344 2804 56384
rect 2668 56008 2708 56048
rect 3244 56848 3284 56888
rect 2956 56008 2996 56048
rect 3628 56848 3668 56888
rect 3340 56512 3380 56552
rect 2572 55420 2612 55460
rect 2860 55084 2900 55124
rect 3052 54832 3092 54872
rect 3052 54664 3092 54704
rect 2956 54328 2996 54368
rect 2956 54160 2996 54200
rect 2188 52648 2228 52688
rect 2572 53740 2612 53780
rect 2092 52312 2132 52352
rect 2380 52312 2420 52352
rect 2572 52312 2612 52352
rect 2092 52144 2132 52184
rect 2572 52144 2612 52184
rect 1900 51724 1940 51764
rect 2092 50548 2132 50588
rect 3820 57016 3860 57056
rect 4588 59032 4628 59072
rect 4588 58192 4628 58232
rect 4780 59872 4820 59912
rect 5740 62980 5780 63020
rect 6028 63904 6068 63944
rect 7276 69868 7316 69908
rect 6892 69196 6932 69236
rect 7084 69112 7124 69152
rect 7468 70792 7508 70832
rect 7468 70540 7508 70580
rect 7660 70624 7700 70664
rect 7372 69280 7412 69320
rect 6892 68860 6932 68900
rect 6892 68440 6932 68480
rect 7084 68020 7124 68060
rect 7276 68944 7316 68984
rect 6796 67516 6836 67556
rect 7084 67096 7124 67136
rect 6796 67012 6836 67052
rect 6892 66508 6932 66548
rect 6796 66340 6836 66380
rect 6700 65752 6740 65792
rect 6412 65416 6452 65456
rect 6604 65332 6644 65372
rect 6412 65248 6452 65288
rect 5932 63064 5972 63104
rect 6028 62896 6068 62936
rect 5836 62140 5876 62180
rect 5740 61888 5780 61928
rect 5644 61048 5684 61088
rect 5548 60376 5588 60416
rect 4492 57772 4532 57812
rect 4396 57016 4436 57056
rect 4204 56932 4244 56972
rect 3724 56512 3764 56552
rect 3436 55588 3476 55628
rect 3340 55084 3380 55124
rect 3340 54916 3380 54956
rect 3436 54748 3476 54788
rect 3436 53320 3476 53360
rect 2764 53236 2804 53276
rect 4396 56428 4436 56468
rect 4300 56260 4340 56300
rect 3688 55924 3728 55964
rect 3770 55924 3810 55964
rect 3852 55924 3892 55964
rect 3934 55924 3974 55964
rect 4016 55924 4056 55964
rect 3916 55336 3956 55376
rect 3820 54832 3860 54872
rect 3688 54412 3728 54452
rect 3770 54412 3810 54452
rect 3852 54412 3892 54452
rect 3934 54412 3974 54452
rect 4016 54412 4056 54452
rect 3724 54160 3764 54200
rect 3628 53908 3668 53948
rect 3628 53488 3668 53528
rect 2764 53068 2804 53108
rect 2668 52060 2708 52100
rect 2380 51724 2420 51764
rect 2956 52900 2996 52940
rect 2860 52312 2900 52352
rect 2764 51640 2804 51680
rect 2764 51136 2804 51176
rect 2668 50800 2708 50840
rect 1900 49876 1940 49916
rect 1708 49372 1748 49412
rect 2668 50296 2708 50336
rect 2476 50044 2516 50084
rect 2284 49372 2324 49412
rect 2380 48868 2420 48908
rect 3820 53992 3860 54032
rect 3916 53908 3956 53948
rect 4396 54916 4436 54956
rect 4396 54160 4436 54200
rect 4492 53992 4532 54032
rect 4204 53320 4244 53360
rect 3724 53068 3764 53108
rect 3916 53068 3956 53108
rect 3436 52900 3476 52940
rect 3148 51640 3188 51680
rect 3052 51052 3092 51092
rect 2956 50716 2996 50756
rect 2860 50044 2900 50084
rect 3052 49960 3092 50000
rect 2956 49456 2996 49496
rect 3340 50968 3380 51008
rect 3688 52900 3728 52940
rect 3770 52900 3810 52940
rect 3852 52900 3892 52940
rect 3934 52900 3974 52940
rect 4016 52900 4056 52940
rect 3724 52732 3764 52772
rect 3628 52480 3668 52520
rect 3820 52480 3860 52520
rect 4108 52060 4148 52100
rect 3628 51724 3668 51764
rect 4300 53068 4340 53108
rect 4396 52732 4436 52772
rect 3688 51388 3728 51428
rect 3770 51388 3810 51428
rect 3852 51388 3892 51428
rect 3934 51388 3974 51428
rect 4016 51388 4056 51428
rect 4012 50968 4052 51008
rect 1996 48616 2036 48656
rect 2284 48532 2324 48572
rect 1708 48112 1748 48152
rect 1804 48028 1844 48068
rect 1996 47944 2036 47984
rect 2668 48532 2708 48572
rect 2860 48196 2900 48236
rect 2476 48112 2516 48152
rect 2380 47272 2420 47312
rect 1996 47188 2036 47228
rect 1900 47104 1940 47144
rect 1516 46768 1556 46808
rect 2572 47944 2612 47984
rect 2284 45760 2324 45800
rect 2476 45760 2516 45800
rect 1708 45676 1748 45716
rect 1516 45424 1556 45464
rect 1324 42652 1364 42692
rect 2092 45256 2132 45296
rect 2092 45004 2132 45044
rect 1900 44416 1940 44456
rect 2380 45676 2420 45716
rect 2764 47860 2804 47900
rect 2668 46264 2708 46304
rect 2668 45760 2708 45800
rect 1996 44164 2036 44204
rect 2188 43996 2228 44036
rect 2476 44164 2516 44204
rect 1900 41224 1940 41264
rect 1420 41140 1460 41180
rect 1420 40468 1460 40508
rect 1708 40468 1748 40508
rect 2476 41476 2516 41516
rect 1324 40384 1364 40424
rect 1516 39880 1556 39920
rect 1420 39712 1460 39752
rect 940 39460 980 39500
rect 76 34840 116 34880
rect 76 34672 116 34712
rect 268 34084 308 34124
rect 172 32824 212 32864
rect 76 29128 116 29168
rect 748 31564 788 31604
rect 748 26608 788 26648
rect 268 21568 308 21608
rect 172 18880 212 18920
rect 76 13168 116 13208
rect 1324 38872 1364 38912
rect 1324 37696 1364 37736
rect 1516 39544 1556 39584
rect 1612 38284 1652 38324
rect 1612 38032 1652 38072
rect 1420 37444 1460 37484
rect 2668 43996 2708 44036
rect 2668 42820 2708 42860
rect 2668 41896 2708 41936
rect 2572 40384 2612 40424
rect 2380 40300 2420 40340
rect 2668 40300 2708 40340
rect 2572 39796 2612 39836
rect 1804 39544 1844 39584
rect 1420 37024 1460 37064
rect 1324 35848 1364 35888
rect 1228 34756 1268 34796
rect 1420 34756 1460 34796
rect 1132 34000 1172 34040
rect 1420 33160 1460 33200
rect 1132 29800 1172 29840
rect 1420 30640 1460 30680
rect 1420 30220 1460 30260
rect 1036 29044 1076 29084
rect 1612 36856 1652 36896
rect 1708 33664 1748 33704
rect 1708 30892 1748 30932
rect 1708 30220 1748 30260
rect 1996 39040 2036 39080
rect 1996 38872 2036 38912
rect 1996 38620 2036 38660
rect 1900 37444 1940 37484
rect 2092 36352 2132 36392
rect 2284 38200 2324 38240
rect 3052 48700 3092 48740
rect 3148 48280 3188 48320
rect 3052 47272 3092 47312
rect 3052 44752 3092 44792
rect 3244 48112 3284 48152
rect 4108 50800 4148 50840
rect 4012 50044 4052 50084
rect 3688 49876 3728 49916
rect 3770 49876 3810 49916
rect 3852 49876 3892 49916
rect 3934 49876 3974 49916
rect 4016 49876 4056 49916
rect 3436 49036 3476 49076
rect 3436 47776 3476 47816
rect 3340 47272 3380 47312
rect 3148 43576 3188 43616
rect 2860 43492 2900 43532
rect 4300 51220 4340 51260
rect 4684 56512 4724 56552
rect 4928 59704 4968 59744
rect 5010 59704 5050 59744
rect 5092 59704 5132 59744
rect 5174 59704 5214 59744
rect 5256 59704 5296 59744
rect 5452 59368 5492 59408
rect 5356 59200 5396 59240
rect 4972 58696 5012 58736
rect 5356 58612 5396 58652
rect 5164 58360 5204 58400
rect 4928 58192 4968 58232
rect 5010 58192 5050 58232
rect 5092 58192 5132 58232
rect 5174 58192 5214 58232
rect 5256 58192 5296 58232
rect 5068 57940 5108 57980
rect 5548 58360 5588 58400
rect 5452 57016 5492 57056
rect 5836 60544 5876 60584
rect 5740 60208 5780 60248
rect 5740 57016 5780 57056
rect 4928 56680 4968 56720
rect 5010 56680 5050 56720
rect 5092 56680 5132 56720
rect 5174 56680 5214 56720
rect 5256 56680 5296 56720
rect 4684 55672 4724 55712
rect 5260 55672 5300 55712
rect 4684 55420 4724 55460
rect 4588 51388 4628 51428
rect 4588 51220 4628 51260
rect 4928 55168 4968 55208
rect 5010 55168 5050 55208
rect 5092 55168 5132 55208
rect 5174 55168 5214 55208
rect 5256 55168 5296 55208
rect 5068 55000 5108 55040
rect 4780 54328 4820 54368
rect 5356 54832 5396 54872
rect 5740 56512 5780 56552
rect 5644 56260 5684 56300
rect 5740 56092 5780 56132
rect 4928 53656 4968 53696
rect 5010 53656 5050 53696
rect 5092 53656 5132 53696
rect 5174 53656 5214 53696
rect 5256 53656 5296 53696
rect 4780 53320 4820 53360
rect 5068 53236 5108 53276
rect 4780 52984 4820 53024
rect 5932 53908 5972 53948
rect 5548 53824 5588 53864
rect 5836 52984 5876 53024
rect 5548 52900 5588 52940
rect 5548 52480 5588 52520
rect 4928 52144 4968 52184
rect 5010 52144 5050 52184
rect 5092 52144 5132 52184
rect 5174 52144 5214 52184
rect 5256 52144 5296 52184
rect 4972 51388 5012 51428
rect 4780 50968 4820 51008
rect 4780 50800 4820 50840
rect 4928 50632 4968 50672
rect 5010 50632 5050 50672
rect 5092 50632 5132 50672
rect 5174 50632 5214 50672
rect 5256 50632 5296 50672
rect 4300 50296 4340 50336
rect 4300 50044 4340 50084
rect 3916 49372 3956 49412
rect 4204 49372 4244 49412
rect 3688 48364 3728 48404
rect 3770 48364 3810 48404
rect 3852 48364 3892 48404
rect 3934 48364 3974 48404
rect 4016 48364 4056 48404
rect 3628 48112 3668 48152
rect 3628 47944 3668 47984
rect 3820 47776 3860 47816
rect 4012 47188 4052 47228
rect 3688 46852 3728 46892
rect 3770 46852 3810 46892
rect 3852 46852 3892 46892
rect 3934 46852 3974 46892
rect 4016 46852 4056 46892
rect 4012 46264 4052 46304
rect 3916 45592 3956 45632
rect 4108 45844 4148 45884
rect 3688 45340 3728 45380
rect 3770 45340 3810 45380
rect 3852 45340 3892 45380
rect 3934 45340 3974 45380
rect 4016 45340 4056 45380
rect 3628 44920 3668 44960
rect 4012 44920 4052 44960
rect 3532 44836 3572 44876
rect 3820 44668 3860 44708
rect 3628 44248 3668 44288
rect 3436 43492 3476 43532
rect 3244 42904 3284 42944
rect 2956 42736 2996 42776
rect 4492 50044 4532 50084
rect 4492 49372 4532 49412
rect 4396 49036 4436 49076
rect 4684 50380 4724 50420
rect 5452 50548 5492 50588
rect 4876 50044 4916 50084
rect 5356 49456 5396 49496
rect 4588 49288 4628 49328
rect 4928 49120 4968 49160
rect 5010 49120 5050 49160
rect 5092 49120 5132 49160
rect 5174 49120 5214 49160
rect 5256 49120 5296 49160
rect 5356 49036 5396 49076
rect 5068 48784 5108 48824
rect 4876 48280 4916 48320
rect 5260 48700 5300 48740
rect 5068 48112 5108 48152
rect 5068 47860 5108 47900
rect 6604 65164 6644 65204
rect 6316 62392 6356 62432
rect 6124 57940 6164 57980
rect 6508 61552 6548 61592
rect 6796 65080 6836 65120
rect 6700 64660 6740 64700
rect 6796 64408 6836 64448
rect 6796 64072 6836 64112
rect 6700 63148 6740 63188
rect 6700 61552 6740 61592
rect 6700 61300 6740 61340
rect 6604 61048 6644 61088
rect 6412 60376 6452 60416
rect 7372 67516 7412 67556
rect 7180 66844 7220 66884
rect 7180 65752 7220 65792
rect 6988 65248 7028 65288
rect 7276 65416 7316 65456
rect 7180 65332 7220 65372
rect 7180 64492 7220 64532
rect 7180 64072 7220 64112
rect 7084 63904 7124 63944
rect 7084 63736 7124 63776
rect 6988 63652 7028 63692
rect 6892 62560 6932 62600
rect 6892 62392 6932 62432
rect 6796 61132 6836 61172
rect 6796 60880 6836 60920
rect 6700 60712 6740 60752
rect 6604 60292 6644 60332
rect 6316 58108 6356 58148
rect 6316 57856 6356 57896
rect 6316 57604 6356 57644
rect 6220 56092 6260 56132
rect 6604 58780 6644 58820
rect 7180 63148 7220 63188
rect 7084 62644 7124 62684
rect 7372 64408 7412 64448
rect 7372 63904 7412 63944
rect 8236 76000 8276 76040
rect 8044 74488 8084 74528
rect 8236 74320 8276 74360
rect 8428 76504 8468 76544
rect 8044 73312 8084 73352
rect 7948 72304 7988 72344
rect 8812 78184 8852 78224
rect 8716 77428 8756 77468
rect 8620 76504 8660 76544
rect 8524 76000 8564 76040
rect 8812 76840 8852 76880
rect 8620 75916 8660 75956
rect 9004 77428 9044 77468
rect 8908 76672 8948 76712
rect 8908 75916 8948 75956
rect 8812 75748 8852 75788
rect 8716 74656 8756 74696
rect 8620 74572 8660 74612
rect 9292 82216 9332 82256
rect 9580 85744 9620 85784
rect 9964 85828 10004 85868
rect 9868 84484 9908 84524
rect 9676 84400 9716 84440
rect 9772 83476 9812 83516
rect 9196 80620 9236 80660
rect 9196 79024 9236 79064
rect 9484 81796 9524 81836
rect 9292 77932 9332 77972
rect 10636 85240 10676 85280
rect 10252 84400 10292 84440
rect 10444 84400 10484 84440
rect 10444 84064 10484 84104
rect 10636 83476 10676 83516
rect 10252 83140 10292 83180
rect 10828 80368 10868 80408
rect 10156 79780 10196 79820
rect 9676 79360 9716 79400
rect 9484 78184 9524 78224
rect 9484 76840 9524 76880
rect 10156 79024 10196 79064
rect 10540 79024 10580 79064
rect 9964 78772 10004 78812
rect 10348 78772 10388 78812
rect 9868 76588 9908 76628
rect 9100 75664 9140 75704
rect 9196 75580 9236 75620
rect 9100 75496 9140 75536
rect 9100 75076 9140 75116
rect 8716 74320 8756 74360
rect 8524 73732 8564 73772
rect 8908 74320 8948 74360
rect 8812 74236 8852 74276
rect 8716 73060 8756 73100
rect 8812 72892 8852 72932
rect 8716 72472 8756 72512
rect 8332 72304 8372 72344
rect 8044 71968 8084 72008
rect 7948 71464 7988 71504
rect 7660 70120 7700 70160
rect 7852 70120 7892 70160
rect 7756 69196 7796 69236
rect 7660 66088 7700 66128
rect 7660 65752 7700 65792
rect 7564 65416 7604 65456
rect 7852 68272 7892 68312
rect 8140 71800 8180 71840
rect 8236 70120 8276 70160
rect 8236 69784 8276 69824
rect 8044 69700 8084 69740
rect 7756 65164 7796 65204
rect 8428 71968 8468 72008
rect 8620 71968 8660 72008
rect 8524 71800 8564 71840
rect 8812 72136 8852 72176
rect 9100 74320 9140 74360
rect 9292 74320 9332 74360
rect 9196 74236 9236 74276
rect 9676 76084 9716 76124
rect 11308 83728 11348 83768
rect 11020 78436 11060 78476
rect 10348 75832 10388 75872
rect 10156 74824 10196 74864
rect 9484 73816 9524 73856
rect 9868 74572 9908 74612
rect 9676 74488 9716 74528
rect 9964 74320 10004 74360
rect 10348 74656 10388 74696
rect 10252 74572 10292 74612
rect 10540 75076 10580 75116
rect 10060 74236 10100 74276
rect 9580 73732 9620 73772
rect 9388 73648 9428 73688
rect 9676 73480 9716 73520
rect 10252 73900 10292 73940
rect 10060 73732 10100 73772
rect 10156 73648 10196 73688
rect 10348 73648 10388 73688
rect 10060 73480 10100 73520
rect 9484 73312 9524 73352
rect 9100 72892 9140 72932
rect 9196 72808 9236 72848
rect 9004 72304 9044 72344
rect 8620 70624 8660 70664
rect 10252 73144 10292 73184
rect 10540 73648 10580 73688
rect 10828 75580 10868 75620
rect 11020 76084 11060 76124
rect 10924 75160 10964 75200
rect 10828 75076 10868 75116
rect 10732 74320 10772 74360
rect 10828 73900 10868 73940
rect 10732 73144 10772 73184
rect 11020 73312 11060 73352
rect 11308 78520 11348 78560
rect 11212 76756 11252 76796
rect 11212 76000 11252 76040
rect 11500 83476 11540 83516
rect 11788 84400 11828 84440
rect 11596 82468 11636 82508
rect 12076 85240 12116 85280
rect 11596 80620 11636 80660
rect 11404 76756 11444 76796
rect 10732 72724 10772 72764
rect 10924 72724 10964 72764
rect 10828 72640 10868 72680
rect 9292 72556 9332 72596
rect 9196 72304 9236 72344
rect 9388 72304 9428 72344
rect 9868 72304 9908 72344
rect 8524 69532 8564 69572
rect 8140 68692 8180 68732
rect 8140 68524 8180 68564
rect 8044 67096 8084 67136
rect 8044 66844 8084 66884
rect 8716 68020 8756 68060
rect 9004 71464 9044 71504
rect 9484 72220 9524 72260
rect 9292 72052 9332 72092
rect 9196 71968 9236 72008
rect 9196 71800 9236 71840
rect 9100 70960 9140 71000
rect 9004 70624 9044 70664
rect 8908 67432 8948 67472
rect 8620 67096 8660 67136
rect 8908 67012 8948 67052
rect 8332 66676 8372 66716
rect 8236 66592 8276 66632
rect 8140 66172 8180 66212
rect 8044 65584 8084 65624
rect 7948 65080 7988 65120
rect 7948 64240 7988 64280
rect 7468 63652 7508 63692
rect 7756 63904 7796 63944
rect 7660 63400 7700 63440
rect 8236 65416 8276 65456
rect 8332 64072 8372 64112
rect 7948 63568 7988 63608
rect 7852 63400 7892 63440
rect 7372 63064 7412 63104
rect 7660 63064 7700 63104
rect 7756 62980 7796 63020
rect 7660 62812 7700 62852
rect 7276 62392 7316 62432
rect 7468 62392 7508 62432
rect 6988 61636 7028 61676
rect 7564 61468 7604 61508
rect 6892 60124 6932 60164
rect 7180 60880 7220 60920
rect 7084 60040 7124 60080
rect 6796 59536 6836 59576
rect 6988 59368 7028 59408
rect 7276 60040 7316 60080
rect 7276 59872 7316 59912
rect 7180 58780 7220 58820
rect 6700 58444 6740 58484
rect 7084 58444 7124 58484
rect 6604 57940 6644 57980
rect 6700 57016 6740 57056
rect 6988 57016 7028 57056
rect 6892 56848 6932 56888
rect 6892 55756 6932 55796
rect 7468 61132 7508 61172
rect 8140 63400 8180 63440
rect 8044 63316 8084 63356
rect 8428 63652 8468 63692
rect 8044 63064 8084 63104
rect 8332 63064 8372 63104
rect 7948 61888 7988 61928
rect 7948 61720 7988 61760
rect 7852 60964 7892 61004
rect 7852 60712 7892 60752
rect 7660 60376 7700 60416
rect 7468 60208 7508 60248
rect 7660 60124 7700 60164
rect 7372 58444 7412 58484
rect 7276 57016 7316 57056
rect 7564 57856 7604 57896
rect 7756 59200 7796 59240
rect 7852 57772 7892 57812
rect 7756 57100 7796 57140
rect 7564 57016 7604 57056
rect 7180 56428 7220 56468
rect 7468 56764 7508 56804
rect 6220 55084 6260 55124
rect 6220 54160 6260 54200
rect 6124 51220 6164 51260
rect 6412 53236 6452 53276
rect 6412 51976 6452 52016
rect 5932 50968 5972 51008
rect 5836 50212 5876 50252
rect 5836 49456 5876 49496
rect 5836 49036 5876 49076
rect 5548 48448 5588 48488
rect 5740 48448 5780 48488
rect 5356 48280 5396 48320
rect 6028 49960 6068 50000
rect 5932 48532 5972 48572
rect 5548 48280 5588 48320
rect 5356 48112 5396 48152
rect 4928 47608 4968 47648
rect 5010 47608 5050 47648
rect 5092 47608 5132 47648
rect 5174 47608 5214 47648
rect 5256 47608 5296 47648
rect 5452 47949 5492 47984
rect 5452 47944 5492 47949
rect 4300 44668 4340 44708
rect 4012 43996 4052 44036
rect 4928 46096 4968 46136
rect 5010 46096 5050 46136
rect 5092 46096 5132 46136
rect 5174 46096 5214 46136
rect 5256 46096 5296 46136
rect 5452 47272 5492 47312
rect 5644 47608 5684 47648
rect 4588 44920 4628 44960
rect 5356 45760 5396 45800
rect 5932 48196 5972 48236
rect 6412 50800 6452 50840
rect 6220 50548 6260 50588
rect 6124 48196 6164 48236
rect 3688 43828 3728 43868
rect 3770 43828 3810 43868
rect 3852 43828 3892 43868
rect 3934 43828 3974 43868
rect 4016 43828 4056 43868
rect 3724 43576 3764 43616
rect 3628 43492 3668 43532
rect 4108 43492 4148 43532
rect 3532 42904 3572 42944
rect 3688 42316 3728 42356
rect 3770 42316 3810 42356
rect 3852 42316 3892 42356
rect 3934 42316 3974 42356
rect 4016 42316 4056 42356
rect 4012 41896 4052 41936
rect 3532 41812 3572 41852
rect 3916 41812 3956 41852
rect 4204 42820 4244 42860
rect 4108 41812 4148 41852
rect 3532 41560 3572 41600
rect 3340 41476 3380 41516
rect 2956 40972 2996 41012
rect 2860 40552 2900 40592
rect 2860 40048 2900 40088
rect 2764 39544 2804 39584
rect 2668 39040 2708 39080
rect 2572 37864 2612 37904
rect 2284 36604 2324 36644
rect 2572 37360 2612 37400
rect 2476 36940 2516 36980
rect 2476 36604 2516 36644
rect 2380 36184 2420 36224
rect 2188 36100 2228 36140
rect 1900 35848 1940 35888
rect 1996 35008 2036 35048
rect 2380 34840 2420 34880
rect 1996 34420 2036 34460
rect 2188 34336 2228 34376
rect 2188 33580 2228 33620
rect 2188 33076 2228 33116
rect 2092 32824 2132 32864
rect 1996 31312 2036 31352
rect 1900 30808 1940 30848
rect 2092 30808 2132 30848
rect 2668 36184 2708 36224
rect 2668 35848 2708 35888
rect 2572 35764 2612 35804
rect 2668 34504 2708 34544
rect 4928 44584 4968 44624
rect 5010 44584 5050 44624
rect 5092 44584 5132 44624
rect 5174 44584 5214 44624
rect 5256 44584 5296 44624
rect 5068 44164 5108 44204
rect 5260 44080 5300 44120
rect 4780 43492 4820 43532
rect 4928 43072 4968 43112
rect 5010 43072 5050 43112
rect 5092 43072 5132 43112
rect 5174 43072 5214 43112
rect 5256 43072 5296 43112
rect 5068 42736 5108 42776
rect 4876 42652 4916 42692
rect 5644 45340 5684 45380
rect 5932 46600 5972 46640
rect 6604 55168 6644 55208
rect 6508 50296 6548 50336
rect 7660 56344 7700 56384
rect 8044 60712 8084 60752
rect 8044 57856 8084 57896
rect 8716 66592 8756 66632
rect 8716 66256 8756 66296
rect 8620 65500 8660 65540
rect 8620 64660 8660 64700
rect 8620 63652 8660 63692
rect 8524 63400 8564 63440
rect 8908 66844 8948 66884
rect 8812 65920 8852 65960
rect 8908 65836 8948 65876
rect 9772 72136 9812 72176
rect 10828 72220 10868 72260
rect 9676 71968 9716 72008
rect 9580 71800 9620 71840
rect 9772 71716 9812 71756
rect 9580 71464 9620 71504
rect 9772 71464 9812 71504
rect 10348 72136 10388 72176
rect 10348 71968 10388 72008
rect 10444 71716 10484 71756
rect 10828 71548 10868 71588
rect 10636 71380 10676 71420
rect 10540 70792 10580 70832
rect 9868 70372 9908 70412
rect 9484 69952 9524 69992
rect 9868 69868 9908 69908
rect 9484 69196 9524 69236
rect 10060 69112 10100 69152
rect 9676 68944 9716 68984
rect 9484 68524 9524 68564
rect 9100 67852 9140 67892
rect 9100 67684 9140 67724
rect 9676 68356 9716 68396
rect 9676 68020 9716 68060
rect 10156 68944 10196 68984
rect 10636 69868 10676 69908
rect 10444 69280 10484 69320
rect 10540 69112 10580 69152
rect 10828 70624 10868 70664
rect 10732 69280 10772 69320
rect 10348 68608 10388 68648
rect 9772 67852 9812 67892
rect 10060 67852 10100 67892
rect 10156 67684 10196 67724
rect 9772 67516 9812 67556
rect 10060 67516 10100 67556
rect 9676 67432 9716 67472
rect 9196 67096 9236 67136
rect 9388 67012 9428 67052
rect 9868 67012 9908 67052
rect 8908 65500 8948 65540
rect 9388 66256 9428 66296
rect 9868 66844 9908 66884
rect 9772 66760 9812 66800
rect 9484 65920 9524 65960
rect 9196 65248 9236 65288
rect 9964 66256 10004 66296
rect 9676 66004 9716 66044
rect 9676 65836 9716 65876
rect 9580 64912 9620 64952
rect 9580 64492 9620 64532
rect 9004 64324 9044 64364
rect 8812 63904 8852 63944
rect 8812 63568 8852 63608
rect 8812 63148 8852 63188
rect 8716 63064 8756 63104
rect 10252 67180 10292 67220
rect 10252 66340 10292 66380
rect 10156 65920 10196 65960
rect 10060 64996 10100 65036
rect 9196 64240 9236 64280
rect 9292 63652 9332 63692
rect 9004 62392 9044 62432
rect 9196 62560 9236 62600
rect 8428 61804 8468 61844
rect 9100 62308 9140 62348
rect 8332 61552 8372 61592
rect 8716 61636 8756 61676
rect 8716 60964 8756 61004
rect 8620 60880 8660 60920
rect 8524 60544 8564 60584
rect 8428 60040 8468 60080
rect 8524 59872 8564 59912
rect 9004 61720 9044 61760
rect 8908 60964 8948 61004
rect 8812 60628 8852 60668
rect 8716 60376 8756 60416
rect 9388 63400 9428 63440
rect 9388 62560 9428 62600
rect 9964 64156 10004 64196
rect 9580 63736 9620 63776
rect 10060 64072 10100 64112
rect 11116 69952 11156 69992
rect 11116 69700 11156 69740
rect 11404 75580 11444 75620
rect 11308 75244 11348 75284
rect 11500 75496 11540 75536
rect 11404 74908 11444 74948
rect 11308 73312 11348 73352
rect 11308 71716 11348 71756
rect 11308 69112 11348 69152
rect 10732 68608 10772 68648
rect 10636 68356 10676 68396
rect 10540 64744 10580 64784
rect 10444 64576 10484 64616
rect 10348 64072 10388 64112
rect 10636 64072 10676 64112
rect 10252 63988 10292 64028
rect 10540 63988 10580 64028
rect 10060 63568 10100 63608
rect 10252 63316 10292 63356
rect 9964 63232 10004 63272
rect 9868 63148 9908 63188
rect 10060 63064 10100 63104
rect 11116 67096 11156 67136
rect 10828 65332 10868 65372
rect 11020 64828 11060 64868
rect 10924 64744 10964 64784
rect 11020 64576 11060 64616
rect 11116 64408 11156 64448
rect 10924 63988 10964 64028
rect 10828 63904 10868 63944
rect 10540 63568 10580 63608
rect 9964 62980 10004 63020
rect 10444 63064 10484 63104
rect 9676 62560 9716 62600
rect 9868 62560 9908 62600
rect 10348 62560 10388 62600
rect 9772 62392 9812 62432
rect 10156 62392 10196 62432
rect 10732 63400 10772 63440
rect 11020 63568 11060 63608
rect 10924 63232 10964 63272
rect 10924 63064 10964 63104
rect 11308 68524 11348 68564
rect 11788 75412 11828 75452
rect 11980 80536 12020 80576
rect 11788 74656 11828 74696
rect 11596 73648 11636 73688
rect 11596 73144 11636 73184
rect 11884 72976 11924 73016
rect 11884 72724 11924 72764
rect 11980 72052 12020 72092
rect 11596 70456 11636 70496
rect 11884 70120 11924 70160
rect 11692 69952 11732 69992
rect 11500 69117 11540 69152
rect 11500 69112 11540 69117
rect 11308 67432 11348 67472
rect 11500 66928 11540 66968
rect 11308 65248 11348 65288
rect 11308 64828 11348 64868
rect 11212 63484 11252 63524
rect 11212 63148 11252 63188
rect 10828 62980 10868 63020
rect 10732 62896 10772 62936
rect 9676 62308 9716 62348
rect 9580 61888 9620 61928
rect 9676 61552 9716 61592
rect 9484 61132 9524 61172
rect 9100 60964 9140 61004
rect 9292 60796 9332 60836
rect 9004 60376 9044 60416
rect 9292 60208 9332 60248
rect 8908 60124 8948 60164
rect 9100 59872 9140 59912
rect 9004 59788 9044 59828
rect 8913 59368 8953 59408
rect 8620 59200 8660 59240
rect 8524 57856 8564 57896
rect 8140 57688 8180 57728
rect 8044 57100 8084 57140
rect 7948 56680 7988 56720
rect 7948 56344 7988 56384
rect 9004 58612 9044 58652
rect 9004 58444 9044 58484
rect 8812 57688 8852 57728
rect 8236 57016 8276 57056
rect 6700 54160 6740 54200
rect 6700 53908 6740 53948
rect 6316 49288 6356 49328
rect 6316 48196 6356 48236
rect 6796 52564 6836 52604
rect 7084 53992 7124 54032
rect 6988 52480 7028 52520
rect 7564 54832 7604 54872
rect 7564 54076 7604 54116
rect 7564 53824 7604 53864
rect 7756 55084 7796 55124
rect 7372 52900 7412 52940
rect 7276 52732 7316 52772
rect 7180 52228 7220 52268
rect 7084 52060 7124 52100
rect 6892 51556 6932 51596
rect 7180 51976 7220 52016
rect 7372 52396 7412 52436
rect 7660 52480 7700 52520
rect 7468 52228 7508 52268
rect 7276 51892 7316 51932
rect 6796 50296 6836 50336
rect 6700 49456 6740 49496
rect 7084 49960 7124 50000
rect 7084 49288 7124 49328
rect 6796 49120 6836 49160
rect 6508 48196 6548 48236
rect 6700 48028 6740 48068
rect 6412 47272 6452 47312
rect 6892 48028 6932 48068
rect 6988 47860 7028 47900
rect 6316 45928 6356 45968
rect 5644 44332 5684 44372
rect 5548 44080 5588 44120
rect 6220 45424 6260 45464
rect 7084 46600 7124 46640
rect 7372 51556 7412 51596
rect 7276 50548 7316 50588
rect 7276 49120 7316 49160
rect 6700 45928 6740 45968
rect 5932 44836 5972 44876
rect 6220 44836 6260 44876
rect 6700 44752 6740 44792
rect 6220 43996 6260 44036
rect 5260 42568 5300 42608
rect 5164 42484 5204 42524
rect 5164 42316 5204 42356
rect 5452 42484 5492 42524
rect 4928 41560 4968 41600
rect 5010 41560 5050 41600
rect 5092 41560 5132 41600
rect 5174 41560 5214 41600
rect 5256 41560 5296 41600
rect 4300 41224 4340 41264
rect 4492 41224 4532 41264
rect 4876 41224 4916 41264
rect 5452 41224 5492 41264
rect 3628 40972 3668 41012
rect 3688 40804 3728 40844
rect 3770 40804 3810 40844
rect 3852 40804 3892 40844
rect 3934 40804 3974 40844
rect 4016 40804 4056 40844
rect 3148 40300 3188 40340
rect 3916 40468 3956 40508
rect 4108 40300 4148 40340
rect 3052 39880 3092 39920
rect 2956 39712 2996 39752
rect 3436 39712 3476 39752
rect 3340 39544 3380 39584
rect 3244 38872 3284 38912
rect 2860 38200 2900 38240
rect 3148 38200 3188 38240
rect 2860 37360 2900 37400
rect 2956 36856 2996 36896
rect 3148 37780 3188 37820
rect 2956 36520 2996 36560
rect 2860 35764 2900 35804
rect 2860 35260 2900 35300
rect 3052 35176 3092 35216
rect 2956 34924 2996 34964
rect 2668 34168 2708 34208
rect 2572 33748 2612 33788
rect 2476 33664 2516 33704
rect 4012 39712 4052 39752
rect 4108 39460 4148 39500
rect 3688 39292 3728 39332
rect 3770 39292 3810 39332
rect 3852 39292 3892 39332
rect 3934 39292 3974 39332
rect 4016 39292 4056 39332
rect 4876 40720 4916 40760
rect 5164 40720 5204 40760
rect 4396 40468 4436 40508
rect 4300 38452 4340 38492
rect 5164 40384 5204 40424
rect 5548 40384 5588 40424
rect 4928 40048 4968 40088
rect 5010 40048 5050 40088
rect 5092 40048 5132 40088
rect 5174 40048 5214 40088
rect 5256 40048 5296 40088
rect 5356 40048 5396 40088
rect 4588 39628 4628 39668
rect 4492 39376 4532 39416
rect 5260 38956 5300 38996
rect 4396 38284 4436 38324
rect 3724 38200 3764 38240
rect 3688 37780 3728 37820
rect 3770 37780 3810 37820
rect 3852 37780 3892 37820
rect 3934 37780 3974 37820
rect 4016 37780 4056 37820
rect 3532 37528 3572 37568
rect 3628 37360 3668 37400
rect 4108 37192 4148 37232
rect 4300 37276 4340 37316
rect 4300 37108 4340 37148
rect 4928 38536 4968 38576
rect 5010 38536 5050 38576
rect 5092 38536 5132 38576
rect 5174 38536 5214 38576
rect 5256 38536 5296 38576
rect 5164 38284 5204 38324
rect 5548 38200 5588 38240
rect 4780 38116 4820 38156
rect 4972 38116 5012 38156
rect 6700 42820 6740 42860
rect 6028 42736 6068 42776
rect 5740 42484 5780 42524
rect 6604 42400 6644 42440
rect 6028 42316 6068 42356
rect 5836 41140 5876 41180
rect 5932 40888 5972 40928
rect 5932 40552 5972 40592
rect 5740 40048 5780 40088
rect 5740 39880 5780 39920
rect 6412 41224 6452 41264
rect 6508 40720 6548 40760
rect 6604 40468 6644 40508
rect 7084 46264 7124 46304
rect 6988 45340 7028 45380
rect 7948 54832 7988 54872
rect 8524 57016 8564 57056
rect 8428 56680 8468 56720
rect 8332 54076 8372 54116
rect 7948 53992 7988 54032
rect 8524 55168 8564 55208
rect 8908 56932 8948 56972
rect 9292 59620 9332 59660
rect 9580 60796 9620 60836
rect 9772 60796 9812 60836
rect 9868 60376 9908 60416
rect 9196 57856 9236 57896
rect 9484 59368 9524 59408
rect 9868 59536 9908 59576
rect 9772 58276 9812 58316
rect 9292 56932 9332 56972
rect 9004 56428 9044 56468
rect 8044 52900 8084 52940
rect 8140 52564 8180 52604
rect 8716 53488 8756 53528
rect 7852 52480 7892 52520
rect 7756 51220 7796 51260
rect 7660 50632 7700 50672
rect 7564 50548 7604 50588
rect 7564 50296 7604 50336
rect 7372 49036 7412 49076
rect 7756 48952 7796 48992
rect 8620 53068 8660 53108
rect 8524 52228 8564 52268
rect 8044 51724 8084 51764
rect 8332 51640 8372 51680
rect 7948 49036 7988 49076
rect 8140 50968 8180 51008
rect 8140 48280 8180 48320
rect 8140 48112 8180 48152
rect 8236 47944 8276 47984
rect 7468 46516 7508 46556
rect 7372 46180 7412 46220
rect 7276 45844 7316 45884
rect 7180 45508 7220 45548
rect 7276 45340 7316 45380
rect 7372 45172 7412 45212
rect 7276 45004 7316 45044
rect 7564 46264 7604 46304
rect 7564 45760 7604 45800
rect 7756 45508 7796 45548
rect 7948 45004 7988 45044
rect 7564 44920 7604 44960
rect 7468 44164 7508 44204
rect 7468 43492 7508 43532
rect 8140 46432 8180 46472
rect 6988 42820 7028 42860
rect 6988 40468 7028 40508
rect 6796 40132 6836 40172
rect 6220 39712 6260 39752
rect 6124 39628 6164 39668
rect 6700 39712 6740 39752
rect 6508 39544 6548 39584
rect 6028 38956 6068 38996
rect 5932 38872 5972 38912
rect 6124 38200 6164 38240
rect 4928 37024 4968 37064
rect 5010 37024 5050 37064
rect 5092 37024 5132 37064
rect 5174 37024 5214 37064
rect 5256 37024 5296 37064
rect 4108 36604 4148 36644
rect 3628 36520 3668 36560
rect 3688 36268 3728 36308
rect 3770 36268 3810 36308
rect 3852 36268 3892 36308
rect 3934 36268 3974 36308
rect 4016 36268 4056 36308
rect 3244 36016 3284 36056
rect 4108 35848 4148 35888
rect 4108 35260 4148 35300
rect 3820 35092 3860 35132
rect 3724 35008 3764 35048
rect 3244 34924 3284 34964
rect 3532 34924 3572 34964
rect 4108 34924 4148 34964
rect 2956 34252 2996 34292
rect 2860 33832 2900 33872
rect 2956 33664 2996 33704
rect 2764 32824 2804 32864
rect 2284 32656 2324 32696
rect 2860 32740 2900 32780
rect 2476 31816 2516 31856
rect 2380 31396 2420 31436
rect 1996 30556 2036 30596
rect 2188 30640 2228 30680
rect 2092 30472 2132 30512
rect 1900 29128 1940 29168
rect 2188 30136 2228 30176
rect 2092 29716 2132 29756
rect 2092 29212 2132 29252
rect 1996 28624 2036 28664
rect 1708 28288 1748 28328
rect 1324 28204 1364 28244
rect 1324 27700 1364 27740
rect 1132 26608 1172 26648
rect 1036 26020 1076 26060
rect 1036 23416 1076 23456
rect 940 2836 980 2876
rect 1036 1240 1076 1280
rect 1516 26104 1556 26144
rect 1516 25684 1556 25724
rect 1324 24928 1364 24968
rect 1324 24508 1364 24548
rect 1420 23752 1460 23792
rect 1324 23668 1364 23708
rect 1420 22828 1460 22868
rect 1324 20476 1364 20516
rect 1324 19720 1364 19760
rect 1516 20728 1556 20768
rect 1804 27448 1844 27488
rect 1804 24928 1844 24968
rect 1804 24760 1844 24800
rect 1708 24088 1748 24128
rect 1708 23500 1748 23540
rect 1708 22156 1748 22196
rect 1708 21568 1748 21608
rect 1612 19888 1652 19928
rect 1708 19804 1748 19844
rect 1996 25600 2036 25640
rect 2476 31060 2516 31100
rect 2476 30472 2516 30512
rect 2668 31480 2708 31520
rect 2860 31480 2900 31520
rect 3244 34168 3284 34208
rect 3148 33916 3188 33956
rect 3436 33748 3476 33788
rect 3340 33664 3380 33704
rect 3052 32740 3092 32780
rect 3340 32824 3380 32864
rect 3244 32656 3284 32696
rect 3688 34756 3728 34796
rect 3770 34756 3810 34796
rect 3852 34756 3892 34796
rect 3934 34756 3974 34796
rect 4016 34756 4056 34796
rect 3820 34336 3860 34376
rect 4300 35176 4340 35216
rect 4204 34336 4244 34376
rect 3724 33916 3764 33956
rect 3916 34252 3956 34292
rect 4204 33496 4244 33536
rect 3688 33244 3728 33284
rect 3770 33244 3810 33284
rect 3852 33244 3892 33284
rect 3934 33244 3974 33284
rect 4016 33244 4056 33284
rect 4204 32992 4244 33032
rect 3532 32740 3572 32780
rect 3724 32740 3764 32780
rect 3244 31984 3284 32024
rect 3052 31480 3092 31520
rect 3436 31480 3476 31520
rect 2860 31312 2900 31352
rect 3052 31312 3092 31352
rect 2956 31144 2996 31184
rect 3340 30976 3380 31016
rect 3244 30892 3284 30932
rect 2764 30724 2804 30764
rect 3148 30724 3188 30764
rect 2284 28960 2324 29000
rect 2284 27700 2324 27740
rect 2188 26104 2228 26144
rect 2188 25852 2228 25892
rect 2188 25432 2228 25472
rect 2476 28960 2516 29000
rect 2668 29128 2708 29168
rect 2668 28960 2708 29000
rect 2572 27784 2612 27824
rect 2476 27364 2516 27404
rect 2476 26776 2516 26816
rect 2380 25768 2420 25808
rect 2476 25516 2516 25556
rect 2380 25264 2420 25304
rect 2476 25012 2516 25052
rect 3052 30640 3092 30680
rect 2956 30556 2996 30596
rect 2860 30388 2900 30428
rect 2956 29800 2996 29840
rect 2956 29548 2996 29588
rect 2956 29044 2996 29084
rect 2860 27784 2900 27824
rect 2860 27448 2900 27488
rect 2764 27364 2804 27404
rect 3340 30472 3380 30512
rect 3436 29632 3476 29672
rect 3436 29044 3476 29084
rect 3148 28876 3188 28916
rect 3244 28372 3284 28412
rect 3436 28120 3476 28160
rect 2956 26440 2996 26480
rect 2860 26104 2900 26144
rect 2764 25516 2804 25556
rect 2860 25348 2900 25388
rect 3148 26692 3188 26732
rect 3148 26188 3188 26228
rect 3436 26440 3476 26480
rect 5164 36772 5204 36812
rect 4684 35848 4724 35888
rect 4588 35596 4628 35636
rect 4492 35344 4532 35384
rect 4492 35008 4532 35048
rect 4396 34336 4436 34376
rect 4396 34168 4436 34208
rect 4396 32740 4436 32780
rect 4396 32320 4436 32360
rect 4204 31984 4244 32024
rect 3724 31900 3764 31940
rect 3688 31732 3728 31772
rect 3770 31732 3810 31772
rect 3852 31732 3892 31772
rect 3934 31732 3974 31772
rect 4016 31732 4056 31772
rect 3724 31396 3764 31436
rect 4300 31732 4340 31772
rect 3628 31060 3668 31100
rect 3916 31144 3956 31184
rect 3724 30976 3764 31016
rect 3820 30808 3860 30848
rect 3628 30472 3668 30512
rect 3688 30220 3728 30260
rect 3770 30220 3810 30260
rect 3852 30220 3892 30260
rect 3934 30220 3974 30260
rect 4016 30220 4056 30260
rect 4204 30640 4244 30680
rect 3628 29800 3668 29840
rect 4204 29800 4244 29840
rect 3628 29128 3668 29168
rect 4204 29128 4244 29168
rect 4012 28876 4052 28916
rect 3688 28708 3728 28748
rect 3770 28708 3810 28748
rect 3852 28708 3892 28748
rect 3934 28708 3974 28748
rect 4016 28708 4056 28748
rect 3628 28456 3668 28496
rect 4108 28456 4148 28496
rect 3724 28120 3764 28160
rect 4108 28288 4148 28328
rect 4588 34840 4628 34880
rect 4972 35848 5012 35888
rect 4928 35512 4968 35552
rect 5010 35512 5050 35552
rect 5092 35512 5132 35552
rect 5174 35512 5214 35552
rect 5256 35512 5296 35552
rect 5164 35344 5204 35384
rect 4780 35008 4820 35048
rect 4684 33328 4724 33368
rect 4492 31984 4532 32024
rect 5068 34336 5108 34376
rect 5260 34672 5300 34712
rect 5068 34168 5108 34208
rect 4928 34000 4968 34040
rect 5010 34000 5050 34040
rect 5092 34000 5132 34040
rect 5174 34000 5214 34040
rect 5256 34000 5296 34040
rect 4928 32488 4968 32528
rect 5010 32488 5050 32528
rect 5092 32488 5132 32528
rect 5174 32488 5214 32528
rect 5256 32488 5296 32528
rect 5452 37444 5492 37484
rect 5548 36604 5588 36644
rect 5452 35344 5492 35384
rect 5452 35176 5492 35216
rect 6028 38116 6068 38156
rect 5836 37444 5876 37484
rect 5836 35932 5876 35972
rect 5836 35260 5876 35300
rect 6028 35260 6068 35300
rect 5740 35176 5780 35216
rect 5548 34336 5588 34376
rect 5644 33916 5684 33956
rect 5644 33748 5684 33788
rect 5548 32404 5588 32444
rect 5068 31480 5108 31520
rect 5356 31480 5396 31520
rect 4780 31396 4820 31436
rect 4492 30808 4532 30848
rect 4684 31144 4724 31184
rect 5356 31312 5396 31352
rect 4588 30724 4628 30764
rect 4588 30388 4628 30428
rect 4396 30052 4436 30092
rect 4300 28120 4340 28160
rect 4108 28036 4148 28076
rect 3820 27700 3860 27740
rect 4012 27700 4052 27740
rect 4108 27448 4148 27488
rect 3688 27196 3728 27236
rect 3770 27196 3810 27236
rect 3852 27196 3892 27236
rect 3934 27196 3974 27236
rect 4016 27196 4056 27236
rect 4300 27448 4340 27488
rect 4204 27280 4244 27320
rect 4204 26944 4244 26984
rect 3724 26776 3764 26816
rect 3724 26608 3764 26648
rect 3244 26104 3284 26144
rect 3148 25516 3188 25556
rect 3148 25264 3188 25304
rect 2668 25012 2708 25052
rect 2476 24424 2516 24464
rect 2284 23752 2324 23792
rect 2188 23668 2228 23708
rect 1996 23332 2036 23372
rect 2092 22912 2132 22952
rect 2284 22912 2324 22952
rect 1996 22828 2036 22868
rect 1900 22576 1940 22616
rect 2092 21568 2132 21608
rect 2092 21400 2132 21440
rect 2668 23920 2708 23960
rect 2572 23836 2612 23876
rect 2476 23752 2516 23792
rect 2476 23332 2516 23372
rect 2668 22996 2708 23036
rect 2572 22744 2612 22784
rect 2476 22240 2516 22280
rect 3148 24508 3188 24548
rect 3052 24424 3092 24464
rect 2860 23752 2900 23792
rect 3244 24340 3284 24380
rect 3340 24256 3380 24296
rect 3532 26104 3572 26144
rect 4684 29296 4724 29336
rect 4972 31144 5012 31184
rect 4928 30976 4968 31016
rect 5010 30976 5050 31016
rect 5092 30976 5132 31016
rect 5174 30976 5214 31016
rect 5256 30976 5296 31016
rect 5068 30808 5108 30848
rect 5068 30304 5108 30344
rect 5548 31312 5588 31352
rect 5452 30220 5492 30260
rect 5644 30052 5684 30092
rect 5548 29800 5588 29840
rect 5356 29716 5396 29756
rect 4928 29464 4968 29504
rect 5010 29464 5050 29504
rect 5092 29464 5132 29504
rect 5174 29464 5214 29504
rect 5256 29464 5296 29504
rect 5356 29128 5396 29168
rect 4780 28708 4820 28748
rect 5452 28540 5492 28580
rect 5356 28204 5396 28244
rect 5548 28456 5588 28496
rect 4684 28036 4724 28076
rect 4928 27952 4968 27992
rect 5010 27952 5050 27992
rect 5092 27952 5132 27992
rect 5174 27952 5214 27992
rect 5256 27952 5296 27992
rect 4780 27616 4820 27656
rect 5260 27616 5300 27656
rect 5452 27616 5492 27656
rect 4780 27280 4820 27320
rect 4492 26776 4532 26816
rect 4396 26440 4436 26480
rect 3532 25852 3572 25892
rect 3688 25684 3728 25724
rect 3770 25684 3810 25724
rect 3852 25684 3892 25724
rect 3934 25684 3974 25724
rect 4016 25684 4056 25724
rect 3820 25264 3860 25304
rect 3688 24172 3728 24212
rect 3770 24172 3810 24212
rect 3852 24172 3892 24212
rect 3934 24172 3974 24212
rect 4016 24172 4056 24212
rect 3820 24004 3860 24044
rect 3532 23920 3572 23960
rect 3148 23752 3188 23792
rect 3052 22240 3092 22280
rect 2956 21904 2996 21944
rect 2764 21652 2804 21692
rect 3148 21736 3188 21776
rect 3532 23668 3572 23708
rect 4204 25684 4244 25724
rect 4204 25264 4244 25304
rect 4300 25180 4340 25220
rect 4204 24844 4244 24884
rect 4492 26104 4532 26144
rect 4204 24676 4244 24716
rect 4396 24508 4436 24548
rect 4396 24088 4436 24128
rect 4300 23920 4340 23960
rect 4108 23416 4148 23456
rect 3436 22912 3476 22952
rect 2860 21400 2900 21440
rect 2764 21064 2804 21104
rect 1804 19720 1844 19760
rect 1804 18544 1844 18584
rect 1324 17956 1364 17996
rect 1516 17704 1556 17744
rect 1612 17116 1652 17156
rect 1420 17032 1460 17072
rect 1804 17452 1844 17492
rect 1228 16780 1268 16820
rect 1516 15856 1556 15896
rect 1324 15184 1364 15224
rect 1612 15604 1652 15644
rect 2476 19804 2516 19844
rect 2668 20728 2708 20768
rect 2572 19384 2612 19424
rect 2572 18712 2612 18752
rect 2956 20896 2996 20936
rect 2956 20308 2996 20348
rect 2764 19468 2804 19508
rect 3052 19468 3092 19508
rect 2956 19384 2996 19424
rect 3340 20980 3380 21020
rect 3148 18880 3188 18920
rect 2668 17620 2708 17660
rect 1900 16444 1940 16484
rect 2284 16444 2324 16484
rect 1708 15520 1748 15560
rect 1612 15184 1652 15224
rect 2572 17116 2612 17156
rect 2956 18040 2996 18080
rect 2860 17620 2900 17660
rect 3052 17620 3092 17660
rect 2956 17452 2996 17492
rect 2860 17284 2900 17324
rect 2956 17116 2996 17156
rect 2860 17032 2900 17072
rect 4012 23080 4052 23120
rect 3916 22996 3956 23036
rect 3688 22660 3728 22700
rect 3770 22660 3810 22700
rect 3852 22660 3892 22700
rect 3934 22660 3974 22700
rect 4016 22660 4056 22700
rect 3532 22324 3572 22364
rect 4108 21904 4148 21944
rect 3532 21736 3572 21776
rect 3724 21652 3764 21692
rect 3436 20896 3476 20936
rect 4204 21568 4244 21608
rect 3688 21148 3728 21188
rect 3770 21148 3810 21188
rect 3852 21148 3892 21188
rect 3934 21148 3974 21188
rect 4016 21148 4056 21188
rect 3724 20896 3764 20936
rect 3532 20812 3572 20852
rect 3436 20728 3476 20768
rect 3916 20812 3956 20852
rect 4684 26776 4724 26816
rect 5260 26692 5300 26732
rect 5644 27700 5684 27740
rect 5932 34672 5972 34712
rect 6897 39712 6937 39752
rect 6796 39040 6836 39080
rect 6892 38956 6932 38996
rect 6508 38788 6548 38828
rect 6700 37864 6740 37904
rect 6700 37444 6740 37484
rect 6220 36520 6260 36560
rect 6220 35176 6260 35216
rect 6124 34336 6164 34376
rect 6028 34252 6068 34292
rect 5932 33916 5972 33956
rect 6604 37360 6644 37400
rect 6604 35848 6644 35888
rect 6508 35344 6548 35384
rect 6604 35260 6644 35300
rect 6412 34588 6452 34628
rect 6316 34336 6356 34376
rect 6316 34168 6356 34208
rect 6220 34000 6260 34040
rect 6220 33832 6260 33872
rect 6124 33664 6164 33704
rect 6988 38284 7028 38324
rect 6988 38032 7028 38072
rect 6892 35848 6932 35888
rect 6892 35344 6932 35384
rect 7276 41056 7316 41096
rect 7180 40720 7220 40760
rect 7180 40384 7220 40424
rect 7180 40132 7220 40172
rect 8140 42736 8180 42776
rect 7564 41644 7604 41684
rect 7660 40552 7700 40592
rect 7276 38956 7316 38996
rect 7180 38536 7220 38576
rect 7276 38032 7316 38072
rect 7564 39712 7604 39752
rect 7756 40384 7796 40424
rect 7468 39544 7508 39584
rect 7660 38956 7700 38996
rect 8140 39712 8180 39752
rect 7948 39376 7988 39416
rect 8044 39040 8084 39080
rect 7948 37864 7988 37904
rect 7276 37528 7316 37568
rect 7083 37444 7123 37484
rect 7180 37024 7220 37064
rect 7084 36604 7124 36644
rect 6988 35176 7028 35216
rect 6796 35092 6836 35132
rect 6892 34756 6932 34796
rect 6700 34672 6740 34712
rect 6796 34252 6836 34292
rect 6604 34168 6644 34208
rect 6508 34000 6548 34040
rect 6604 33664 6644 33704
rect 6028 33580 6068 33620
rect 6124 33160 6164 33200
rect 5836 32404 5876 32444
rect 5932 32236 5972 32276
rect 5932 31732 5972 31772
rect 5836 30892 5876 30932
rect 5836 30724 5876 30764
rect 5836 30472 5876 30512
rect 5836 29464 5876 29504
rect 6220 32572 6260 32612
rect 6508 32404 6548 32444
rect 6412 32068 6452 32108
rect 6316 31564 6356 31604
rect 6124 30640 6164 30680
rect 6124 29800 6164 29840
rect 5932 28624 5972 28664
rect 5836 28456 5876 28496
rect 5932 28036 5972 28076
rect 5932 27868 5972 27908
rect 5740 26944 5780 26984
rect 4928 26440 4968 26480
rect 5010 26440 5050 26480
rect 5092 26440 5132 26480
rect 5174 26440 5214 26480
rect 5256 26440 5296 26480
rect 5548 26440 5588 26480
rect 5068 26272 5108 26312
rect 5452 26272 5492 26312
rect 4780 25936 4820 25976
rect 4972 25600 5012 25640
rect 4684 25432 4724 25472
rect 4780 25264 4820 25304
rect 5260 26104 5300 26144
rect 5164 25516 5204 25556
rect 5260 25432 5300 25472
rect 5164 25348 5204 25388
rect 5068 25096 5108 25136
rect 4928 24928 4968 24968
rect 5010 24928 5050 24968
rect 5092 24928 5132 24968
rect 5174 24928 5214 24968
rect 5256 24928 5296 24968
rect 5452 25180 5492 25220
rect 4876 24760 4916 24800
rect 5356 24760 5396 24800
rect 5356 24424 5396 24464
rect 4588 24088 4628 24128
rect 5260 24088 5300 24128
rect 4928 23416 4968 23456
rect 5010 23416 5050 23456
rect 5092 23416 5132 23456
rect 5174 23416 5214 23456
rect 5256 23416 5296 23456
rect 5452 23752 5492 23792
rect 5356 22828 5396 22868
rect 4492 22240 4532 22280
rect 4492 20056 4532 20096
rect 3436 19972 3476 20012
rect 4396 19972 4436 20012
rect 3340 18712 3380 18752
rect 3340 18124 3380 18164
rect 3244 17788 3284 17828
rect 3244 17284 3284 17324
rect 5452 22240 5492 22280
rect 4684 22072 4724 22112
rect 4780 21988 4820 22028
rect 4684 20896 4724 20936
rect 4928 21904 4968 21944
rect 5010 21904 5050 21944
rect 5092 21904 5132 21944
rect 5174 21904 5214 21944
rect 5256 21904 5296 21944
rect 5164 21736 5204 21776
rect 5356 21652 5396 21692
rect 5164 21603 5204 21608
rect 5164 21568 5204 21603
rect 5644 25432 5684 25472
rect 5932 26692 5972 26732
rect 6700 32824 6740 32864
rect 7084 33916 7124 33956
rect 6892 33580 6932 33620
rect 7084 33076 7124 33116
rect 7276 36604 7316 36644
rect 7276 34252 7316 34292
rect 7276 33916 7316 33956
rect 7276 33664 7316 33704
rect 7276 33412 7316 33452
rect 7468 37024 7508 37064
rect 7468 36688 7508 36728
rect 7564 36604 7604 36644
rect 7564 36436 7604 36476
rect 7564 35764 7604 35804
rect 7468 34588 7508 34628
rect 7564 33916 7604 33956
rect 7468 33832 7508 33872
rect 7468 33664 7508 33704
rect 7564 33412 7604 33452
rect 7372 33244 7412 33284
rect 6796 32656 6836 32696
rect 6892 31816 6932 31856
rect 6892 31564 6932 31604
rect 6700 31312 6740 31352
rect 7180 32908 7220 32948
rect 7084 31144 7124 31184
rect 7084 30556 7124 30596
rect 6412 30220 6452 30260
rect 6988 30220 7028 30260
rect 6412 29800 6452 29840
rect 6316 29380 6356 29420
rect 7852 37528 7892 37568
rect 7756 37192 7796 37232
rect 7852 37108 7892 37148
rect 8428 49372 8468 49412
rect 8620 51640 8660 51680
rect 8620 51220 8660 51260
rect 9580 57856 9620 57896
rect 9580 57520 9620 57560
rect 9676 57100 9716 57140
rect 10060 59788 10100 59828
rect 9964 58696 10004 58736
rect 9964 58360 10004 58400
rect 9868 57436 9908 57476
rect 9292 56260 9332 56300
rect 9196 56092 9236 56132
rect 9196 54832 9236 54872
rect 9484 56176 9524 56216
rect 9580 56008 9620 56048
rect 9676 55672 9716 55712
rect 10252 62224 10292 62264
rect 10444 60460 10484 60500
rect 10156 59200 10196 59240
rect 10348 59872 10388 59912
rect 10156 58108 10196 58148
rect 10252 57772 10292 57812
rect 10444 59368 10484 59408
rect 10444 58360 10484 58400
rect 11212 62896 11252 62936
rect 10924 61636 10964 61676
rect 11212 61552 11252 61592
rect 10924 61048 10964 61088
rect 11116 61048 11156 61088
rect 10924 60712 10964 60752
rect 10924 60124 10964 60164
rect 10732 60049 10772 60080
rect 10732 60040 10772 60049
rect 10828 59956 10868 59996
rect 10924 59872 10964 59912
rect 10732 59368 10772 59408
rect 10636 58192 10676 58232
rect 10156 57100 10196 57140
rect 9964 55672 10004 55712
rect 9868 55504 9908 55544
rect 9868 55252 9908 55292
rect 9868 55084 9908 55124
rect 10156 55084 10196 55124
rect 8716 50212 8756 50252
rect 8812 49960 8852 50000
rect 8716 49540 8756 49580
rect 8620 49456 8660 49496
rect 9100 53355 9140 53360
rect 9100 53320 9140 53355
rect 9292 53488 9332 53528
rect 9580 53908 9620 53948
rect 9196 53236 9236 53276
rect 9772 53320 9812 53360
rect 9388 51724 9428 51764
rect 9292 51640 9332 51680
rect 9196 51304 9236 51344
rect 9292 51052 9332 51092
rect 8908 49456 8948 49496
rect 8908 48784 8948 48824
rect 9100 48784 9140 48824
rect 9388 48784 9428 48824
rect 9004 48196 9044 48236
rect 8908 48112 8948 48152
rect 9004 47776 9044 47816
rect 8620 46432 8660 46472
rect 8908 46180 8948 46220
rect 8812 46012 8852 46052
rect 8812 45172 8852 45212
rect 9004 45004 9044 45044
rect 8812 43492 8852 43532
rect 8428 43324 8468 43364
rect 9004 43240 9044 43280
rect 8908 43156 8948 43196
rect 8812 42064 8852 42104
rect 9964 54160 10004 54200
rect 10060 53992 10100 54032
rect 9964 53236 10004 53276
rect 9580 51640 9620 51680
rect 9388 48028 9428 48068
rect 9484 47944 9524 47984
rect 9292 47776 9332 47816
rect 9196 45928 9236 45968
rect 9196 44920 9236 44960
rect 9484 46432 9524 46472
rect 9388 46180 9428 46220
rect 9580 46264 9620 46304
rect 9676 46180 9716 46220
rect 9676 45844 9716 45884
rect 9676 44416 9716 44456
rect 9484 43996 9524 44036
rect 9292 43912 9332 43952
rect 10156 53824 10196 53864
rect 10348 57436 10388 57476
rect 10348 55924 10388 55964
rect 10540 56092 10580 56132
rect 10636 55924 10676 55964
rect 10444 54832 10484 54872
rect 10348 54160 10388 54200
rect 10348 53992 10388 54032
rect 10348 53068 10388 53108
rect 10732 55504 10772 55544
rect 11212 60712 11252 60752
rect 11404 63232 11444 63272
rect 11788 69280 11828 69320
rect 11692 68860 11732 68900
rect 11788 68692 11828 68732
rect 11788 67768 11828 67808
rect 11692 67180 11732 67220
rect 11788 66928 11828 66968
rect 11788 66760 11828 66800
rect 11788 66592 11828 66632
rect 11692 66172 11732 66212
rect 11692 66004 11732 66044
rect 11596 62812 11636 62852
rect 12364 83056 12404 83096
rect 12364 76840 12404 76880
rect 12940 84400 12980 84440
rect 13516 85576 13556 85616
rect 13708 84484 13748 84524
rect 13324 84400 13364 84440
rect 13900 84400 13940 84440
rect 14092 84736 14132 84776
rect 13324 84232 13364 84272
rect 13996 84232 14036 84272
rect 13996 83560 14036 83600
rect 13708 83476 13748 83516
rect 13132 83308 13172 83348
rect 13900 83308 13940 83348
rect 13516 83140 13556 83180
rect 13036 81880 13076 81920
rect 12844 76840 12884 76880
rect 12556 74656 12596 74696
rect 12268 73648 12308 73688
rect 12172 72976 12212 73016
rect 12364 72724 12404 72764
rect 12172 71464 12212 71504
rect 12172 70456 12212 70496
rect 12172 69868 12212 69908
rect 12076 69784 12116 69824
rect 11980 69700 12020 69740
rect 11980 68692 12020 68732
rect 12076 68440 12116 68480
rect 12076 68104 12116 68144
rect 11884 66508 11924 66548
rect 11884 66172 11924 66212
rect 11884 65332 11924 65372
rect 11884 64660 11924 64700
rect 12076 66928 12116 66968
rect 12172 66760 12212 66800
rect 12172 66508 12212 66548
rect 11788 62812 11828 62852
rect 11020 58864 11060 58904
rect 11020 58696 11060 58736
rect 11212 60124 11252 60164
rect 11308 59284 11348 59324
rect 11212 58864 11252 58904
rect 11116 58360 11156 58400
rect 11020 57940 11060 57980
rect 11308 58528 11348 58568
rect 11308 56932 11348 56972
rect 11212 56764 11252 56804
rect 11116 56596 11156 56636
rect 11020 56260 11060 56300
rect 11308 55672 11348 55712
rect 11020 55504 11060 55544
rect 9868 51556 9908 51596
rect 10060 50968 10100 51008
rect 9868 49456 9908 49496
rect 9868 48028 9908 48068
rect 9964 46432 10004 46472
rect 10252 51640 10292 51680
rect 10444 50968 10484 51008
rect 10540 50548 10580 50588
rect 10252 50296 10292 50336
rect 10828 54916 10868 54956
rect 10828 54496 10868 54536
rect 11308 54832 11348 54872
rect 11500 61552 11540 61592
rect 11692 62224 11732 62264
rect 11596 60796 11636 60836
rect 11692 60376 11732 60416
rect 11692 59872 11732 59912
rect 11596 59032 11636 59072
rect 11500 57436 11540 57476
rect 12076 63904 12116 63944
rect 12076 63232 12116 63272
rect 11980 62224 12020 62264
rect 12460 72136 12500 72176
rect 12364 71800 12404 71840
rect 12460 71632 12500 71672
rect 12364 66676 12404 66716
rect 12556 71464 12596 71504
rect 12652 71044 12692 71084
rect 12940 76756 12980 76796
rect 14476 84736 14516 84776
rect 14380 84316 14420 84356
rect 14284 83476 14324 83516
rect 14284 83308 14324 83348
rect 14764 84400 14804 84440
rect 14668 83308 14708 83348
rect 14572 83224 14612 83264
rect 15052 84316 15092 84356
rect 15436 84400 15476 84440
rect 15052 83308 15092 83348
rect 14188 82552 14228 82592
rect 14572 81880 14612 81920
rect 13132 71968 13172 72008
rect 13036 70624 13076 70664
rect 13612 71968 13652 72008
rect 13132 69700 13172 69740
rect 13036 68944 13076 68984
rect 12844 68860 12884 68900
rect 12748 68020 12788 68060
rect 12748 67348 12788 67388
rect 12556 66844 12596 66884
rect 12460 66004 12500 66044
rect 12364 65584 12404 65624
rect 12556 65500 12596 65540
rect 12364 65332 12404 65372
rect 12556 65332 12596 65372
rect 12364 65164 12404 65204
rect 12364 64828 12404 64868
rect 12268 64240 12308 64280
rect 12268 63904 12308 63944
rect 11884 60796 11924 60836
rect 12076 60964 12116 61004
rect 11980 60712 12020 60752
rect 11788 59200 11828 59240
rect 11692 57856 11732 57896
rect 11404 54664 11444 54704
rect 11308 54412 11348 54452
rect 11596 57016 11636 57056
rect 11596 56764 11636 56804
rect 11212 54160 11252 54200
rect 10732 53236 10772 53276
rect 10924 53068 10964 53108
rect 11116 53320 11156 53360
rect 11884 58696 11924 58736
rect 12076 59452 12116 59492
rect 11980 58528 12020 58568
rect 11884 57856 11924 57896
rect 12556 64408 12596 64448
rect 12460 63904 12500 63944
rect 13036 68356 13076 68396
rect 13516 69700 13556 69740
rect 13804 71464 13844 71504
rect 13804 71044 13844 71084
rect 13708 69280 13748 69320
rect 13324 69028 13364 69068
rect 13708 68776 13748 68816
rect 12940 66928 12980 66968
rect 12844 66424 12884 66464
rect 13036 66592 13076 66632
rect 13132 66508 13172 66548
rect 13708 68188 13748 68228
rect 13324 68020 13364 68060
rect 13804 68020 13844 68060
rect 13324 66928 13364 66968
rect 13804 67348 13844 67388
rect 14284 72304 14324 72344
rect 13996 71380 14036 71420
rect 14476 70624 14516 70664
rect 14380 70204 14420 70244
rect 14572 69700 14612 69740
rect 14284 69112 14324 69152
rect 14092 67348 14132 67388
rect 13900 67180 13940 67220
rect 14188 66928 14228 66968
rect 13228 66424 13268 66464
rect 12844 66088 12884 66128
rect 13612 66088 13652 66128
rect 13036 66004 13076 66044
rect 13228 66004 13268 66044
rect 13708 66004 13748 66044
rect 13324 65920 13364 65960
rect 14188 65920 14228 65960
rect 14380 65920 14420 65960
rect 13612 65836 13652 65876
rect 12748 65752 12788 65792
rect 13324 65500 13364 65540
rect 12748 65248 12788 65288
rect 12748 64912 12788 64952
rect 13132 65416 13172 65456
rect 13228 65416 13268 65456
rect 13036 65332 13076 65372
rect 13420 65248 13460 65288
rect 13036 64996 13076 65036
rect 13516 64996 13556 65036
rect 12748 64492 12788 64532
rect 12940 64576 12980 64616
rect 13036 64492 13076 64532
rect 12844 64408 12884 64448
rect 12940 63988 12980 64028
rect 12556 63736 12596 63776
rect 12460 62728 12500 62768
rect 12460 62392 12500 62432
rect 12556 62224 12596 62264
rect 13324 64408 13364 64448
rect 13228 64240 13268 64280
rect 13516 64576 13556 64616
rect 13516 64324 13556 64364
rect 13132 63400 13172 63440
rect 13228 63064 13268 63104
rect 12364 61048 12404 61088
rect 12748 61048 12788 61088
rect 12364 60899 12404 60920
rect 12364 60880 12404 60899
rect 12652 60880 12692 60920
rect 12556 60292 12596 60332
rect 12460 60124 12500 60164
rect 12364 59452 12404 59492
rect 12364 59032 12404 59072
rect 12172 57604 12212 57644
rect 12364 57184 12404 57224
rect 12268 56680 12308 56720
rect 12076 56596 12116 56636
rect 12844 60880 12884 60920
rect 13036 60880 13076 60920
rect 12748 60040 12788 60080
rect 12844 59956 12884 59996
rect 13228 60376 13268 60416
rect 13708 65584 13748 65624
rect 13900 65332 13940 65372
rect 13804 64912 13844 64952
rect 13708 64492 13748 64532
rect 14476 65080 14516 65120
rect 14284 64828 14324 64868
rect 14476 64828 14516 64868
rect 14092 64744 14132 64784
rect 14188 64660 14228 64700
rect 13804 64324 13844 64364
rect 13804 63904 13844 63944
rect 13708 62560 13748 62600
rect 13420 61552 13460 61592
rect 13516 60880 13556 60920
rect 13036 59452 13076 59492
rect 12940 59368 12980 59408
rect 12556 59032 12596 59072
rect 12556 58612 12596 58652
rect 12556 58108 12596 58148
rect 12839 58612 12879 58652
rect 12940 58528 12980 58568
rect 13036 58360 13076 58400
rect 13324 59452 13364 59492
rect 13228 58360 13268 58400
rect 12460 57100 12500 57140
rect 12940 57940 12980 57980
rect 11980 56260 12020 56300
rect 11884 56008 11924 56048
rect 11692 55252 11732 55292
rect 12364 55252 12404 55292
rect 12076 54664 12116 54704
rect 11788 54328 11828 54368
rect 12268 54328 12308 54368
rect 11404 54076 11444 54116
rect 11404 52564 11444 52604
rect 11980 53992 12020 54032
rect 11788 53656 11828 53696
rect 11596 53236 11636 53276
rect 11212 51640 11252 51680
rect 11500 51640 11540 51680
rect 10444 50212 10484 50252
rect 10636 50212 10676 50252
rect 10348 49540 10388 49580
rect 10636 47692 10676 47732
rect 9868 46264 9908 46304
rect 10060 46264 10100 46304
rect 10060 46096 10100 46136
rect 9964 45676 10004 45716
rect 10060 44248 10100 44288
rect 9868 44164 9908 44204
rect 9868 43912 9908 43952
rect 9772 43828 9812 43868
rect 9388 43492 9428 43532
rect 9196 42400 9236 42440
rect 8812 41560 8852 41600
rect 9004 41728 9044 41768
rect 9004 41560 9044 41600
rect 8332 38956 8372 38996
rect 8716 38872 8756 38912
rect 8524 38200 8564 38240
rect 9100 41308 9140 41348
rect 9004 40720 9044 40760
rect 9004 40468 9044 40508
rect 8908 40384 8948 40424
rect 8908 39712 8948 39752
rect 9388 41728 9428 41768
rect 9292 41560 9332 41600
rect 9484 41560 9524 41600
rect 10348 46516 10388 46556
rect 10540 46432 10580 46472
rect 10444 46096 10484 46136
rect 10348 45676 10388 45716
rect 11020 50800 11060 50840
rect 11116 49456 11156 49496
rect 11116 46768 11156 46808
rect 11500 50968 11540 51008
rect 11980 53152 12020 53192
rect 11980 52900 12020 52940
rect 12172 53488 12212 53528
rect 11692 51052 11732 51092
rect 11596 50296 11636 50336
rect 11404 50212 11444 50252
rect 11308 49624 11348 49664
rect 11596 49624 11636 49664
rect 11788 50968 11828 51008
rect 11500 48784 11540 48824
rect 11500 47188 11540 47228
rect 11404 46684 11444 46724
rect 10732 46516 10772 46556
rect 10924 46432 10964 46472
rect 10924 46180 10964 46220
rect 10828 44920 10868 44960
rect 11212 44920 11252 44960
rect 12556 54851 12596 54872
rect 12556 54832 12596 54851
rect 12556 53908 12596 53948
rect 12364 53488 12404 53528
rect 12364 52564 12404 52604
rect 12268 52060 12308 52100
rect 13132 56680 13172 56720
rect 13324 57688 13364 57728
rect 13324 57436 13364 57476
rect 13324 56764 13364 56804
rect 12748 53992 12788 54032
rect 12748 52984 12788 53024
rect 12652 52648 12692 52688
rect 12940 54328 12980 54368
rect 12364 51892 12404 51932
rect 12652 51808 12692 51848
rect 12172 51052 12212 51092
rect 12268 50548 12308 50588
rect 12076 49792 12116 49832
rect 11884 48616 11924 48656
rect 11788 47020 11828 47060
rect 12172 49540 12212 49580
rect 12076 46012 12116 46052
rect 11884 45340 11924 45380
rect 11404 45088 11444 45128
rect 11308 44416 11348 44456
rect 10636 44164 10676 44204
rect 12076 45088 12116 45128
rect 12364 47188 12404 47228
rect 12364 47020 12404 47060
rect 12364 46684 12404 46724
rect 12268 46516 12308 46556
rect 12268 45340 12308 45380
rect 12748 50968 12788 51008
rect 12844 50296 12884 50336
rect 12748 49708 12788 49748
rect 13132 53908 13172 53948
rect 13228 52900 13268 52940
rect 13036 52648 13076 52688
rect 13228 52312 13268 52352
rect 13132 52228 13172 52268
rect 13036 52144 13076 52184
rect 13612 58780 13652 58820
rect 13516 58612 13556 58652
rect 13612 58528 13652 58568
rect 13516 57772 13556 57812
rect 13900 61636 13940 61676
rect 13996 60964 14036 61004
rect 14380 64660 14420 64700
rect 14284 63820 14324 63860
rect 15628 81292 15668 81332
rect 15820 79024 15860 79064
rect 15340 75664 15380 75704
rect 15052 72304 15092 72344
rect 15148 71800 15188 71840
rect 15052 70792 15092 70832
rect 14860 70624 14900 70664
rect 15052 70624 15092 70664
rect 14764 69280 14804 69320
rect 14764 69112 14804 69152
rect 15052 69784 15092 69824
rect 15916 72220 15956 72260
rect 15820 71716 15860 71756
rect 15244 70540 15284 70580
rect 15532 70624 15572 70664
rect 15820 71044 15860 71084
rect 16396 84400 16436 84440
rect 16588 84400 16628 84440
rect 16876 85828 16916 85868
rect 16204 71884 16244 71924
rect 16204 71716 16244 71756
rect 16108 71548 16148 71588
rect 16012 70960 16052 71000
rect 15916 70624 15956 70664
rect 15916 70372 15956 70412
rect 15724 70288 15764 70328
rect 15340 70120 15380 70160
rect 15532 69868 15572 69908
rect 15244 69448 15284 69488
rect 15148 69364 15188 69404
rect 15052 69196 15092 69236
rect 14956 69112 14996 69152
rect 14956 68440 14996 68480
rect 14860 67684 14900 67724
rect 15052 68020 15092 68060
rect 14764 66928 14804 66968
rect 15340 69280 15380 69320
rect 15340 68272 15380 68312
rect 15148 67684 15188 67724
rect 15436 67684 15476 67724
rect 15628 68944 15668 68984
rect 15628 68104 15668 68144
rect 14956 66340 14996 66380
rect 14860 65416 14900 65456
rect 14860 65164 14900 65204
rect 14764 64828 14804 64868
rect 14860 64660 14900 64700
rect 14668 64324 14708 64364
rect 14764 64156 14804 64196
rect 14668 63904 14708 63944
rect 15532 67516 15572 67556
rect 15820 68440 15860 68480
rect 15724 67684 15764 67724
rect 15436 67432 15476 67472
rect 15628 67432 15668 67472
rect 15628 67264 15668 67304
rect 15340 64660 15380 64700
rect 16012 69978 16052 69992
rect 16012 69952 16052 69978
rect 16204 71044 16244 71084
rect 17932 83812 17972 83852
rect 18124 83476 18164 83516
rect 18412 83812 18452 83852
rect 18316 83728 18356 83768
rect 18316 83476 18356 83516
rect 18508 83476 18548 83516
rect 19084 84988 19124 85028
rect 19660 84988 19700 85028
rect 18808 84652 18848 84692
rect 18890 84652 18930 84692
rect 18972 84652 19012 84692
rect 19054 84652 19094 84692
rect 19136 84652 19176 84692
rect 18892 83728 18932 83768
rect 18700 83476 18740 83516
rect 19084 83476 19124 83516
rect 19276 83476 19316 83516
rect 18796 83308 18836 83348
rect 19276 83308 19316 83348
rect 18808 83140 18848 83180
rect 18890 83140 18930 83180
rect 18972 83140 19012 83180
rect 19054 83140 19094 83180
rect 19136 83140 19176 83180
rect 19468 83476 19508 83516
rect 20048 83896 20088 83936
rect 20130 83896 20170 83936
rect 20212 83896 20252 83936
rect 20294 83896 20334 83936
rect 20376 83896 20416 83936
rect 17356 82552 17396 82592
rect 17740 82552 17780 82592
rect 18700 82048 18740 82088
rect 18124 81880 18164 81920
rect 18508 81880 18548 81920
rect 16780 72304 16820 72344
rect 16588 71632 16628 71672
rect 16396 71548 16436 71588
rect 16396 70120 16436 70160
rect 16300 70036 16340 70076
rect 16588 69952 16628 69992
rect 16108 69700 16148 69740
rect 16300 69616 16340 69656
rect 16012 69364 16052 69404
rect 17164 71800 17204 71840
rect 18316 71884 18356 71924
rect 17548 71380 17588 71420
rect 18124 70876 18164 70916
rect 17644 70456 17684 70496
rect 17164 70036 17204 70076
rect 17068 69952 17108 69992
rect 16684 69532 16724 69572
rect 16396 68608 16436 68648
rect 16300 68440 16340 68480
rect 15916 67516 15956 67556
rect 15820 66928 15860 66968
rect 16300 67768 16340 67808
rect 16108 67600 16148 67640
rect 16012 66508 16052 66548
rect 16204 67516 16244 67556
rect 16012 66088 16052 66128
rect 17068 67768 17108 67808
rect 16876 67684 16916 67724
rect 16972 67600 17012 67640
rect 16492 67432 16532 67472
rect 16300 66508 16340 66548
rect 16876 67432 16916 67472
rect 16876 66928 16916 66968
rect 17068 66676 17108 66716
rect 16588 66340 16628 66380
rect 16780 66340 16820 66380
rect 16588 66088 16628 66128
rect 16876 66172 16916 66212
rect 16684 66004 16724 66044
rect 15820 65668 15860 65708
rect 15724 65416 15764 65456
rect 15532 64408 15572 64448
rect 14860 63736 14900 63776
rect 14188 61132 14228 61172
rect 15052 62560 15092 62600
rect 14668 62224 14708 62264
rect 15052 62224 15092 62264
rect 14380 61468 14420 61508
rect 14380 61048 14420 61088
rect 14956 61636 14996 61676
rect 14572 61048 14612 61088
rect 14476 60964 14516 61004
rect 14572 60880 14612 60920
rect 14380 60460 14420 60500
rect 14380 60040 14420 60080
rect 13900 59956 13940 59996
rect 13804 59536 13844 59576
rect 13804 58360 13844 58400
rect 13804 57688 13844 57728
rect 13900 57184 13940 57224
rect 13900 56932 13940 56972
rect 13804 56680 13844 56720
rect 13708 55336 13748 55376
rect 13708 55084 13748 55124
rect 13516 54748 13556 54788
rect 13420 54328 13460 54368
rect 13420 53992 13460 54032
rect 13324 51892 13364 51932
rect 13132 51808 13172 51848
rect 13324 50968 13364 51008
rect 13228 50464 13268 50504
rect 13612 53908 13652 53948
rect 13804 53992 13844 54032
rect 13516 52228 13556 52268
rect 13804 52648 13844 52688
rect 13804 52312 13844 52352
rect 13708 52228 13748 52268
rect 13612 51892 13652 51932
rect 12940 49456 12980 49496
rect 12844 49372 12884 49412
rect 12844 49204 12884 49244
rect 13516 49624 13556 49664
rect 13516 49456 13556 49496
rect 13516 49120 13556 49160
rect 12748 47272 12788 47312
rect 12652 46264 12692 46304
rect 12460 44416 12500 44456
rect 10444 42064 10484 42104
rect 10828 41896 10868 41936
rect 10060 41812 10100 41852
rect 9964 40468 10004 40508
rect 9868 40384 9908 40424
rect 9772 40132 9812 40172
rect 9964 40048 10004 40088
rect 10540 41476 10580 41516
rect 10444 41308 10484 41348
rect 11116 42064 11156 42104
rect 11116 41896 11156 41936
rect 11596 41476 11636 41516
rect 10924 41140 10964 41180
rect 10636 40720 10676 40760
rect 10444 40384 10484 40424
rect 10636 40384 10676 40424
rect 11500 41224 11540 41264
rect 11500 40468 11540 40508
rect 11020 40216 11060 40256
rect 10060 39964 10100 40004
rect 9292 39544 9332 39584
rect 9100 39040 9140 39080
rect 9196 38956 9236 38996
rect 8812 38536 8852 38576
rect 8716 36856 8756 36896
rect 8716 36520 8756 36560
rect 7756 35512 7796 35552
rect 7756 34336 7796 34376
rect 7756 34000 7796 34040
rect 7660 32908 7700 32948
rect 7564 32656 7604 32696
rect 7756 32656 7796 32696
rect 8140 35512 8180 35552
rect 8044 35344 8084 35384
rect 7948 34672 7988 34712
rect 7948 34252 7988 34292
rect 7948 33160 7988 33200
rect 8140 34336 8180 34376
rect 8908 38200 8948 38240
rect 9004 37192 9044 37232
rect 8524 34336 8564 34376
rect 8332 33916 8372 33956
rect 8236 33664 8276 33704
rect 8332 33160 8372 33200
rect 8044 32908 8084 32948
rect 7949 32740 7989 32780
rect 7852 32572 7892 32612
rect 7756 32488 7796 32528
rect 7564 32236 7604 32276
rect 7660 32152 7700 32192
rect 7372 31984 7412 32024
rect 7276 31396 7316 31436
rect 7276 31144 7316 31184
rect 6988 29128 7028 29168
rect 6412 28960 6452 29000
rect 6604 28960 6644 29000
rect 6412 28708 6452 28748
rect 6316 28288 6356 28328
rect 6316 28036 6356 28076
rect 6892 28456 6932 28496
rect 6700 28288 6740 28328
rect 6412 26860 6452 26900
rect 6220 26692 6260 26732
rect 6028 25852 6068 25892
rect 5836 25516 5876 25556
rect 5836 25348 5876 25388
rect 5740 24928 5780 24968
rect 5932 24508 5972 24548
rect 5644 24172 5684 24212
rect 6412 25264 6452 25304
rect 6316 25012 6356 25052
rect 6124 24424 6164 24464
rect 6220 24340 6260 24380
rect 6028 24088 6068 24128
rect 5836 23836 5876 23876
rect 5740 23752 5780 23792
rect 6316 23836 6356 23876
rect 6124 23668 6164 23708
rect 6028 22996 6068 23036
rect 5740 22240 5780 22280
rect 6124 22240 6164 22280
rect 6220 22156 6260 22196
rect 6412 22324 6452 22364
rect 6796 28120 6836 28160
rect 6796 27280 6836 27320
rect 6796 26860 6836 26900
rect 6604 25684 6644 25724
rect 6700 25264 6740 25304
rect 6892 26776 6932 26816
rect 7084 28204 7124 28244
rect 7372 29128 7412 29168
rect 7084 26104 7124 26144
rect 6796 25180 6836 25220
rect 6988 25180 7028 25220
rect 6892 25012 6932 25052
rect 6604 23836 6644 23876
rect 6700 23752 6740 23792
rect 6604 22828 6644 22868
rect 6983 24760 7023 24800
rect 7084 24760 7124 24800
rect 7084 24340 7124 24380
rect 7276 26776 7316 26816
rect 7564 27952 7604 27992
rect 7468 26272 7508 26312
rect 7372 26104 7412 26144
rect 7276 25264 7316 25304
rect 7372 24424 7412 24464
rect 7180 24256 7220 24296
rect 7564 25852 7604 25892
rect 8236 32404 8276 32444
rect 8524 33076 8564 33116
rect 8428 32908 8468 32948
rect 7852 32152 7892 32192
rect 8332 32236 8372 32276
rect 8812 34084 8852 34124
rect 8716 33664 8756 33704
rect 8716 32152 8756 32192
rect 8140 31396 8180 31436
rect 8332 31396 8372 31436
rect 8044 31144 8084 31184
rect 7948 29296 7988 29336
rect 7852 28204 7892 28244
rect 7756 27028 7796 27068
rect 8236 31312 8276 31352
rect 8140 28120 8180 28160
rect 8044 27952 8084 27992
rect 7756 26692 7796 26732
rect 7756 26104 7796 26144
rect 7756 25852 7796 25892
rect 7660 25516 7700 25556
rect 7276 23836 7316 23876
rect 6892 22996 6932 23036
rect 7084 23248 7124 23288
rect 7564 23920 7604 23960
rect 7468 23668 7508 23708
rect 7084 22828 7124 22868
rect 6796 22240 6836 22280
rect 6700 22156 6740 22196
rect 5548 21820 5588 21860
rect 5932 21820 5972 21860
rect 5548 21568 5588 21608
rect 5740 21568 5780 21608
rect 5356 21148 5396 21188
rect 5356 20896 5396 20936
rect 5068 20812 5108 20852
rect 5164 20728 5204 20768
rect 5356 20728 5396 20768
rect 5932 21484 5972 21524
rect 6028 21400 6068 21440
rect 6028 20896 6068 20936
rect 5836 20728 5876 20768
rect 5644 20476 5684 20516
rect 4928 20392 4968 20432
rect 5010 20392 5050 20432
rect 5092 20392 5132 20432
rect 5174 20392 5214 20432
rect 5256 20392 5296 20432
rect 5356 20392 5396 20432
rect 4876 20140 4916 20180
rect 4684 19888 4724 19928
rect 5260 19972 5300 20012
rect 3688 19636 3728 19676
rect 3770 19636 3810 19676
rect 3852 19636 3892 19676
rect 3934 19636 3974 19676
rect 4016 19636 4056 19676
rect 4204 19300 4244 19340
rect 4300 18544 4340 18584
rect 4108 18292 4148 18332
rect 3532 18124 3572 18164
rect 3688 18124 3728 18164
rect 3770 18124 3810 18164
rect 3852 18124 3892 18164
rect 3934 18124 3974 18164
rect 4016 18124 4056 18164
rect 3628 17956 3668 17996
rect 3724 17704 3764 17744
rect 3724 16780 3764 16820
rect 4012 16780 4052 16820
rect 4300 16780 4340 16820
rect 3688 16612 3728 16652
rect 3770 16612 3810 16652
rect 3852 16612 3892 16652
rect 3934 16612 3974 16652
rect 4016 16612 4056 16652
rect 4108 16444 4148 16484
rect 2860 16360 2900 16400
rect 3340 16360 3380 16400
rect 2764 16192 2804 16232
rect 2476 15688 2516 15728
rect 2764 15688 2804 15728
rect 1900 15268 1940 15308
rect 1516 14260 1556 14300
rect 1228 13504 1268 13544
rect 1804 14176 1844 14216
rect 1228 13252 1268 13292
rect 1324 12496 1364 12536
rect 1420 11152 1460 11192
rect 1612 13000 1652 13040
rect 1708 12832 1748 12872
rect 2092 14596 2132 14636
rect 1996 14428 2036 14468
rect 2284 14008 2324 14048
rect 2092 12748 2132 12788
rect 1996 11908 2036 11948
rect 1708 11824 1748 11864
rect 1996 11740 2036 11780
rect 1612 10900 1652 10940
rect 1900 11488 1940 11528
rect 3148 16192 3188 16232
rect 3052 15688 3092 15728
rect 3148 15520 3188 15560
rect 3340 16192 3380 16232
rect 3532 16192 3572 16232
rect 4300 16192 4340 16232
rect 4300 15772 4340 15812
rect 5260 19216 5300 19256
rect 5548 20056 5588 20096
rect 5452 19720 5492 19760
rect 5740 19636 5780 19676
rect 5644 19468 5684 19508
rect 4928 18880 4968 18920
rect 5010 18880 5050 18920
rect 5092 18880 5132 18920
rect 5174 18880 5214 18920
rect 5256 18880 5296 18920
rect 4780 18796 4820 18836
rect 4684 18040 4724 18080
rect 5356 18544 5396 18584
rect 3975 15688 4015 15728
rect 4396 15688 4436 15728
rect 3340 15436 3380 15476
rect 3532 15436 3572 15476
rect 3820 15520 3860 15560
rect 4396 15436 4436 15476
rect 3436 15268 3476 15308
rect 3688 15100 3728 15140
rect 3770 15100 3810 15140
rect 3852 15100 3892 15140
rect 3934 15100 3974 15140
rect 4016 15100 4056 15140
rect 2956 14596 2996 14636
rect 2860 14512 2900 14552
rect 3340 14512 3380 14552
rect 3532 14512 3572 14552
rect 2668 14008 2708 14048
rect 2572 13504 2612 13544
rect 3244 14008 3284 14048
rect 2860 13504 2900 13544
rect 2476 13168 2516 13208
rect 2764 13168 2804 13208
rect 2380 12664 2420 12704
rect 2188 12580 2228 12620
rect 2668 12664 2708 12704
rect 2956 12664 2996 12704
rect 2764 12580 2804 12620
rect 2188 11908 2228 11948
rect 2380 11404 2420 11444
rect 1612 10228 1652 10268
rect 1900 10060 1940 10100
rect 1900 9808 1940 9848
rect 1324 9472 1364 9512
rect 1324 9304 1364 9344
rect 1228 8800 1268 8840
rect 1516 9220 1556 9260
rect 1420 8884 1460 8924
rect 1516 8128 1556 8168
rect 2188 11068 2228 11108
rect 2092 9892 2132 9932
rect 2092 9388 2132 9428
rect 2284 10144 2324 10184
rect 1708 8716 1748 8756
rect 1900 8464 1940 8504
rect 1804 8296 1844 8336
rect 1516 7960 1556 8000
rect 1324 7456 1364 7496
rect 1324 6112 1364 6152
rect 1228 5356 1268 5396
rect 1612 7876 1652 7916
rect 1708 7456 1748 7496
rect 1612 7372 1652 7412
rect 1708 6784 1748 6824
rect 3052 12580 3092 12620
rect 3244 12580 3284 12620
rect 3148 12496 3188 12536
rect 3052 12412 3092 12452
rect 2476 10564 2516 10604
rect 2476 10396 2516 10436
rect 3820 14344 3860 14384
rect 4204 14680 4244 14720
rect 4300 14344 4340 14384
rect 3436 14008 3476 14048
rect 5260 17536 5300 17576
rect 5644 19048 5684 19088
rect 5644 18880 5684 18920
rect 5548 18712 5588 18752
rect 5548 18544 5588 18584
rect 6316 21568 6356 21608
rect 6220 19888 6260 19928
rect 6124 19216 6164 19256
rect 6028 19132 6068 19172
rect 5932 19048 5972 19088
rect 5740 18376 5780 18416
rect 5644 17704 5684 17744
rect 5356 17452 5396 17492
rect 4928 17368 4968 17408
rect 5010 17368 5050 17408
rect 5092 17368 5132 17408
rect 5174 17368 5214 17408
rect 5256 17368 5296 17408
rect 4780 17116 4820 17156
rect 5164 17116 5204 17156
rect 4972 17032 5012 17072
rect 5356 17032 5396 17072
rect 4588 16612 4628 16652
rect 3820 14008 3860 14048
rect 3724 13840 3764 13880
rect 3688 13588 3728 13628
rect 3770 13588 3810 13628
rect 3852 13588 3892 13628
rect 3934 13588 3974 13628
rect 4016 13588 4056 13628
rect 4780 16360 4820 16400
rect 4684 14764 4724 14804
rect 4588 13420 4628 13460
rect 4684 13336 4724 13376
rect 4492 13252 4532 13292
rect 4108 13168 4148 13208
rect 4300 13084 4340 13124
rect 3628 12580 3668 12620
rect 3916 12496 3956 12536
rect 4588 13084 4628 13124
rect 3724 12412 3764 12452
rect 4396 12244 4436 12284
rect 3688 12076 3728 12116
rect 3770 12076 3810 12116
rect 3852 12076 3892 12116
rect 3934 12076 3974 12116
rect 4016 12076 4056 12116
rect 4492 11992 4532 12032
rect 2860 9976 2900 10016
rect 3052 11152 3092 11192
rect 2956 9808 2996 9848
rect 2668 9136 2708 9176
rect 2380 8800 2420 8840
rect 2764 9052 2804 9092
rect 3052 9472 3092 9512
rect 2860 8632 2900 8672
rect 3052 9052 3092 9092
rect 2476 8464 2516 8504
rect 2668 8380 2708 8420
rect 2860 8128 2900 8168
rect 2092 7708 2132 7748
rect 1996 7624 2036 7664
rect 2860 7456 2900 7496
rect 2764 7036 2804 7076
rect 2668 6952 2708 6992
rect 3052 8128 3092 8168
rect 3340 11152 3380 11192
rect 6124 18544 6164 18584
rect 6028 18460 6068 18500
rect 5932 18376 5972 18416
rect 5836 16948 5876 16988
rect 5548 16612 5588 16652
rect 6028 17284 6068 17324
rect 6028 16612 6068 16652
rect 4928 15856 4968 15896
rect 5010 15856 5050 15896
rect 5092 15856 5132 15896
rect 5174 15856 5214 15896
rect 5256 15856 5296 15896
rect 5260 15268 5300 15308
rect 5164 14932 5204 14972
rect 4928 14344 4968 14384
rect 5010 14344 5050 14384
rect 5092 14344 5132 14384
rect 5174 14344 5214 14384
rect 5256 14344 5296 14384
rect 4972 14092 5012 14132
rect 5932 16192 5972 16232
rect 5932 15772 5972 15812
rect 5836 14596 5876 14636
rect 5836 14176 5876 14216
rect 5452 14008 5492 14048
rect 5068 13420 5108 13460
rect 5644 13252 5684 13292
rect 4928 12832 4968 12872
rect 5010 12832 5050 12872
rect 5092 12832 5132 12872
rect 5174 12832 5214 12872
rect 5256 12832 5296 12872
rect 5356 11992 5396 12032
rect 5836 13168 5876 13208
rect 6316 19216 6356 19256
rect 6508 21820 6548 21860
rect 6988 21988 7028 22028
rect 6796 21904 6836 21944
rect 6700 21736 6740 21776
rect 6700 21316 6740 21356
rect 6604 19636 6644 19676
rect 6796 20392 6836 20432
rect 6796 19804 6836 19844
rect 6796 19636 6836 19676
rect 6508 19300 6548 19340
rect 6700 19300 6740 19340
rect 6604 19216 6644 19256
rect 6700 19132 6740 19172
rect 6412 18544 6452 18584
rect 6604 18796 6644 18836
rect 6316 16780 6356 16820
rect 6796 18712 6836 18752
rect 7180 21652 7220 21692
rect 7180 21400 7220 21440
rect 8140 26692 8180 26732
rect 8332 29800 8372 29840
rect 8524 30640 8564 30680
rect 8620 30472 8660 30512
rect 9004 34336 9044 34376
rect 8812 30976 8852 31016
rect 8812 30640 8852 30680
rect 8812 30472 8852 30512
rect 8908 30304 8948 30344
rect 8716 29716 8756 29756
rect 8620 29212 8660 29252
rect 8332 28288 8372 28328
rect 8620 27616 8660 27656
rect 8812 29464 8852 29504
rect 8332 26944 8372 26984
rect 8812 26104 8852 26144
rect 7948 25180 7988 25220
rect 7852 24508 7892 24548
rect 7756 23752 7796 23792
rect 7660 23500 7700 23540
rect 7660 22240 7700 22280
rect 7372 21820 7412 21860
rect 7564 21820 7604 21860
rect 8044 23920 8084 23960
rect 8428 25012 8468 25052
rect 8236 24424 8276 24464
rect 8140 23836 8180 23876
rect 8140 23500 8180 23540
rect 8332 23752 8372 23792
rect 8140 22828 8180 22868
rect 8428 23584 8468 23624
rect 8716 25012 8756 25052
rect 8620 23752 8660 23792
rect 8812 24256 8852 24296
rect 10636 39712 10676 39752
rect 10156 39040 10196 39080
rect 10348 38704 10388 38744
rect 9676 38620 9716 38660
rect 9772 37696 9812 37736
rect 9676 37612 9716 37652
rect 10252 37864 10292 37904
rect 10636 39208 10676 39248
rect 11500 38200 11540 38240
rect 10348 37696 10388 37736
rect 10444 37696 10484 37736
rect 9964 37444 10004 37484
rect 9772 37360 9812 37400
rect 9676 36688 9716 36728
rect 9580 36184 9620 36224
rect 9580 35932 9620 35972
rect 9388 35512 9428 35552
rect 9196 31564 9236 31604
rect 9292 31396 9332 31436
rect 9004 30220 9044 30260
rect 10156 36940 10196 36980
rect 10060 36856 10100 36896
rect 10060 36604 10100 36644
rect 10060 36352 10100 36392
rect 9676 35512 9716 35552
rect 9580 34084 9620 34124
rect 9772 33832 9812 33872
rect 10060 35848 10100 35888
rect 10060 35008 10100 35048
rect 10060 34336 10100 34376
rect 10444 37444 10484 37484
rect 11692 39124 11732 39164
rect 11692 38200 11732 38240
rect 11404 37780 11444 37820
rect 12172 43324 12212 43364
rect 12076 41896 12116 41936
rect 11884 39712 11924 39752
rect 11596 37780 11636 37820
rect 11308 37696 11348 37736
rect 10924 37276 10964 37316
rect 10732 36940 10772 36980
rect 10828 36856 10868 36896
rect 10348 36688 10388 36728
rect 10348 36352 10388 36392
rect 10252 36016 10292 36056
rect 10252 34924 10292 34964
rect 9964 33832 10004 33872
rect 9580 33664 9620 33704
rect 9388 31060 9428 31100
rect 9196 30976 9236 31016
rect 9388 30724 9428 30764
rect 9484 30640 9524 30680
rect 9196 29968 9236 30008
rect 9196 29800 9236 29840
rect 9388 30304 9428 30344
rect 9004 28372 9044 28412
rect 9292 28120 9332 28160
rect 9292 27868 9332 27908
rect 9100 27700 9140 27740
rect 9004 26104 9044 26144
rect 9100 25768 9140 25808
rect 9196 25684 9236 25724
rect 9292 24760 9332 24800
rect 9484 29632 9524 29672
rect 9676 30892 9716 30932
rect 9676 30724 9716 30764
rect 9580 29128 9620 29168
rect 9484 27616 9524 27656
rect 9964 33160 10004 33200
rect 9964 32320 10004 32360
rect 9868 31312 9908 31352
rect 9964 30976 10004 31016
rect 9580 26776 9620 26816
rect 9484 25684 9524 25724
rect 9388 24340 9428 24380
rect 8812 23752 8852 23792
rect 9100 23668 9140 23708
rect 8524 22996 8564 23036
rect 8428 22828 8468 22868
rect 8524 22576 8564 22616
rect 8332 22240 8372 22280
rect 7660 21652 7700 21692
rect 7948 21652 7988 21692
rect 7564 21400 7604 21440
rect 7084 20896 7124 20936
rect 6988 20812 7028 20852
rect 6988 20560 7028 20600
rect 7084 19720 7124 19760
rect 6988 19216 7028 19256
rect 7372 21064 7412 21104
rect 7276 20560 7316 20600
rect 7756 21232 7796 21272
rect 7852 20812 7892 20852
rect 7468 20056 7508 20096
rect 7564 19972 7604 20012
rect 7372 19300 7412 19340
rect 7180 18880 7220 18920
rect 6796 18544 6836 18584
rect 7084 18544 7124 18584
rect 6316 16108 6356 16148
rect 6508 16276 6548 16316
rect 6508 16108 6548 16148
rect 6412 15940 6452 15980
rect 6220 14764 6260 14804
rect 6508 14008 6548 14048
rect 6220 13252 6260 13292
rect 6508 13252 6548 13292
rect 6028 12832 6068 12872
rect 6220 12832 6260 12872
rect 6316 12748 6356 12788
rect 4972 11824 5012 11864
rect 5644 11824 5684 11864
rect 4108 11488 4148 11528
rect 4012 11152 4052 11192
rect 3436 10984 3476 11024
rect 3688 10564 3728 10604
rect 3770 10564 3810 10604
rect 3852 10564 3892 10604
rect 3934 10564 3974 10604
rect 4016 10564 4056 10604
rect 5644 11572 5684 11612
rect 5932 11488 5972 11528
rect 4684 11320 4724 11360
rect 4928 11320 4968 11360
rect 5010 11320 5050 11360
rect 5092 11320 5132 11360
rect 5174 11320 5214 11360
rect 5256 11320 5296 11360
rect 3244 9640 3284 9680
rect 3244 9472 3284 9512
rect 3436 9472 3476 9512
rect 3820 10144 3860 10184
rect 4396 10312 4436 10352
rect 3724 9976 3764 10016
rect 4204 10144 4244 10184
rect 4492 9976 4532 10016
rect 4108 9724 4148 9764
rect 4012 9556 4052 9596
rect 3820 9472 3860 9512
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 5356 11236 5396 11276
rect 4780 11152 4820 11192
rect 4684 10060 4724 10100
rect 4588 9808 4628 9848
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 4300 9472 4340 9512
rect 4780 9640 4820 9680
rect 5073 9556 5113 9596
rect 4204 9136 4244 9176
rect 3340 8632 3380 8672
rect 3468 8632 3508 8672
rect 3244 8464 3284 8504
rect 3724 8800 3764 8840
rect 4108 8716 4148 8756
rect 4012 8632 4052 8672
rect 3916 8380 3956 8420
rect 3244 7792 3284 7832
rect 3436 7876 3476 7916
rect 2092 6784 2132 6824
rect 2668 6784 2708 6824
rect 2860 6784 2900 6824
rect 2284 6700 2324 6740
rect 2956 6700 2996 6740
rect 3057 6700 3097 6740
rect 2188 6532 2228 6572
rect 2572 6448 2612 6488
rect 2380 6364 2420 6404
rect 2668 6364 2708 6404
rect 1900 5440 1940 5480
rect 1132 1156 1172 1196
rect 1420 4432 1460 4472
rect 1804 4768 1844 4808
rect 1708 4600 1748 4640
rect 1996 4348 2036 4388
rect 1420 3424 1460 3464
rect 1612 3256 1652 3296
rect 1708 3172 1748 3212
rect 1900 3004 1940 3044
rect 1804 2920 1844 2960
rect 1612 2500 1652 2540
rect 1516 1744 1556 1784
rect 2188 5860 2228 5900
rect 2284 5776 2324 5816
rect 2284 4096 2324 4136
rect 2284 3424 2324 3464
rect 2188 3340 2228 3380
rect 2092 2164 2132 2204
rect 1900 2080 1940 2120
rect 1996 1744 2036 1784
rect 1516 1072 1556 1112
rect 1804 988 1844 1028
rect 1324 652 1364 692
rect 1900 148 1940 188
rect 2572 5272 2612 5312
rect 2668 4852 2708 4892
rect 2476 4180 2516 4220
rect 2476 3928 2516 3968
rect 3148 6616 3188 6656
rect 4108 8044 4148 8084
rect 3628 7960 3668 8000
rect 4588 7624 4628 7664
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 3724 7288 3764 7328
rect 3340 7204 3380 7244
rect 3340 6784 3380 6824
rect 3340 6532 3380 6572
rect 3244 6448 3284 6488
rect 2956 5608 2996 5648
rect 2860 5272 2900 5312
rect 2572 3844 2612 3884
rect 2476 3508 2516 3548
rect 2668 3760 2708 3800
rect 2572 3004 2612 3044
rect 3532 7120 3572 7160
rect 3532 6448 3572 6488
rect 4300 7204 4340 7244
rect 4972 9472 5012 9512
rect 5260 9472 5300 9512
rect 5548 10984 5588 11024
rect 5452 10312 5492 10352
rect 5356 8632 5396 8672
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 4876 8044 4916 8084
rect 4780 7540 4820 7580
rect 5260 7792 5300 7832
rect 6316 11992 6356 12032
rect 6220 11488 6260 11528
rect 6028 11404 6068 11444
rect 6124 11236 6164 11276
rect 6412 11236 6452 11276
rect 6316 10732 6356 10772
rect 6124 10648 6164 10688
rect 7084 18292 7124 18332
rect 6892 17956 6932 17996
rect 6892 17032 6932 17072
rect 6892 16780 6932 16820
rect 7084 17956 7124 17996
rect 7084 16108 7124 16148
rect 6700 15352 6740 15392
rect 6796 15184 6836 15224
rect 6700 14512 6740 14552
rect 6988 15352 7028 15392
rect 7084 13840 7124 13880
rect 6988 12580 7028 12620
rect 7084 12412 7124 12452
rect 7084 11908 7124 11948
rect 6988 11572 7028 11612
rect 6700 11236 6740 11276
rect 6604 10732 6644 10772
rect 6508 10564 6548 10604
rect 5548 10144 5588 10184
rect 5932 10144 5972 10184
rect 6412 10312 6452 10352
rect 6028 9892 6068 9932
rect 6316 9892 6356 9932
rect 5836 9640 5876 9680
rect 5548 8548 5588 8588
rect 5740 7876 5780 7916
rect 5452 7540 5492 7580
rect 6604 8632 6644 8672
rect 5932 8128 5972 8168
rect 6028 7792 6068 7832
rect 5740 7120 5780 7160
rect 5548 7036 5588 7076
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 4593 6700 4633 6740
rect 3820 6448 3860 6488
rect 3052 5104 3092 5144
rect 3052 4600 3092 4640
rect 3436 4768 3476 4808
rect 3244 4600 3284 4640
rect 3148 3928 3188 3968
rect 2956 3088 2996 3128
rect 2860 2584 2900 2624
rect 2380 2416 2420 2456
rect 2284 1408 2324 1448
rect 2476 1828 2516 1868
rect 2092 820 2132 860
rect 2284 736 2324 776
rect 2188 652 2228 692
rect 2668 400 2708 440
rect 3052 2752 3092 2792
rect 3436 4096 3476 4136
rect 3244 2836 3284 2876
rect 3148 1240 3188 1280
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 4492 6448 4532 6488
rect 4876 6532 4916 6572
rect 4396 6028 4436 6068
rect 4396 5692 4436 5732
rect 4588 5692 4628 5732
rect 5356 6028 5396 6068
rect 4780 5608 4820 5648
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 5164 4936 5204 4976
rect 4588 4852 4628 4892
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 3628 4264 3668 4304
rect 4588 3928 4628 3968
rect 3628 3676 3668 3716
rect 3532 3004 3572 3044
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 4204 3004 4244 3044
rect 3532 2836 3572 2876
rect 4204 2584 4244 2624
rect 4396 2332 4436 2372
rect 4204 1912 4244 1952
rect 3340 1660 3380 1700
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 2956 232 2996 272
rect 3916 1240 3956 1280
rect 3724 316 3764 356
rect 3532 232 3572 272
rect 4108 1156 4148 1196
rect 4300 1828 4340 1868
rect 4204 568 4244 608
rect 4492 2248 4532 2288
rect 4876 4852 4916 4892
rect 6124 7036 6164 7076
rect 7084 11236 7124 11276
rect 7084 10060 7124 10100
rect 7084 9220 7124 9260
rect 7276 18124 7316 18164
rect 7276 17032 7316 17072
rect 7660 19216 7700 19256
rect 7564 17956 7604 17996
rect 7660 17032 7700 17072
rect 7468 15940 7508 15980
rect 7372 15856 7412 15896
rect 7564 15604 7604 15644
rect 7660 15184 7700 15224
rect 7564 15100 7604 15140
rect 7372 14512 7412 14552
rect 7276 13168 7316 13208
rect 7276 11656 7316 11696
rect 6892 8632 6932 8672
rect 6700 8296 6740 8336
rect 6700 8128 6740 8168
rect 6604 7876 6644 7916
rect 6508 7792 6548 7832
rect 6604 7288 6644 7328
rect 6028 5692 6068 5732
rect 6316 5692 6356 5732
rect 6124 5272 6164 5312
rect 6028 5188 6068 5228
rect 5548 4852 5588 4892
rect 5740 4768 5780 4808
rect 5932 4600 5972 4640
rect 4876 3928 4916 3968
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 4972 3592 5012 3632
rect 4684 2584 4724 2624
rect 5068 3424 5108 3464
rect 5356 3592 5396 3632
rect 5164 3172 5204 3212
rect 5164 2920 5204 2960
rect 5740 3760 5780 3800
rect 6508 5692 6548 5732
rect 6604 5608 6644 5648
rect 6700 5104 6740 5144
rect 6220 5020 6260 5060
rect 6124 4012 6164 4052
rect 6412 4852 6452 4892
rect 6124 3760 6164 3800
rect 5644 3424 5684 3464
rect 6316 3760 6356 3800
rect 6220 3424 6260 3464
rect 5068 2668 5108 2708
rect 4972 2584 5012 2624
rect 5260 2584 5300 2624
rect 5164 2416 5204 2456
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 4972 1912 5012 1952
rect 5260 2080 5300 2120
rect 5452 2584 5492 2624
rect 5932 2584 5972 2624
rect 5548 2332 5588 2372
rect 5452 2248 5492 2288
rect 4492 1660 4532 1700
rect 4396 1492 4436 1532
rect 4684 1408 4724 1448
rect 4492 64 4532 104
rect 5356 1408 5396 1448
rect 5740 2248 5780 2288
rect 5548 1408 5588 1448
rect 6796 5020 6836 5060
rect 7180 8464 7220 8504
rect 7084 8296 7124 8336
rect 7468 13840 7508 13880
rect 7468 12412 7508 12452
rect 7468 12160 7508 12200
rect 7660 14848 7700 14888
rect 7660 12580 7700 12620
rect 7852 14764 7892 14804
rect 8140 17956 8180 17996
rect 8044 16360 8084 16400
rect 8044 15856 8084 15896
rect 8428 19972 8468 20012
rect 8332 19216 8372 19256
rect 8236 15856 8276 15896
rect 8044 15016 8084 15056
rect 8140 14848 8180 14888
rect 8044 13252 8084 13292
rect 7852 12916 7892 12956
rect 7948 12412 7988 12452
rect 8044 12244 8084 12284
rect 7948 11908 7988 11948
rect 7852 11656 7892 11696
rect 8140 11488 8180 11528
rect 7468 10648 7508 10688
rect 7372 10060 7412 10100
rect 7660 10144 7700 10184
rect 7372 9304 7412 9344
rect 7948 10480 7988 10520
rect 8812 23584 8852 23624
rect 8716 22912 8756 22952
rect 8908 22240 8948 22280
rect 9484 23752 9524 23792
rect 9484 23164 9524 23204
rect 8908 22072 8948 22112
rect 9388 22072 9428 22112
rect 8812 21232 8852 21272
rect 9388 21568 9428 21608
rect 9196 21484 9236 21524
rect 8716 20392 8756 20432
rect 8716 19972 8756 20012
rect 8524 17956 8564 17996
rect 8812 18796 8852 18836
rect 8812 18376 8852 18416
rect 8908 17788 8948 17828
rect 8524 17704 8564 17744
rect 8812 17620 8852 17660
rect 8716 17200 8756 17240
rect 8428 17116 8468 17156
rect 8428 16612 8468 16652
rect 8908 15940 8948 15980
rect 8428 15268 8468 15308
rect 8428 14848 8468 14888
rect 8716 14764 8756 14804
rect 8620 14008 8660 14048
rect 8428 13336 8468 13376
rect 8524 13168 8564 13208
rect 8332 12832 8372 12872
rect 8716 13924 8756 13964
rect 8620 11908 8660 11948
rect 8812 11824 8852 11864
rect 8332 10144 8372 10184
rect 8716 11488 8756 11528
rect 8620 9640 8660 9680
rect 7468 8548 7508 8588
rect 7276 7960 7316 8000
rect 7468 7960 7508 8000
rect 7660 9220 7700 9260
rect 7180 7792 7220 7832
rect 7084 7624 7124 7664
rect 6988 7036 7028 7076
rect 7468 6952 7508 6992
rect 6988 6448 7028 6488
rect 6988 5776 7028 5816
rect 7084 5692 7124 5732
rect 6988 5356 7028 5396
rect 6988 5188 7028 5228
rect 8140 9136 8180 9176
rect 8428 9136 8468 9176
rect 8332 8800 8372 8840
rect 8236 8632 8276 8672
rect 8620 9220 8660 9260
rect 8524 8464 8564 8504
rect 8044 8128 8084 8168
rect 7852 7960 7892 8000
rect 8044 7876 8084 7916
rect 8236 7036 8276 7076
rect 8812 9892 8852 9932
rect 8716 8212 8756 8252
rect 8332 6784 8372 6824
rect 8524 7540 8564 7580
rect 8908 7876 8948 7916
rect 9100 20056 9140 20096
rect 9100 19384 9140 19424
rect 9388 19552 9428 19592
rect 9196 18880 9236 18920
rect 9100 17536 9140 17576
rect 9100 17116 9140 17156
rect 9100 12580 9140 12620
rect 9100 9472 9140 9512
rect 9580 20728 9620 20768
rect 9580 20560 9620 20600
rect 9868 29632 9908 29672
rect 9964 29296 10004 29336
rect 9868 28288 9908 28328
rect 10156 34168 10196 34208
rect 10540 36520 10580 36560
rect 11020 36688 11060 36728
rect 10828 36604 10868 36644
rect 10540 36016 10580 36056
rect 10732 36016 10772 36056
rect 10636 35848 10676 35888
rect 10540 35680 10580 35720
rect 10732 35764 10772 35804
rect 11212 37024 11252 37064
rect 11596 37360 11636 37400
rect 11788 37192 11828 37232
rect 11596 36604 11636 36644
rect 11308 36436 11348 36476
rect 11308 36184 11348 36224
rect 10924 36016 10964 36056
rect 10828 35512 10868 35552
rect 10540 35092 10580 35132
rect 10444 35008 10484 35048
rect 10348 33580 10388 33620
rect 10636 34924 10676 34964
rect 10828 35008 10868 35048
rect 10732 34336 10772 34376
rect 11020 35932 11060 35972
rect 11020 35680 11060 35720
rect 10924 34504 10964 34544
rect 10444 33076 10484 33116
rect 10348 30892 10388 30932
rect 11116 35176 11156 35216
rect 11116 34924 11156 34964
rect 11116 34588 11156 34628
rect 10924 34084 10964 34124
rect 11308 35680 11348 35720
rect 11308 35512 11348 35552
rect 11596 35764 11636 35804
rect 11500 35680 11540 35720
rect 11788 36688 11828 36728
rect 13132 48700 13172 48740
rect 13228 48532 13268 48572
rect 13036 46432 13076 46472
rect 12844 44080 12884 44120
rect 13420 48784 13460 48824
rect 13804 48700 13844 48740
rect 13708 48616 13748 48656
rect 13612 48532 13652 48572
rect 13420 47860 13460 47900
rect 13324 46264 13364 46304
rect 13516 47272 13556 47312
rect 14380 59536 14420 59576
rect 14188 59368 14228 59408
rect 14092 58864 14132 58904
rect 14092 57940 14132 57980
rect 14092 55336 14132 55376
rect 14092 54832 14132 54872
rect 13996 53824 14036 53864
rect 13996 53488 14036 53528
rect 14860 61384 14900 61424
rect 14956 61300 14996 61340
rect 14764 61216 14804 61256
rect 14956 61132 14996 61172
rect 14764 60040 14804 60080
rect 14668 59956 14708 59996
rect 14476 57772 14516 57812
rect 14284 57268 14324 57308
rect 14380 57184 14420 57224
rect 14284 57100 14324 57140
rect 14284 56596 14324 56636
rect 13996 53152 14036 53192
rect 13996 52648 14036 52688
rect 14764 57520 14804 57560
rect 14956 59284 14996 59324
rect 14860 57184 14900 57224
rect 14860 57016 14900 57056
rect 14668 56680 14708 56720
rect 14572 56596 14612 56636
rect 14476 56344 14516 56384
rect 14380 55924 14420 55964
rect 14380 55672 14420 55712
rect 14668 55924 14708 55964
rect 14380 54916 14420 54956
rect 14860 55840 14900 55880
rect 15724 64324 15764 64364
rect 15724 64072 15764 64112
rect 15724 63904 15764 63944
rect 15340 63820 15380 63860
rect 15244 62728 15284 62768
rect 16204 64408 16244 64448
rect 16012 64156 16052 64196
rect 15916 64072 15956 64112
rect 15916 63904 15956 63944
rect 15340 62224 15380 62264
rect 15244 61804 15284 61844
rect 15532 62392 15572 62432
rect 15244 61300 15284 61340
rect 16204 63820 16244 63860
rect 16780 65332 16820 65372
rect 16396 65248 16436 65288
rect 16684 65080 16724 65120
rect 17548 69700 17588 69740
rect 17740 69700 17780 69740
rect 18028 70036 18068 70076
rect 17932 69868 17972 69908
rect 17644 69364 17684 69404
rect 17644 69196 17684 69236
rect 17548 68188 17588 68228
rect 17836 69364 17876 69404
rect 17740 67600 17780 67640
rect 17644 67516 17684 67556
rect 17356 66676 17396 66716
rect 17548 66760 17588 66800
rect 18220 69784 18260 69824
rect 18028 68104 18068 68144
rect 18028 67936 18068 67976
rect 18604 71632 18644 71672
rect 18604 70624 18644 70664
rect 18412 69280 18452 69320
rect 20044 82552 20084 82592
rect 20048 82384 20088 82424
rect 20130 82384 20170 82424
rect 20212 82384 20252 82424
rect 20294 82384 20334 82424
rect 20376 82384 20416 82424
rect 19660 82048 19700 82088
rect 18796 81964 18836 82004
rect 19276 81880 19316 81920
rect 18808 81628 18848 81668
rect 18890 81628 18930 81668
rect 18972 81628 19012 81668
rect 19054 81628 19094 81668
rect 19136 81628 19176 81668
rect 20048 80872 20088 80912
rect 20130 80872 20170 80912
rect 20212 80872 20252 80912
rect 20294 80872 20334 80912
rect 20376 80872 20416 80912
rect 18808 80116 18848 80156
rect 18890 80116 18930 80156
rect 18972 80116 19012 80156
rect 19054 80116 19094 80156
rect 19136 80116 19176 80156
rect 20048 79360 20088 79400
rect 20130 79360 20170 79400
rect 20212 79360 20252 79400
rect 20294 79360 20334 79400
rect 20376 79360 20416 79400
rect 18808 78604 18848 78644
rect 18890 78604 18930 78644
rect 18972 78604 19012 78644
rect 19054 78604 19094 78644
rect 19136 78604 19176 78644
rect 20812 78520 20852 78560
rect 20048 77848 20088 77888
rect 20130 77848 20170 77888
rect 20212 77848 20252 77888
rect 20294 77848 20334 77888
rect 20376 77848 20416 77888
rect 18808 77092 18848 77132
rect 18890 77092 18930 77132
rect 18972 77092 19012 77132
rect 19054 77092 19094 77132
rect 19136 77092 19176 77132
rect 20524 76504 20564 76544
rect 20048 76336 20088 76376
rect 20130 76336 20170 76376
rect 20212 76336 20252 76376
rect 20294 76336 20334 76376
rect 20376 76336 20416 76376
rect 18808 75580 18848 75620
rect 18890 75580 18930 75620
rect 18972 75580 19012 75620
rect 19054 75580 19094 75620
rect 19136 75580 19176 75620
rect 20048 74824 20088 74864
rect 20130 74824 20170 74864
rect 20212 74824 20252 74864
rect 20294 74824 20334 74864
rect 20376 74824 20416 74864
rect 18808 74068 18848 74108
rect 18890 74068 18930 74108
rect 18972 74068 19012 74108
rect 19054 74068 19094 74108
rect 19136 74068 19176 74108
rect 20048 73312 20088 73352
rect 20130 73312 20170 73352
rect 20212 73312 20252 73352
rect 20294 73312 20334 73352
rect 20376 73312 20416 73352
rect 18808 72556 18848 72596
rect 18890 72556 18930 72596
rect 18972 72556 19012 72596
rect 19054 72556 19094 72596
rect 19136 72556 19176 72596
rect 20048 71800 20088 71840
rect 20130 71800 20170 71840
rect 20212 71800 20252 71840
rect 20294 71800 20334 71840
rect 20376 71800 20416 71840
rect 18796 71632 18836 71672
rect 19372 71464 19412 71504
rect 18808 71044 18848 71084
rect 18890 71044 18930 71084
rect 18972 71044 19012 71084
rect 19054 71044 19094 71084
rect 19136 71044 19176 71084
rect 19372 70792 19412 70832
rect 18892 70624 18932 70664
rect 18796 70456 18836 70496
rect 18700 70120 18740 70160
rect 18700 69952 18740 69992
rect 18988 70036 19028 70076
rect 19084 69952 19124 69992
rect 19468 70624 19508 70664
rect 19372 70036 19412 70076
rect 18988 69784 19028 69824
rect 19756 70456 19796 70496
rect 20044 70540 20084 70580
rect 20048 70288 20088 70328
rect 20130 70288 20170 70328
rect 20212 70288 20252 70328
rect 20294 70288 20334 70328
rect 20376 70288 20416 70328
rect 20044 70036 20084 70076
rect 19084 69700 19124 69740
rect 19276 69616 19316 69656
rect 18808 69532 18848 69572
rect 18890 69532 18930 69572
rect 18972 69532 19012 69572
rect 19054 69532 19094 69572
rect 19136 69532 19176 69572
rect 18700 69364 18740 69404
rect 18892 69364 18932 69404
rect 19276 69364 19316 69404
rect 18604 69196 18644 69236
rect 18316 68944 18356 68984
rect 18988 69196 19028 69236
rect 20236 69952 20276 69992
rect 19372 69112 19412 69152
rect 19180 69028 19220 69068
rect 19276 68944 19316 68984
rect 19660 69616 19700 69656
rect 19852 69448 19892 69488
rect 19948 69280 19988 69320
rect 19756 69112 19796 69152
rect 18796 68776 18836 68816
rect 20048 68776 20088 68816
rect 20130 68776 20170 68816
rect 20212 68776 20252 68816
rect 20294 68776 20334 68816
rect 20376 68776 20416 68816
rect 18700 68440 18740 68480
rect 18412 68188 18452 68228
rect 18892 68188 18932 68228
rect 19276 68440 19316 68480
rect 18604 68104 18644 68144
rect 18220 68020 18260 68060
rect 17932 66760 17972 66800
rect 17452 66172 17492 66212
rect 17260 66088 17300 66128
rect 17452 65500 17492 65540
rect 17932 65500 17972 65540
rect 16780 64072 16820 64112
rect 16396 63904 16436 63944
rect 16492 63736 16532 63776
rect 16012 62392 16052 62432
rect 16012 62140 16052 62180
rect 15820 61720 15860 61760
rect 15724 61636 15764 61676
rect 15820 61552 15860 61592
rect 15436 61468 15476 61508
rect 15436 61300 15476 61340
rect 15724 61384 15764 61424
rect 15628 61300 15668 61340
rect 15340 61132 15380 61172
rect 15916 61216 15956 61256
rect 15628 61048 15668 61088
rect 15244 59200 15284 59240
rect 15148 58528 15188 58568
rect 15628 60544 15668 60584
rect 15532 58696 15572 58736
rect 15436 58612 15476 58652
rect 16012 61048 16052 61088
rect 16300 63316 16340 63356
rect 16492 63064 16532 63104
rect 16396 62728 16436 62768
rect 15820 60880 15860 60920
rect 15820 60628 15860 60668
rect 15820 59872 15860 59912
rect 16012 58948 16052 58988
rect 16780 63736 16820 63776
rect 16588 62560 16628 62600
rect 16492 62140 16532 62180
rect 16396 60880 16436 60920
rect 16300 60208 16340 60248
rect 16300 59368 16340 59408
rect 16108 58780 16148 58820
rect 16012 58612 16052 58652
rect 16108 58528 16148 58568
rect 16300 58528 16340 58568
rect 15340 57772 15380 57812
rect 16012 57856 16052 57896
rect 15916 57520 15956 57560
rect 15340 57352 15380 57392
rect 15052 56260 15092 56300
rect 15244 56176 15284 56216
rect 14764 54916 14804 54956
rect 15052 55084 15092 55124
rect 15148 54748 15188 54788
rect 15052 54496 15092 54536
rect 15052 54160 15092 54200
rect 14764 53824 14804 53864
rect 14380 53488 14420 53528
rect 14188 51808 14228 51848
rect 13996 50968 14036 51008
rect 13996 50380 14036 50420
rect 13996 49624 14036 49664
rect 13996 48784 14036 48824
rect 14284 50968 14324 51008
rect 14188 47776 14228 47816
rect 13996 47188 14036 47228
rect 13612 46516 13652 46556
rect 13708 46348 13748 46388
rect 13324 45340 13364 45380
rect 13324 44920 13364 44960
rect 13324 43576 13364 43616
rect 13516 44584 13556 44624
rect 13804 44920 13844 44960
rect 13708 44584 13748 44624
rect 13708 44248 13748 44288
rect 13900 44668 13940 44708
rect 13996 44248 14036 44288
rect 12940 41896 12980 41936
rect 12556 41728 12596 41768
rect 12940 41392 12980 41432
rect 12364 41224 12404 41264
rect 13228 40636 13268 40676
rect 13036 40468 13076 40508
rect 12748 40300 12788 40340
rect 12844 39544 12884 39584
rect 12748 39208 12788 39248
rect 12940 38956 12980 38996
rect 12748 37948 12788 37988
rect 12652 37696 12692 37736
rect 12172 37444 12212 37484
rect 12172 37276 12212 37316
rect 12076 36940 12116 36980
rect 12556 37360 12596 37400
rect 12268 36856 12308 36896
rect 11788 35848 11828 35888
rect 12268 36100 12308 36140
rect 12076 35848 12116 35888
rect 12652 37024 12692 37064
rect 13228 39544 13268 39584
rect 13132 38956 13172 38996
rect 13036 38200 13076 38240
rect 13420 38872 13460 38912
rect 12940 37948 12980 37988
rect 13804 43576 13844 43616
rect 13900 43408 13940 43448
rect 13516 38200 13556 38240
rect 13132 37864 13172 37904
rect 13324 37864 13364 37904
rect 13516 37864 13556 37904
rect 13036 37276 13076 37316
rect 12844 37192 12884 37232
rect 13036 36856 13076 36896
rect 12844 36772 12884 36812
rect 12940 36688 12980 36728
rect 12748 36604 12788 36644
rect 12460 36520 12500 36560
rect 12844 36100 12884 36140
rect 12652 36016 12692 36056
rect 11788 35596 11828 35636
rect 11212 33832 11252 33872
rect 11212 33664 11252 33704
rect 11404 35176 11444 35216
rect 11500 35092 11540 35132
rect 11404 35008 11444 35048
rect 11500 34924 11540 34964
rect 11404 33664 11444 33704
rect 11884 35260 11924 35300
rect 11596 34504 11636 34544
rect 11596 34336 11636 34376
rect 11788 35176 11828 35216
rect 12076 35176 12116 35216
rect 12556 35848 12596 35888
rect 12940 35932 12980 35972
rect 12748 35680 12788 35720
rect 13612 37612 13652 37652
rect 13324 37024 13364 37064
rect 13228 36856 13268 36896
rect 13900 38200 13940 38240
rect 13900 37864 13940 37904
rect 13804 37024 13844 37064
rect 14188 45088 14228 45128
rect 14188 44248 14228 44288
rect 14572 53404 14612 53444
rect 14476 50800 14516 50840
rect 14476 50296 14516 50336
rect 14572 49624 14612 49664
rect 14572 49120 14612 49160
rect 14572 48532 14612 48572
rect 14476 47944 14516 47984
rect 14476 47776 14516 47816
rect 15148 52984 15188 53024
rect 14764 51808 14804 51848
rect 15244 51808 15284 51848
rect 15148 51052 15188 51092
rect 15244 50968 15284 51008
rect 14956 50800 14996 50840
rect 14764 49708 14804 49748
rect 15628 56428 15668 56468
rect 15532 56260 15572 56300
rect 15532 54832 15572 54872
rect 15916 56260 15956 56300
rect 15820 55504 15860 55544
rect 15532 54412 15572 54452
rect 15820 53992 15860 54032
rect 15436 50380 15476 50420
rect 15052 49540 15092 49580
rect 15148 49372 15188 49412
rect 14860 47944 14900 47984
rect 14668 46264 14708 46304
rect 14668 44920 14708 44960
rect 14572 40636 14612 40676
rect 14572 39544 14612 39584
rect 14476 39208 14516 39248
rect 14380 39040 14420 39080
rect 14092 38200 14132 38240
rect 14188 37948 14228 37988
rect 14668 38704 14708 38744
rect 15724 53320 15764 53360
rect 15628 53236 15668 53276
rect 15820 53068 15860 53108
rect 16012 55420 16052 55460
rect 16588 61048 16628 61088
rect 16684 60880 16724 60920
rect 16588 59452 16628 59492
rect 16588 58780 16628 58820
rect 16396 57604 16436 57644
rect 16300 57268 16340 57308
rect 16972 63652 17012 63692
rect 16972 60880 17012 60920
rect 17836 65248 17876 65288
rect 17452 64408 17492 64448
rect 17932 64408 17972 64448
rect 17351 63904 17391 63944
rect 18220 65416 18260 65456
rect 18028 64324 18068 64364
rect 17644 63988 17684 64028
rect 18604 65332 18644 65372
rect 18412 64912 18452 64952
rect 17548 63316 17588 63356
rect 18028 63736 18068 63776
rect 17932 63316 17972 63356
rect 17932 63064 17972 63104
rect 17452 61384 17492 61424
rect 17164 61300 17204 61340
rect 16876 59200 16916 59240
rect 16780 58192 16820 58232
rect 16876 57520 16916 57560
rect 16300 56344 16340 56384
rect 16492 56344 16532 56384
rect 16300 55588 16340 55628
rect 16876 57016 16916 57056
rect 16876 56512 16916 56552
rect 17260 59368 17300 59408
rect 17356 59116 17396 59156
rect 17644 60880 17684 60920
rect 17548 60544 17588 60584
rect 17644 60460 17684 60500
rect 17836 60628 17876 60668
rect 17740 60376 17780 60416
rect 17548 59368 17588 59408
rect 17740 59284 17780 59324
rect 17644 59200 17684 59240
rect 17644 57856 17684 57896
rect 17164 57604 17204 57644
rect 17260 56932 17300 56972
rect 17068 56680 17108 56720
rect 16588 55924 16628 55964
rect 16972 55924 17012 55964
rect 16108 54748 16148 54788
rect 16396 55168 16436 55208
rect 16300 55000 16340 55040
rect 16300 53320 16340 53360
rect 16204 52564 16244 52604
rect 15724 52312 15764 52352
rect 16012 52312 16052 52352
rect 15820 51808 15860 51848
rect 15628 51724 15668 51764
rect 15532 49540 15572 49580
rect 15436 49372 15476 49412
rect 15820 51052 15860 51092
rect 16012 51976 16052 52016
rect 15916 50968 15956 51008
rect 16204 51976 16244 52016
rect 16204 51724 16244 51764
rect 16204 51052 16244 51092
rect 15820 50044 15860 50084
rect 16012 50212 16052 50252
rect 15916 49540 15956 49580
rect 15724 49456 15764 49496
rect 14860 46264 14900 46304
rect 15244 46768 15284 46808
rect 15244 45760 15284 45800
rect 15244 44920 15284 44960
rect 15052 43828 15092 43868
rect 14860 42316 14900 42356
rect 15244 44248 15284 44288
rect 15148 39460 15188 39500
rect 14860 39208 14900 39248
rect 14476 37780 14516 37820
rect 14380 37528 14420 37568
rect 13996 36688 14036 36728
rect 13900 36604 13940 36644
rect 13324 36268 13364 36308
rect 13228 36016 13268 36056
rect 13708 36268 13748 36308
rect 13228 35680 13268 35720
rect 13228 35428 13268 35468
rect 13420 35848 13460 35888
rect 12748 35260 12788 35300
rect 12172 35092 12212 35132
rect 12556 35092 12596 35132
rect 11980 34504 12020 34544
rect 11692 34084 11732 34124
rect 11884 34084 11924 34124
rect 11692 33916 11732 33956
rect 11788 33832 11828 33872
rect 10636 31396 10676 31436
rect 10636 31228 10676 31268
rect 10540 30976 10580 31016
rect 10444 30724 10484 30764
rect 10348 30556 10388 30596
rect 10444 29968 10484 30008
rect 10540 29800 10580 29840
rect 10828 30640 10868 30680
rect 10732 30556 10772 30596
rect 11020 31984 11060 32024
rect 11212 32320 11252 32360
rect 11692 33328 11732 33368
rect 11500 31564 11540 31604
rect 11212 31312 11252 31352
rect 11404 31480 11444 31520
rect 11308 31144 11348 31184
rect 10924 30472 10964 30512
rect 10540 29632 10580 29672
rect 10252 29380 10292 29420
rect 10540 29380 10580 29420
rect 10156 29128 10196 29168
rect 10156 28120 10196 28160
rect 10348 28540 10388 28580
rect 10636 29296 10676 29336
rect 10924 30136 10964 30176
rect 10924 29800 10964 29840
rect 11212 30892 11252 30932
rect 11212 30724 11252 30764
rect 11308 30556 11348 30596
rect 11500 30472 11540 30512
rect 11116 29968 11156 30008
rect 11116 29464 11156 29504
rect 11020 29212 11060 29252
rect 10924 29128 10964 29168
rect 10828 28960 10868 29000
rect 10636 28876 10676 28916
rect 9772 26860 9812 26900
rect 9964 27112 10004 27152
rect 10156 27448 10196 27488
rect 10060 26860 10100 26900
rect 10252 27196 10292 27236
rect 9964 26272 10004 26312
rect 10060 26020 10100 26060
rect 9772 25264 9812 25304
rect 9964 25768 10004 25808
rect 9868 24760 9908 24800
rect 9868 24592 9908 24632
rect 9868 22912 9908 22952
rect 9772 22408 9812 22448
rect 9868 21316 9908 21356
rect 10060 23080 10100 23120
rect 10348 26692 10388 26732
rect 10252 26524 10292 26564
rect 10540 27616 10580 27656
rect 11596 29968 11636 30008
rect 11596 29464 11636 29504
rect 11308 29044 11348 29084
rect 11692 29128 11732 29168
rect 11500 28624 11540 28664
rect 11212 28540 11252 28580
rect 11116 28120 11156 28160
rect 10732 27448 10772 27488
rect 10636 26776 10676 26816
rect 10252 25768 10292 25808
rect 10252 25264 10292 25304
rect 9964 20560 10004 20600
rect 9868 20308 9908 20348
rect 9580 18544 9620 18584
rect 9484 18208 9524 18248
rect 9676 18040 9716 18080
rect 9292 17620 9332 17660
rect 9676 17620 9716 17660
rect 9388 17116 9428 17156
rect 9484 17032 9524 17072
rect 9484 16528 9524 16568
rect 10540 24340 10580 24380
rect 11020 27700 11060 27740
rect 10924 27532 10964 27572
rect 10924 27280 10964 27320
rect 11308 27196 11348 27236
rect 10828 26776 10868 26816
rect 10828 26608 10868 26648
rect 11116 26860 11156 26900
rect 11500 26944 11540 26984
rect 11884 33664 11924 33704
rect 11884 31564 11924 31604
rect 12076 34420 12116 34460
rect 12076 33664 12116 33704
rect 12652 35008 12692 35048
rect 12556 34420 12596 34460
rect 12460 34336 12500 34376
rect 12268 34000 12308 34040
rect 12172 33412 12212 33452
rect 12172 33244 12212 33284
rect 12076 32824 12116 32864
rect 12076 32320 12116 32360
rect 11980 30724 12020 30764
rect 13324 35344 13364 35384
rect 13516 35344 13556 35384
rect 13420 35260 13460 35300
rect 13036 35176 13076 35216
rect 13132 35092 13172 35132
rect 12940 35008 12980 35048
rect 13516 35008 13556 35048
rect 13420 34924 13460 34964
rect 13324 34840 13364 34880
rect 12940 34504 12980 34544
rect 13036 34420 13076 34460
rect 12844 34168 12884 34208
rect 12940 34084 12980 34124
rect 12748 34000 12788 34040
rect 12748 33832 12788 33872
rect 12556 33412 12596 33452
rect 12268 32656 12308 32696
rect 12172 30892 12212 30932
rect 11884 29632 11924 29672
rect 11980 29296 12020 29336
rect 12172 29464 12212 29504
rect 12172 29296 12212 29336
rect 12076 29128 12116 29168
rect 12460 32320 12500 32360
rect 12364 32152 12404 32192
rect 12460 30724 12500 30764
rect 12364 30640 12404 30680
rect 12460 29884 12500 29924
rect 12364 29632 12404 29672
rect 12268 28960 12308 29000
rect 11980 28876 12020 28916
rect 11884 28540 11924 28580
rect 11788 28120 11828 28160
rect 11884 27868 11924 27908
rect 11692 27448 11732 27488
rect 11596 26776 11636 26816
rect 11020 26524 11060 26564
rect 11404 26524 11444 26564
rect 11212 26272 11252 26312
rect 11500 26188 11540 26228
rect 11404 25432 11444 25472
rect 10924 25264 10964 25304
rect 11116 24760 11156 24800
rect 11116 24340 11156 24380
rect 10444 23164 10484 23204
rect 10444 22660 10484 22700
rect 10444 21652 10484 21692
rect 10156 19804 10196 19844
rect 10348 21148 10388 21188
rect 10732 23668 10772 23708
rect 10636 21064 10676 21104
rect 10636 20476 10676 20516
rect 10828 21232 10868 21272
rect 11596 24676 11636 24716
rect 11308 24256 11348 24296
rect 11212 23752 11252 23792
rect 11308 23668 11348 23708
rect 11788 27364 11828 27404
rect 12076 28624 12116 28664
rect 12172 28540 12212 28580
rect 11980 26944 12020 26984
rect 12172 27616 12212 27656
rect 12460 27868 12500 27908
rect 12268 27448 12308 27488
rect 12364 27364 12404 27404
rect 12172 26944 12212 26984
rect 11980 25936 12020 25976
rect 11884 24928 11924 24968
rect 11692 24172 11732 24212
rect 11692 23920 11732 23960
rect 12460 26944 12500 26984
rect 12268 26440 12308 26480
rect 12364 26188 12404 26228
rect 12364 24340 12404 24380
rect 12460 24088 12500 24128
rect 13228 34504 13268 34544
rect 13516 34168 13556 34208
rect 13420 33832 13460 33872
rect 13804 35428 13844 35468
rect 13708 34840 13748 34880
rect 14188 35848 14228 35888
rect 14476 35932 14516 35972
rect 14092 35008 14132 35048
rect 14284 35176 14324 35216
rect 14188 34924 14228 34964
rect 13804 34504 13844 34544
rect 14188 34504 14228 34544
rect 13708 34336 13748 34376
rect 13804 34168 13844 34208
rect 13708 34000 13748 34040
rect 13420 33664 13460 33704
rect 13228 32824 13268 32864
rect 13612 33664 13652 33704
rect 13900 34000 13940 34040
rect 14003 34000 14043 34040
rect 13516 33412 13556 33452
rect 13516 33244 13556 33284
rect 13420 32992 13460 33032
rect 13900 33412 13940 33452
rect 13132 32740 13172 32780
rect 14476 35008 14516 35048
rect 14380 34588 14420 34628
rect 14572 34420 14612 34460
rect 14380 34168 14420 34208
rect 14572 34168 14612 34208
rect 14092 33412 14132 33452
rect 13996 33244 14036 33284
rect 13996 33076 14036 33116
rect 14188 32992 14228 33032
rect 15244 39040 15284 39080
rect 15052 37948 15092 37988
rect 14860 35848 14900 35888
rect 14764 35176 14804 35216
rect 14764 34000 14804 34040
rect 14476 33664 14516 33704
rect 13996 32824 14036 32864
rect 12652 32236 12692 32276
rect 13516 32236 13556 32276
rect 12844 32152 12884 32192
rect 13036 32152 13076 32192
rect 12940 31564 12980 31604
rect 12748 31480 12788 31520
rect 12940 31144 12980 31184
rect 12748 31060 12788 31100
rect 13420 32152 13460 32192
rect 13228 31564 13268 31604
rect 12748 30472 12788 30512
rect 13228 31144 13268 31184
rect 13324 31060 13364 31100
rect 13228 30724 13268 30764
rect 13132 30472 13172 30512
rect 13132 29716 13172 29756
rect 13036 29632 13076 29672
rect 12748 28540 12788 28580
rect 12652 28372 12692 28412
rect 12748 28288 12788 28328
rect 12652 24592 12692 24632
rect 13132 29464 13172 29504
rect 13516 31312 13556 31352
rect 13420 30724 13460 30764
rect 13804 30640 13844 30680
rect 13708 30052 13748 30092
rect 13612 29296 13652 29336
rect 13228 28540 13268 28580
rect 13228 27616 13268 27656
rect 11500 23752 11540 23792
rect 11884 23752 11924 23792
rect 12076 23752 12116 23792
rect 12076 23248 12116 23288
rect 11500 23164 11540 23204
rect 11692 23080 11732 23120
rect 11596 22240 11636 22280
rect 11788 22492 11828 22532
rect 12076 22912 12116 22952
rect 11980 22660 12020 22700
rect 11884 22324 11924 22364
rect 12172 22408 12212 22448
rect 12076 22324 12116 22364
rect 12172 22156 12212 22196
rect 11308 21652 11348 21692
rect 11404 21484 11444 21524
rect 11308 21064 11348 21104
rect 10828 20560 10868 20600
rect 10252 19636 10292 19676
rect 10060 18460 10100 18500
rect 9964 18208 10004 18248
rect 10156 17956 10196 17996
rect 10348 19048 10388 19088
rect 10060 17872 10100 17912
rect 10252 17788 10292 17828
rect 10156 17704 10196 17744
rect 9676 16444 9716 16484
rect 9388 16108 9428 16148
rect 9292 14680 9332 14720
rect 9868 16276 9908 16316
rect 9772 16192 9812 16232
rect 10060 16192 10100 16232
rect 9964 15184 10004 15224
rect 9292 14176 9332 14216
rect 9484 14092 9524 14132
rect 9580 13840 9620 13880
rect 9388 13756 9428 13796
rect 9004 7540 9044 7580
rect 8620 7036 8660 7076
rect 8716 6616 8756 6656
rect 8044 6196 8084 6236
rect 8428 6196 8468 6236
rect 8524 5944 8564 5984
rect 6700 2332 6740 2372
rect 6604 2164 6644 2204
rect 7084 4516 7124 4556
rect 6892 4432 6932 4472
rect 7660 5020 7700 5060
rect 7756 4936 7796 4976
rect 7372 4684 7412 4724
rect 7852 4600 7892 4640
rect 7756 4516 7796 4556
rect 7468 4432 7508 4472
rect 7468 3508 7508 3548
rect 7660 3928 7700 3968
rect 8236 3928 8276 3968
rect 8428 5188 8468 5228
rect 8236 3592 8276 3632
rect 7756 3508 7796 3548
rect 7660 3340 7700 3380
rect 6988 2080 7028 2120
rect 7564 3256 7604 3296
rect 8140 3424 8180 3464
rect 7852 3172 7892 3212
rect 8044 3172 8084 3212
rect 6220 1324 6260 1364
rect 6124 1156 6164 1196
rect 6220 1072 6260 1112
rect 5932 904 5972 944
rect 5836 820 5876 860
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 4876 568 4916 608
rect 5068 568 5108 608
rect 5452 484 5492 524
rect 5260 148 5300 188
rect 5644 400 5684 440
rect 6028 232 6068 272
rect 6412 988 6452 1028
rect 6316 904 6356 944
rect 6412 736 6452 776
rect 6508 568 6548 608
rect 6796 1408 6836 1448
rect 8428 2752 8468 2792
rect 7852 1828 7892 1868
rect 8236 1828 8276 1868
rect 7852 1408 7892 1448
rect 7180 1324 7220 1364
rect 6700 1240 6740 1280
rect 7372 1240 7412 1280
rect 7756 1240 7796 1280
rect 6796 904 6836 944
rect 6604 400 6644 440
rect 6604 148 6644 188
rect 7180 1156 7220 1196
rect 6988 736 7028 776
rect 6892 400 6932 440
rect 7756 988 7796 1028
rect 7372 568 7412 608
rect 7564 568 7604 608
rect 7564 400 7604 440
rect 8044 1324 8084 1364
rect 7948 1156 7988 1196
rect 8428 1492 8468 1532
rect 8620 4600 8660 4640
rect 8620 4012 8660 4052
rect 8620 3424 8660 3464
rect 8908 6868 8948 6908
rect 9004 6532 9044 6572
rect 8812 4852 8852 4892
rect 9196 7876 9236 7916
rect 9196 7120 9236 7160
rect 9196 6532 9236 6572
rect 8812 1828 8852 1868
rect 8140 1240 8180 1280
rect 8524 1156 8564 1196
rect 8140 568 8180 608
rect 8716 1240 8756 1280
rect 8620 652 8660 692
rect 9004 1660 9044 1700
rect 9004 1156 9044 1196
rect 8812 820 8852 860
rect 9196 1492 9236 1532
rect 9484 12244 9524 12284
rect 9388 11572 9428 11612
rect 9772 13084 9812 13124
rect 10636 19804 10676 19844
rect 10924 18796 10964 18836
rect 11404 20056 11444 20096
rect 11212 19468 11252 19508
rect 11212 19132 11252 19172
rect 11116 18796 11156 18836
rect 11020 18712 11060 18752
rect 10636 18544 10676 18584
rect 11212 18628 11252 18668
rect 10540 17788 10580 17828
rect 10540 17368 10580 17408
rect 10156 15940 10196 15980
rect 10060 14932 10100 14972
rect 10348 16192 10388 16232
rect 10732 18208 10772 18248
rect 10252 13756 10292 13796
rect 9964 12580 10004 12620
rect 9868 11824 9908 11864
rect 9676 11320 9716 11360
rect 9388 7036 9428 7076
rect 9388 2752 9428 2792
rect 9388 2332 9428 2372
rect 9580 8548 9620 8588
rect 9580 7960 9620 8000
rect 9868 11152 9908 11192
rect 10444 14932 10484 14972
rect 10924 17116 10964 17156
rect 11596 18460 11636 18500
rect 11596 18124 11636 18164
rect 11404 17788 11444 17828
rect 11212 17368 11252 17408
rect 11020 16864 11060 16904
rect 11308 17116 11348 17156
rect 11596 17704 11636 17744
rect 11500 17452 11540 17492
rect 11500 17200 11540 17240
rect 11020 16024 11060 16064
rect 11020 14680 11060 14720
rect 10732 12580 10772 12620
rect 11020 13189 11060 13217
rect 11020 13177 11060 13189
rect 11692 15436 11732 15476
rect 12076 21484 12116 21524
rect 11884 19972 11924 20012
rect 12748 23920 12788 23960
rect 12364 23836 12404 23876
rect 12364 23080 12404 23120
rect 12652 23752 12692 23792
rect 13900 29800 13940 29840
rect 13420 27448 13460 27488
rect 13420 26944 13460 26984
rect 13516 26608 13556 26648
rect 13132 25852 13172 25892
rect 13708 24088 13748 24128
rect 13132 23920 13172 23960
rect 13516 23836 13556 23876
rect 12556 23416 12596 23456
rect 12556 23248 12596 23288
rect 12268 20728 12308 20768
rect 12556 22072 12596 22112
rect 12460 21736 12500 21776
rect 12652 21652 12692 21692
rect 12844 23248 12884 23288
rect 12940 22996 12980 23036
rect 13132 23584 13172 23624
rect 13516 23584 13556 23624
rect 13420 23164 13460 23204
rect 13132 22660 13172 22700
rect 13132 22408 13172 22448
rect 13036 22240 13076 22280
rect 12844 22156 12884 22196
rect 13324 22240 13364 22280
rect 13228 22156 13268 22196
rect 13132 21904 13172 21944
rect 12556 21400 12596 21440
rect 12748 21568 12788 21608
rect 12844 21400 12884 21440
rect 12652 20728 12692 20768
rect 12268 20140 12308 20180
rect 12268 19972 12308 20012
rect 12172 19888 12212 19928
rect 11884 15520 11924 15560
rect 10924 12076 10964 12116
rect 10540 11656 10580 11696
rect 10444 11488 10484 11528
rect 10828 11404 10868 11444
rect 10156 11152 10196 11192
rect 10252 11068 10292 11108
rect 10156 10984 10196 11024
rect 10060 10900 10100 10940
rect 9964 10144 10004 10184
rect 9772 9556 9812 9596
rect 9868 9472 9908 9512
rect 10060 8800 10100 8840
rect 9964 8632 10004 8672
rect 10156 8716 10196 8756
rect 10636 11068 10676 11108
rect 10444 10984 10484 11024
rect 10732 10816 10772 10856
rect 10348 10144 10388 10184
rect 10348 9640 10388 9680
rect 10540 10312 10580 10352
rect 10540 10144 10580 10184
rect 10348 9136 10388 9176
rect 10503 8716 10543 8756
rect 10060 8464 10100 8504
rect 10060 8212 10100 8252
rect 9676 7876 9716 7916
rect 9772 7036 9812 7076
rect 10348 8464 10388 8504
rect 10252 7456 10292 7496
rect 10252 6868 10292 6908
rect 10156 5860 10196 5900
rect 9868 5608 9908 5648
rect 9772 5104 9812 5144
rect 9676 4600 9716 4640
rect 9964 5524 10004 5564
rect 9772 4096 9812 4136
rect 10252 5608 10292 5648
rect 10732 10396 10772 10436
rect 10828 9640 10868 9680
rect 10444 8212 10484 8252
rect 10444 7036 10484 7076
rect 10924 8548 10964 8588
rect 10924 8296 10964 8336
rect 11212 12076 11252 12116
rect 11212 11824 11252 11864
rect 11308 11404 11348 11444
rect 11212 11320 11252 11360
rect 11116 10144 11156 10184
rect 11020 8128 11060 8168
rect 10924 7876 10964 7916
rect 11692 14512 11732 14552
rect 11692 11320 11732 11360
rect 11500 11236 11540 11276
rect 11692 11152 11732 11192
rect 11500 11068 11540 11108
rect 11404 10984 11444 11024
rect 11404 10144 11444 10184
rect 11308 10060 11348 10100
rect 11212 8716 11252 8756
rect 11116 7540 11156 7580
rect 11020 7456 11060 7496
rect 11404 8128 11444 8168
rect 11297 7456 11337 7496
rect 11212 7288 11252 7328
rect 11404 7288 11444 7328
rect 10924 7036 10964 7076
rect 11212 7036 11252 7076
rect 10636 6700 10676 6740
rect 10732 6448 10772 6488
rect 11116 6616 11156 6656
rect 10924 6448 10964 6488
rect 11500 7204 11540 7244
rect 12172 17704 12212 17744
rect 12364 19888 12404 19928
rect 12652 20140 12692 20180
rect 12556 19804 12596 19844
rect 12556 19132 12596 19172
rect 12460 18964 12500 19004
rect 12748 18880 12788 18920
rect 12652 18796 12692 18836
rect 12364 16780 12404 16820
rect 12748 18628 12788 18668
rect 12748 18124 12788 18164
rect 12652 18040 12692 18080
rect 12556 17956 12596 17996
rect 12268 15772 12308 15812
rect 12076 15436 12116 15476
rect 12172 14764 12212 14804
rect 12076 10732 12116 10772
rect 11980 10648 12020 10688
rect 11884 10564 11924 10604
rect 12076 10564 12116 10604
rect 11980 10480 12020 10520
rect 11884 10396 11924 10436
rect 11980 10144 12020 10184
rect 11788 9556 11828 9596
rect 11788 8800 11828 8840
rect 11692 7036 11732 7076
rect 11884 8464 11924 8504
rect 11884 8044 11924 8084
rect 11212 6532 11252 6572
rect 11356 6364 11396 6404
rect 10732 6280 10772 6320
rect 11020 6280 11060 6320
rect 11212 6280 11252 6320
rect 10540 5944 10580 5984
rect 10156 5104 10196 5144
rect 10156 4768 10196 4808
rect 10060 4096 10100 4136
rect 10156 3928 10196 3968
rect 9676 3844 9716 3884
rect 10540 5524 10580 5564
rect 10828 5356 10868 5396
rect 9868 3172 9908 3212
rect 10444 4096 10484 4136
rect 10636 4096 10676 4136
rect 10156 3256 10196 3296
rect 9964 2752 10004 2792
rect 10156 3004 10196 3044
rect 10060 2584 10100 2624
rect 9580 2332 9620 2372
rect 9484 1660 9524 1700
rect 9484 1492 9524 1532
rect 9196 904 9236 944
rect 9100 736 9140 776
rect 9100 568 9140 608
rect 8908 316 8948 356
rect 9868 1912 9908 1952
rect 10732 3592 10772 3632
rect 10924 4348 10964 4388
rect 10828 3508 10868 3548
rect 10540 3256 10580 3296
rect 10924 3424 10964 3464
rect 10828 3256 10868 3296
rect 10732 3172 10772 3212
rect 10444 2668 10484 2708
rect 10924 2668 10964 2708
rect 11308 5944 11348 5984
rect 11212 4768 11252 4808
rect 11788 6616 11828 6656
rect 11630 6364 11670 6404
rect 11692 6196 11732 6236
rect 11596 6112 11636 6152
rect 11596 4264 11636 4304
rect 11500 4180 11540 4220
rect 11212 3592 11252 3632
rect 11116 3508 11156 3548
rect 11212 3256 11252 3296
rect 11116 3172 11156 3212
rect 10444 2500 10484 2540
rect 10060 1996 10100 2036
rect 10540 1996 10580 2036
rect 10540 1576 10580 1616
rect 9868 1492 9908 1532
rect 10156 1156 10196 1196
rect 10732 1408 10772 1448
rect 10636 1324 10676 1364
rect 10060 904 10100 944
rect 9964 400 10004 440
rect 10252 820 10292 860
rect 10924 2080 10964 2120
rect 10924 1660 10964 1700
rect 10828 1156 10868 1196
rect 10732 484 10772 524
rect 10828 400 10868 440
rect 11308 3088 11348 3128
rect 11308 2668 11348 2708
rect 12268 13336 12308 13376
rect 12460 11656 12500 11696
rect 12748 17788 12788 17828
rect 13036 18712 13076 18752
rect 12940 17956 12980 17996
rect 12748 16696 12788 16736
rect 12748 15520 12788 15560
rect 12652 15268 12692 15308
rect 12844 15436 12884 15476
rect 13612 23248 13652 23288
rect 13612 23080 13652 23120
rect 13516 21904 13556 21944
rect 13708 22828 13748 22868
rect 13708 22240 13748 22280
rect 13228 21568 13268 21608
rect 13420 21568 13460 21608
rect 13420 21400 13460 21440
rect 13324 19300 13364 19340
rect 13132 17536 13172 17576
rect 13132 15856 13172 15896
rect 12844 14848 12884 14888
rect 12748 14680 12788 14720
rect 12652 12244 12692 12284
rect 12556 10732 12596 10772
rect 12460 10312 12500 10352
rect 12364 10144 12404 10184
rect 12748 10564 12788 10604
rect 12652 10144 12692 10184
rect 12556 8968 12596 9008
rect 12460 8800 12500 8840
rect 12556 8212 12596 8252
rect 12268 7876 12308 7916
rect 13036 14680 13076 14720
rect 12940 14512 12980 14552
rect 13228 14848 13268 14888
rect 13612 21568 13652 21608
rect 13708 21400 13748 21440
rect 13516 20728 13556 20768
rect 13612 19300 13652 19340
rect 13516 19216 13556 19256
rect 13516 17704 13556 17744
rect 13708 18964 13748 19004
rect 14380 32152 14420 32192
rect 14188 31732 14228 31772
rect 14380 31564 14420 31604
rect 14956 34000 14996 34040
rect 14668 33664 14708 33704
rect 15436 49120 15476 49160
rect 15628 49120 15668 49160
rect 15820 49120 15860 49160
rect 15820 48196 15860 48236
rect 16204 50632 16244 50672
rect 16204 48868 16244 48908
rect 16012 46768 16052 46808
rect 16108 46180 16148 46220
rect 15724 46096 15764 46136
rect 15532 45340 15572 45380
rect 15436 44920 15476 44960
rect 15436 44416 15476 44456
rect 15532 43156 15572 43196
rect 15436 37864 15476 37904
rect 15340 36184 15380 36224
rect 15532 35176 15572 35216
rect 15532 34672 15572 34712
rect 16012 45592 16052 45632
rect 15724 44416 15764 44456
rect 15820 44164 15860 44204
rect 15820 43408 15860 43448
rect 15820 43156 15860 43196
rect 15724 39712 15764 39752
rect 16108 44584 16148 44624
rect 16204 44332 16244 44372
rect 16876 55588 16916 55628
rect 16972 55504 17012 55544
rect 16588 55168 16628 55208
rect 16780 55336 16820 55376
rect 16684 54832 16724 54872
rect 16588 54244 16628 54284
rect 16780 54160 16820 54200
rect 16684 53824 16724 53864
rect 16588 53068 16628 53108
rect 16972 53824 17012 53864
rect 16876 53488 16916 53528
rect 17548 57016 17588 57056
rect 17356 56260 17396 56300
rect 17452 55252 17492 55292
rect 17260 54916 17300 54956
rect 17356 54832 17396 54872
rect 17164 54076 17204 54116
rect 17452 54076 17492 54116
rect 17356 53488 17396 53528
rect 17260 53404 17300 53444
rect 17068 53068 17108 53108
rect 16780 52060 16820 52100
rect 16972 51976 17012 52016
rect 16780 50968 16820 51008
rect 16684 50380 16724 50420
rect 16396 49708 16436 49748
rect 16396 49456 16436 49496
rect 16396 47440 16436 47480
rect 16588 50044 16628 50084
rect 16588 49708 16628 49748
rect 16588 49456 16628 49496
rect 17068 51052 17108 51092
rect 17068 50380 17108 50420
rect 17452 52900 17492 52940
rect 17260 52060 17300 52100
rect 17260 51220 17300 51260
rect 17260 50464 17300 50504
rect 17068 50212 17108 50252
rect 16972 50128 17012 50168
rect 16876 49708 16916 49748
rect 17164 50128 17204 50168
rect 16876 47944 16916 47984
rect 16780 47440 16820 47480
rect 16972 47272 17012 47312
rect 16108 43408 16148 43448
rect 16012 41476 16052 41516
rect 16300 39628 16340 39668
rect 16300 39124 16340 39164
rect 15820 37864 15860 37904
rect 15724 33664 15764 33704
rect 16012 33496 16052 33536
rect 16204 33664 16244 33704
rect 14764 32656 14804 32696
rect 14668 32152 14708 32192
rect 14668 31984 14708 32024
rect 14572 31816 14612 31856
rect 14476 31480 14516 31520
rect 15148 32152 15188 32192
rect 14860 31984 14900 32024
rect 14860 31816 14900 31856
rect 14572 31060 14612 31100
rect 14572 30640 14612 30680
rect 14476 29800 14516 29840
rect 14380 29548 14420 29588
rect 14188 28288 14228 28328
rect 14284 27616 14324 27656
rect 14188 27028 14228 27068
rect 14764 30640 14804 30680
rect 14668 30220 14708 30260
rect 14668 30052 14708 30092
rect 14764 29800 14804 29840
rect 14476 27448 14516 27488
rect 14092 25516 14132 25556
rect 14092 24844 14132 24884
rect 13996 23920 14036 23960
rect 13996 23752 14036 23792
rect 14380 25180 14420 25220
rect 14380 24592 14420 24632
rect 14188 24088 14228 24128
rect 14380 23920 14420 23960
rect 14284 23752 14324 23792
rect 13996 22492 14036 22532
rect 14092 22324 14132 22364
rect 14092 21820 14132 21860
rect 13996 20728 14036 20768
rect 13996 20560 14036 20600
rect 14284 22996 14324 23036
rect 14188 20140 14228 20180
rect 14092 19972 14132 20012
rect 13996 19888 14036 19928
rect 13996 19300 14036 19340
rect 14380 22576 14420 22616
rect 14380 20980 14420 21020
rect 14764 27616 14804 27656
rect 14668 27532 14708 27572
rect 14572 26524 14612 26564
rect 14668 26104 14708 26144
rect 14572 26020 14612 26060
rect 14668 25600 14708 25640
rect 14572 25516 14612 25556
rect 14572 23920 14612 23960
rect 14572 23752 14612 23792
rect 14476 20560 14516 20600
rect 14380 20056 14420 20096
rect 14476 19804 14516 19844
rect 14380 19636 14420 19676
rect 14284 19300 14324 19340
rect 13900 19048 13940 19088
rect 13804 18712 13844 18752
rect 13804 18544 13844 18584
rect 14188 19216 14228 19256
rect 13516 17032 13556 17072
rect 13420 15856 13460 15896
rect 13708 15520 13748 15560
rect 13612 15268 13652 15308
rect 14188 16864 14228 16904
rect 13996 15772 14036 15812
rect 14092 15688 14132 15728
rect 13132 13840 13172 13880
rect 13132 13168 13172 13208
rect 13324 14428 13364 14468
rect 13516 14428 13556 14468
rect 13420 13336 13460 13376
rect 13612 13252 13652 13292
rect 13420 13168 13460 13208
rect 14284 15268 14324 15308
rect 13996 14848 14036 14888
rect 13804 13672 13844 13712
rect 13900 13252 13940 13292
rect 13036 12244 13076 12284
rect 12940 11740 12980 11780
rect 13420 12832 13460 12872
rect 13324 11572 13364 11612
rect 13036 10984 13076 11024
rect 12940 10816 12980 10856
rect 12844 8716 12884 8756
rect 12748 8632 12788 8672
rect 12940 8212 12980 8252
rect 12652 7960 12692 8000
rect 12556 7876 12596 7916
rect 12268 6616 12308 6656
rect 11980 5356 12020 5396
rect 11884 5104 11924 5144
rect 11788 5020 11828 5060
rect 12172 6448 12212 6488
rect 12268 5524 12308 5564
rect 12268 5104 12308 5144
rect 12556 6616 12596 6656
rect 12748 7456 12788 7496
rect 12940 7960 12980 8000
rect 13420 10984 13460 11024
rect 13324 10144 13364 10184
rect 13228 9304 13268 9344
rect 13132 7120 13172 7160
rect 13036 6700 13076 6740
rect 12844 6448 12884 6488
rect 13132 6448 13172 6488
rect 12460 5608 12500 5648
rect 12556 5524 12596 5564
rect 12460 5188 12500 5228
rect 13036 6364 13076 6404
rect 12940 5608 12980 5648
rect 12556 5020 12596 5060
rect 12076 4936 12116 4976
rect 12172 4852 12212 4892
rect 11788 4096 11828 4136
rect 11980 4096 12020 4136
rect 11308 2164 11348 2204
rect 11212 1912 11252 1952
rect 12844 5020 12884 5060
rect 12748 4936 12788 4976
rect 13036 4936 13076 4976
rect 13420 7792 13460 7832
rect 13324 6952 13364 6992
rect 13708 12832 13748 12872
rect 13612 12244 13652 12284
rect 13804 11572 13844 11612
rect 13708 10564 13748 10604
rect 13708 10312 13748 10352
rect 13612 9472 13652 9512
rect 13708 9220 13748 9260
rect 13612 8212 13652 8252
rect 13612 7120 13652 7160
rect 13612 6868 13652 6908
rect 13516 6448 13556 6488
rect 13324 6364 13364 6404
rect 14188 14092 14228 14132
rect 14188 13336 14228 13376
rect 14092 12244 14132 12284
rect 14572 18880 14612 18920
rect 14764 20728 14804 20768
rect 14764 20560 14804 20600
rect 14956 31480 14996 31520
rect 15340 32320 15380 32360
rect 15436 32152 15476 32192
rect 15244 31480 15284 31520
rect 15340 31228 15380 31268
rect 15244 31144 15284 31184
rect 15148 30640 15188 30680
rect 15820 32152 15860 32192
rect 15916 32068 15956 32108
rect 15052 30472 15092 30512
rect 14956 28288 14996 28328
rect 15244 30556 15284 30596
rect 15244 29968 15284 30008
rect 15340 29716 15380 29756
rect 15244 29548 15284 29588
rect 14956 26188 14996 26228
rect 14956 25516 14996 25556
rect 14956 25264 14996 25304
rect 15148 26104 15188 26144
rect 15628 30595 15668 30596
rect 15628 30556 15668 30595
rect 15724 30472 15764 30512
rect 15820 30220 15860 30260
rect 15724 30052 15764 30092
rect 15628 29800 15668 29840
rect 15916 29800 15956 29840
rect 15820 29632 15860 29672
rect 15244 25600 15284 25640
rect 15148 25516 15188 25556
rect 15532 28876 15572 28916
rect 15436 27952 15476 27992
rect 15532 27616 15572 27656
rect 15724 27616 15764 27656
rect 15628 27532 15668 27572
rect 16108 33328 16148 33368
rect 16204 32908 16244 32948
rect 16108 31900 16148 31940
rect 16780 45760 16820 45800
rect 16492 44836 16532 44876
rect 16876 45172 16916 45212
rect 17068 45340 17108 45380
rect 17068 44248 17108 44288
rect 17452 52060 17492 52100
rect 18316 63904 18356 63944
rect 18220 63736 18260 63776
rect 18220 63316 18260 63356
rect 18412 63232 18452 63272
rect 18316 63064 18356 63104
rect 18220 60712 18260 60752
rect 18124 60460 18164 60500
rect 17836 58108 17876 58148
rect 17836 57100 17876 57140
rect 18124 59284 18164 59324
rect 18028 59116 18068 59156
rect 18316 60376 18356 60416
rect 18316 59200 18356 59240
rect 17932 56932 17972 56972
rect 17836 56848 17876 56888
rect 17740 56260 17780 56300
rect 18220 58192 18260 58232
rect 18124 58108 18164 58148
rect 18028 56848 18068 56888
rect 18028 56260 18068 56300
rect 18124 56176 18164 56216
rect 18124 55504 18164 55544
rect 17644 55084 17684 55124
rect 17644 54496 17684 54536
rect 17932 54916 17972 54956
rect 17548 51976 17588 52016
rect 17740 51808 17780 51848
rect 17644 51220 17684 51260
rect 17452 50968 17492 51008
rect 17548 50464 17588 50504
rect 17452 50380 17492 50420
rect 17548 50044 17588 50084
rect 17356 49120 17396 49160
rect 17260 47272 17300 47312
rect 17164 44164 17204 44204
rect 16972 42400 17012 42440
rect 17164 42148 17204 42188
rect 16588 34924 16628 34964
rect 16492 33496 16532 33536
rect 16300 32320 16340 32360
rect 16108 31144 16148 31184
rect 16204 31060 16244 31100
rect 16204 30220 16244 30260
rect 16588 32656 16628 32696
rect 16780 31900 16820 31940
rect 16588 30976 16628 31016
rect 16300 29548 16340 29588
rect 16588 30472 16628 30512
rect 16684 29884 16724 29924
rect 16492 29380 16532 29420
rect 16300 29296 16340 29336
rect 16684 29296 16724 29336
rect 16492 29212 16532 29252
rect 16396 29044 16436 29084
rect 15916 27532 15956 27572
rect 16204 27700 16244 27740
rect 16108 26944 16148 26984
rect 15436 26104 15476 26144
rect 14956 24592 14996 24632
rect 15148 24256 15188 24296
rect 15340 25264 15380 25304
rect 15916 26608 15956 26648
rect 15820 26188 15860 26228
rect 16012 25852 16052 25892
rect 16204 26104 16244 26144
rect 16780 29128 16820 29168
rect 16684 28876 16724 28916
rect 16588 27448 16628 27488
rect 16588 26944 16628 26984
rect 16108 25516 16148 25556
rect 15436 25180 15476 25220
rect 15340 24592 15380 24632
rect 15052 23757 15092 23792
rect 15052 23752 15092 23757
rect 14956 23416 14996 23456
rect 15244 23668 15284 23708
rect 15532 24256 15572 24296
rect 15628 24004 15668 24044
rect 15532 23668 15572 23708
rect 15244 23416 15284 23456
rect 15244 23164 15284 23204
rect 14956 21652 14996 21692
rect 14956 20728 14996 20768
rect 15532 23416 15572 23456
rect 15436 23248 15476 23288
rect 15532 23080 15572 23120
rect 15436 22996 15476 23036
rect 15532 22912 15572 22952
rect 15436 21316 15476 21356
rect 15724 23836 15764 23876
rect 16108 24760 16148 24800
rect 15916 23836 15956 23876
rect 15820 23752 15860 23792
rect 16108 23584 16148 23624
rect 16108 23416 16148 23456
rect 15820 23248 15860 23288
rect 15628 22744 15668 22784
rect 15916 22744 15956 22784
rect 15724 21568 15764 21608
rect 15628 20728 15668 20768
rect 14860 18292 14900 18332
rect 15244 18292 15284 18332
rect 14956 18124 14996 18164
rect 14956 17956 14996 17996
rect 15244 17872 15284 17912
rect 14668 17620 14708 17660
rect 14572 16948 14612 16988
rect 14572 16780 14612 16820
rect 15148 17536 15188 17576
rect 15244 17032 15284 17072
rect 14956 16948 14996 16988
rect 14860 16864 14900 16904
rect 15052 16780 15092 16820
rect 15148 16444 15188 16484
rect 14380 13336 14420 13376
rect 14092 11488 14132 11528
rect 13996 10060 14036 10100
rect 13900 8044 13940 8084
rect 13804 7792 13844 7832
rect 13804 7120 13844 7160
rect 12460 4768 12500 4808
rect 12364 4600 12404 4640
rect 12556 4096 12596 4136
rect 13036 4516 13076 4556
rect 12364 3340 12404 3380
rect 12940 2668 12980 2708
rect 12844 2332 12884 2372
rect 11500 1660 11540 1700
rect 11692 1324 11732 1364
rect 11116 1240 11156 1280
rect 12268 1828 12308 1868
rect 12940 1828 12980 1868
rect 12844 1744 12884 1784
rect 12364 1660 12404 1700
rect 11980 1408 12020 1448
rect 11116 904 11156 944
rect 11212 736 11252 776
rect 11788 904 11828 944
rect 11596 484 11636 524
rect 12172 1240 12212 1280
rect 12076 232 12116 272
rect 13132 4432 13172 4472
rect 12748 1492 12788 1532
rect 12748 1240 12788 1280
rect 12556 1072 12596 1112
rect 13900 6364 13940 6404
rect 13804 5104 13844 5144
rect 13804 4936 13844 4976
rect 13708 4684 13748 4724
rect 13708 4096 13748 4136
rect 13420 3424 13460 3464
rect 13228 3088 13268 3128
rect 13228 2668 13268 2708
rect 13228 2500 13268 2540
rect 13804 3592 13844 3632
rect 14380 11152 14420 11192
rect 14380 10984 14420 11024
rect 14188 10900 14228 10940
rect 14284 10480 14324 10520
rect 14284 10144 14324 10184
rect 14188 9640 14228 9680
rect 14188 8800 14228 8840
rect 14572 14512 14612 14552
rect 15052 15268 15092 15308
rect 14956 14512 14996 14552
rect 15244 15352 15284 15392
rect 15628 19552 15668 19592
rect 15820 20728 15860 20768
rect 15820 19804 15860 19844
rect 15724 18964 15764 19004
rect 15628 18880 15668 18920
rect 15436 18796 15476 18836
rect 15436 17788 15476 17828
rect 15628 18208 15668 18248
rect 16108 22828 16148 22868
rect 16300 25432 16340 25472
rect 16492 25180 16532 25220
rect 16684 25852 16724 25892
rect 16780 24760 16820 24800
rect 17644 49372 17684 49412
rect 17644 48784 17684 48824
rect 17548 44584 17588 44624
rect 17932 50548 17972 50588
rect 18412 58276 18452 58316
rect 18808 68020 18848 68060
rect 18890 68020 18930 68060
rect 18972 68020 19012 68060
rect 19054 68020 19094 68060
rect 19136 68020 19176 68060
rect 18988 67852 19028 67892
rect 19276 67516 19316 67556
rect 19564 68104 19604 68144
rect 19468 67600 19508 67640
rect 19660 67600 19700 67640
rect 19852 67600 19892 67640
rect 19756 67348 19796 67388
rect 19372 66760 19412 66800
rect 18808 66508 18848 66548
rect 18890 66508 18930 66548
rect 18972 66508 19012 66548
rect 19054 66508 19094 66548
rect 19136 66508 19176 66548
rect 18808 64996 18848 65036
rect 18890 64996 18930 65036
rect 18972 64996 19012 65036
rect 19054 64996 19094 65036
rect 19136 64996 19176 65036
rect 18808 63484 18848 63524
rect 18890 63484 18930 63524
rect 18972 63484 19012 63524
rect 19054 63484 19094 63524
rect 19136 63484 19176 63524
rect 18700 63232 18740 63272
rect 18604 60292 18644 60332
rect 18808 61972 18848 62012
rect 18890 61972 18930 62012
rect 18972 61972 19012 62012
rect 19054 61972 19094 62012
rect 19136 61972 19176 62012
rect 20236 67516 20276 67556
rect 20044 67432 20084 67472
rect 20048 67264 20088 67304
rect 20130 67264 20170 67304
rect 20212 67264 20252 67304
rect 20294 67264 20334 67304
rect 20376 67264 20416 67304
rect 19948 66760 19988 66800
rect 20048 65752 20088 65792
rect 20130 65752 20170 65792
rect 20212 65752 20252 65792
rect 20294 65752 20334 65792
rect 20376 65752 20416 65792
rect 19660 64660 19700 64700
rect 20048 64240 20088 64280
rect 20130 64240 20170 64280
rect 20212 64240 20252 64280
rect 20294 64240 20334 64280
rect 20376 64240 20416 64280
rect 19948 62980 19988 63020
rect 19468 60880 19508 60920
rect 18808 60460 18848 60500
rect 18890 60460 18930 60500
rect 18972 60460 19012 60500
rect 19054 60460 19094 60500
rect 19136 60460 19176 60500
rect 19084 60124 19124 60164
rect 18700 59872 18740 59912
rect 19276 59872 19316 59912
rect 19276 59452 19316 59492
rect 19084 59116 19124 59156
rect 18808 58948 18848 58988
rect 18890 58948 18930 58988
rect 18972 58948 19012 58988
rect 19054 58948 19094 58988
rect 19136 58948 19176 58988
rect 18700 58192 18740 58232
rect 19276 57940 19316 57980
rect 18808 57436 18848 57476
rect 18890 57436 18930 57476
rect 18972 57436 19012 57476
rect 19054 57436 19094 57476
rect 19136 57436 19176 57476
rect 18892 57184 18932 57224
rect 18604 57100 18644 57140
rect 19180 56428 19220 56468
rect 18604 56176 18644 56216
rect 18316 54748 18356 54788
rect 18808 55924 18848 55964
rect 18890 55924 18930 55964
rect 18972 55924 19012 55964
rect 19054 55924 19094 55964
rect 19136 55924 19176 55964
rect 19372 55756 19412 55796
rect 19660 60124 19700 60164
rect 19852 59116 19892 59156
rect 19852 57520 19892 57560
rect 19564 57184 19604 57224
rect 19564 57016 19604 57056
rect 19564 55672 19604 55712
rect 18508 54496 18548 54536
rect 18316 54244 18356 54284
rect 18220 53236 18260 53276
rect 17836 50128 17876 50168
rect 18316 51892 18356 51932
rect 18412 51808 18452 51848
rect 17932 49792 17972 49832
rect 19276 54580 19316 54620
rect 18808 54412 18848 54452
rect 18890 54412 18930 54452
rect 18972 54412 19012 54452
rect 19054 54412 19094 54452
rect 19136 54412 19176 54452
rect 19180 54244 19220 54284
rect 19084 53992 19124 54032
rect 18700 53320 18740 53360
rect 18808 52900 18848 52940
rect 18890 52900 18930 52940
rect 18972 52900 19012 52940
rect 19054 52900 19094 52940
rect 19136 52900 19176 52940
rect 19468 53572 19508 53612
rect 19852 54748 19892 54788
rect 19660 54496 19700 54536
rect 19852 54328 19892 54368
rect 19852 54076 19892 54116
rect 18604 50464 18644 50504
rect 18796 51892 18836 51932
rect 19276 52144 19316 52184
rect 19372 52060 19412 52100
rect 18796 51724 18836 51764
rect 18808 51388 18848 51428
rect 18890 51388 18930 51428
rect 18972 51388 19012 51428
rect 19054 51388 19094 51428
rect 19136 51388 19176 51428
rect 19180 51052 19220 51092
rect 19180 50800 19220 50840
rect 19372 50800 19412 50840
rect 19276 50464 19316 50504
rect 18220 50128 18260 50168
rect 18124 49792 18164 49832
rect 18028 49540 18068 49580
rect 18124 49372 18164 49412
rect 18508 49792 18548 49832
rect 18808 49876 18848 49916
rect 18890 49876 18930 49916
rect 18972 49876 19012 49916
rect 19054 49876 19094 49916
rect 19136 49876 19176 49916
rect 19756 53320 19796 53360
rect 20048 62728 20088 62768
rect 20130 62728 20170 62768
rect 20212 62728 20252 62768
rect 20294 62728 20334 62768
rect 20376 62728 20416 62768
rect 20716 74488 20756 74528
rect 20716 63400 20756 63440
rect 20524 62476 20564 62516
rect 20716 61720 20756 61760
rect 20048 61216 20088 61256
rect 20130 61216 20170 61256
rect 20212 61216 20252 61256
rect 20294 61216 20334 61256
rect 20376 61216 20416 61256
rect 20048 59704 20088 59744
rect 20130 59704 20170 59744
rect 20212 59704 20252 59744
rect 20294 59704 20334 59744
rect 20376 59704 20416 59744
rect 20620 59704 20660 59744
rect 20048 58192 20088 58232
rect 20130 58192 20170 58232
rect 20212 58192 20252 58232
rect 20294 58192 20334 58232
rect 20376 58192 20416 58232
rect 20044 57940 20084 57980
rect 20048 56680 20088 56720
rect 20130 56680 20170 56720
rect 20212 56680 20252 56720
rect 20294 56680 20334 56720
rect 20376 56680 20416 56720
rect 20048 55168 20088 55208
rect 20130 55168 20170 55208
rect 20212 55168 20252 55208
rect 20294 55168 20334 55208
rect 20376 55168 20416 55208
rect 20236 55000 20276 55040
rect 20044 54748 20084 54788
rect 20044 53824 20084 53864
rect 20048 53656 20088 53696
rect 20130 53656 20170 53696
rect 20212 53656 20252 53696
rect 20294 53656 20334 53696
rect 20376 53656 20416 53696
rect 19756 52732 19796 52772
rect 19756 52396 19796 52436
rect 19660 52312 19700 52352
rect 19660 52060 19700 52100
rect 19564 51976 19604 52016
rect 19564 50800 19604 50840
rect 19468 50044 19508 50084
rect 18988 49708 19028 49748
rect 18700 49456 18740 49496
rect 18412 48868 18452 48908
rect 18316 48784 18356 48824
rect 17836 47944 17876 47984
rect 17740 47776 17780 47816
rect 18028 47776 18068 47816
rect 17932 47020 17972 47060
rect 17836 45340 17876 45380
rect 17740 44920 17780 44960
rect 17644 44500 17684 44540
rect 17452 43744 17492 43784
rect 17740 44080 17780 44120
rect 17740 43492 17780 43532
rect 17932 45172 17972 45212
rect 18316 47776 18356 47816
rect 18220 47188 18260 47228
rect 18412 47020 18452 47060
rect 18316 46852 18356 46892
rect 18604 48616 18644 48656
rect 19180 48952 19220 48992
rect 19372 49624 19412 49664
rect 20044 52396 20084 52436
rect 20048 52144 20088 52184
rect 20130 52144 20170 52184
rect 20212 52144 20252 52184
rect 20294 52144 20334 52184
rect 20376 52144 20416 52184
rect 20044 51976 20084 52016
rect 19948 51640 19988 51680
rect 19948 51304 19988 51344
rect 19756 50464 19796 50504
rect 20140 50968 20180 51008
rect 19948 50632 19988 50672
rect 20048 50632 20088 50672
rect 20130 50632 20170 50672
rect 20212 50632 20252 50672
rect 20294 50632 20334 50672
rect 20376 50632 20416 50672
rect 19852 50380 19892 50420
rect 19660 50296 19700 50336
rect 19852 50128 19892 50168
rect 19660 49624 19700 49664
rect 20044 50296 20084 50336
rect 18808 48364 18848 48404
rect 18890 48364 18930 48404
rect 18972 48364 19012 48404
rect 19054 48364 19094 48404
rect 19136 48364 19176 48404
rect 19276 47524 19316 47564
rect 19276 47356 19316 47396
rect 18700 46852 18740 46892
rect 18808 46852 18848 46892
rect 18890 46852 18930 46892
rect 18972 46852 19012 46892
rect 19054 46852 19094 46892
rect 19136 46852 19176 46892
rect 18988 46684 19028 46724
rect 18220 45676 18260 45716
rect 18124 45088 18164 45128
rect 18508 46432 18548 46472
rect 18508 45172 18548 45212
rect 18316 44836 18356 44876
rect 18124 44500 18164 44540
rect 18316 44248 18356 44288
rect 18220 44164 18260 44204
rect 17548 42820 17588 42860
rect 17452 32656 17492 32696
rect 18028 42904 18068 42944
rect 17932 42232 17972 42272
rect 17740 40384 17780 40424
rect 17740 31312 17780 31352
rect 17836 31228 17876 31268
rect 18028 41980 18068 42020
rect 17740 30724 17780 30764
rect 17644 30220 17684 30260
rect 17356 30052 17396 30092
rect 17548 29800 17588 29840
rect 17164 29296 17204 29336
rect 16972 29212 17012 29252
rect 17220 29044 17260 29084
rect 17740 29464 17780 29504
rect 17644 29380 17684 29420
rect 17548 29044 17588 29084
rect 17740 29128 17780 29168
rect 17068 27616 17108 27656
rect 17164 27448 17204 27488
rect 17260 27280 17300 27320
rect 17068 26608 17108 26648
rect 16972 26188 17012 26228
rect 17356 26692 17396 26732
rect 17452 26524 17492 26564
rect 17164 25432 17204 25472
rect 16972 24760 17012 24800
rect 16876 24592 16916 24632
rect 16492 24424 16532 24464
rect 16300 23584 16340 23624
rect 16396 23332 16436 23372
rect 16012 22072 16052 22112
rect 16204 22660 16244 22700
rect 16204 21820 16244 21860
rect 16012 21484 16052 21524
rect 16108 21400 16148 21440
rect 16012 21316 16052 21356
rect 15916 18712 15956 18752
rect 15724 17956 15764 17996
rect 15820 17872 15860 17912
rect 15436 17200 15476 17240
rect 15436 14848 15476 14888
rect 15724 15268 15764 15308
rect 15532 14680 15572 14720
rect 14668 13756 14708 13796
rect 15148 13336 15188 13376
rect 15052 13000 15092 13040
rect 15340 13840 15380 13880
rect 15244 12580 15284 12620
rect 14956 11656 14996 11696
rect 14860 11488 14900 11528
rect 15436 13756 15476 13796
rect 14956 10984 14996 11024
rect 15052 10900 15092 10940
rect 14668 10816 14708 10856
rect 14668 10228 14708 10268
rect 14668 9892 14708 9932
rect 14572 9472 14612 9512
rect 14572 8380 14612 8420
rect 14476 8044 14516 8084
rect 14092 7708 14132 7748
rect 14380 7456 14420 7496
rect 14284 7372 14324 7412
rect 14860 9472 14900 9512
rect 14860 9304 14900 9344
rect 15628 13336 15668 13376
rect 15532 13168 15572 13208
rect 15148 8212 15188 8252
rect 15340 8884 15380 8924
rect 15436 8716 15476 8756
rect 14956 7120 14996 7160
rect 14380 6868 14420 6908
rect 14188 5524 14228 5564
rect 14764 5356 14804 5396
rect 14188 5188 14228 5228
rect 14188 4180 14228 4220
rect 15724 13168 15764 13208
rect 15628 12580 15668 12620
rect 15724 10396 15764 10436
rect 16012 17704 16052 17744
rect 15916 17536 15956 17576
rect 15916 17116 15956 17156
rect 16204 20728 16244 20768
rect 16396 22576 16436 22616
rect 16396 22240 16436 22280
rect 17356 24760 17396 24800
rect 17260 24088 17300 24128
rect 18028 30472 18068 30512
rect 17932 30304 17972 30344
rect 18892 45928 18932 45968
rect 18892 45760 18932 45800
rect 18700 45676 18740 45716
rect 18988 45676 19028 45716
rect 19756 48952 19796 48992
rect 20048 49120 20088 49160
rect 20130 49120 20170 49160
rect 20212 49120 20252 49160
rect 20294 49120 20334 49160
rect 20376 49120 20416 49160
rect 19948 48952 19988 48992
rect 19948 48448 19988 48488
rect 19852 48280 19892 48320
rect 19852 48028 19892 48068
rect 19468 47944 19508 47984
rect 19468 47524 19508 47564
rect 19852 47188 19892 47228
rect 20140 47776 20180 47816
rect 20048 47608 20088 47648
rect 20130 47608 20170 47648
rect 20212 47608 20252 47648
rect 20294 47608 20334 47648
rect 20376 47608 20416 47648
rect 19948 46936 19988 46976
rect 19468 46684 19508 46724
rect 19852 46516 19892 46556
rect 19276 45760 19316 45800
rect 18796 45508 18836 45548
rect 19084 45508 19124 45548
rect 18808 45340 18848 45380
rect 18890 45340 18930 45380
rect 18972 45340 19012 45380
rect 19054 45340 19094 45380
rect 19136 45340 19176 45380
rect 18892 45172 18932 45212
rect 18988 45088 19028 45128
rect 18988 44920 19028 44960
rect 18892 44752 18932 44792
rect 18808 43828 18848 43868
rect 18890 43828 18930 43868
rect 18972 43828 19012 43868
rect 19054 43828 19094 43868
rect 19136 43828 19176 43868
rect 19180 43660 19220 43700
rect 18988 43492 19028 43532
rect 19372 45508 19412 45548
rect 19564 45844 19604 45884
rect 20044 46264 20084 46304
rect 20048 46096 20088 46136
rect 20130 46096 20170 46136
rect 20212 46096 20252 46136
rect 20294 46096 20334 46136
rect 20376 46096 20416 46136
rect 19660 45676 19700 45716
rect 19660 45508 19700 45548
rect 19852 45004 19892 45044
rect 19756 44920 19796 44960
rect 19852 44752 19892 44792
rect 19756 44500 19796 44540
rect 19372 44248 19412 44288
rect 19180 42568 19220 42608
rect 18796 42484 18836 42524
rect 18508 41980 18548 42020
rect 18508 41728 18548 41768
rect 18316 40972 18356 41012
rect 18316 35008 18356 35048
rect 18316 33496 18356 33536
rect 18220 33328 18260 33368
rect 18412 31228 18452 31268
rect 18412 30220 18452 30260
rect 17836 28372 17876 28412
rect 17836 27784 17876 27824
rect 17740 27700 17780 27740
rect 17644 26692 17684 26732
rect 18124 29884 18164 29924
rect 18316 29884 18356 29924
rect 18124 29632 18164 29672
rect 18412 29800 18452 29840
rect 18124 29212 18164 29252
rect 18028 29128 18068 29168
rect 18124 27784 18164 27824
rect 18316 27952 18356 27992
rect 18220 27532 18260 27572
rect 18028 27196 18068 27236
rect 17932 26776 17972 26816
rect 17836 25180 17876 25220
rect 17068 23920 17108 23960
rect 17836 23920 17876 23960
rect 16780 23500 16820 23540
rect 16684 23416 16724 23456
rect 16588 21820 16628 21860
rect 16492 21736 16532 21776
rect 16396 21400 16436 21440
rect 16972 22660 17012 22700
rect 17644 23668 17684 23708
rect 17836 23500 17876 23540
rect 17836 23332 17876 23372
rect 17452 23248 17492 23288
rect 17356 22576 17396 22616
rect 17452 22492 17492 22532
rect 16588 21484 16628 21524
rect 16300 20476 16340 20516
rect 16876 20728 16916 20768
rect 16780 20644 16820 20684
rect 16300 18964 16340 19004
rect 16204 18712 16244 18752
rect 16204 17116 16244 17156
rect 16204 16864 16244 16904
rect 16300 16444 16340 16484
rect 16972 20560 17012 20600
rect 16876 19972 16916 20012
rect 17164 21400 17204 21440
rect 17164 20812 17204 20852
rect 17356 20812 17396 20852
rect 17740 22072 17780 22112
rect 17548 21400 17588 21440
rect 17548 20644 17588 20684
rect 17164 20476 17204 20516
rect 17068 20056 17108 20096
rect 16876 19720 16916 19760
rect 16876 19300 16916 19340
rect 17356 20308 17396 20348
rect 17836 20644 17876 20684
rect 17740 20476 17780 20516
rect 18412 27112 18452 27152
rect 18220 25180 18260 25220
rect 18988 42484 19028 42524
rect 18808 42316 18848 42356
rect 18890 42316 18930 42356
rect 18972 42316 19012 42356
rect 19054 42316 19094 42356
rect 19136 42316 19176 42356
rect 19276 42148 19316 42188
rect 18892 42064 18932 42104
rect 18700 41812 18740 41852
rect 19756 42652 19796 42692
rect 19660 42232 19700 42272
rect 20048 44584 20088 44624
rect 20130 44584 20170 44624
rect 20212 44584 20252 44624
rect 20294 44584 20334 44624
rect 20376 44584 20416 44624
rect 19948 44248 19988 44288
rect 19948 43576 19988 43616
rect 19948 43240 19988 43280
rect 20048 43072 20088 43112
rect 20130 43072 20170 43112
rect 20212 43072 20252 43112
rect 20294 43072 20334 43112
rect 20376 43072 20416 43112
rect 19852 42148 19892 42188
rect 19372 41560 19412 41600
rect 18892 41392 18932 41432
rect 19084 41392 19124 41432
rect 19372 41308 19412 41348
rect 19276 41140 19316 41180
rect 18988 41056 19028 41096
rect 18892 40972 18932 41012
rect 18808 40804 18848 40844
rect 18890 40804 18930 40844
rect 18972 40804 19012 40844
rect 19054 40804 19094 40844
rect 19136 40804 19176 40844
rect 19084 40636 19124 40676
rect 19468 40972 19508 41012
rect 19468 40636 19508 40676
rect 19660 41728 19700 41768
rect 19660 41476 19700 41516
rect 19564 40552 19604 40592
rect 19660 40468 19700 40508
rect 18988 40132 19028 40172
rect 19564 39964 19604 40004
rect 19852 41812 19892 41852
rect 19948 41644 19988 41684
rect 20048 41560 20088 41600
rect 20130 41560 20170 41600
rect 20212 41560 20252 41600
rect 20294 41560 20334 41600
rect 20376 41560 20416 41600
rect 19852 40972 19892 41012
rect 20044 41224 20084 41264
rect 19948 40468 19988 40508
rect 19852 40216 19892 40256
rect 20048 40048 20088 40088
rect 20130 40048 20170 40088
rect 20212 40048 20252 40088
rect 20294 40048 20334 40088
rect 20376 40048 20416 40088
rect 19948 39880 19988 39920
rect 19372 39712 19412 39752
rect 19564 39712 19604 39752
rect 18808 39292 18848 39332
rect 18890 39292 18930 39332
rect 18972 39292 19012 39332
rect 19054 39292 19094 39332
rect 19136 39292 19176 39332
rect 19372 39460 19412 39500
rect 19756 39628 19796 39668
rect 20524 39544 20564 39584
rect 19660 39376 19700 39416
rect 19276 38872 19316 38912
rect 18700 38452 18740 38492
rect 19276 38368 19316 38408
rect 18808 37780 18848 37820
rect 18890 37780 18930 37820
rect 18972 37780 19012 37820
rect 19054 37780 19094 37820
rect 19136 37780 19176 37820
rect 18700 37528 18740 37568
rect 19564 38200 19604 38240
rect 19564 38032 19604 38072
rect 18988 37276 19028 37316
rect 18892 37192 18932 37232
rect 19180 36856 19220 36896
rect 19564 37444 19604 37484
rect 20048 38536 20088 38576
rect 20130 38536 20170 38576
rect 20212 38536 20252 38576
rect 20294 38536 20334 38576
rect 20376 38536 20416 38576
rect 19948 37612 19988 37652
rect 19660 37276 19700 37316
rect 19468 37192 19508 37232
rect 19756 37108 19796 37148
rect 20048 37024 20088 37064
rect 20130 37024 20170 37064
rect 20212 37024 20252 37064
rect 20294 37024 20334 37064
rect 20376 37024 20416 37064
rect 19372 36604 19412 36644
rect 18892 36436 18932 36476
rect 18808 36268 18848 36308
rect 18890 36268 18930 36308
rect 18972 36268 19012 36308
rect 19054 36268 19094 36308
rect 19136 36268 19176 36308
rect 19276 36184 19316 36224
rect 19180 36016 19220 36056
rect 19180 35260 19220 35300
rect 18978 35008 19018 35048
rect 18808 34756 18848 34796
rect 18890 34756 18930 34796
rect 18972 34756 19012 34796
rect 19054 34756 19094 34796
rect 19136 34756 19176 34796
rect 18700 33328 18740 33368
rect 18808 33244 18848 33284
rect 18890 33244 18930 33284
rect 18972 33244 19012 33284
rect 19054 33244 19094 33284
rect 19136 33244 19176 33284
rect 18808 31732 18848 31772
rect 18890 31732 18930 31772
rect 18972 31732 19012 31772
rect 19054 31732 19094 31772
rect 19136 31732 19176 31772
rect 19372 35092 19412 35132
rect 19564 36772 19604 36812
rect 19660 36604 19700 36644
rect 19564 36268 19604 36308
rect 19564 35008 19604 35048
rect 19468 34840 19508 34880
rect 19564 34588 19604 34628
rect 19372 34000 19412 34040
rect 20908 75832 20948 75872
rect 20812 59788 20852 59828
rect 21388 75160 21428 75200
rect 21004 73144 21044 73184
rect 21100 63736 21140 63776
rect 21004 62644 21044 62684
rect 21004 59032 21044 59072
rect 20908 56764 20948 56804
rect 20716 48532 20756 48572
rect 20620 36016 20660 36056
rect 19948 35596 19988 35636
rect 20048 35512 20088 35552
rect 20130 35512 20170 35552
rect 20212 35512 20252 35552
rect 20294 35512 20334 35552
rect 20376 35512 20416 35552
rect 21292 62392 21332 62432
rect 21196 61048 21236 61088
rect 21196 39880 21236 39920
rect 21388 61552 21428 61592
rect 21292 38788 21332 38828
rect 21100 36268 21140 36308
rect 21388 35764 21428 35804
rect 21388 35512 21428 35552
rect 21004 35260 21044 35300
rect 19756 35176 19796 35216
rect 19756 34504 19796 34544
rect 19852 34168 19892 34208
rect 20048 34000 20088 34040
rect 20130 34000 20170 34040
rect 20212 34000 20252 34040
rect 20294 34000 20334 34040
rect 20376 34000 20416 34040
rect 20048 32488 20088 32528
rect 20130 32488 20170 32528
rect 20212 32488 20252 32528
rect 20294 32488 20334 32528
rect 20376 32488 20416 32528
rect 19660 32236 19700 32276
rect 19276 31564 19316 31604
rect 19468 31312 19508 31352
rect 18700 30976 18740 31016
rect 19276 30976 19316 31016
rect 18604 30640 18644 30680
rect 18796 30892 18836 30932
rect 18700 30472 18740 30512
rect 18604 29464 18644 29504
rect 18028 23836 18068 23876
rect 18124 23752 18164 23792
rect 18028 23500 18068 23540
rect 18028 21400 18068 21440
rect 18220 23248 18260 23288
rect 18124 21064 18164 21104
rect 18124 20728 18164 20768
rect 19276 30472 19316 30512
rect 19084 30388 19124 30428
rect 18808 30220 18848 30260
rect 18890 30220 18930 30260
rect 18972 30220 19012 30260
rect 19054 30220 19094 30260
rect 19136 30220 19176 30260
rect 20044 31144 20084 31184
rect 19948 30976 19988 31016
rect 20048 30976 20088 31016
rect 20130 30976 20170 31016
rect 20212 30976 20252 31016
rect 20294 30976 20334 31016
rect 20376 30976 20416 31016
rect 19660 30220 19700 30260
rect 19468 29968 19508 30008
rect 19084 29632 19124 29672
rect 19564 29800 19604 29840
rect 19564 29464 19604 29504
rect 19948 30640 19988 30680
rect 19852 29968 19892 30008
rect 19948 29716 19988 29756
rect 20236 30640 20276 30680
rect 20620 30472 20660 30512
rect 20524 30388 20564 30428
rect 20044 29632 20084 29672
rect 20048 29464 20088 29504
rect 20130 29464 20170 29504
rect 20212 29464 20252 29504
rect 20294 29464 20334 29504
rect 20376 29464 20416 29504
rect 20140 29296 20180 29336
rect 19660 29212 19700 29252
rect 19948 29128 19988 29168
rect 18808 28708 18848 28748
rect 18890 28708 18930 28748
rect 18972 28708 19012 28748
rect 19054 28708 19094 28748
rect 19136 28708 19176 28748
rect 18700 27532 18740 27572
rect 20044 28456 20084 28496
rect 19468 27868 19508 27908
rect 19756 27952 19796 27992
rect 19948 28288 19988 28328
rect 19852 27784 19892 27824
rect 18808 27196 18848 27236
rect 18890 27196 18930 27236
rect 18972 27196 19012 27236
rect 19054 27196 19094 27236
rect 19136 27196 19176 27236
rect 19276 27196 19316 27236
rect 19468 27280 19508 27320
rect 18700 26776 18740 26816
rect 19372 26776 19412 26816
rect 19660 27196 19700 27236
rect 20048 27952 20088 27992
rect 20130 27952 20170 27992
rect 20212 27952 20252 27992
rect 20294 27952 20334 27992
rect 20376 27952 20416 27992
rect 19948 27448 19988 27488
rect 20140 27700 20180 27740
rect 20044 27364 20084 27404
rect 19852 27196 19892 27236
rect 19084 26440 19124 26480
rect 19276 26440 19316 26480
rect 19564 26608 19604 26648
rect 18808 25684 18848 25724
rect 18890 25684 18930 25724
rect 18972 25684 19012 25724
rect 19054 25684 19094 25724
rect 19136 25684 19176 25724
rect 18808 24172 18848 24212
rect 18890 24172 18930 24212
rect 18972 24172 19012 24212
rect 19054 24172 19094 24212
rect 19136 24172 19176 24212
rect 19756 26776 19796 26816
rect 19948 26692 19988 26732
rect 18604 23332 18644 23372
rect 18412 23248 18452 23288
rect 18700 23080 18740 23120
rect 19372 23920 19412 23960
rect 19180 23836 19220 23876
rect 19276 23584 19316 23624
rect 19852 23668 19892 23708
rect 19564 23584 19604 23624
rect 19852 23500 19892 23540
rect 18604 22072 18644 22112
rect 18508 21736 18548 21776
rect 18808 22660 18848 22700
rect 18890 22660 18930 22700
rect 18972 22660 19012 22700
rect 19054 22660 19094 22700
rect 19136 22660 19176 22700
rect 19276 21652 19316 21692
rect 18988 21568 19028 21608
rect 18808 21148 18848 21188
rect 18890 21148 18930 21188
rect 18972 21148 19012 21188
rect 19054 21148 19094 21188
rect 19136 21148 19176 21188
rect 18508 20812 18548 20852
rect 18028 20644 18068 20684
rect 16492 17536 16532 17576
rect 16876 17536 16916 17576
rect 16684 17368 16724 17408
rect 17068 17032 17108 17072
rect 16780 16948 16820 16988
rect 16204 16360 16244 16400
rect 16396 16276 16436 16316
rect 16684 16276 16724 16316
rect 16876 16864 16916 16904
rect 16108 14092 16148 14132
rect 16012 13840 16052 13880
rect 15916 13672 15956 13712
rect 16204 13672 16244 13712
rect 15916 13252 15956 13292
rect 16588 15520 16628 15560
rect 16588 15268 16628 15308
rect 16492 14848 16532 14888
rect 16492 14512 16532 14552
rect 16396 13252 16436 13292
rect 15916 12496 15956 12536
rect 16300 12496 16340 12536
rect 16108 11908 16148 11948
rect 15916 11152 15956 11192
rect 15628 8884 15668 8924
rect 15532 8632 15572 8672
rect 16012 10396 16052 10436
rect 15820 9052 15860 9092
rect 15436 7120 15476 7160
rect 15436 6952 15476 6992
rect 16012 9472 16052 9512
rect 15244 5356 15284 5396
rect 15724 5440 15764 5480
rect 15532 5020 15572 5060
rect 14956 4180 14996 4220
rect 14764 4096 14804 4136
rect 14188 3340 14228 3380
rect 13996 2920 14036 2960
rect 14572 3256 14612 3296
rect 14860 3172 14900 3212
rect 14188 2584 14228 2624
rect 15052 2752 15092 2792
rect 15244 4096 15284 4136
rect 15916 5020 15956 5060
rect 15820 4096 15860 4136
rect 15244 3424 15284 3464
rect 15436 2920 15476 2960
rect 15532 2752 15572 2792
rect 14668 2416 14708 2456
rect 13708 2332 13748 2372
rect 13900 1828 13940 1868
rect 14284 1828 14324 1868
rect 13324 1576 13364 1616
rect 14284 1408 14324 1448
rect 13900 1240 13940 1280
rect 13708 820 13748 860
rect 13420 736 13460 776
rect 13516 652 13556 692
rect 14092 736 14132 776
rect 14476 904 14516 944
rect 15244 1828 15284 1868
rect 14956 1072 14996 1112
rect 14860 988 14900 1028
rect 14956 904 14996 944
rect 15436 1408 15476 1448
rect 15148 1156 15188 1196
rect 15436 988 15476 1028
rect 15244 820 15284 860
rect 15052 484 15092 524
rect 14956 316 14996 356
rect 15628 1828 15668 1868
rect 15628 1240 15668 1280
rect 15532 316 15572 356
rect 16108 7960 16148 8000
rect 16396 11740 16436 11780
rect 16300 10984 16340 11024
rect 16492 11152 16532 11192
rect 16300 8632 16340 8672
rect 16204 6700 16244 6740
rect 16780 14680 16820 14720
rect 16684 14176 16724 14216
rect 17356 19804 17396 19844
rect 17740 20056 17780 20096
rect 18124 20476 18164 20516
rect 18028 20224 18068 20264
rect 18412 20392 18452 20432
rect 18316 20308 18356 20348
rect 18316 20140 18356 20180
rect 17836 19972 17876 20012
rect 17452 19216 17492 19256
rect 17356 19048 17396 19088
rect 17260 16108 17300 16148
rect 17068 15268 17108 15308
rect 17260 14764 17300 14804
rect 17164 14680 17204 14720
rect 17548 18628 17588 18668
rect 17644 17704 17684 17744
rect 17836 16864 17876 16904
rect 17836 16360 17876 16400
rect 17740 16192 17780 16232
rect 17548 16108 17588 16148
rect 18028 16192 18068 16232
rect 17548 14764 17588 14804
rect 17644 14680 17684 14720
rect 18220 14680 18260 14720
rect 17356 14260 17396 14300
rect 17164 13840 17204 13880
rect 17068 13420 17108 13460
rect 17068 13252 17108 13292
rect 16972 11488 17012 11528
rect 17356 13420 17396 13460
rect 17068 10312 17108 10352
rect 16684 8212 16724 8252
rect 16780 8128 16820 8168
rect 16396 7960 16436 8000
rect 16396 7792 16436 7832
rect 16300 5860 16340 5900
rect 16204 5440 16244 5480
rect 16108 4936 16148 4976
rect 16108 4180 16148 4220
rect 16972 9724 17012 9764
rect 17260 12580 17300 12620
rect 17644 13924 17684 13964
rect 17260 10060 17300 10100
rect 17260 9724 17300 9764
rect 17164 8800 17204 8840
rect 17068 8716 17108 8756
rect 16972 8128 17012 8168
rect 17260 8212 17300 8252
rect 16684 7120 16724 7160
rect 16588 6868 16628 6908
rect 16492 5020 16532 5060
rect 16012 1828 16052 1868
rect 16012 988 16052 1028
rect 15724 736 15764 776
rect 15820 484 15860 524
rect 15820 316 15860 356
rect 16396 1828 16436 1868
rect 16876 6448 16916 6488
rect 16684 5188 16724 5228
rect 17164 7876 17204 7916
rect 17164 7288 17204 7328
rect 16972 5356 17012 5396
rect 17260 5524 17300 5564
rect 17260 5356 17300 5396
rect 16780 4936 16820 4976
rect 16684 2752 16724 2792
rect 16300 988 16340 1028
rect 16204 820 16244 860
rect 16972 4936 17012 4976
rect 16876 2584 16916 2624
rect 17644 12328 17684 12368
rect 17452 11572 17492 11612
rect 17548 11488 17588 11528
rect 17836 11572 17876 11612
rect 17740 9640 17780 9680
rect 17644 9388 17684 9428
rect 17740 8884 17780 8924
rect 17548 8632 17588 8672
rect 17452 8128 17492 8168
rect 17548 7960 17588 8000
rect 17644 7288 17684 7328
rect 17644 6784 17684 6824
rect 18700 20560 18740 20600
rect 18604 19804 18644 19844
rect 18808 19636 18848 19676
rect 18890 19636 18930 19676
rect 18972 19636 19012 19676
rect 19054 19636 19094 19676
rect 19136 19636 19176 19676
rect 18700 19300 18740 19340
rect 18604 19048 18644 19088
rect 18508 18712 18548 18752
rect 18892 19048 18932 19088
rect 18508 17620 18548 17660
rect 18808 18124 18848 18164
rect 18890 18124 18930 18164
rect 18972 18124 19012 18164
rect 19054 18124 19094 18164
rect 19136 18124 19176 18164
rect 19084 17620 19124 17660
rect 18892 17536 18932 17576
rect 19276 17536 19316 17576
rect 18508 16864 18548 16904
rect 18316 13336 18356 13376
rect 18028 10984 18068 11024
rect 18028 10564 18068 10604
rect 18412 11488 18452 11528
rect 18700 17116 18740 17156
rect 18604 14176 18644 14216
rect 18808 16612 18848 16652
rect 18890 16612 18930 16652
rect 18972 16612 19012 16652
rect 19054 16612 19094 16652
rect 19136 16612 19176 16652
rect 18808 15100 18848 15140
rect 18890 15100 18930 15140
rect 18972 15100 19012 15140
rect 19054 15100 19094 15140
rect 19136 15100 19176 15140
rect 19756 23080 19796 23120
rect 21388 29968 21428 30008
rect 20048 26440 20088 26480
rect 20130 26440 20170 26480
rect 20212 26440 20252 26480
rect 20294 26440 20334 26480
rect 20376 26440 20416 26480
rect 20048 24928 20088 24968
rect 20130 24928 20170 24968
rect 20212 24928 20252 24968
rect 20294 24928 20334 24968
rect 20376 24928 20416 24968
rect 20044 23584 20084 23624
rect 20048 23416 20088 23456
rect 20130 23416 20170 23456
rect 20212 23416 20252 23456
rect 20294 23416 20334 23456
rect 20376 23416 20416 23456
rect 20048 21904 20088 21944
rect 20130 21904 20170 21944
rect 20212 21904 20252 21944
rect 20294 21904 20334 21944
rect 20376 21904 20416 21944
rect 20048 20392 20088 20432
rect 20130 20392 20170 20432
rect 20212 20392 20252 20432
rect 20294 20392 20334 20432
rect 20376 20392 20416 20432
rect 20048 18880 20088 18920
rect 20130 18880 20170 18920
rect 20212 18880 20252 18920
rect 20294 18880 20334 18920
rect 20376 18880 20416 18920
rect 19372 17452 19412 17492
rect 20048 17368 20088 17408
rect 20130 17368 20170 17408
rect 20212 17368 20252 17408
rect 20294 17368 20334 17408
rect 20376 17368 20416 17408
rect 20048 15856 20088 15896
rect 20130 15856 20170 15896
rect 20212 15856 20252 15896
rect 20294 15856 20334 15896
rect 20376 15856 20416 15896
rect 18796 14512 18836 14552
rect 18700 14092 18740 14132
rect 20048 14344 20088 14384
rect 20130 14344 20170 14384
rect 20212 14344 20252 14384
rect 20294 14344 20334 14384
rect 20376 14344 20416 14384
rect 19180 14176 19220 14216
rect 19276 14092 19316 14132
rect 18988 13840 19028 13880
rect 18808 13588 18848 13628
rect 18890 13588 18930 13628
rect 18972 13588 19012 13628
rect 19054 13588 19094 13628
rect 19136 13588 19176 13628
rect 18808 12076 18848 12116
rect 18890 12076 18930 12116
rect 18972 12076 19012 12116
rect 19054 12076 19094 12116
rect 19136 12076 19176 12116
rect 20048 12832 20088 12872
rect 20130 12832 20170 12872
rect 20212 12832 20252 12872
rect 20294 12832 20334 12872
rect 20376 12832 20416 12872
rect 19564 12496 19604 12536
rect 18316 10984 18356 11024
rect 18508 10984 18548 11024
rect 18412 10144 18452 10184
rect 18316 9472 18356 9512
rect 18316 9052 18356 9092
rect 18124 8884 18164 8924
rect 18700 10564 18740 10604
rect 18808 10564 18848 10604
rect 18890 10564 18930 10604
rect 18972 10564 19012 10604
rect 19054 10564 19094 10604
rect 19136 10564 19176 10604
rect 18700 10396 18740 10436
rect 20048 11320 20088 11360
rect 20130 11320 20170 11360
rect 20212 11320 20252 11360
rect 20294 11320 20334 11360
rect 20376 11320 20416 11360
rect 19276 9472 19316 9512
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 18700 8800 18740 8840
rect 19468 10396 19508 10436
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 19372 7960 19412 8000
rect 18796 7876 18836 7916
rect 19180 7876 19220 7916
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 18508 6280 18548 6320
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 18892 5272 18932 5312
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 18412 4936 18452 4976
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 21292 24508 21332 24548
rect 20620 24004 20660 24044
rect 20620 23416 20660 23456
rect 20620 18544 20660 18584
rect 20620 16024 20660 16064
rect 21388 18040 21428 18080
rect 21292 15352 21332 15392
rect 21388 8632 21428 8672
rect 21388 8128 21428 8168
rect 20524 1828 20564 1868
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 17356 1240 17396 1280
rect 17548 1240 17588 1280
rect 18124 1240 18164 1280
rect 18508 1240 18548 1280
rect 19276 1240 19316 1280
rect 19468 1240 19508 1280
rect 17932 988 17972 1028
rect 17740 820 17780 860
rect 18316 904 18356 944
rect 19084 1156 19124 1196
rect 18892 1072 18932 1112
rect 18700 568 18740 608
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
<< metal3 >>
rect 2179 85912 2188 85952
rect 2228 85912 15140 85952
rect 15100 85868 15140 85912
rect 3715 85828 3724 85868
rect 3764 85828 9964 85868
rect 10004 85828 10013 85868
rect 15100 85828 16876 85868
rect 16916 85828 16925 85868
rect 0 85784 80 85804
rect 0 85744 268 85784
rect 308 85744 317 85784
rect 4291 85744 4300 85784
rect 4340 85744 9580 85784
rect 9620 85744 9629 85784
rect 0 85724 80 85744
rect 15715 85616 15773 85617
rect 13507 85576 13516 85616
rect 13556 85576 15724 85616
rect 15764 85576 15773 85616
rect 15715 85575 15773 85576
rect 0 85448 80 85468
rect 4771 85448 4829 85449
rect 0 85408 4780 85448
rect 4820 85408 4829 85448
rect 0 85388 80 85408
rect 4771 85407 4829 85408
rect 2659 85240 2668 85280
rect 2708 85240 3148 85280
rect 3188 85240 3197 85280
rect 10627 85240 10636 85280
rect 10676 85240 12076 85280
rect 12116 85240 12125 85280
rect 0 85112 80 85132
rect 1315 85112 1373 85113
rect 0 85072 1324 85112
rect 1364 85072 1373 85112
rect 0 85052 80 85072
rect 1315 85071 1373 85072
rect 19075 84988 19084 85028
rect 19124 84988 19660 85028
rect 19700 84988 19709 85028
rect 8227 84944 8285 84945
rect 15907 84944 15965 84945
rect 8227 84904 8236 84944
rect 8276 84904 8716 84944
rect 8756 84904 8765 84944
rect 9091 84904 9100 84944
rect 9140 84904 15916 84944
rect 15956 84904 15965 84944
rect 8227 84903 8285 84904
rect 15907 84903 15965 84904
rect 4195 84820 4204 84860
rect 4244 84820 4684 84860
rect 4724 84820 4733 84860
rect 0 84777 80 84796
rect 0 84776 125 84777
rect 0 84736 76 84776
rect 116 84736 125 84776
rect 14083 84736 14092 84776
rect 14132 84736 14476 84776
rect 14516 84736 14525 84776
rect 0 84735 125 84736
rect 0 84716 80 84735
rect 3679 84652 3688 84692
rect 3728 84652 3770 84692
rect 3810 84652 3852 84692
rect 3892 84652 3934 84692
rect 3974 84652 4016 84692
rect 4056 84652 4065 84692
rect 18799 84652 18808 84692
rect 18848 84652 18890 84692
rect 18930 84652 18972 84692
rect 19012 84652 19054 84692
rect 19094 84652 19136 84692
rect 19176 84652 19185 84692
rect 2947 84568 2956 84608
rect 2996 84568 3436 84608
rect 3476 84568 3485 84608
rect 5539 84524 5597 84525
rect 7363 84524 7421 84525
rect 12355 84524 12413 84525
rect 5539 84484 5548 84524
rect 5588 84484 6028 84524
rect 6068 84484 6077 84524
rect 6595 84484 6604 84524
rect 6644 84484 7372 84524
rect 7412 84484 7421 84524
rect 9859 84484 9868 84524
rect 9908 84484 12364 84524
rect 12404 84484 12413 84524
rect 5539 84483 5597 84484
rect 7363 84483 7421 84484
rect 12355 84483 12413 84484
rect 12835 84524 12893 84525
rect 12835 84484 12844 84524
rect 12884 84484 13708 84524
rect 13748 84484 13757 84524
rect 12835 84483 12893 84484
rect 0 84440 80 84460
rect 5827 84440 5885 84441
rect 0 84400 2092 84440
rect 2132 84400 2141 84440
rect 5251 84400 5260 84440
rect 5300 84400 5644 84440
rect 5684 84400 5693 84440
rect 5742 84400 5836 84440
rect 5876 84400 5885 84440
rect 0 84380 80 84400
rect 5827 84399 5885 84400
rect 6115 84440 6173 84441
rect 6403 84440 6461 84441
rect 6691 84440 6749 84441
rect 7171 84440 7229 84441
rect 9667 84440 9725 84441
rect 10243 84440 10301 84441
rect 6115 84400 6124 84440
rect 6164 84400 6220 84440
rect 6260 84400 6269 84440
rect 6403 84400 6412 84440
rect 6452 84400 6546 84440
rect 6691 84400 6700 84440
rect 6740 84400 6796 84440
rect 6836 84400 6845 84440
rect 6979 84400 6988 84440
rect 7028 84400 7180 84440
rect 7220 84400 7229 84440
rect 9582 84400 9676 84440
rect 9716 84400 9725 84440
rect 10158 84400 10252 84440
rect 10292 84400 10301 84440
rect 6115 84399 6173 84400
rect 6403 84399 6461 84400
rect 6691 84399 6749 84400
rect 7171 84399 7229 84400
rect 9667 84399 9725 84400
rect 10243 84399 10301 84400
rect 10435 84440 10493 84441
rect 11779 84440 11837 84441
rect 12931 84440 12989 84441
rect 13315 84440 13373 84441
rect 14083 84440 14141 84441
rect 16387 84440 16445 84441
rect 16867 84440 16925 84441
rect 10435 84400 10444 84440
rect 10484 84400 10578 84440
rect 11694 84400 11788 84440
rect 11828 84400 11837 84440
rect 12846 84400 12940 84440
rect 12980 84400 12989 84440
rect 13230 84400 13324 84440
rect 13364 84400 13373 84440
rect 13891 84400 13900 84440
rect 13940 84400 14092 84440
rect 14132 84400 14141 84440
rect 14755 84400 14764 84440
rect 14804 84400 15436 84440
rect 15476 84400 15485 84440
rect 16302 84400 16396 84440
rect 16436 84400 16445 84440
rect 16579 84400 16588 84440
rect 16628 84400 16876 84440
rect 16916 84400 16925 84440
rect 10435 84399 10493 84400
rect 11779 84399 11837 84400
rect 12931 84399 12989 84400
rect 13315 84399 13373 84400
rect 14083 84399 14141 84400
rect 16387 84399 16445 84400
rect 16867 84399 16925 84400
rect 3235 84356 3293 84357
rect 3150 84316 3244 84356
rect 3284 84316 3293 84356
rect 8323 84316 8332 84356
rect 8372 84316 8812 84356
rect 8852 84316 8861 84356
rect 14371 84316 14380 84356
rect 14420 84316 15052 84356
rect 15092 84316 15101 84356
rect 3235 84315 3293 84316
rect 1219 84272 1277 84273
rect 1219 84232 1228 84272
rect 1268 84232 5548 84272
rect 5588 84232 5597 84272
rect 13315 84232 13324 84272
rect 13364 84232 13996 84272
rect 14036 84232 14045 84272
rect 1219 84231 1277 84232
rect 3619 84148 3628 84188
rect 3668 84148 8332 84188
rect 8372 84148 8381 84188
rect 0 84104 80 84124
rect 0 84064 1324 84104
rect 1364 84064 1373 84104
rect 5059 84064 5068 84104
rect 5108 84064 10444 84104
rect 10484 84064 10493 84104
rect 0 84044 80 84064
rect 1795 83980 1804 84020
rect 1844 83980 6412 84020
rect 6452 83980 6461 84020
rect 4919 83896 4928 83936
rect 4968 83896 5010 83936
rect 5050 83896 5092 83936
rect 5132 83896 5174 83936
rect 5214 83896 5256 83936
rect 5296 83896 5305 83936
rect 20039 83896 20048 83936
rect 20088 83896 20130 83936
rect 20170 83896 20212 83936
rect 20252 83896 20294 83936
rect 20334 83896 20376 83936
rect 20416 83896 20425 83936
rect 2179 83812 2188 83852
rect 2228 83812 5548 83852
rect 5588 83812 5597 83852
rect 6211 83812 6220 83852
rect 6260 83812 7180 83852
rect 7220 83812 7229 83852
rect 17923 83812 17932 83852
rect 17972 83812 18412 83852
rect 18452 83812 18461 83852
rect 0 83768 80 83788
rect 0 83728 76 83768
rect 116 83728 125 83768
rect 3043 83728 3052 83768
rect 3092 83728 4300 83768
rect 4340 83728 4349 83768
rect 6979 83728 6988 83768
rect 7028 83728 7756 83768
rect 7796 83728 7805 83768
rect 8131 83728 8140 83768
rect 8180 83728 8428 83768
rect 8468 83728 8477 83768
rect 11299 83728 11308 83768
rect 11348 83728 11357 83768
rect 18307 83728 18316 83768
rect 18356 83728 18892 83768
rect 18932 83728 18941 83768
rect 0 83708 80 83728
rect 11308 83684 11348 83728
rect 5635 83644 5644 83684
rect 5684 83644 11348 83684
rect 1708 83560 13996 83600
rect 14036 83560 14045 83600
rect 1708 83516 1748 83560
rect 2947 83516 3005 83517
rect 4387 83516 4445 83517
rect 6019 83516 6077 83517
rect 7747 83516 7805 83517
rect 9763 83516 9821 83517
rect 11011 83516 11069 83517
rect 11683 83516 11741 83517
rect 18307 83516 18365 83517
rect 18595 83516 18653 83517
rect 19075 83516 19133 83517
rect 19555 83516 19613 83517
rect 1699 83476 1708 83516
rect 1748 83476 1757 83516
rect 2851 83476 2860 83516
rect 2900 83476 2956 83516
rect 2996 83476 3005 83516
rect 4302 83476 4396 83516
rect 4436 83476 4445 83516
rect 5731 83476 5740 83516
rect 5780 83476 6028 83516
rect 6068 83476 6077 83516
rect 7662 83476 7756 83516
rect 7796 83476 7805 83516
rect 9678 83476 9772 83516
rect 9812 83476 9821 83516
rect 10627 83476 10636 83516
rect 10676 83476 11020 83516
rect 11060 83476 11069 83516
rect 11491 83476 11500 83516
rect 11540 83476 11692 83516
rect 11732 83476 11741 83516
rect 13699 83476 13708 83516
rect 13748 83476 14284 83516
rect 14324 83476 14333 83516
rect 18115 83476 18124 83516
rect 18164 83476 18316 83516
rect 18356 83476 18365 83516
rect 18480 83476 18508 83516
rect 18548 83476 18604 83516
rect 18644 83476 18700 83516
rect 18740 83476 18749 83516
rect 18990 83476 19084 83516
rect 19124 83476 19133 83516
rect 19267 83476 19276 83516
rect 19316 83476 19468 83516
rect 19508 83476 19564 83516
rect 19604 83476 19613 83516
rect 2947 83475 3005 83476
rect 4387 83475 4445 83476
rect 6019 83475 6077 83476
rect 7747 83475 7805 83476
rect 9763 83475 9821 83476
rect 11011 83475 11069 83476
rect 11683 83475 11741 83476
rect 18307 83475 18365 83476
rect 18595 83475 18653 83476
rect 19075 83475 19133 83476
rect 19555 83475 19613 83476
rect 0 83432 80 83452
rect 7075 83432 7133 83433
rect 0 83392 7084 83432
rect 7124 83392 7133 83432
rect 7363 83392 7372 83432
rect 7412 83392 8524 83432
rect 8564 83392 8573 83432
rect 0 83372 80 83392
rect 7075 83391 7133 83392
rect 2563 83348 2621 83349
rect 13123 83348 13181 83349
rect 13987 83348 14045 83349
rect 14467 83348 14525 83349
rect 14659 83348 14717 83349
rect 15043 83348 15101 83349
rect 2563 83308 2572 83348
rect 2612 83308 3628 83348
rect 3668 83308 3677 83348
rect 4963 83308 4972 83348
rect 5012 83308 9004 83348
rect 9044 83308 9053 83348
rect 13038 83308 13132 83348
rect 13172 83308 13181 83348
rect 13891 83308 13900 83348
rect 13940 83308 13996 83348
rect 14036 83308 14045 83348
rect 14275 83308 14284 83348
rect 14324 83308 14476 83348
rect 14516 83308 14525 83348
rect 14574 83308 14668 83348
rect 14708 83308 14717 83348
rect 14958 83308 15052 83348
rect 15092 83308 15101 83348
rect 18787 83308 18796 83348
rect 18836 83308 19276 83348
rect 19316 83308 19325 83348
rect 2563 83307 2621 83308
rect 13123 83307 13181 83308
rect 13987 83307 14045 83308
rect 14467 83307 14525 83308
rect 14659 83307 14717 83308
rect 15043 83307 15101 83308
rect 7651 83264 7709 83265
rect 6787 83224 6796 83264
rect 6836 83224 7660 83264
rect 7700 83224 7709 83264
rect 8131 83224 8140 83264
rect 8180 83224 14572 83264
rect 14612 83224 14621 83264
rect 7651 83223 7709 83224
rect 10819 83180 10877 83181
rect 3679 83140 3688 83180
rect 3728 83140 3770 83180
rect 3810 83140 3852 83180
rect 3892 83140 3934 83180
rect 3974 83140 4016 83180
rect 4056 83140 4065 83180
rect 7459 83140 7468 83180
rect 7508 83140 8044 83180
rect 8084 83140 8093 83180
rect 10243 83140 10252 83180
rect 10292 83140 10828 83180
rect 10868 83140 10877 83180
rect 10819 83139 10877 83140
rect 12739 83180 12797 83181
rect 12739 83140 12748 83180
rect 12788 83140 13516 83180
rect 13556 83140 13565 83180
rect 18799 83140 18808 83180
rect 18848 83140 18890 83180
rect 18930 83140 18972 83180
rect 19012 83140 19054 83180
rect 19094 83140 19136 83180
rect 19176 83140 19185 83180
rect 12739 83139 12797 83140
rect 0 83096 80 83116
rect 1891 83096 1949 83097
rect 0 83056 1900 83096
rect 1940 83056 1949 83096
rect 6499 83056 6508 83096
rect 6548 83056 12364 83096
rect 12404 83056 12413 83096
rect 0 83036 80 83056
rect 1891 83055 1949 83056
rect 6883 82804 6892 82844
rect 6932 82804 7276 82844
rect 7316 82804 7325 82844
rect 0 82760 80 82780
rect 2467 82760 2525 82761
rect 0 82720 2476 82760
rect 2516 82720 2525 82760
rect 4099 82720 4108 82760
rect 4148 82720 7948 82760
rect 7988 82720 7997 82760
rect 0 82700 80 82720
rect 2467 82719 2525 82720
rect 1891 82676 1949 82677
rect 4108 82676 4148 82720
rect 1891 82636 1900 82676
rect 1940 82636 4148 82676
rect 1891 82635 1949 82636
rect 14179 82592 14237 82593
rect 17347 82592 17405 82593
rect 17731 82592 17789 82593
rect 2563 82552 2572 82592
rect 2612 82552 3148 82592
rect 3188 82552 4108 82592
rect 4148 82552 4157 82592
rect 14094 82552 14188 82592
rect 14228 82552 14237 82592
rect 17262 82552 17356 82592
rect 17396 82552 17405 82592
rect 17646 82552 17740 82592
rect 17780 82552 17789 82592
rect 14179 82551 14237 82552
rect 17347 82551 17405 82552
rect 17731 82551 17789 82552
rect 19459 82592 19517 82593
rect 19459 82552 19468 82592
rect 19508 82552 20044 82592
rect 20084 82552 20093 82592
rect 19459 82551 19517 82552
rect 4675 82468 4684 82508
rect 4724 82468 11596 82508
rect 11636 82468 11645 82508
rect 0 82424 80 82444
rect 4291 82424 4349 82425
rect 0 82384 4300 82424
rect 4340 82384 4349 82424
rect 4919 82384 4928 82424
rect 4968 82384 5010 82424
rect 5050 82384 5092 82424
rect 5132 82384 5174 82424
rect 5214 82384 5256 82424
rect 5296 82384 5305 82424
rect 20039 82384 20048 82424
rect 20088 82384 20130 82424
rect 20170 82384 20212 82424
rect 20252 82384 20294 82424
rect 20334 82384 20376 82424
rect 20416 82384 20425 82424
rect 0 82364 80 82384
rect 4291 82383 4349 82384
rect 1699 82216 1708 82256
rect 1748 82216 2476 82256
rect 2516 82216 2525 82256
rect 8899 82216 8908 82256
rect 8948 82216 9292 82256
rect 9332 82216 9341 82256
rect 0 82088 80 82108
rect 0 82048 1132 82088
rect 1172 82048 1181 82088
rect 3427 82048 3436 82088
rect 3476 82048 3724 82088
rect 3764 82048 3773 82088
rect 18691 82048 18700 82088
rect 18740 82048 19660 82088
rect 19700 82048 19709 82088
rect 0 82028 80 82048
rect 18403 82004 18461 82005
rect 1219 81964 1228 82004
rect 1268 81964 1804 82004
rect 1844 81964 1853 82004
rect 18403 81964 18412 82004
rect 18452 81964 18796 82004
rect 18836 81964 18845 82004
rect 18403 81963 18461 81964
rect 18115 81920 18173 81921
rect 18499 81920 18557 81921
rect 19267 81920 19325 81921
rect 3811 81880 3820 81920
rect 3860 81880 3869 81920
rect 6595 81880 6604 81920
rect 6644 81880 6653 81920
rect 13027 81880 13036 81920
rect 13076 81880 13085 81920
rect 14563 81880 14572 81920
rect 14612 81880 14621 81920
rect 18030 81880 18124 81920
rect 18164 81880 18173 81920
rect 18414 81880 18508 81920
rect 18548 81880 18557 81920
rect 19182 81880 19276 81920
rect 19316 81880 19325 81920
rect 0 81752 80 81772
rect 3820 81752 3860 81880
rect 6604 81836 6644 81880
rect 7555 81836 7613 81837
rect 13036 81836 13076 81880
rect 4099 81796 4108 81836
rect 4148 81796 4972 81836
rect 5012 81796 5021 81836
rect 6604 81796 7564 81836
rect 7604 81796 7613 81836
rect 9475 81796 9484 81836
rect 9524 81796 13076 81836
rect 13891 81836 13949 81837
rect 14572 81836 14612 81880
rect 18115 81879 18173 81880
rect 18499 81879 18557 81880
rect 19267 81879 19325 81880
rect 13891 81796 13900 81836
rect 13940 81796 14612 81836
rect 0 81712 2540 81752
rect 3427 81712 3436 81752
rect 3476 81712 3860 81752
rect 4972 81752 5012 81796
rect 7555 81795 7613 81796
rect 13891 81795 13949 81796
rect 4972 81712 6316 81752
rect 6356 81712 7372 81752
rect 7412 81712 7421 81752
rect 0 81692 80 81712
rect 2500 81500 2540 81712
rect 3679 81628 3688 81668
rect 3728 81628 3770 81668
rect 3810 81628 3852 81668
rect 3892 81628 3934 81668
rect 3974 81628 4016 81668
rect 4056 81628 4065 81668
rect 18799 81628 18808 81668
rect 18848 81628 18890 81668
rect 18930 81628 18972 81668
rect 19012 81628 19054 81668
rect 19094 81628 19136 81668
rect 19176 81628 19185 81668
rect 2500 81460 4012 81500
rect 4052 81460 4061 81500
rect 0 81416 80 81436
rect 0 81376 3148 81416
rect 3188 81376 3197 81416
rect 0 81356 80 81376
rect 7363 81292 7372 81332
rect 7412 81292 15628 81332
rect 15668 81292 15677 81332
rect 1219 81124 1228 81164
rect 1268 81124 1516 81164
rect 1556 81124 1565 81164
rect 0 81080 80 81100
rect 1603 81080 1661 81081
rect 0 81040 1612 81080
rect 1652 81040 1661 81080
rect 6979 81040 6988 81080
rect 7028 81040 7564 81080
rect 7604 81040 7613 81080
rect 0 81020 80 81040
rect 1603 81039 1661 81040
rect 4919 80872 4928 80912
rect 4968 80872 5010 80912
rect 5050 80872 5092 80912
rect 5132 80872 5174 80912
rect 5214 80872 5256 80912
rect 5296 80872 5305 80912
rect 20039 80872 20048 80912
rect 20088 80872 20130 80912
rect 20170 80872 20212 80912
rect 20252 80872 20294 80912
rect 20334 80872 20376 80912
rect 20416 80872 20425 80912
rect 0 80744 80 80764
rect 2755 80744 2813 80745
rect 0 80704 2668 80744
rect 2708 80704 2764 80744
rect 2804 80704 2813 80744
rect 0 80684 80 80704
rect 2755 80703 2813 80704
rect 1411 80620 1420 80660
rect 1460 80620 2860 80660
rect 2900 80620 2909 80660
rect 4963 80620 4972 80660
rect 5012 80620 5740 80660
rect 5780 80620 6796 80660
rect 6836 80620 6845 80660
rect 9187 80620 9196 80660
rect 9236 80620 11596 80660
rect 11636 80620 11645 80660
rect 1603 80576 1661 80577
rect 1518 80536 1612 80576
rect 1652 80536 1661 80576
rect 1603 80535 1661 80536
rect 2275 80576 2333 80577
rect 2467 80576 2525 80577
rect 2275 80536 2284 80576
rect 2324 80536 2476 80576
rect 2516 80536 6220 80576
rect 6260 80536 6269 80576
rect 8995 80536 9004 80576
rect 9044 80536 11980 80576
rect 12020 80536 12029 80576
rect 2275 80535 2333 80536
rect 2467 80535 2525 80536
rect 5443 80492 5501 80493
rect 1516 80452 1900 80492
rect 1940 80452 1949 80492
rect 4579 80452 4588 80492
rect 4628 80452 4972 80492
rect 5012 80452 5021 80492
rect 5443 80452 5452 80492
rect 5492 80452 6028 80492
rect 6068 80452 6077 80492
rect 0 80408 80 80428
rect 1516 80409 1556 80452
rect 5443 80451 5501 80452
rect 1507 80408 1565 80409
rect 6787 80408 6845 80409
rect 0 80368 1516 80408
rect 1556 80368 1565 80408
rect 1795 80368 1804 80408
rect 1844 80368 2572 80408
rect 2612 80368 3724 80408
rect 3764 80368 3773 80408
rect 5923 80368 5932 80408
rect 5972 80368 6796 80408
rect 6836 80368 10828 80408
rect 10868 80368 10877 80408
rect 0 80348 80 80368
rect 1507 80367 1565 80368
rect 6787 80367 6845 80368
rect 5155 80284 5164 80324
rect 5204 80284 5452 80324
rect 5492 80284 5501 80324
rect 3679 80116 3688 80156
rect 3728 80116 3770 80156
rect 3810 80116 3852 80156
rect 3892 80116 3934 80156
rect 3974 80116 4016 80156
rect 4056 80116 4065 80156
rect 18799 80116 18808 80156
rect 18848 80116 18890 80156
rect 18930 80116 18972 80156
rect 19012 80116 19054 80156
rect 19094 80116 19136 80156
rect 19176 80116 19185 80156
rect 0 80072 80 80092
rect 0 80032 3340 80072
rect 3380 80032 6412 80072
rect 6452 80032 6461 80072
rect 0 80012 80 80032
rect 835 79988 893 79989
rect 835 79948 844 79988
rect 884 79948 5548 79988
rect 5588 79948 5597 79988
rect 835 79947 893 79948
rect 5347 79820 5405 79821
rect 4099 79780 4108 79820
rect 4148 79780 5356 79820
rect 5396 79780 10156 79820
rect 10196 79780 10205 79820
rect 5347 79779 5405 79780
rect 0 79736 80 79756
rect 2275 79736 2333 79737
rect 4675 79736 4733 79737
rect 0 79696 364 79736
rect 404 79696 413 79736
rect 2275 79696 2284 79736
rect 2324 79696 2668 79736
rect 2708 79696 2717 79736
rect 4195 79696 4204 79736
rect 4244 79696 4684 79736
rect 4724 79696 4733 79736
rect 0 79676 80 79696
rect 2275 79695 2333 79696
rect 4675 79695 4733 79696
rect 8995 79652 9053 79653
rect 3715 79612 3724 79652
rect 3764 79612 4300 79652
rect 4340 79612 9004 79652
rect 9044 79612 9053 79652
rect 8995 79611 9053 79612
rect 12163 79568 12221 79569
rect 172 79528 12172 79568
rect 12212 79528 12221 79568
rect 0 79400 80 79420
rect 172 79400 212 79528
rect 12163 79527 12221 79528
rect 3139 79400 3197 79401
rect 0 79360 212 79400
rect 1219 79360 1228 79400
rect 1268 79360 1420 79400
rect 1460 79360 1469 79400
rect 3054 79360 3148 79400
rect 3188 79360 3197 79400
rect 4919 79360 4928 79400
rect 4968 79360 5010 79400
rect 5050 79360 5092 79400
rect 5132 79360 5174 79400
rect 5214 79360 5256 79400
rect 5296 79360 5305 79400
rect 5539 79360 5548 79400
rect 5588 79360 9676 79400
rect 9716 79360 9725 79400
rect 20039 79360 20048 79400
rect 20088 79360 20130 79400
rect 20170 79360 20212 79400
rect 20252 79360 20294 79400
rect 20334 79360 20376 79400
rect 20416 79360 20425 79400
rect 0 79340 80 79360
rect 3139 79359 3197 79360
rect 5443 79276 5452 79316
rect 5492 79276 7276 79316
rect 7316 79276 8044 79316
rect 8084 79276 8093 79316
rect 5923 79192 5932 79232
rect 5972 79192 7180 79232
rect 7220 79192 7229 79232
rect 7363 79192 7372 79232
rect 7412 79192 7948 79232
rect 7988 79192 7997 79232
rect 2371 79108 2380 79148
rect 2420 79108 2860 79148
rect 2900 79108 3188 79148
rect 5251 79108 5260 79148
rect 5300 79108 5548 79148
rect 5588 79108 5597 79148
rect 0 79064 80 79084
rect 3148 79064 3188 79108
rect 0 79024 2668 79064
rect 2708 79024 2717 79064
rect 3139 79024 3148 79064
rect 3188 79024 5452 79064
rect 5492 79024 5501 79064
rect 5827 79024 5836 79064
rect 5876 79024 6988 79064
rect 7028 79024 7037 79064
rect 7459 79024 7468 79064
rect 7508 79024 9196 79064
rect 9236 79024 10156 79064
rect 10196 79024 10540 79064
rect 10580 79024 15820 79064
rect 15860 79024 15869 79064
rect 0 79004 80 79024
rect 1891 78980 1949 78981
rect 1806 78940 1900 78980
rect 1940 78940 1949 78980
rect 1891 78939 1949 78940
rect 2500 78940 4204 78980
rect 4244 78940 8908 78980
rect 8948 78940 8957 78980
rect 1507 78896 1565 78897
rect 2500 78896 2540 78940
rect 1507 78856 1516 78896
rect 1556 78856 2540 78896
rect 2659 78856 2668 78896
rect 2708 78856 4492 78896
rect 4532 78856 4876 78896
rect 4916 78856 4925 78896
rect 5827 78856 5836 78896
rect 5876 78856 8140 78896
rect 8180 78856 8189 78896
rect 1507 78855 1565 78856
rect 6979 78772 6988 78812
rect 7028 78772 7852 78812
rect 7892 78772 7901 78812
rect 9955 78772 9964 78812
rect 10004 78772 10348 78812
rect 10388 78772 10397 78812
rect 0 78728 80 78748
rect 0 78688 212 78728
rect 0 78668 80 78688
rect 172 78560 212 78688
rect 3679 78604 3688 78644
rect 3728 78604 3770 78644
rect 3810 78604 3852 78644
rect 3892 78604 3934 78644
rect 3974 78604 4016 78644
rect 4056 78604 4065 78644
rect 18799 78604 18808 78644
rect 18848 78604 18890 78644
rect 18930 78604 18972 78644
rect 19012 78604 19054 78644
rect 19094 78604 19136 78644
rect 19176 78604 19185 78644
rect 21424 78560 21504 78580
rect 172 78520 5260 78560
rect 5300 78520 5309 78560
rect 8323 78520 8332 78560
rect 8372 78520 11308 78560
rect 11348 78520 11357 78560
rect 20803 78520 20812 78560
rect 20852 78520 21504 78560
rect 21424 78500 21504 78520
rect 3907 78436 3916 78476
rect 3956 78436 11020 78476
rect 11060 78436 11069 78476
rect 0 78392 80 78412
rect 0 78352 2572 78392
rect 2612 78352 2621 78392
rect 5347 78352 5356 78392
rect 5396 78352 5644 78392
rect 5684 78352 5693 78392
rect 0 78332 80 78352
rect 3139 78224 3197 78225
rect 3139 78184 3148 78224
rect 3188 78184 3340 78224
rect 3380 78184 3389 78224
rect 7171 78184 7180 78224
rect 7220 78184 7468 78224
rect 7508 78184 7948 78224
rect 7988 78184 7997 78224
rect 8803 78184 8812 78224
rect 8852 78184 9484 78224
rect 9524 78184 9533 78224
rect 3139 78183 3197 78184
rect 7459 78140 7517 78141
rect 1795 78100 1804 78140
rect 1844 78100 2668 78140
rect 2708 78100 2717 78140
rect 4867 78100 4876 78140
rect 4916 78100 7468 78140
rect 7508 78100 7517 78140
rect 7459 78099 7517 78100
rect 0 78056 80 78076
rect 0 78016 2956 78056
rect 2996 78016 3148 78056
rect 3188 78016 3197 78056
rect 4291 78016 4300 78056
rect 4340 78016 4972 78056
rect 5012 78016 5021 78056
rect 0 77996 80 78016
rect 4195 77972 4253 77973
rect 3331 77932 3340 77972
rect 3380 77932 4204 77972
rect 4244 77932 9292 77972
rect 9332 77932 9341 77972
rect 4195 77931 4253 77932
rect 21187 77888 21245 77889
rect 21424 77888 21504 77908
rect 4919 77848 4928 77888
rect 4968 77848 5010 77888
rect 5050 77848 5092 77888
rect 5132 77848 5174 77888
rect 5214 77848 5256 77888
rect 5296 77848 5305 77888
rect 20039 77848 20048 77888
rect 20088 77848 20130 77888
rect 20170 77848 20212 77888
rect 20252 77848 20294 77888
rect 20334 77848 20376 77888
rect 20416 77848 20425 77888
rect 21187 77848 21196 77888
rect 21236 77848 21504 77888
rect 21187 77847 21245 77848
rect 21424 77828 21504 77848
rect 0 77720 80 77740
rect 3331 77720 3389 77721
rect 0 77680 3340 77720
rect 3380 77680 3389 77720
rect 6019 77680 6028 77720
rect 6068 77680 6604 77720
rect 6644 77680 6653 77720
rect 0 77660 80 77680
rect 3331 77679 3389 77680
rect 3427 77596 3436 77636
rect 3476 77596 4204 77636
rect 4244 77596 4253 77636
rect 2947 77552 3005 77553
rect 2862 77512 2956 77552
rect 2996 77512 3005 77552
rect 2947 77511 3005 77512
rect 4771 77552 4829 77553
rect 4771 77512 4780 77552
rect 4820 77512 5260 77552
rect 5300 77512 6028 77552
rect 6068 77512 6077 77552
rect 6403 77512 6412 77552
rect 6452 77512 6892 77552
rect 6932 77512 6941 77552
rect 7843 77512 7852 77552
rect 7892 77512 8524 77552
rect 8564 77512 8573 77552
rect 4771 77511 4829 77512
rect 3427 77468 3485 77469
rect 3342 77428 3436 77468
rect 3476 77428 3485 77468
rect 8323 77428 8332 77468
rect 8372 77428 8716 77468
rect 8756 77428 9004 77468
rect 9044 77428 9053 77468
rect 3427 77427 3485 77428
rect 0 77384 80 77404
rect 0 77344 212 77384
rect 0 77324 80 77344
rect 172 77216 212 77344
rect 7459 77260 7468 77300
rect 7508 77260 8428 77300
rect 8468 77260 8477 77300
rect 21424 77217 21504 77236
rect 21379 77216 21504 77217
rect 172 77176 6700 77216
rect 6740 77176 6749 77216
rect 7267 77176 7276 77216
rect 7316 77176 8332 77216
rect 8372 77176 8381 77216
rect 21379 77176 21388 77216
rect 21428 77176 21504 77216
rect 21379 77175 21504 77176
rect 21424 77156 21504 77175
rect 3679 77092 3688 77132
rect 3728 77092 3770 77132
rect 3810 77092 3852 77132
rect 3892 77092 3934 77132
rect 3974 77092 4016 77132
rect 4056 77092 4065 77132
rect 18799 77092 18808 77132
rect 18848 77092 18890 77132
rect 18930 77092 18972 77132
rect 19012 77092 19054 77132
rect 19094 77092 19136 77132
rect 19176 77092 19185 77132
rect 0 77048 80 77068
rect 0 77008 7276 77048
rect 7316 77008 7325 77048
rect 0 76988 80 77008
rect 6499 76964 6557 76965
rect 6414 76924 6508 76964
rect 6548 76924 6557 76964
rect 6499 76923 6557 76924
rect 4579 76880 4637 76881
rect 4494 76840 4588 76880
rect 4628 76840 4637 76880
rect 6307 76840 6316 76880
rect 6356 76840 7084 76880
rect 7124 76840 7133 76880
rect 8803 76840 8812 76880
rect 8852 76840 9484 76880
rect 9524 76840 9533 76880
rect 12355 76840 12364 76880
rect 12404 76840 12844 76880
rect 12884 76840 12893 76880
rect 4579 76839 4637 76840
rect 2275 76756 2284 76796
rect 2324 76756 2476 76796
rect 2516 76756 3340 76796
rect 3380 76756 4492 76796
rect 4532 76756 5644 76796
rect 5684 76756 5693 76796
rect 6211 76756 6220 76796
rect 6260 76756 7756 76796
rect 7796 76756 7948 76796
rect 7988 76756 11212 76796
rect 11252 76756 11261 76796
rect 11395 76756 11404 76796
rect 11444 76756 12940 76796
rect 12980 76756 12989 76796
rect 0 76712 80 76732
rect 1987 76712 2045 76713
rect 0 76672 1996 76712
rect 2036 76672 2045 76712
rect 4099 76672 4108 76712
rect 4148 76672 4396 76712
rect 4436 76672 4445 76712
rect 5347 76672 5356 76712
rect 5396 76672 6124 76712
rect 6164 76672 6508 76712
rect 6548 76672 6557 76712
rect 8227 76672 8236 76712
rect 8276 76672 8908 76712
rect 8948 76672 8957 76712
rect 0 76652 80 76672
rect 1987 76671 2045 76672
rect 8803 76628 8861 76629
rect 5644 76588 6028 76628
rect 6068 76588 8812 76628
rect 8852 76588 9868 76628
rect 9908 76588 9917 76628
rect 3523 76544 3581 76545
rect 5644 76544 5684 76588
rect 8803 76587 8861 76588
rect 21424 76544 21504 76564
rect 3438 76504 3532 76544
rect 3572 76504 3581 76544
rect 5635 76504 5644 76544
rect 5684 76504 5693 76544
rect 5827 76504 5836 76544
rect 5876 76504 6220 76544
rect 6260 76504 6269 76544
rect 6595 76504 6604 76544
rect 6644 76504 6653 76544
rect 8419 76504 8428 76544
rect 8468 76504 8620 76544
rect 8660 76504 8669 76544
rect 20515 76504 20524 76544
rect 20564 76504 21504 76544
rect 3523 76503 3581 76504
rect 0 76376 80 76396
rect 0 76336 172 76376
rect 212 76336 221 76376
rect 4919 76336 4928 76376
rect 4968 76336 5010 76376
rect 5050 76336 5092 76376
rect 5132 76336 5174 76376
rect 5214 76336 5256 76376
rect 5296 76336 5305 76376
rect 0 76316 80 76336
rect 2179 76252 2188 76292
rect 2228 76252 3244 76292
rect 3284 76252 3293 76292
rect 5443 76252 5452 76292
rect 5492 76252 5501 76292
rect 5452 76208 5492 76252
rect 6604 76208 6644 76504
rect 21424 76484 21504 76504
rect 6691 76420 6700 76460
rect 6740 76420 6749 76460
rect 6700 76292 6740 76420
rect 20039 76336 20048 76376
rect 20088 76336 20130 76376
rect 20170 76336 20212 76376
rect 20252 76336 20294 76376
rect 20334 76336 20376 76376
rect 20416 76336 20425 76376
rect 6700 76252 6836 76292
rect 5452 76168 5740 76208
rect 5780 76168 5789 76208
rect 6604 76168 6700 76208
rect 6740 76168 6749 76208
rect 6796 76124 6836 76252
rect 7747 76168 7756 76208
rect 7796 76168 7805 76208
rect 6595 76084 6604 76124
rect 6644 76084 6836 76124
rect 0 76040 80 76060
rect 355 76040 413 76041
rect 1795 76040 1853 76041
rect 0 76000 364 76040
rect 404 76000 413 76040
rect 1603 76000 1612 76040
rect 1652 76000 1804 76040
rect 1844 76000 1853 76040
rect 4387 76000 4396 76040
rect 4436 76000 5068 76040
rect 5108 76000 5117 76040
rect 6499 76000 6508 76040
rect 6548 76000 6988 76040
rect 7028 76000 7037 76040
rect 7171 76000 7180 76040
rect 7220 76000 7468 76040
rect 7508 76000 7517 76040
rect 0 75980 80 76000
rect 355 75999 413 76000
rect 1795 75999 1853 76000
rect 4579 75956 4637 75957
rect 1795 75916 1804 75956
rect 1844 75916 2188 75956
rect 2228 75916 2237 75956
rect 2563 75916 2572 75956
rect 2612 75916 4588 75956
rect 4628 75916 4637 75956
rect 4579 75915 4637 75916
rect 4771 75956 4829 75957
rect 4771 75916 4780 75956
rect 4820 75916 5452 75956
rect 5492 75916 5501 75956
rect 4771 75915 4829 75916
rect 7756 75872 7796 76168
rect 9667 76084 9676 76124
rect 9716 76084 11020 76124
rect 11060 76084 11069 76124
rect 8227 76000 8236 76040
rect 8276 76000 8524 76040
rect 8564 76000 8573 76040
rect 11203 76000 11212 76040
rect 11252 76000 11261 76040
rect 8515 75956 8573 75957
rect 8515 75916 8524 75956
rect 8564 75916 8620 75956
rect 8660 75916 8908 75956
rect 8948 75916 8957 75956
rect 8515 75915 8573 75916
rect 11212 75872 11252 76000
rect 21424 75872 21504 75892
rect 4963 75832 4972 75872
rect 5012 75832 7372 75872
rect 7412 75832 7421 75872
rect 7555 75832 7564 75872
rect 7604 75832 7796 75872
rect 10339 75832 10348 75872
rect 10388 75832 11252 75872
rect 20899 75832 20908 75872
rect 20948 75832 21504 75872
rect 21424 75812 21504 75832
rect 5539 75748 5548 75788
rect 5588 75748 8812 75788
rect 8852 75748 8861 75788
rect 0 75704 80 75724
rect 7459 75704 7517 75705
rect 0 75664 7361 75704
rect 7401 75664 7410 75704
rect 7459 75664 7468 75704
rect 7508 75664 7564 75704
rect 7604 75664 7613 75704
rect 9091 75664 9100 75704
rect 9140 75664 15340 75704
rect 15380 75664 15389 75704
rect 0 75644 80 75664
rect 7459 75663 7517 75664
rect 6499 75620 6557 75621
rect 9571 75620 9629 75621
rect 3679 75580 3688 75620
rect 3728 75580 3770 75620
rect 3810 75580 3852 75620
rect 3892 75580 3934 75620
rect 3974 75580 4016 75620
rect 4056 75580 4065 75620
rect 4867 75580 4876 75620
rect 4916 75580 5644 75620
rect 5684 75580 5693 75620
rect 6414 75580 6508 75620
rect 6548 75580 6557 75620
rect 6979 75580 6988 75620
rect 7028 75580 7468 75620
rect 7508 75580 7517 75620
rect 9187 75580 9196 75620
rect 9236 75580 9580 75620
rect 9620 75580 9629 75620
rect 6499 75579 6557 75580
rect 9571 75579 9629 75580
rect 10627 75620 10685 75621
rect 10627 75580 10636 75620
rect 10676 75580 10828 75620
rect 10868 75580 11404 75620
rect 11444 75580 11453 75620
rect 18799 75580 18808 75620
rect 18848 75580 18890 75620
rect 18930 75580 18972 75620
rect 19012 75580 19054 75620
rect 19094 75580 19136 75620
rect 19176 75580 19185 75620
rect 10627 75579 10685 75580
rect 2500 75496 4780 75536
rect 4820 75496 4829 75536
rect 5443 75496 5452 75536
rect 5492 75496 5501 75536
rect 9091 75496 9100 75536
rect 9140 75496 11500 75536
rect 11540 75496 11549 75536
rect 2500 75452 2540 75496
rect 5452 75452 5492 75496
rect 11299 75452 11357 75453
rect 1891 75412 1900 75452
rect 1940 75412 2092 75452
rect 2132 75412 2540 75452
rect 3715 75412 3724 75452
rect 3764 75412 5356 75452
rect 5396 75412 5405 75452
rect 5452 75412 11308 75452
rect 11348 75412 11788 75452
rect 11828 75412 11837 75452
rect 11299 75411 11357 75412
rect 0 75368 80 75388
rect 0 75328 5644 75368
rect 5684 75328 5693 75368
rect 0 75308 80 75328
rect 3139 75284 3197 75285
rect 9187 75284 9245 75285
rect 3043 75244 3052 75284
rect 3092 75244 3148 75284
rect 3188 75244 9196 75284
rect 9236 75244 9245 75284
rect 3139 75243 3197 75244
rect 9187 75243 9245 75244
rect 10435 75284 10493 75285
rect 10435 75244 10444 75284
rect 10484 75244 11308 75284
rect 11348 75244 11357 75284
rect 10435 75243 10493 75244
rect 11011 75200 11069 75201
rect 21424 75200 21504 75220
rect 2371 75160 2380 75200
rect 2420 75160 2764 75200
rect 2804 75160 2813 75200
rect 5251 75160 5260 75200
rect 5300 75160 6220 75200
rect 6260 75160 6269 75200
rect 10915 75160 10924 75200
rect 10964 75160 11020 75200
rect 11060 75160 11069 75200
rect 21379 75160 21388 75200
rect 21428 75160 21504 75200
rect 11011 75159 11069 75160
rect 21424 75140 21504 75160
rect 6019 75116 6077 75117
rect 451 75076 460 75116
rect 500 75076 940 75116
rect 980 75076 4052 75116
rect 5934 75076 6028 75116
rect 6068 75076 6077 75116
rect 9091 75076 9100 75116
rect 9140 75076 9149 75116
rect 10531 75076 10540 75116
rect 10580 75076 10828 75116
rect 10868 75076 10877 75116
rect 0 75032 80 75052
rect 0 74992 2540 75032
rect 0 74972 80 74992
rect 2500 74864 2540 74992
rect 1411 74824 1420 74864
rect 1460 74824 1804 74864
rect 1844 74824 1853 74864
rect 2500 74824 2572 74864
rect 2612 74824 2621 74864
rect 4012 74780 4052 75076
rect 6019 75075 6077 75076
rect 9100 75032 9140 75076
rect 4099 74992 4108 75032
rect 4148 74992 4396 75032
rect 4436 74992 9140 75032
rect 8899 74948 8957 74949
rect 4771 74908 4780 74948
rect 4820 74908 8908 74948
rect 8948 74908 8957 74948
rect 8899 74907 8957 74908
rect 9187 74948 9245 74949
rect 9187 74908 9196 74948
rect 9236 74908 11404 74948
rect 11444 74908 11453 74948
rect 9187 74907 9245 74908
rect 4919 74824 4928 74864
rect 4968 74824 5010 74864
rect 5050 74824 5092 74864
rect 5132 74824 5174 74864
rect 5214 74824 5256 74864
rect 5296 74824 5305 74864
rect 5827 74824 5836 74864
rect 5876 74824 10156 74864
rect 10196 74824 10205 74864
rect 20039 74824 20048 74864
rect 20088 74824 20130 74864
rect 20170 74824 20212 74864
rect 20252 74824 20294 74864
rect 20334 74824 20376 74864
rect 20416 74824 20425 74864
rect 10147 74780 10205 74781
rect 1699 74740 1708 74780
rect 1748 74740 2860 74780
rect 2900 74740 2909 74780
rect 4012 74740 5452 74780
rect 5492 74740 5740 74780
rect 5780 74740 5789 74780
rect 6316 74740 10156 74780
rect 10196 74740 10205 74780
rect 0 74696 80 74716
rect 6316 74696 6356 74740
rect 10147 74739 10205 74740
rect 9379 74696 9437 74697
rect 0 74656 6356 74696
rect 7555 74656 7564 74696
rect 7604 74656 8716 74696
rect 8756 74656 9388 74696
rect 9428 74656 9437 74696
rect 10339 74656 10348 74696
rect 10388 74656 11788 74696
rect 11828 74656 12556 74696
rect 12596 74656 12605 74696
rect 0 74636 80 74656
rect 9379 74655 9437 74656
rect 8803 74612 8861 74613
rect 9283 74612 9341 74613
rect 2659 74572 2668 74612
rect 2708 74572 3052 74612
rect 3092 74572 3101 74612
rect 5356 74572 5548 74612
rect 5588 74572 5597 74612
rect 8611 74572 8620 74612
rect 8660 74572 8812 74612
rect 8852 74572 9292 74612
rect 9332 74572 9341 74612
rect 9859 74572 9868 74612
rect 9908 74572 10252 74612
rect 10292 74572 10301 74612
rect 1411 74488 1420 74528
rect 1460 74488 2540 74528
rect 2851 74488 2860 74528
rect 2900 74488 3244 74528
rect 3284 74488 3293 74528
rect 4099 74488 4108 74528
rect 4148 74488 4157 74528
rect 2500 74444 2540 74488
rect 4108 74444 4148 74488
rect 2500 74404 2764 74444
rect 2804 74404 3052 74444
rect 3092 74404 4148 74444
rect 0 74360 80 74380
rect 5356 74360 5396 74572
rect 8803 74571 8861 74572
rect 9283 74571 9341 74572
rect 6019 74528 6077 74529
rect 21424 74528 21504 74548
rect 5443 74488 5452 74528
rect 5492 74488 6028 74528
rect 6068 74488 6077 74528
rect 8035 74488 8044 74528
rect 8084 74488 9676 74528
rect 9716 74488 9725 74528
rect 20707 74488 20716 74528
rect 20756 74488 21504 74528
rect 6019 74487 6077 74488
rect 21424 74468 21504 74488
rect 8803 74444 8861 74445
rect 6403 74404 6412 74444
rect 6452 74404 8812 74444
rect 8852 74404 8861 74444
rect 8803 74403 8861 74404
rect 6979 74360 7037 74361
rect 8899 74360 8957 74361
rect 10627 74360 10685 74361
rect 0 74320 556 74360
rect 596 74320 605 74360
rect 1603 74320 1612 74360
rect 1652 74320 3532 74360
rect 3572 74320 3581 74360
rect 3628 74320 3724 74360
rect 3764 74320 3773 74360
rect 5356 74320 5492 74360
rect 5539 74320 5548 74360
rect 5588 74320 6988 74360
rect 7028 74320 7037 74360
rect 8227 74320 8236 74360
rect 8276 74320 8716 74360
rect 8756 74320 8765 74360
rect 8899 74320 8908 74360
rect 8948 74320 9100 74360
rect 9140 74320 9149 74360
rect 9283 74320 9292 74360
rect 9332 74320 9964 74360
rect 10004 74320 10013 74360
rect 10627 74320 10636 74360
rect 10676 74320 10732 74360
rect 10772 74320 10781 74360
rect 0 74300 80 74320
rect 1219 74236 1228 74276
rect 1268 74236 1708 74276
rect 1748 74236 1757 74276
rect 2755 74236 2764 74276
rect 2804 74236 3436 74276
rect 3476 74236 3485 74276
rect 3628 74192 3668 74320
rect 4099 74276 4157 74277
rect 5452 74276 5492 74320
rect 6979 74319 7037 74320
rect 8899 74319 8957 74320
rect 10627 74319 10685 74320
rect 4099 74236 4108 74276
rect 4148 74236 4300 74276
rect 4340 74236 4349 74276
rect 5443 74236 5452 74276
rect 5492 74236 5501 74276
rect 6403 74236 6412 74276
rect 6452 74236 6892 74276
rect 6932 74236 6941 74276
rect 7843 74236 7852 74276
rect 7892 74236 8812 74276
rect 8852 74236 9196 74276
rect 9236 74236 10060 74276
rect 10100 74236 10109 74276
rect 4099 74235 4157 74236
rect 2851 74152 2860 74192
rect 2900 74152 3668 74192
rect 6787 74152 6796 74192
rect 6836 74152 7468 74192
rect 7508 74152 7756 74192
rect 7796 74152 7805 74192
rect 3679 74068 3688 74108
rect 3728 74068 3770 74108
rect 3810 74068 3852 74108
rect 3892 74068 3934 74108
rect 3974 74068 4016 74108
rect 4056 74068 4065 74108
rect 6883 74068 6892 74108
rect 6932 74068 7372 74108
rect 7412 74068 7421 74108
rect 18799 74068 18808 74108
rect 18848 74068 18890 74108
rect 18930 74068 18972 74108
rect 19012 74068 19054 74108
rect 19094 74068 19136 74108
rect 19176 74068 19185 74108
rect 0 74024 80 74044
rect 0 73984 1324 74024
rect 1364 73984 1373 74024
rect 0 73964 80 73984
rect 1987 73900 1996 73940
rect 2036 73900 2188 73940
rect 2228 73900 2237 73940
rect 5347 73900 5356 73940
rect 5396 73900 5836 73940
rect 5876 73900 6796 73940
rect 6836 73900 6845 73940
rect 10243 73900 10252 73940
rect 10292 73900 10828 73940
rect 10868 73900 10877 73940
rect 2467 73856 2525 73857
rect 9955 73856 10013 73857
rect 1516 73816 1900 73856
rect 1940 73816 1949 73856
rect 2275 73816 2284 73856
rect 2324 73816 2476 73856
rect 2516 73816 2525 73856
rect 9475 73816 9484 73856
rect 9524 73816 9964 73856
rect 10004 73816 10013 73856
rect 0 73688 80 73708
rect 1516 73688 1556 73816
rect 2467 73815 2525 73816
rect 9955 73815 10013 73816
rect 16291 73856 16349 73857
rect 21424 73856 21504 73876
rect 16291 73816 16300 73856
rect 16340 73816 21504 73856
rect 16291 73815 16349 73816
rect 21424 73796 21504 73816
rect 2563 73732 2572 73772
rect 2612 73732 5260 73772
rect 5300 73732 6412 73772
rect 6452 73732 6461 73772
rect 8515 73732 8524 73772
rect 8564 73732 9580 73772
rect 9620 73732 10060 73772
rect 10100 73732 10109 73772
rect 6979 73688 7037 73689
rect 0 73648 1556 73688
rect 1603 73648 1612 73688
rect 1652 73648 2380 73688
rect 2420 73648 2429 73688
rect 6499 73648 6508 73688
rect 6548 73648 6557 73688
rect 6979 73648 6988 73688
rect 7028 73648 7180 73688
rect 7220 73648 7229 73688
rect 9379 73648 9388 73688
rect 9428 73648 10156 73688
rect 10196 73648 10205 73688
rect 10339 73648 10348 73688
rect 10388 73648 10540 73688
rect 10580 73648 10589 73688
rect 11320 73648 11596 73688
rect 11636 73648 12268 73688
rect 12308 73648 12317 73688
rect 0 73628 80 73648
rect 6508 73604 6548 73648
rect 6979 73647 7037 73648
rect 11320 73604 11360 73648
rect 3139 73564 3148 73604
rect 3188 73564 3380 73604
rect 6508 73564 11360 73604
rect 3340 73520 3380 73564
rect 6499 73520 6557 73521
rect 1315 73480 1324 73520
rect 1364 73480 1804 73520
rect 1844 73480 1853 73520
rect 3331 73480 3340 73520
rect 3380 73480 3389 73520
rect 6414 73480 6508 73520
rect 6548 73480 6557 73520
rect 9667 73480 9676 73520
rect 9716 73480 10060 73520
rect 10100 73480 10109 73520
rect 6499 73479 6557 73480
rect 1507 73396 1516 73436
rect 1556 73396 2540 73436
rect 2947 73396 2956 73436
rect 2996 73396 3148 73436
rect 3188 73396 3197 73436
rect 6307 73396 6316 73436
rect 6356 73396 7281 73436
rect 7321 73396 7660 73436
rect 7700 73396 7709 73436
rect 0 73352 80 73372
rect 2500 73352 2540 73396
rect 0 73312 1132 73352
rect 1172 73312 1181 73352
rect 2500 73312 4684 73352
rect 4724 73312 4733 73352
rect 4919 73312 4928 73352
rect 4968 73312 5010 73352
rect 5050 73312 5092 73352
rect 5132 73312 5174 73352
rect 5214 73312 5256 73352
rect 5296 73312 5305 73352
rect 6595 73312 6604 73352
rect 6644 73312 7180 73352
rect 7220 73312 7229 73352
rect 8035 73312 8044 73352
rect 8084 73312 9484 73352
rect 9524 73312 11020 73352
rect 11060 73312 11308 73352
rect 11348 73312 11357 73352
rect 20039 73312 20048 73352
rect 20088 73312 20130 73352
rect 20170 73312 20212 73352
rect 20252 73312 20294 73352
rect 20334 73312 20376 73352
rect 20416 73312 20425 73352
rect 0 73292 80 73312
rect 6499 73228 6508 73268
rect 6548 73228 7084 73268
rect 7124 73228 7133 73268
rect 21424 73184 21504 73204
rect 3043 73144 3052 73184
rect 3092 73144 3101 73184
rect 6595 73144 6604 73184
rect 6644 73144 6653 73184
rect 10243 73144 10252 73184
rect 10292 73144 10732 73184
rect 10772 73144 10781 73184
rect 11320 73144 11596 73184
rect 11636 73144 11645 73184
rect 20995 73144 21004 73184
rect 21044 73144 21504 73184
rect 0 73016 80 73036
rect 1699 73016 1757 73017
rect 2275 73016 2333 73017
rect 0 72976 212 73016
rect 1219 72976 1228 73016
rect 1268 72976 1708 73016
rect 1748 72976 2284 73016
rect 2324 72976 2333 73016
rect 0 72956 80 72976
rect 172 72848 212 72976
rect 1699 72975 1757 72976
rect 2275 72975 2333 72976
rect 2467 73016 2525 73017
rect 3052 73016 3092 73144
rect 3523 73100 3581 73101
rect 3438 73060 3532 73100
rect 3572 73060 3581 73100
rect 3523 73059 3581 73060
rect 3139 73016 3197 73017
rect 6604 73016 6644 73144
rect 8620 73060 8716 73100
rect 8756 73060 8765 73100
rect 8620 73016 8660 73060
rect 2467 72976 2476 73016
rect 2516 72976 2610 73016
rect 3052 72976 3148 73016
rect 3188 72976 3197 73016
rect 4483 72976 4492 73016
rect 4532 72976 4541 73016
rect 6604 72976 8660 73016
rect 2467 72975 2525 72976
rect 3139 72975 3197 72976
rect 4492 72932 4532 72976
rect 11320 72932 11360 73144
rect 21424 73124 21504 73144
rect 11875 72976 11884 73016
rect 11924 72976 12172 73016
rect 12212 72976 12221 73016
rect 259 72892 268 72932
rect 308 72892 1036 72932
rect 1076 72892 4532 72932
rect 8803 72892 8812 72932
rect 8852 72892 9100 72932
rect 9140 72892 9149 72932
rect 10924 72892 11360 72932
rect 172 72808 9196 72848
rect 9236 72808 9245 72848
rect 10723 72764 10781 72765
rect 10924 72764 10964 72892
rect 355 72724 364 72764
rect 404 72724 1748 72764
rect 2851 72724 2860 72764
rect 2900 72724 3436 72764
rect 3476 72724 3485 72764
rect 5923 72724 5932 72764
rect 5972 72724 6316 72764
rect 6356 72724 6365 72764
rect 10638 72724 10732 72764
rect 10772 72724 10781 72764
rect 10915 72724 10924 72764
rect 10964 72724 10973 72764
rect 11875 72724 11884 72764
rect 11924 72724 12364 72764
rect 12404 72724 12413 72764
rect 0 72680 80 72700
rect 1708 72680 1748 72724
rect 10723 72723 10781 72724
rect 0 72640 1612 72680
rect 1652 72640 1661 72680
rect 1708 72640 6892 72680
rect 6932 72640 10828 72680
rect 10868 72640 10877 72680
rect 0 72620 80 72640
rect 3523 72596 3581 72597
rect 3331 72556 3340 72596
rect 3380 72556 3532 72596
rect 3572 72556 3581 72596
rect 3679 72556 3688 72596
rect 3728 72556 3770 72596
rect 3810 72556 3852 72596
rect 3892 72556 3934 72596
rect 3974 72556 4016 72596
rect 4056 72556 4065 72596
rect 5731 72556 5740 72596
rect 5780 72556 5972 72596
rect 3523 72555 3581 72556
rect 451 72512 509 72513
rect 451 72472 460 72512
rect 500 72472 5836 72512
rect 5876 72472 5885 72512
rect 451 72471 509 72472
rect 5932 72428 5972 72556
rect 7756 72556 9292 72596
rect 9332 72556 9341 72596
rect 18799 72556 18808 72596
rect 18848 72556 18890 72596
rect 18930 72556 18972 72596
rect 19012 72556 19054 72596
rect 19094 72556 19136 72596
rect 19176 72556 19185 72596
rect 7756 72513 7796 72556
rect 7747 72512 7805 72513
rect 8899 72512 8957 72513
rect 21424 72512 21504 72532
rect 6115 72472 6124 72512
rect 6164 72472 7756 72512
rect 7796 72472 7805 72512
rect 8707 72472 8716 72512
rect 8756 72472 8908 72512
rect 8948 72472 8957 72512
rect 7747 72471 7805 72472
rect 8899 72471 8957 72472
rect 11320 72472 21504 72512
rect 8419 72428 8477 72429
rect 11320 72428 11360 72472
rect 21424 72452 21504 72472
rect 1036 72388 2956 72428
rect 2996 72388 3005 72428
rect 3235 72388 3244 72428
rect 3284 72388 4588 72428
rect 4628 72388 4637 72428
rect 5923 72388 5932 72428
rect 5972 72388 7180 72428
rect 7220 72388 7229 72428
rect 8419 72388 8428 72428
rect 8468 72388 11360 72428
rect 0 72344 80 72364
rect 1036 72344 1076 72388
rect 8419 72387 8477 72388
rect 8803 72344 8861 72345
rect 0 72304 1076 72344
rect 1123 72304 1132 72344
rect 1172 72304 6932 72344
rect 7939 72304 7948 72344
rect 7988 72304 8332 72344
rect 8372 72304 8381 72344
rect 8803 72304 8812 72344
rect 8852 72304 9004 72344
rect 9044 72304 9053 72344
rect 9187 72304 9196 72344
rect 9236 72304 9245 72344
rect 9379 72304 9388 72344
rect 9428 72304 9868 72344
rect 9908 72304 9917 72344
rect 14275 72304 14284 72344
rect 14324 72304 15052 72344
rect 15092 72304 16780 72344
rect 16820 72304 16829 72344
rect 0 72284 80 72304
rect 6019 72260 6077 72261
rect 6211 72260 6269 72261
rect 3244 72220 6028 72260
rect 6068 72220 6220 72260
rect 6260 72220 6269 72260
rect 1411 72136 1420 72176
rect 1460 72136 1900 72176
rect 1940 72136 2092 72176
rect 2132 72136 2141 72176
rect 3244 72092 3284 72220
rect 6019 72219 6077 72220
rect 6211 72219 6269 72220
rect 5635 72136 5644 72176
rect 5684 72136 6412 72176
rect 6452 72136 6461 72176
rect 1507 72052 1516 72092
rect 1556 72052 2284 72092
rect 2324 72052 2476 72092
rect 2516 72052 2525 72092
rect 2947 72052 2956 72092
rect 2996 72052 3244 72092
rect 3284 72052 3293 72092
rect 5443 72052 5452 72092
rect 5492 72052 6316 72092
rect 6356 72052 6365 72092
rect 0 72008 80 72028
rect 3043 72008 3101 72009
rect 5635 72008 5693 72009
rect 6211 72008 6269 72009
rect 0 71968 2324 72008
rect 0 71948 80 71968
rect 2284 71840 2324 71968
rect 3043 71968 3052 72008
rect 3092 71968 3724 72008
rect 3764 71968 3773 72008
rect 4579 71968 4588 72008
rect 4628 71968 5644 72008
rect 5684 71968 5693 72008
rect 6126 71968 6220 72008
rect 6260 71968 6269 72008
rect 3043 71967 3101 71968
rect 5635 71967 5693 71968
rect 6211 71967 6269 71968
rect 6595 72008 6653 72009
rect 6595 71968 6604 72008
rect 6644 71968 6796 72008
rect 6836 71968 6845 72008
rect 6595 71967 6653 71968
rect 2467 71924 2525 71925
rect 6892 71924 6932 72304
rect 8803 72303 8861 72304
rect 9196 72260 9236 72304
rect 9196 72220 9484 72260
rect 9524 72220 9533 72260
rect 10819 72220 10828 72260
rect 10868 72220 15916 72260
rect 15956 72220 15965 72260
rect 12451 72176 12509 72177
rect 8803 72136 8812 72176
rect 8852 72136 9772 72176
rect 9812 72136 9821 72176
rect 10339 72136 10348 72176
rect 10388 72136 10397 72176
rect 12366 72136 12460 72176
rect 12500 72136 12509 72176
rect 9091 72092 9149 72093
rect 10348 72092 10388 72136
rect 12451 72135 12509 72136
rect 15235 72092 15293 72093
rect 6979 72052 6988 72092
rect 7028 72052 9100 72092
rect 9140 72052 9149 72092
rect 9283 72052 9292 72092
rect 9332 72052 10388 72092
rect 11971 72052 11980 72092
rect 12020 72052 15244 72092
rect 15284 72052 15293 72092
rect 9091 72051 9149 72052
rect 15235 72051 15293 72052
rect 13795 72008 13853 72009
rect 8035 71968 8044 72008
rect 8084 71968 8428 72008
rect 8468 71968 8620 72008
rect 8660 71968 9196 72008
rect 9236 71968 9245 72008
rect 9667 71968 9676 72008
rect 9716 71968 10348 72008
rect 10388 71968 10397 72008
rect 13123 71968 13132 72008
rect 13172 71968 13612 72008
rect 13652 71968 13661 72008
rect 13795 71968 13804 72008
rect 13844 71968 21332 72008
rect 13795 71967 13853 71968
rect 2382 71884 2476 71924
rect 2516 71884 3916 71924
rect 3956 71884 3965 71924
rect 4771 71884 4780 71924
rect 4820 71884 6836 71924
rect 6892 71884 16204 71924
rect 16244 71884 18316 71924
rect 18356 71884 18365 71924
rect 2467 71883 2525 71884
rect 6595 71840 6653 71841
rect 2284 71800 3628 71840
rect 3668 71800 3677 71840
rect 4919 71800 4928 71840
rect 4968 71800 5010 71840
rect 5050 71800 5092 71840
rect 5132 71800 5174 71840
rect 5214 71800 5256 71840
rect 5296 71800 5305 71840
rect 6403 71800 6412 71840
rect 6452 71800 6604 71840
rect 6644 71800 6653 71840
rect 6796 71840 6836 71884
rect 11587 71840 11645 71841
rect 12355 71840 12413 71841
rect 21292 71840 21332 71968
rect 21424 71840 21504 71860
rect 6796 71800 8140 71840
rect 8180 71800 8524 71840
rect 8564 71800 8573 71840
rect 9187 71800 9196 71840
rect 9236 71800 9580 71840
rect 9620 71800 9629 71840
rect 11587 71800 11596 71840
rect 11636 71800 12364 71840
rect 12404 71800 12413 71840
rect 15139 71800 15148 71840
rect 15188 71800 17164 71840
rect 17204 71800 17213 71840
rect 20039 71800 20048 71840
rect 20088 71800 20130 71840
rect 20170 71800 20212 71840
rect 20252 71800 20294 71840
rect 20334 71800 20376 71840
rect 20416 71800 20425 71840
rect 21292 71800 21504 71840
rect 6595 71799 6653 71800
rect 11587 71799 11645 71800
rect 12355 71799 12413 71800
rect 21424 71780 21504 71800
rect 3331 71756 3389 71757
rect 3331 71716 3340 71756
rect 3380 71716 7756 71756
rect 7796 71716 9772 71756
rect 9812 71716 9821 71756
rect 10435 71716 10444 71756
rect 10484 71716 11308 71756
rect 11348 71716 15764 71756
rect 15811 71716 15820 71756
rect 15860 71716 16204 71756
rect 16244 71716 16253 71756
rect 3331 71715 3389 71716
rect 0 71672 80 71692
rect 15724 71672 15764 71716
rect 0 71632 12460 71672
rect 12500 71632 12509 71672
rect 15724 71632 16588 71672
rect 16628 71632 18604 71672
rect 18644 71632 18796 71672
rect 18836 71632 18845 71672
rect 0 71612 80 71632
rect 4675 71548 4684 71588
rect 4724 71548 5932 71588
rect 5972 71548 6836 71588
rect 7075 71548 7084 71588
rect 7124 71548 10828 71588
rect 10868 71548 10877 71588
rect 11320 71548 12596 71588
rect 16099 71548 16108 71588
rect 16148 71548 16396 71588
rect 16436 71548 16445 71588
rect 1891 71504 1949 71505
rect 1891 71464 1900 71504
rect 1940 71464 2860 71504
rect 2900 71464 3532 71504
rect 3572 71464 3581 71504
rect 3907 71464 3916 71504
rect 3956 71464 4108 71504
rect 4148 71464 4157 71504
rect 5059 71464 5068 71504
rect 5108 71464 5447 71504
rect 5487 71464 5496 71504
rect 5539 71464 5548 71504
rect 5588 71464 6700 71504
rect 6740 71464 6749 71504
rect 1891 71463 1949 71464
rect 3523 71420 3581 71421
rect 6796 71420 6836 71548
rect 11320 71504 11360 71548
rect 12163 71504 12221 71505
rect 12556 71504 12596 71548
rect 19363 71504 19421 71505
rect 7939 71464 7948 71504
rect 7988 71464 9004 71504
rect 9044 71464 9580 71504
rect 9620 71464 9629 71504
rect 9763 71464 9772 71504
rect 9812 71464 11360 71504
rect 12078 71464 12172 71504
rect 12212 71464 12221 71504
rect 12547 71464 12556 71504
rect 12596 71464 13804 71504
rect 13844 71464 13853 71504
rect 19278 71464 19372 71504
rect 19412 71464 19421 71504
rect 12163 71463 12221 71464
rect 19363 71463 19421 71464
rect 12172 71420 12212 71463
rect 2179 71380 2188 71420
rect 2228 71380 2668 71420
rect 2708 71380 2717 71420
rect 3523 71380 3532 71420
rect 3572 71380 5260 71420
rect 5300 71380 5309 71420
rect 5731 71380 5740 71420
rect 5780 71380 6028 71420
rect 6068 71380 6508 71420
rect 6548 71380 6557 71420
rect 6796 71380 10636 71420
rect 10676 71380 10685 71420
rect 12172 71380 13996 71420
rect 14036 71380 17548 71420
rect 17588 71380 17597 71420
rect 3523 71379 3581 71380
rect 0 71336 80 71356
rect 0 71296 6220 71336
rect 6260 71296 6269 71336
rect 6595 71296 6604 71336
rect 6644 71296 6988 71336
rect 7028 71296 7037 71336
rect 7363 71296 7372 71336
rect 7412 71296 7660 71336
rect 7700 71296 7709 71336
rect 0 71276 80 71296
rect 2083 71252 2141 71253
rect 15811 71252 15869 71253
rect 2083 71212 2092 71252
rect 2132 71212 2668 71252
rect 2708 71212 2717 71252
rect 3043 71212 3052 71252
rect 3092 71212 3628 71252
rect 3668 71212 15820 71252
rect 15860 71212 15869 71252
rect 2083 71211 2141 71212
rect 15811 71211 15869 71212
rect 9859 71168 9917 71169
rect 21424 71168 21504 71188
rect 2851 71128 2860 71168
rect 2900 71128 5876 71168
rect 6883 71128 6892 71168
rect 6932 71128 7180 71168
rect 7220 71128 7229 71168
rect 9859 71128 9868 71168
rect 9908 71128 21504 71168
rect 5836 71084 5876 71128
rect 9859 71127 9917 71128
rect 21424 71108 21504 71128
rect 3679 71044 3688 71084
rect 3728 71044 3770 71084
rect 3810 71044 3852 71084
rect 3892 71044 3934 71084
rect 3974 71044 4016 71084
rect 4056 71044 4065 71084
rect 5836 71044 12652 71084
rect 12692 71044 13804 71084
rect 13844 71044 13853 71084
rect 15811 71044 15820 71084
rect 15860 71044 16204 71084
rect 16244 71044 16253 71084
rect 18799 71044 18808 71084
rect 18848 71044 18890 71084
rect 18930 71044 18972 71084
rect 19012 71044 19054 71084
rect 19094 71044 19136 71084
rect 19176 71044 19185 71084
rect 0 71000 80 71020
rect 16003 71000 16061 71001
rect 0 70960 9100 71000
rect 9140 70960 9149 71000
rect 15918 70960 16012 71000
rect 16052 70960 16061 71000
rect 0 70940 80 70960
rect 16003 70959 16061 70960
rect 2500 70876 18124 70916
rect 18164 70876 18173 70916
rect 2500 70832 2540 70876
rect 1324 70792 2540 70832
rect 3139 70832 3197 70833
rect 10531 70832 10589 70833
rect 15619 70832 15677 70833
rect 3139 70792 3148 70832
rect 3188 70792 3724 70832
rect 3764 70792 3773 70832
rect 5251 70792 5260 70832
rect 5300 70792 5740 70832
rect 5780 70792 5789 70832
rect 6691 70792 6700 70832
rect 6740 70792 7084 70832
rect 7124 70792 7133 70832
rect 7267 70792 7276 70832
rect 7316 70792 7468 70832
rect 7508 70792 7517 70832
rect 10446 70792 10540 70832
rect 10580 70792 10589 70832
rect 15043 70792 15052 70832
rect 15092 70792 15101 70832
rect 15619 70792 15628 70832
rect 15668 70792 19372 70832
rect 19412 70792 19421 70832
rect 0 70664 80 70684
rect 1324 70664 1364 70792
rect 3139 70791 3197 70792
rect 10531 70791 10589 70792
rect 1411 70748 1469 70749
rect 4099 70748 4157 70749
rect 1411 70708 1420 70748
rect 1460 70708 2956 70748
rect 2996 70708 3005 70748
rect 4003 70708 4012 70748
rect 4052 70708 4108 70748
rect 4148 70708 4157 70748
rect 1411 70707 1469 70708
rect 4099 70707 4157 70708
rect 6979 70748 7037 70749
rect 15052 70748 15092 70792
rect 15619 70791 15677 70792
rect 6979 70708 6988 70748
rect 7028 70708 7180 70748
rect 7220 70708 7229 70748
rect 15052 70708 15956 70748
rect 6979 70707 7037 70708
rect 0 70624 1364 70664
rect 2179 70664 2237 70665
rect 4771 70664 4829 70665
rect 8131 70664 8189 70665
rect 9283 70664 9341 70665
rect 15916 70664 15956 70708
rect 2179 70624 2188 70664
rect 2228 70624 2572 70664
rect 2612 70624 2621 70664
rect 2851 70624 2860 70664
rect 2900 70624 3532 70664
rect 3572 70624 3581 70664
rect 4771 70624 4780 70664
rect 4820 70624 5164 70664
rect 5204 70624 5356 70664
rect 5396 70624 5405 70664
rect 7075 70624 7084 70664
rect 7124 70624 7660 70664
rect 7700 70624 7709 70664
rect 8131 70624 8140 70664
rect 8180 70624 8620 70664
rect 8660 70624 8669 70664
rect 8995 70624 9004 70664
rect 9044 70624 9292 70664
rect 9332 70624 9341 70664
rect 10819 70624 10828 70664
rect 10868 70624 13036 70664
rect 13076 70624 13085 70664
rect 14467 70624 14476 70664
rect 14516 70624 14860 70664
rect 14900 70624 14909 70664
rect 15043 70624 15052 70664
rect 15092 70624 15532 70664
rect 15572 70624 15581 70664
rect 15907 70624 15916 70664
rect 15956 70624 15965 70664
rect 18595 70624 18604 70664
rect 18644 70624 18892 70664
rect 18932 70624 18941 70664
rect 19459 70624 19468 70664
rect 19508 70624 19517 70664
rect 0 70604 80 70624
rect 2179 70623 2237 70624
rect 4771 70623 4829 70624
rect 8131 70623 8189 70624
rect 9283 70623 9341 70624
rect 14860 70580 14900 70624
rect 19468 70580 19508 70624
rect 1219 70540 1228 70580
rect 1268 70540 2380 70580
rect 2420 70540 2429 70580
rect 6019 70540 6028 70580
rect 6068 70540 6077 70580
rect 6787 70540 6796 70580
rect 6836 70540 7468 70580
rect 7508 70540 7517 70580
rect 14860 70540 15244 70580
rect 15284 70540 15293 70580
rect 19468 70540 20044 70580
rect 20084 70540 20093 70580
rect 6028 70496 6068 70540
rect 7747 70496 7805 70497
rect 21424 70496 21504 70516
rect 6028 70456 7756 70496
rect 7796 70456 7805 70496
rect 11587 70456 11596 70496
rect 11636 70456 12172 70496
rect 12212 70456 12221 70496
rect 14476 70456 17644 70496
rect 17684 70456 17693 70496
rect 18787 70456 18796 70496
rect 18836 70456 19756 70496
rect 19796 70456 19805 70496
rect 20140 70456 21504 70496
rect 7747 70455 7805 70456
rect 9955 70412 10013 70413
rect 9859 70372 9868 70412
rect 9908 70372 9964 70412
rect 10004 70372 10013 70412
rect 9955 70371 10013 70372
rect 0 70328 80 70348
rect 0 70288 2540 70328
rect 4919 70288 4928 70328
rect 4968 70288 5010 70328
rect 5050 70288 5092 70328
rect 5132 70288 5174 70328
rect 5214 70288 5256 70328
rect 5296 70288 5305 70328
rect 0 70268 80 70288
rect 2500 70244 2540 70288
rect 2500 70204 14380 70244
rect 14420 70204 14429 70244
rect 14476 70160 14516 70456
rect 15811 70412 15869 70413
rect 20140 70412 20180 70456
rect 21424 70436 21504 70456
rect 15811 70372 15820 70412
rect 15860 70372 15916 70412
rect 15956 70372 15965 70412
rect 16300 70372 20180 70412
rect 15811 70371 15869 70372
rect 15619 70328 15677 70329
rect 15619 70288 15628 70328
rect 15668 70288 15724 70328
rect 15764 70288 15773 70328
rect 15619 70287 15677 70288
rect 14947 70244 15005 70245
rect 16300 70244 16340 70372
rect 20039 70288 20048 70328
rect 20088 70288 20130 70328
rect 20170 70288 20212 70328
rect 20252 70288 20294 70328
rect 20334 70288 20376 70328
rect 20416 70288 20425 70328
rect 14947 70204 14956 70244
rect 14996 70204 16340 70244
rect 14947 70203 15005 70204
rect 19651 70160 19709 70161
rect 5923 70120 5932 70160
rect 5972 70120 7660 70160
rect 7700 70120 7709 70160
rect 7843 70120 7852 70160
rect 7892 70120 8236 70160
rect 8276 70120 11884 70160
rect 11924 70120 14516 70160
rect 15331 70120 15340 70160
rect 15380 70120 16396 70160
rect 16436 70120 16445 70160
rect 18691 70120 18700 70160
rect 18740 70120 19660 70160
rect 19700 70120 19709 70160
rect 19651 70119 19709 70120
rect 2851 70076 2909 70077
rect 2766 70036 2860 70076
rect 2900 70036 2909 70076
rect 4675 70036 4684 70076
rect 4724 70036 5644 70076
rect 5684 70036 6892 70076
rect 6932 70036 6941 70076
rect 16291 70036 16300 70076
rect 16340 70036 17164 70076
rect 17204 70036 18028 70076
rect 18068 70036 18988 70076
rect 19028 70036 19037 70076
rect 19363 70036 19372 70076
rect 19412 70036 20044 70076
rect 20084 70036 20093 70076
rect 2851 70035 2909 70036
rect 0 69992 80 70012
rect 1315 69992 1373 69993
rect 4291 69992 4349 69993
rect 11683 69992 11741 69993
rect 12547 69992 12605 69993
rect 0 69952 1172 69992
rect 1230 69952 1324 69992
rect 1364 69952 1373 69992
rect 2467 69952 2476 69992
rect 2516 69952 2668 69992
rect 2708 69952 3052 69992
rect 3092 69952 4108 69992
rect 4148 69952 4157 69992
rect 4291 69952 4300 69992
rect 4340 69952 4434 69992
rect 4579 69952 4588 69992
rect 4628 69952 6316 69992
rect 6356 69952 6365 69992
rect 6499 69952 6508 69992
rect 6548 69952 6796 69992
rect 6836 69952 6845 69992
rect 9475 69952 9484 69992
rect 9524 69952 11116 69992
rect 11156 69952 11165 69992
rect 11598 69952 11692 69992
rect 11732 69952 12556 69992
rect 12596 69952 12605 69992
rect 16003 69952 16012 69992
rect 16052 69952 16588 69992
rect 16628 69952 17068 69992
rect 17108 69952 17117 69992
rect 17620 69952 18700 69992
rect 18740 69952 18749 69992
rect 19075 69952 19084 69992
rect 19124 69952 20236 69992
rect 20276 69952 20285 69992
rect 0 69932 80 69952
rect 1132 69908 1172 69952
rect 1315 69951 1373 69952
rect 4291 69951 4349 69952
rect 11683 69951 11741 69952
rect 12547 69951 12605 69952
rect 1132 69868 4244 69908
rect 2659 69740 2717 69741
rect 3139 69740 3197 69741
rect 2574 69700 2668 69740
rect 2708 69700 2717 69740
rect 2851 69700 2860 69740
rect 2900 69700 3148 69740
rect 3188 69700 3197 69740
rect 2659 69699 2717 69700
rect 3139 69699 3197 69700
rect 3427 69740 3485 69741
rect 4204 69740 4244 69868
rect 4300 69824 4340 69951
rect 5731 69908 5789 69909
rect 11875 69908 11933 69909
rect 17620 69908 17660 69952
rect 5731 69868 5740 69908
rect 5780 69868 6124 69908
rect 6164 69868 6173 69908
rect 6883 69868 6892 69908
rect 6932 69868 7276 69908
rect 7316 69868 7325 69908
rect 9859 69868 9868 69908
rect 9908 69868 10636 69908
rect 10676 69868 10685 69908
rect 11875 69868 11884 69908
rect 11924 69868 12172 69908
rect 12212 69868 12221 69908
rect 15523 69868 15532 69908
rect 15572 69868 17660 69908
rect 17923 69868 17932 69908
rect 17972 69868 20180 69908
rect 5731 69867 5789 69868
rect 11875 69867 11933 69868
rect 11491 69824 11549 69825
rect 20140 69824 20180 69868
rect 21424 69824 21504 69844
rect 4300 69784 8236 69824
rect 8276 69784 8285 69824
rect 11491 69784 11500 69824
rect 11540 69784 12076 69824
rect 12116 69784 12125 69824
rect 15043 69784 15052 69824
rect 15092 69784 18220 69824
rect 18260 69784 18269 69824
rect 18979 69784 18988 69824
rect 19028 69784 19700 69824
rect 20140 69784 21504 69824
rect 11491 69783 11549 69784
rect 3427 69700 3436 69740
rect 3476 69700 3724 69740
rect 3764 69700 3773 69740
rect 4204 69700 8044 69740
rect 8084 69700 8093 69740
rect 11107 69700 11116 69740
rect 11156 69700 11980 69740
rect 12020 69700 13132 69740
rect 13172 69700 13516 69740
rect 13556 69700 13565 69740
rect 14563 69700 14572 69740
rect 14612 69700 16108 69740
rect 16148 69700 17548 69740
rect 17588 69700 17740 69740
rect 17780 69700 17789 69740
rect 19075 69700 19084 69740
rect 19124 69700 19133 69740
rect 3427 69699 3485 69700
rect 0 69656 80 69676
rect 16003 69656 16061 69657
rect 19084 69656 19124 69700
rect 19660 69656 19700 69784
rect 21424 69764 21504 69784
rect 0 69616 5548 69656
rect 5588 69616 5597 69656
rect 6307 69616 6316 69656
rect 6356 69616 6604 69656
rect 6644 69616 6653 69656
rect 16003 69616 16012 69656
rect 16052 69616 16300 69656
rect 16340 69616 16349 69656
rect 19084 69616 19276 69656
rect 19316 69616 19325 69656
rect 19651 69616 19660 69656
rect 19700 69616 19709 69656
rect 0 69596 80 69616
rect 16003 69615 16061 69616
rect 4771 69572 4829 69573
rect 10147 69572 10205 69573
rect 3679 69532 3688 69572
rect 3728 69532 3770 69572
rect 3810 69532 3852 69572
rect 3892 69532 3934 69572
rect 3974 69532 4016 69572
rect 4056 69532 4065 69572
rect 4771 69532 4780 69572
rect 4820 69532 8524 69572
rect 8564 69532 8573 69572
rect 10147 69532 10156 69572
rect 10196 69532 16684 69572
rect 16724 69532 16733 69572
rect 18799 69532 18808 69572
rect 18848 69532 18890 69572
rect 18930 69532 18972 69572
rect 19012 69532 19054 69572
rect 19094 69532 19136 69572
rect 19176 69532 19185 69572
rect 4771 69531 4829 69532
rect 10147 69531 10205 69532
rect 16012 69489 16052 69532
rect 16003 69488 16061 69489
rect 16771 69488 16829 69489
rect 2500 69448 15244 69488
rect 15284 69448 15293 69488
rect 16003 69448 16012 69488
rect 16052 69448 16092 69488
rect 16771 69448 16780 69488
rect 16820 69448 19852 69488
rect 19892 69448 19901 69488
rect 0 69320 80 69340
rect 2500 69320 2540 69448
rect 16003 69447 16061 69448
rect 16771 69447 16829 69448
rect 3235 69404 3293 69405
rect 3235 69364 3244 69404
rect 3284 69364 3628 69404
rect 3668 69364 3677 69404
rect 5923 69364 5932 69404
rect 5972 69364 8852 69404
rect 15139 69364 15148 69404
rect 15188 69364 16012 69404
rect 16052 69364 16061 69404
rect 17635 69364 17644 69404
rect 17684 69364 17836 69404
rect 17876 69364 18700 69404
rect 18740 69364 18749 69404
rect 18883 69364 18892 69404
rect 18932 69364 19276 69404
rect 19316 69364 19325 69404
rect 3235 69363 3293 69364
rect 8812 69321 8852 69364
rect 8803 69320 8861 69321
rect 9187 69320 9245 69321
rect 0 69280 2540 69320
rect 4675 69280 4684 69320
rect 4724 69280 5452 69320
rect 5492 69280 6220 69320
rect 6260 69280 6269 69320
rect 6691 69280 6700 69320
rect 6740 69280 7372 69320
rect 7412 69280 7421 69320
rect 8803 69280 8812 69320
rect 8852 69280 9196 69320
rect 9236 69280 9245 69320
rect 0 69260 80 69280
rect 8803 69279 8861 69280
rect 9187 69279 9245 69280
rect 9667 69320 9725 69321
rect 10339 69320 10397 69321
rect 13603 69320 13661 69321
rect 9667 69280 9676 69320
rect 9716 69280 10348 69320
rect 10388 69280 10444 69320
rect 10484 69280 10493 69320
rect 10723 69280 10732 69320
rect 10772 69280 11788 69320
rect 11828 69280 11837 69320
rect 13603 69280 13612 69320
rect 13652 69280 13708 69320
rect 13748 69280 13757 69320
rect 14755 69280 14764 69320
rect 14804 69280 15340 69320
rect 15380 69280 15389 69320
rect 18403 69280 18412 69320
rect 18452 69280 19948 69320
rect 19988 69280 19997 69320
rect 9667 69279 9725 69280
rect 10339 69279 10397 69280
rect 13603 69279 13661 69280
rect 2755 69236 2813 69237
rect 19363 69236 19421 69237
rect 1123 69196 1132 69236
rect 1172 69196 2476 69236
rect 2516 69196 2525 69236
rect 2755 69196 2764 69236
rect 2804 69196 6892 69236
rect 6932 69196 7756 69236
rect 7796 69196 7805 69236
rect 9475 69196 9484 69236
rect 9524 69196 15052 69236
rect 15092 69196 15101 69236
rect 17635 69196 17644 69236
rect 17684 69196 18604 69236
rect 18644 69196 18653 69236
rect 18979 69196 18988 69236
rect 19028 69196 19372 69236
rect 19412 69196 19421 69236
rect 2755 69195 2813 69196
rect 19363 69195 19421 69196
rect 9763 69152 9821 69153
rect 11011 69152 11069 69153
rect 21424 69152 21504 69172
rect 6403 69112 6412 69152
rect 6452 69112 7084 69152
rect 7124 69112 7133 69152
rect 9763 69112 9772 69152
rect 9812 69112 10060 69152
rect 10100 69112 10109 69152
rect 10531 69112 10540 69152
rect 10580 69112 11020 69152
rect 11060 69112 11069 69152
rect 11299 69112 11308 69152
rect 11348 69112 11500 69152
rect 11540 69112 11549 69152
rect 14275 69112 14284 69152
rect 14324 69112 14764 69152
rect 14804 69112 14956 69152
rect 14996 69112 15005 69152
rect 19363 69112 19372 69152
rect 19412 69112 19756 69152
rect 19796 69112 19805 69152
rect 20140 69112 21504 69152
rect 9763 69111 9821 69112
rect 11011 69111 11069 69112
rect 5251 69028 5260 69068
rect 5300 69028 5452 69068
rect 5492 69028 5501 69068
rect 13315 69028 13324 69068
rect 13364 69028 19180 69068
rect 19220 69028 19229 69068
rect 0 68984 80 69004
rect 2755 68984 2813 68985
rect 7267 68984 7325 68985
rect 0 68944 2764 68984
rect 2804 68944 2813 68984
rect 2947 68944 2956 68984
rect 2996 68944 3436 68984
rect 3476 68944 7028 68984
rect 7182 68944 7276 68984
rect 7316 68944 7325 68984
rect 9667 68944 9676 68984
rect 9716 68944 10156 68984
rect 10196 68944 10205 68984
rect 13027 68944 13036 68984
rect 13076 68944 15628 68984
rect 15668 68944 15677 68984
rect 18307 68944 18316 68984
rect 18356 68944 19276 68984
rect 19316 68944 19325 68984
rect 0 68924 80 68944
rect 2755 68943 2813 68944
rect 6988 68900 7028 68944
rect 7267 68943 7325 68944
rect 20140 68900 20180 69112
rect 21424 69092 21504 69112
rect 2563 68860 2572 68900
rect 2612 68860 6892 68900
rect 6932 68860 6941 68900
rect 6988 68860 11692 68900
rect 11732 68860 12844 68900
rect 12884 68860 12893 68900
rect 18796 68860 20180 68900
rect 18796 68816 18836 68860
rect 4919 68776 4928 68816
rect 4968 68776 5010 68816
rect 5050 68776 5092 68816
rect 5132 68776 5174 68816
rect 5214 68776 5256 68816
rect 5296 68776 5305 68816
rect 5731 68776 5740 68816
rect 5780 68776 13708 68816
rect 13748 68776 13757 68816
rect 18787 68776 18796 68816
rect 18836 68776 18845 68816
rect 20039 68776 20048 68816
rect 20088 68776 20130 68816
rect 20170 68776 20212 68816
rect 20252 68776 20294 68816
rect 20334 68776 20376 68816
rect 20416 68776 20425 68816
rect 3811 68692 3820 68732
rect 3860 68692 6124 68732
rect 6164 68692 6173 68732
rect 8131 68692 8140 68732
rect 8180 68692 11788 68732
rect 11828 68692 11980 68732
rect 12020 68692 12029 68732
rect 0 68648 80 68668
rect 5539 68648 5597 68649
rect 0 68608 5164 68648
rect 5204 68608 5213 68648
rect 5539 68608 5548 68648
rect 5588 68608 5740 68648
rect 5780 68608 5789 68648
rect 10339 68608 10348 68648
rect 10388 68608 10397 68648
rect 10723 68608 10732 68648
rect 10772 68608 16396 68648
rect 16436 68608 16445 68648
rect 0 68588 80 68608
rect 5539 68607 5597 68608
rect 3427 68564 3485 68565
rect 3619 68564 3677 68565
rect 4867 68564 4925 68565
rect 10348 68564 10388 68608
rect 3139 68524 3148 68564
rect 3188 68524 3436 68564
rect 3476 68524 3628 68564
rect 3668 68524 3677 68564
rect 4099 68524 4108 68564
rect 4148 68524 4684 68564
rect 4724 68524 4733 68564
rect 4867 68524 4876 68564
rect 4916 68524 8140 68564
rect 8180 68524 9484 68564
rect 9524 68524 9533 68564
rect 10348 68524 11308 68564
rect 11348 68524 11357 68564
rect 3427 68523 3485 68524
rect 3619 68523 3677 68524
rect 4867 68523 4925 68524
rect 21424 68480 21504 68500
rect 1027 68440 1036 68480
rect 1076 68440 2380 68480
rect 2420 68440 2429 68480
rect 2500 68440 3820 68480
rect 3860 68440 3869 68480
rect 4195 68440 4204 68480
rect 4244 68440 4253 68480
rect 4483 68440 4492 68480
rect 4532 68440 6220 68480
rect 6260 68440 6269 68480
rect 6883 68440 6892 68480
rect 6932 68440 12076 68480
rect 12116 68440 12125 68480
rect 14947 68440 14956 68480
rect 14996 68440 15820 68480
rect 15860 68440 16300 68480
rect 16340 68440 16349 68480
rect 18691 68440 18700 68480
rect 18740 68440 19276 68480
rect 19316 68440 19325 68480
rect 20620 68440 21504 68480
rect 2380 68396 2420 68440
rect 2500 68396 2540 68440
rect 2380 68356 2540 68396
rect 4204 68396 4244 68440
rect 17155 68396 17213 68397
rect 20620 68396 20660 68440
rect 21424 68420 21504 68440
rect 4204 68356 5108 68396
rect 9667 68356 9676 68396
rect 9716 68356 10636 68396
rect 10676 68356 13036 68396
rect 13076 68356 13085 68396
rect 17155 68356 17164 68396
rect 17204 68356 20660 68396
rect 0 68312 80 68332
rect 4771 68312 4829 68313
rect 0 68272 4780 68312
rect 4820 68272 4829 68312
rect 0 68252 80 68272
rect 4771 68271 4829 68272
rect 4099 68228 4157 68229
rect 2179 68188 2188 68228
rect 2228 68188 2380 68228
rect 2420 68188 2429 68228
rect 3811 68188 3820 68228
rect 3860 68188 4108 68228
rect 4148 68188 4157 68228
rect 5068 68228 5108 68356
rect 17155 68355 17213 68356
rect 7075 68312 7133 68313
rect 8611 68312 8669 68313
rect 7075 68272 7084 68312
rect 7124 68272 7852 68312
rect 7892 68272 8620 68312
rect 8660 68272 15340 68312
rect 15380 68272 15389 68312
rect 7075 68271 7133 68272
rect 8611 68271 8669 68272
rect 5068 68188 6700 68228
rect 6740 68188 6749 68228
rect 11320 68188 13708 68228
rect 13748 68188 13757 68228
rect 17539 68188 17548 68228
rect 17588 68188 18412 68228
rect 18452 68188 18892 68228
rect 18932 68188 18941 68228
rect 4099 68187 4157 68188
rect 1699 68144 1757 68145
rect 11320 68144 11360 68188
rect 18892 68144 18932 68188
rect 1699 68104 1708 68144
rect 1748 68104 11360 68144
rect 12067 68104 12076 68144
rect 12116 68104 15628 68144
rect 15668 68104 15677 68144
rect 18019 68104 18028 68144
rect 18068 68104 18604 68144
rect 18644 68104 18653 68144
rect 18892 68104 19564 68144
rect 19604 68104 19613 68144
rect 1699 68103 1757 68104
rect 7939 68060 7997 68061
rect 3679 68020 3688 68060
rect 3728 68020 3770 68060
rect 3810 68020 3852 68060
rect 3892 68020 3934 68060
rect 3974 68020 4016 68060
rect 4056 68020 4065 68060
rect 4195 68020 4204 68060
rect 4244 68020 4492 68060
rect 4532 68020 4541 68060
rect 5539 68020 5548 68060
rect 5588 68020 7084 68060
rect 7124 68020 7133 68060
rect 7939 68020 7948 68060
rect 7988 68020 8716 68060
rect 8756 68020 9676 68060
rect 9716 68020 9725 68060
rect 12739 68020 12748 68060
rect 12788 68020 13324 68060
rect 13364 68020 13373 68060
rect 13795 68020 13804 68060
rect 13844 68020 15052 68060
rect 15092 68020 15101 68060
rect 18211 68020 18220 68060
rect 18260 68020 18740 68060
rect 18799 68020 18808 68060
rect 18848 68020 18890 68060
rect 18930 68020 18972 68060
rect 19012 68020 19054 68060
rect 19094 68020 19136 68060
rect 19176 68020 19185 68060
rect 7939 68019 7997 68020
rect 0 67976 80 67996
rect 18700 67976 18740 68020
rect 0 67936 18028 67976
rect 18068 67936 18077 67976
rect 18700 67936 19028 67976
rect 0 67916 80 67936
rect 15139 67892 15197 67893
rect 18988 67892 19028 67936
rect 4579 67852 4588 67892
rect 4628 67852 4876 67892
rect 4916 67852 4925 67892
rect 5251 67852 5260 67892
rect 5300 67852 6700 67892
rect 6740 67852 6749 67892
rect 9091 67852 9100 67892
rect 9140 67852 9772 67892
rect 9812 67852 9821 67892
rect 10051 67852 10060 67892
rect 10100 67852 15148 67892
rect 15188 67852 15197 67892
rect 18979 67852 18988 67892
rect 19028 67852 19037 67892
rect 15139 67851 15197 67852
rect 20131 67808 20189 67809
rect 21424 67808 21504 67828
rect 1795 67768 1804 67808
rect 1844 67768 2476 67808
rect 2516 67768 2860 67808
rect 2900 67768 2909 67808
rect 5452 67768 5932 67808
rect 5972 67768 5981 67808
rect 9100 67768 11788 67808
rect 11828 67768 11837 67808
rect 15148 67768 16300 67808
rect 16340 67768 17068 67808
rect 17108 67768 17117 67808
rect 20131 67768 20140 67808
rect 20180 67768 21504 67808
rect 1603 67724 1661 67725
rect 5452 67724 5492 67768
rect 9100 67724 9140 67768
rect 10147 67724 10205 67725
rect 15148 67724 15188 67768
rect 20131 67767 20189 67768
rect 21424 67748 21504 67768
rect 1603 67684 1612 67724
rect 1652 67684 5492 67724
rect 5548 67684 9100 67724
rect 9140 67684 9149 67724
rect 10062 67684 10156 67724
rect 10196 67684 10205 67724
rect 14851 67684 14860 67724
rect 14900 67684 15148 67724
rect 15188 67684 15197 67724
rect 15427 67684 15436 67724
rect 15476 67684 15724 67724
rect 15764 67684 15773 67724
rect 15820 67684 16876 67724
rect 16916 67684 16925 67724
rect 1603 67683 1661 67684
rect 0 67640 80 67660
rect 5548 67640 5588 67684
rect 10147 67683 10205 67684
rect 13219 67640 13277 67641
rect 15820 67640 15860 67684
rect 0 67600 1132 67640
rect 1172 67600 1181 67640
rect 1987 67600 1996 67640
rect 2036 67600 2476 67640
rect 2516 67600 2525 67640
rect 2572 67600 3628 67640
rect 3668 67600 3677 67640
rect 4483 67600 4492 67640
rect 4532 67600 5588 67640
rect 5731 67600 5740 67640
rect 5780 67600 13228 67640
rect 13268 67600 15860 67640
rect 16099 67600 16108 67640
rect 16148 67600 16972 67640
rect 17012 67600 17021 67640
rect 17731 67600 17740 67640
rect 17780 67600 19468 67640
rect 19508 67600 19517 67640
rect 19651 67600 19660 67640
rect 19700 67600 19852 67640
rect 19892 67600 19901 67640
rect 0 67580 80 67600
rect 2572 67556 2612 67600
rect 13219 67599 13277 67600
rect 15331 67556 15389 67557
rect 2563 67516 2572 67556
rect 2612 67516 2621 67556
rect 2851 67516 2860 67556
rect 2900 67516 3244 67556
rect 3284 67516 3293 67556
rect 3436 67516 3532 67556
rect 3572 67516 6028 67556
rect 6068 67516 6077 67556
rect 6787 67516 6796 67556
rect 6836 67516 7372 67556
rect 7412 67516 7421 67556
rect 9763 67516 9772 67556
rect 9812 67516 10060 67556
rect 10100 67516 10109 67556
rect 15331 67516 15340 67556
rect 15380 67516 15532 67556
rect 15572 67516 15916 67556
rect 15956 67516 15965 67556
rect 16195 67516 16204 67556
rect 16244 67516 17644 67556
rect 17684 67516 17693 67556
rect 19267 67516 19276 67556
rect 19316 67516 20236 67556
rect 20276 67516 20285 67556
rect 3436 67472 3476 67516
rect 15331 67515 15389 67516
rect 3811 67472 3869 67473
rect 11395 67472 11453 67473
rect 3427 67432 3436 67472
rect 3476 67432 3485 67472
rect 3811 67432 3820 67472
rect 3860 67432 4108 67472
rect 4148 67432 4157 67472
rect 8899 67432 8908 67472
rect 8948 67432 9676 67472
rect 9716 67432 9725 67472
rect 11280 67432 11308 67472
rect 11348 67432 11404 67472
rect 11444 67432 11455 67472
rect 15427 67432 15436 67472
rect 15476 67432 15628 67472
rect 15668 67432 15677 67472
rect 16483 67432 16492 67472
rect 16532 67432 16876 67472
rect 16916 67432 16925 67472
rect 19756 67432 20044 67472
rect 20084 67432 20093 67472
rect 3811 67431 3869 67432
rect 11395 67431 11453 67432
rect 19756 67388 19796 67432
rect 547 67348 556 67388
rect 596 67348 2956 67388
rect 2996 67348 12748 67388
rect 12788 67348 12797 67388
rect 13795 67348 13804 67388
rect 13844 67348 14092 67388
rect 14132 67348 14141 67388
rect 19747 67348 19756 67388
rect 19796 67348 19805 67388
rect 0 67304 80 67324
rect 3427 67304 3485 67305
rect 0 67264 3436 67304
rect 3476 67264 3485 67304
rect 4919 67264 4928 67304
rect 4968 67264 5010 67304
rect 5050 67264 5092 67304
rect 5132 67264 5174 67304
rect 5214 67264 5256 67304
rect 5296 67264 5305 67304
rect 6019 67264 6028 67304
rect 6068 67264 15628 67304
rect 15668 67264 15677 67304
rect 20039 67264 20048 67304
rect 20088 67264 20130 67304
rect 20170 67264 20212 67304
rect 20252 67264 20294 67304
rect 20334 67264 20376 67304
rect 20416 67264 20425 67304
rect 0 67244 80 67264
rect 3427 67263 3485 67264
rect 13507 67220 13565 67221
rect 2860 67180 5356 67220
rect 5396 67180 5405 67220
rect 6115 67180 6124 67220
rect 6164 67180 10252 67220
rect 10292 67180 10301 67220
rect 11683 67180 11692 67220
rect 11732 67180 11741 67220
rect 13507 67180 13516 67220
rect 13556 67180 13900 67220
rect 13940 67180 13949 67220
rect 67 67136 125 67137
rect 67 67096 76 67136
rect 116 67096 2572 67136
rect 2612 67096 2621 67136
rect 67 67095 125 67096
rect 2860 67052 2900 67180
rect 9187 67136 9245 67137
rect 11692 67136 11732 67180
rect 13507 67179 13565 67180
rect 6595 67096 6604 67136
rect 6644 67096 7084 67136
rect 7124 67096 7133 67136
rect 8035 67096 8044 67136
rect 8084 67096 8620 67136
rect 8660 67096 8669 67136
rect 9102 67096 9196 67136
rect 9236 67096 9245 67136
rect 11107 67096 11116 67136
rect 11156 67096 11732 67136
rect 12451 67136 12509 67137
rect 21424 67136 21504 67156
rect 12451 67096 12460 67136
rect 12500 67096 21504 67136
rect 9187 67095 9245 67096
rect 12451 67095 12509 67096
rect 21424 67076 21504 67096
rect 844 67012 2900 67052
rect 2947 67012 2956 67052
rect 2996 67012 3148 67052
rect 3188 67012 3197 67052
rect 3523 67012 3532 67052
rect 3572 67012 6796 67052
rect 6836 67012 6845 67052
rect 8899 67012 8908 67052
rect 8948 67012 9388 67052
rect 9428 67012 9437 67052
rect 9859 67012 9868 67052
rect 9908 67012 13364 67052
rect 0 66968 80 66988
rect 844 66968 884 67012
rect 2755 66968 2813 66969
rect 13324 66968 13364 67012
rect 0 66928 884 66968
rect 931 66928 940 66968
rect 980 66928 1708 66968
rect 1748 66928 1757 66968
rect 2755 66928 2764 66968
rect 2804 66928 11360 66968
rect 11491 66928 11500 66968
rect 11540 66928 11788 66968
rect 11828 66928 11837 66968
rect 12067 66928 12076 66968
rect 12116 66928 12940 66968
rect 12980 66928 12989 66968
rect 13315 66928 13324 66968
rect 13364 66928 14188 66968
rect 14228 66928 14764 66968
rect 14804 66928 15820 66968
rect 15860 66928 16876 66968
rect 16916 66928 16925 66968
rect 0 66908 80 66928
rect 2755 66927 2813 66928
rect 355 66884 413 66885
rect 11320 66884 11360 66928
rect 355 66844 364 66884
rect 404 66844 1228 66884
rect 1268 66844 5740 66884
rect 5780 66844 5789 66884
rect 7171 66844 7180 66884
rect 7220 66844 8044 66884
rect 8084 66844 8908 66884
rect 8948 66844 9868 66884
rect 9908 66844 9917 66884
rect 11320 66844 12556 66884
rect 12596 66844 12605 66884
rect 355 66843 413 66844
rect 739 66800 797 66801
rect 2947 66800 3005 66801
rect 4771 66800 4829 66801
rect 17539 66800 17597 66801
rect 19939 66800 19997 66801
rect 739 66760 748 66800
rect 788 66760 2956 66800
rect 2996 66760 3005 66800
rect 739 66759 797 66760
rect 2947 66759 3005 66760
rect 3052 66760 3436 66800
rect 3476 66760 3485 66800
rect 4483 66760 4492 66800
rect 4532 66760 4780 66800
rect 4820 66760 5356 66800
rect 5396 66760 5405 66800
rect 6595 66760 6604 66800
rect 6644 66760 9772 66800
rect 9812 66760 9821 66800
rect 11779 66760 11788 66800
rect 11828 66760 12172 66800
rect 12212 66760 12221 66800
rect 17454 66760 17548 66800
rect 17588 66760 17597 66800
rect 17923 66760 17932 66800
rect 17972 66760 19372 66800
rect 19412 66760 19421 66800
rect 19854 66760 19948 66800
rect 19988 66760 19997 66800
rect 3052 66716 3092 66760
rect 4771 66759 4829 66760
rect 17539 66759 17597 66760
rect 19939 66759 19997 66760
rect 7459 66716 7517 66717
rect 2947 66676 2956 66716
rect 2996 66676 3092 66716
rect 4387 66676 4396 66716
rect 4436 66676 4972 66716
rect 5012 66676 5021 66716
rect 5443 66676 5452 66716
rect 5492 66676 7468 66716
rect 7508 66676 7517 66716
rect 8323 66676 8332 66716
rect 8372 66676 12364 66716
rect 12404 66676 12413 66716
rect 17059 66676 17068 66716
rect 17108 66676 17356 66716
rect 17396 66676 17405 66716
rect 7459 66675 7517 66676
rect 0 66632 80 66652
rect 1123 66632 1181 66633
rect 6019 66632 6077 66633
rect 6307 66632 6365 66633
rect 12643 66632 12701 66633
rect 0 66592 1132 66632
rect 1172 66592 1181 66632
rect 5923 66592 5932 66632
rect 5972 66592 6028 66632
rect 6068 66592 6077 66632
rect 6222 66592 6316 66632
rect 6356 66592 6365 66632
rect 8227 66592 8236 66632
rect 8276 66592 8716 66632
rect 8756 66592 8765 66632
rect 11320 66592 11788 66632
rect 11828 66592 11837 66632
rect 12643 66592 12652 66632
rect 12692 66592 13036 66632
rect 13076 66592 13085 66632
rect 0 66572 80 66592
rect 1123 66591 1181 66592
rect 6019 66591 6077 66592
rect 6307 66591 6365 66592
rect 4579 66548 4637 66549
rect 2083 66508 2092 66548
rect 2132 66508 2284 66548
rect 2324 66508 2333 66548
rect 3679 66508 3688 66548
rect 3728 66508 3770 66548
rect 3810 66508 3852 66548
rect 3892 66508 3934 66548
rect 3974 66508 4016 66548
rect 4056 66508 4065 66548
rect 4579 66508 4588 66548
rect 4628 66508 6892 66548
rect 6932 66508 6941 66548
rect 4579 66507 4637 66508
rect 11320 66464 11360 66592
rect 12643 66591 12701 66592
rect 13123 66548 13181 66549
rect 11875 66508 11884 66548
rect 11924 66508 12172 66548
rect 12212 66508 12221 66548
rect 13038 66508 13132 66548
rect 13172 66508 13181 66548
rect 16003 66508 16012 66548
rect 16052 66508 16300 66548
rect 16340 66508 16349 66548
rect 18799 66508 18808 66548
rect 18848 66508 18890 66548
rect 18930 66508 18972 66548
rect 19012 66508 19054 66548
rect 19094 66508 19136 66548
rect 19176 66508 19185 66548
rect 13123 66507 13181 66508
rect 13027 66464 13085 66465
rect 16099 66464 16157 66465
rect 21424 66464 21504 66484
rect 2500 66424 11360 66464
rect 12835 66424 12844 66464
rect 12884 66424 13036 66464
rect 13076 66424 13085 66464
rect 13219 66424 13228 66464
rect 13268 66424 13277 66464
rect 16099 66424 16108 66464
rect 16148 66424 21504 66464
rect 0 66296 80 66316
rect 2500 66296 2540 66424
rect 13027 66423 13085 66424
rect 6883 66380 6941 66381
rect 13228 66380 13268 66424
rect 16099 66423 16157 66424
rect 21424 66404 21504 66424
rect 4291 66340 4300 66380
rect 4340 66340 6508 66380
rect 6548 66340 6557 66380
rect 6787 66340 6796 66380
rect 6836 66340 6892 66380
rect 6932 66340 6941 66380
rect 10243 66340 10252 66380
rect 10292 66340 13268 66380
rect 13795 66380 13853 66381
rect 13795 66340 13804 66380
rect 13844 66340 14956 66380
rect 14996 66340 15005 66380
rect 16579 66340 16588 66380
rect 16628 66340 16780 66380
rect 16820 66340 16829 66380
rect 6883 66339 6941 66340
rect 13795 66339 13853 66340
rect 4579 66296 4637 66297
rect 0 66256 2540 66296
rect 2668 66256 4588 66296
rect 4628 66256 4637 66296
rect 5539 66256 5548 66296
rect 5588 66256 8716 66296
rect 8756 66256 8765 66296
rect 9379 66256 9388 66296
rect 9428 66256 9964 66296
rect 10004 66256 10013 66296
rect 0 66236 80 66256
rect 2668 66212 2708 66256
rect 4579 66255 4637 66256
rect 2563 66172 2572 66212
rect 2612 66172 2708 66212
rect 3715 66172 3724 66212
rect 3764 66172 4492 66212
rect 4532 66172 4541 66212
rect 5059 66172 5068 66212
rect 5108 66172 8140 66212
rect 8180 66172 8189 66212
rect 11683 66172 11692 66212
rect 11732 66172 11884 66212
rect 11924 66172 11933 66212
rect 16867 66172 16876 66212
rect 16916 66172 17452 66212
rect 17492 66172 17501 66212
rect 8035 66128 8093 66129
rect 16003 66128 16061 66129
rect 3619 66088 3628 66128
rect 3668 66088 3916 66128
rect 3956 66088 3965 66128
rect 4099 66088 4108 66128
rect 4148 66088 6028 66128
rect 6068 66088 6316 66128
rect 6356 66088 6508 66128
rect 6548 66088 6557 66128
rect 7651 66088 7660 66128
rect 7700 66088 8044 66128
rect 8084 66088 8093 66128
rect 12835 66088 12844 66128
rect 12884 66088 13612 66128
rect 13652 66088 13661 66128
rect 15918 66088 16012 66128
rect 16052 66088 16061 66128
rect 16579 66088 16588 66128
rect 16628 66088 17260 66128
rect 17300 66088 17309 66128
rect 8035 66087 8093 66088
rect 16003 66087 16061 66088
rect 5539 66044 5597 66045
rect 16012 66044 16052 66087
rect 3523 66004 3532 66044
rect 3572 66004 4780 66044
rect 4820 66004 5164 66044
rect 5204 66004 5213 66044
rect 5443 66004 5452 66044
rect 5492 66004 5548 66044
rect 5588 66004 5597 66044
rect 9667 66004 9676 66044
rect 9716 66004 9725 66044
rect 11683 66004 11692 66044
rect 11732 66004 12460 66044
rect 12500 66004 13036 66044
rect 13076 66004 13085 66044
rect 13219 66004 13228 66044
rect 13268 66004 13708 66044
rect 13748 66004 13757 66044
rect 16012 66004 16684 66044
rect 16724 66004 16733 66044
rect 5539 66003 5597 66004
rect 0 65960 80 65980
rect 2851 65960 2909 65961
rect 9676 65960 9716 66004
rect 10339 65960 10397 65961
rect 14371 65960 14429 65961
rect 0 65920 2540 65960
rect 2659 65920 2668 65960
rect 2708 65920 2860 65960
rect 2900 65920 2909 65960
rect 4963 65920 4972 65960
rect 5012 65920 5021 65960
rect 5356 65920 6220 65960
rect 6260 65920 6269 65960
rect 8803 65920 8812 65960
rect 8852 65920 9484 65960
rect 9524 65920 9716 65960
rect 10147 65920 10156 65960
rect 10196 65920 10348 65960
rect 10388 65920 10397 65960
rect 13315 65920 13324 65960
rect 13364 65920 14188 65960
rect 14228 65920 14237 65960
rect 14286 65920 14380 65960
rect 14420 65920 14429 65960
rect 0 65900 80 65920
rect 2500 65876 2540 65920
rect 2851 65919 2909 65920
rect 4972 65876 5012 65920
rect 5356 65876 5396 65920
rect 10339 65919 10397 65920
rect 14371 65919 14429 65920
rect 13603 65876 13661 65877
rect 2500 65836 5012 65876
rect 5347 65836 5356 65876
rect 5396 65836 5405 65876
rect 8899 65836 8908 65876
rect 8948 65836 9676 65876
rect 9716 65836 9725 65876
rect 13518 65836 13612 65876
rect 13652 65836 13661 65876
rect 13603 65835 13661 65836
rect 7843 65792 7901 65793
rect 13411 65792 13469 65793
rect 21424 65792 21504 65812
rect 2179 65752 2188 65792
rect 2228 65752 4204 65792
rect 4244 65752 4253 65792
rect 4919 65752 4928 65792
rect 4968 65752 5010 65792
rect 5050 65752 5092 65792
rect 5132 65752 5174 65792
rect 5214 65752 5256 65792
rect 5296 65752 5305 65792
rect 5923 65752 5932 65792
rect 5972 65752 5981 65792
rect 6691 65752 6700 65792
rect 6740 65752 7180 65792
rect 7220 65752 7229 65792
rect 7651 65752 7660 65792
rect 7700 65752 7852 65792
rect 7892 65752 7901 65792
rect 12739 65752 12748 65792
rect 12788 65752 13420 65792
rect 13460 65752 13469 65792
rect 20039 65752 20048 65792
rect 20088 65752 20130 65792
rect 20170 65752 20212 65792
rect 20252 65752 20294 65792
rect 20334 65752 20376 65792
rect 20416 65752 20425 65792
rect 20524 65752 21504 65792
rect 5932 65708 5972 65752
rect 7843 65751 7901 65752
rect 13411 65751 13469 65752
rect 3331 65668 3340 65708
rect 3380 65668 3532 65708
rect 3572 65668 3581 65708
rect 4003 65668 4012 65708
rect 4052 65668 5972 65708
rect 6019 65708 6077 65709
rect 6019 65668 6028 65708
rect 6068 65668 15820 65708
rect 15860 65668 15869 65708
rect 6019 65667 6077 65668
rect 0 65624 80 65644
rect 3139 65624 3197 65625
rect 0 65584 2092 65624
rect 2132 65584 2141 65624
rect 3054 65584 3148 65624
rect 3188 65584 3197 65624
rect 0 65564 80 65584
rect 3139 65583 3197 65584
rect 3427 65624 3485 65625
rect 17443 65624 17501 65625
rect 20524 65624 20564 65752
rect 21424 65732 21504 65752
rect 3427 65584 3436 65624
rect 3476 65584 8044 65624
rect 8084 65584 8093 65624
rect 12355 65584 12364 65624
rect 12404 65584 13708 65624
rect 13748 65584 13757 65624
rect 17443 65584 17452 65624
rect 17492 65584 20564 65624
rect 3427 65583 3485 65584
rect 17443 65583 17501 65584
rect 547 65540 605 65541
rect 17635 65540 17693 65541
rect 547 65500 556 65540
rect 596 65500 3340 65540
rect 3380 65500 3389 65540
rect 6211 65500 6220 65540
rect 6260 65500 8620 65540
rect 8660 65500 8908 65540
rect 8948 65500 8957 65540
rect 12547 65500 12556 65540
rect 12596 65500 13324 65540
rect 13364 65500 13373 65540
rect 15724 65500 17452 65540
rect 17492 65500 17501 65540
rect 17635 65500 17644 65540
rect 17684 65500 17932 65540
rect 17972 65500 17981 65540
rect 547 65499 605 65500
rect 2083 65456 2141 65457
rect 15724 65456 15764 65500
rect 17635 65499 17693 65500
rect 15907 65456 15965 65457
rect 1603 65416 1612 65456
rect 1652 65416 2092 65456
rect 2132 65416 2141 65456
rect 3427 65416 3436 65456
rect 3476 65416 6412 65456
rect 6452 65416 6461 65456
rect 7267 65416 7276 65456
rect 7316 65416 7564 65456
rect 7604 65416 8236 65456
rect 8276 65416 8285 65456
rect 13123 65416 13132 65456
rect 13172 65416 13228 65456
rect 13268 65416 13277 65456
rect 14851 65416 14860 65456
rect 14900 65416 15724 65456
rect 15764 65416 15773 65456
rect 15907 65416 15916 65456
rect 15956 65416 18220 65456
rect 18260 65416 18269 65456
rect 2083 65415 2141 65416
rect 15907 65415 15965 65416
rect 1603 65372 1661 65373
rect 1795 65372 1853 65373
rect 9475 65372 9533 65373
rect 1603 65332 1612 65372
rect 1652 65332 1708 65372
rect 1748 65332 1804 65372
rect 1844 65332 1872 65372
rect 2572 65332 2956 65372
rect 2996 65332 3005 65372
rect 3523 65332 3532 65372
rect 3572 65332 4300 65372
rect 4340 65332 4349 65372
rect 4483 65332 4492 65372
rect 4532 65332 6604 65372
rect 6644 65332 6653 65372
rect 7171 65332 7180 65372
rect 7220 65332 9484 65372
rect 9524 65332 9533 65372
rect 10819 65332 10828 65372
rect 10868 65332 11884 65372
rect 11924 65332 12364 65372
rect 12404 65332 12413 65372
rect 12547 65332 12556 65372
rect 12596 65332 13036 65372
rect 13076 65332 13900 65372
rect 13940 65332 13949 65372
rect 16771 65332 16780 65372
rect 16820 65332 18604 65372
rect 18644 65332 18653 65372
rect 1603 65331 1661 65332
rect 1795 65331 1853 65332
rect 0 65288 80 65308
rect 2572 65288 2612 65332
rect 9475 65331 9533 65332
rect 6307 65288 6365 65289
rect 0 65248 1804 65288
rect 1844 65248 1853 65288
rect 2563 65248 2572 65288
rect 2612 65248 2621 65288
rect 4771 65248 4780 65288
rect 4820 65248 5164 65288
rect 5204 65248 5213 65288
rect 6307 65248 6316 65288
rect 6356 65248 6412 65288
rect 6452 65248 6461 65288
rect 6979 65248 6988 65288
rect 7028 65248 9196 65288
rect 9236 65248 9245 65288
rect 11299 65248 11308 65288
rect 11348 65248 12748 65288
rect 12788 65248 13420 65288
rect 13460 65248 13469 65288
rect 16387 65248 16396 65288
rect 16436 65248 17836 65288
rect 17876 65248 17885 65288
rect 0 65228 80 65248
rect 6307 65247 6365 65248
rect 5539 65204 5597 65205
rect 163 65164 172 65204
rect 212 65164 3532 65204
rect 3572 65164 3581 65204
rect 5539 65164 5548 65204
rect 5588 65164 5740 65204
rect 5780 65164 5789 65204
rect 6595 65164 6604 65204
rect 6644 65164 7756 65204
rect 7796 65164 11360 65204
rect 12355 65164 12364 65204
rect 12404 65164 14860 65204
rect 14900 65164 14909 65204
rect 5539 65163 5597 65164
rect 11320 65120 11360 65164
rect 21424 65120 21504 65140
rect 2083 65080 2092 65120
rect 2132 65080 2476 65120
rect 2516 65080 4780 65120
rect 4820 65080 4829 65120
rect 5539 65080 5548 65120
rect 5588 65080 6796 65120
rect 6836 65080 7948 65120
rect 7988 65080 7997 65120
rect 11320 65080 14476 65120
rect 14516 65080 14525 65120
rect 16675 65080 16684 65120
rect 16724 65080 21504 65120
rect 21424 65060 21504 65080
rect 1315 64996 1324 65036
rect 1364 64996 1516 65036
rect 1556 64996 1565 65036
rect 1795 64996 1804 65036
rect 1844 64996 2572 65036
rect 2612 64996 2621 65036
rect 3679 64996 3688 65036
rect 3728 64996 3770 65036
rect 3810 64996 3852 65036
rect 3892 64996 3934 65036
rect 3974 64996 4016 65036
rect 4056 64996 4065 65036
rect 5164 64996 10060 65036
rect 10100 64996 10109 65036
rect 13027 64996 13036 65036
rect 13076 64996 13516 65036
rect 13556 64996 13565 65036
rect 18799 64996 18808 65036
rect 18848 64996 18890 65036
rect 18930 64996 18972 65036
rect 19012 64996 19054 65036
rect 19094 64996 19136 65036
rect 19176 64996 19185 65036
rect 0 64952 80 64972
rect 5164 64952 5204 64996
rect 0 64912 5204 64952
rect 5251 64912 5260 64952
rect 5300 64912 9580 64952
rect 9620 64912 9629 64952
rect 12739 64912 12748 64952
rect 12788 64912 13804 64952
rect 13844 64912 18412 64952
rect 18452 64912 18461 64952
rect 0 64892 80 64912
rect 931 64868 989 64869
rect 5923 64868 5981 64869
rect 13123 64868 13181 64869
rect 931 64828 940 64868
rect 980 64828 5932 64868
rect 5972 64828 5981 64868
rect 11011 64828 11020 64868
rect 11060 64828 11308 64868
rect 11348 64828 11357 64868
rect 12355 64828 12364 64868
rect 12404 64828 13132 64868
rect 13172 64828 14284 64868
rect 14324 64828 14333 64868
rect 14467 64828 14476 64868
rect 14516 64828 14764 64868
rect 14804 64828 14813 64868
rect 931 64827 989 64828
rect 5923 64827 5981 64828
rect 13123 64827 13181 64828
rect 2500 64744 10540 64784
rect 10580 64744 10924 64784
rect 10964 64744 10973 64784
rect 11320 64744 14092 64784
rect 14132 64744 14141 64784
rect 1315 64700 1373 64701
rect 2500 64700 2540 64744
rect 8611 64700 8669 64701
rect 1315 64660 1324 64700
rect 1364 64660 2540 64700
rect 2659 64660 2668 64700
rect 2708 64660 2956 64700
rect 2996 64660 3005 64700
rect 3436 64660 4012 64700
rect 4052 64660 4061 64700
rect 4771 64660 4780 64700
rect 4820 64660 6700 64700
rect 6740 64660 6749 64700
rect 8526 64660 8620 64700
rect 8660 64660 8669 64700
rect 1315 64659 1373 64660
rect 0 64616 80 64636
rect 3436 64616 3476 64660
rect 8611 64659 8669 64660
rect 9475 64700 9533 64701
rect 11320 64700 11360 64744
rect 9475 64660 9484 64700
rect 9524 64660 11360 64700
rect 11875 64660 11884 64700
rect 11924 64660 14188 64700
rect 14228 64660 14380 64700
rect 14420 64660 14429 64700
rect 14851 64660 14860 64700
rect 14900 64660 15340 64700
rect 15380 64660 19660 64700
rect 19700 64660 19709 64700
rect 9475 64659 9533 64660
rect 0 64576 1324 64616
rect 1364 64576 1373 64616
rect 2755 64576 2764 64616
rect 2804 64576 3476 64616
rect 3523 64576 3532 64616
rect 3572 64576 9620 64616
rect 10435 64576 10444 64616
rect 10484 64576 11020 64616
rect 11060 64576 11069 64616
rect 12931 64576 12940 64616
rect 12980 64576 13516 64616
rect 13556 64576 13565 64616
rect 0 64556 80 64576
rect 9580 64532 9620 64576
rect 2275 64492 2284 64532
rect 2324 64492 7180 64532
rect 7220 64492 7229 64532
rect 9571 64492 9580 64532
rect 9620 64492 12748 64532
rect 12788 64492 12797 64532
rect 13027 64492 13036 64532
rect 13076 64492 13708 64532
rect 13748 64492 13757 64532
rect 13804 64492 20180 64532
rect 11107 64448 11165 64449
rect 13603 64448 13661 64449
rect 13804 64448 13844 64492
rect 5347 64408 5356 64448
rect 5396 64408 6028 64448
rect 6068 64408 6077 64448
rect 6787 64408 6796 64448
rect 6836 64408 7372 64448
rect 7412 64408 7421 64448
rect 11022 64408 11116 64448
rect 11156 64408 11165 64448
rect 11107 64407 11165 64408
rect 12268 64408 12556 64448
rect 12596 64408 12844 64448
rect 12884 64408 13324 64448
rect 13364 64408 13373 64448
rect 13603 64408 13612 64448
rect 13652 64408 13844 64448
rect 15523 64408 15532 64448
rect 15572 64408 16204 64448
rect 16244 64408 16253 64448
rect 17443 64408 17452 64448
rect 17492 64408 17932 64448
rect 17972 64408 17981 64448
rect 5923 64364 5981 64365
rect 2092 64324 2764 64364
rect 2804 64324 3244 64364
rect 3284 64324 3293 64364
rect 5838 64324 5932 64364
rect 5972 64324 5981 64364
rect 0 64280 80 64300
rect 2092 64280 2132 64324
rect 5923 64323 5981 64324
rect 7948 64324 9004 64364
rect 9044 64324 9236 64364
rect 2659 64280 2717 64281
rect 7948 64280 7988 64324
rect 9196 64280 9236 64324
rect 12268 64280 12308 64408
rect 13603 64407 13661 64408
rect 20140 64364 20180 64492
rect 21424 64448 21504 64468
rect 21196 64408 21504 64448
rect 21196 64364 21236 64408
rect 21424 64388 21504 64408
rect 13507 64324 13516 64364
rect 13556 64324 13804 64364
rect 13844 64324 13853 64364
rect 14659 64324 14668 64364
rect 14708 64324 15476 64364
rect 15715 64324 15724 64364
rect 15764 64324 18028 64364
rect 18068 64324 18077 64364
rect 20140 64324 21236 64364
rect 15436 64281 15476 64324
rect 13411 64280 13469 64281
rect 15427 64280 15485 64281
rect 0 64240 2132 64280
rect 2574 64240 2668 64280
rect 2708 64240 2717 64280
rect 4919 64240 4928 64280
rect 4968 64240 5010 64280
rect 5050 64240 5092 64280
rect 5132 64240 5174 64280
rect 5214 64240 5256 64280
rect 5296 64240 5305 64280
rect 7908 64240 7948 64280
rect 7988 64240 7997 64280
rect 9187 64240 9196 64280
rect 9236 64240 9245 64280
rect 12259 64240 12268 64280
rect 12308 64240 12317 64280
rect 12364 64240 13228 64280
rect 13268 64240 13420 64280
rect 13460 64240 13469 64280
rect 15396 64240 15436 64280
rect 15476 64240 15485 64280
rect 20039 64240 20048 64280
rect 20088 64240 20130 64280
rect 20170 64240 20212 64280
rect 20252 64240 20294 64280
rect 20334 64240 20376 64280
rect 20416 64240 20425 64280
rect 0 64220 80 64240
rect 2659 64239 2717 64240
rect 12364 64197 12404 64240
rect 13411 64239 13469 64240
rect 15427 64239 15485 64240
rect 11107 64196 11165 64197
rect 12355 64196 12413 64197
rect 1891 64156 1900 64196
rect 1940 64156 2540 64196
rect 9955 64156 9964 64196
rect 10004 64156 11116 64196
rect 11156 64156 11360 64196
rect 2500 64028 2540 64156
rect 11107 64155 11165 64156
rect 4099 64112 4157 64113
rect 5539 64112 5597 64113
rect 6019 64112 6077 64113
rect 6883 64112 6941 64113
rect 7555 64112 7613 64113
rect 8323 64112 8381 64113
rect 10627 64112 10685 64113
rect 3811 64072 3820 64112
rect 3860 64072 4108 64112
rect 4148 64072 4157 64112
rect 5443 64072 5452 64112
rect 5492 64072 5548 64112
rect 5588 64072 5597 64112
rect 5827 64072 5836 64112
rect 5876 64072 6028 64112
rect 6068 64072 6077 64112
rect 6787 64072 6796 64112
rect 6836 64072 6892 64112
rect 6932 64072 6941 64112
rect 7171 64072 7180 64112
rect 7220 64072 7564 64112
rect 7604 64072 7613 64112
rect 8238 64072 8332 64112
rect 8372 64072 8381 64112
rect 10051 64072 10060 64112
rect 10100 64072 10348 64112
rect 10388 64072 10397 64112
rect 10542 64072 10636 64112
rect 10676 64072 10685 64112
rect 11320 64112 11360 64156
rect 12355 64156 12364 64196
rect 12404 64156 12413 64196
rect 14755 64156 14764 64196
rect 14804 64156 16012 64196
rect 16052 64156 16061 64196
rect 12355 64155 12413 64156
rect 11320 64072 15724 64112
rect 15764 64072 15773 64112
rect 15907 64072 15916 64112
rect 15956 64072 16780 64112
rect 16820 64072 16829 64112
rect 4099 64071 4157 64072
rect 5539 64071 5597 64072
rect 6019 64071 6077 64072
rect 6883 64071 6941 64072
rect 7555 64071 7613 64072
rect 8323 64071 8381 64072
rect 10627 64071 10685 64072
rect 10147 64028 10205 64029
rect 13027 64028 13085 64029
rect 2500 63988 6068 64028
rect 0 63944 80 63964
rect 1411 63944 1469 63945
rect 6028 63944 6068 63988
rect 10147 63988 10156 64028
rect 10196 63988 10252 64028
rect 10292 63988 10301 64028
rect 10531 63988 10540 64028
rect 10580 63988 10924 64028
rect 10964 63988 10973 64028
rect 12931 63988 12940 64028
rect 12980 63988 13036 64028
rect 13076 63988 17644 64028
rect 17684 63988 17693 64028
rect 10147 63987 10205 63988
rect 13027 63987 13085 63988
rect 9091 63944 9149 63945
rect 10915 63944 10973 63945
rect 0 63904 1420 63944
rect 1460 63904 3148 63944
rect 3188 63904 3197 63944
rect 4579 63904 4588 63944
rect 4628 63904 5548 63944
rect 5588 63904 5740 63944
rect 5780 63904 5789 63944
rect 6019 63904 6028 63944
rect 6068 63904 7084 63944
rect 7124 63904 7133 63944
rect 7363 63904 7372 63944
rect 7412 63904 7756 63944
rect 7796 63904 7805 63944
rect 8803 63904 8812 63944
rect 8852 63904 9100 63944
rect 9140 63904 10828 63944
rect 10868 63904 10924 63944
rect 10964 63904 10992 63944
rect 12067 63904 12076 63944
rect 12116 63904 12268 63944
rect 12308 63904 12460 63944
rect 12500 63904 12509 63944
rect 13795 63904 13804 63944
rect 13844 63904 14668 63944
rect 14708 63904 15724 63944
rect 15764 63904 15773 63944
rect 15907 63904 15916 63944
rect 15956 63904 16396 63944
rect 16436 63904 16445 63944
rect 17342 63904 17351 63944
rect 17391 63904 18316 63944
rect 18356 63904 18365 63944
rect 0 63884 80 63904
rect 1411 63903 1469 63904
rect 9091 63903 9149 63904
rect 10915 63903 10973 63904
rect 2500 63820 14284 63860
rect 14324 63820 14333 63860
rect 15331 63820 15340 63860
rect 15380 63820 16204 63860
rect 16244 63820 16253 63860
rect 2500 63776 2540 63820
rect 21424 63776 21504 63796
rect 1123 63736 1132 63776
rect 1172 63736 2540 63776
rect 7075 63736 7084 63776
rect 7124 63736 9580 63776
rect 9620 63736 9629 63776
rect 12547 63736 12556 63776
rect 12596 63736 14860 63776
rect 14900 63736 14909 63776
rect 16483 63736 16492 63776
rect 16532 63736 16780 63776
rect 16820 63736 16829 63776
rect 18019 63736 18028 63776
rect 18068 63736 18220 63776
rect 18260 63736 18269 63776
rect 21091 63736 21100 63776
rect 21140 63736 21504 63776
rect 21424 63716 21504 63736
rect 8035 63692 8093 63693
rect 16963 63692 17021 63693
rect 6979 63652 6988 63692
rect 7028 63652 7468 63692
rect 7508 63652 7517 63692
rect 8035 63652 8044 63692
rect 8084 63652 8428 63692
rect 8468 63652 8477 63692
rect 8611 63652 8620 63692
rect 8660 63652 9292 63692
rect 9332 63652 9341 63692
rect 16878 63652 16972 63692
rect 17012 63652 17021 63692
rect 8035 63651 8093 63652
rect 16963 63651 17021 63652
rect 0 63608 80 63628
rect 0 63568 7948 63608
rect 7988 63568 7997 63608
rect 8803 63568 8812 63608
rect 8852 63568 10060 63608
rect 10100 63568 10109 63608
rect 10531 63568 10540 63608
rect 10580 63568 11020 63608
rect 11060 63568 11069 63608
rect 0 63548 80 63568
rect 7459 63524 7517 63525
rect 11107 63524 11165 63525
rect 3679 63484 3688 63524
rect 3728 63484 3770 63524
rect 3810 63484 3852 63524
rect 3892 63484 3934 63524
rect 3974 63484 4016 63524
rect 4056 63484 4065 63524
rect 7459 63484 7468 63524
rect 7508 63484 11060 63524
rect 7459 63483 7517 63484
rect 1987 63440 2045 63441
rect 7555 63440 7613 63441
rect 1987 63400 1996 63440
rect 2036 63400 2540 63440
rect 1987 63399 2045 63400
rect 2500 63356 2540 63400
rect 7555 63400 7564 63440
rect 7604 63400 7660 63440
rect 7700 63400 7709 63440
rect 7843 63400 7852 63440
rect 7892 63400 7901 63440
rect 8131 63400 8140 63440
rect 8180 63400 8524 63440
rect 8564 63400 8573 63440
rect 9379 63400 9388 63440
rect 9428 63400 10732 63440
rect 10772 63400 10781 63440
rect 7555 63399 7613 63400
rect 3139 63356 3197 63357
rect 7852 63356 7892 63400
rect 8323 63356 8381 63357
rect 11020 63356 11060 63484
rect 11107 63484 11116 63524
rect 11156 63484 11212 63524
rect 11252 63484 11261 63524
rect 18799 63484 18808 63524
rect 18848 63484 18890 63524
rect 18930 63484 18972 63524
rect 19012 63484 19054 63524
rect 19094 63484 19136 63524
rect 19176 63484 19185 63524
rect 11107 63483 11165 63484
rect 12643 63440 12701 63441
rect 19843 63440 19901 63441
rect 12643 63400 12652 63440
rect 12692 63400 13132 63440
rect 13172 63400 13181 63440
rect 19843 63400 19852 63440
rect 19892 63400 20716 63440
rect 20756 63400 20765 63440
rect 12643 63399 12701 63400
rect 19843 63399 19901 63400
rect 2500 63316 3148 63356
rect 3188 63316 3197 63356
rect 3331 63316 3340 63356
rect 3380 63316 3724 63356
rect 3764 63316 7892 63356
rect 8035 63316 8044 63356
rect 8084 63316 8332 63356
rect 8372 63316 10252 63356
rect 10292 63316 10301 63356
rect 11020 63316 16300 63356
rect 16340 63316 16349 63356
rect 17539 63316 17548 63356
rect 17588 63316 17932 63356
rect 17972 63316 18220 63356
rect 18260 63316 18269 63356
rect 3139 63315 3197 63316
rect 8323 63315 8381 63316
rect 0 63272 80 63292
rect 10051 63272 10109 63273
rect 0 63232 2132 63272
rect 2947 63232 2956 63272
rect 2996 63232 3532 63272
rect 3572 63232 3581 63272
rect 5932 63232 9964 63272
rect 10004 63232 10060 63272
rect 10100 63232 10128 63272
rect 10915 63232 10924 63272
rect 10964 63232 11348 63272
rect 11395 63232 11404 63272
rect 11444 63232 12076 63272
rect 12116 63232 12125 63272
rect 18403 63232 18412 63272
rect 18452 63232 18700 63272
rect 18740 63232 18749 63272
rect 0 63212 80 63232
rect 1699 63020 1757 63021
rect 1411 62980 1420 63020
rect 1460 62980 1708 63020
rect 1748 62980 1757 63020
rect 2092 63020 2132 63232
rect 2371 63148 2380 63188
rect 2420 63148 3340 63188
rect 3380 63148 3389 63188
rect 2851 63104 2909 63105
rect 3139 63104 3197 63105
rect 5932 63104 5972 63232
rect 10051 63231 10109 63232
rect 11308 63188 11348 63232
rect 6691 63148 6700 63188
rect 6740 63148 7180 63188
rect 7220 63148 8812 63188
rect 8852 63148 8861 63188
rect 9859 63148 9868 63188
rect 9908 63148 11212 63188
rect 11252 63148 11261 63188
rect 11308 63148 16532 63188
rect 11320 63104 11360 63148
rect 16492 63104 16532 63148
rect 21283 63104 21341 63105
rect 21424 63104 21504 63124
rect 2851 63064 2860 63104
rect 2900 63064 2956 63104
rect 2996 63064 3005 63104
rect 3139 63064 3148 63104
rect 3188 63064 5932 63104
rect 5972 63064 5981 63104
rect 7363 63064 7372 63104
rect 7412 63064 7660 63104
rect 7700 63064 8044 63104
rect 8084 63064 8093 63104
rect 8323 63064 8332 63104
rect 8372 63064 8716 63104
rect 8756 63064 8765 63104
rect 10051 63064 10060 63104
rect 10100 63064 10109 63104
rect 10435 63064 10444 63104
rect 10484 63064 10924 63104
rect 10964 63064 10973 63104
rect 11212 63064 11360 63104
rect 13219 63064 13228 63104
rect 13268 63064 13277 63104
rect 16483 63064 16492 63104
rect 16532 63064 16541 63104
rect 17923 63064 17932 63104
rect 17972 63064 18316 63104
rect 18356 63064 18365 63104
rect 21283 63064 21292 63104
rect 21332 63064 21504 63104
rect 2851 63063 2909 63064
rect 3139 63063 3197 63064
rect 2947 63020 3005 63021
rect 4483 63020 4541 63021
rect 7843 63020 7901 63021
rect 9955 63020 10013 63021
rect 2092 62980 2708 63020
rect 1699 62979 1757 62980
rect 0 62936 80 62956
rect 1603 62936 1661 62937
rect 2668 62936 2708 62980
rect 2947 62980 2956 63020
rect 2996 62980 3052 63020
rect 3092 62980 3101 63020
rect 4398 62980 4492 63020
rect 4532 62980 4541 63020
rect 5731 62980 5740 63020
rect 5780 62980 7756 63020
rect 7796 62980 7852 63020
rect 7892 62980 7920 63020
rect 9870 62980 9964 63020
rect 10004 62980 10013 63020
rect 10060 63020 10100 63064
rect 10060 62980 10828 63020
rect 10868 62980 10877 63020
rect 2947 62979 3005 62980
rect 4483 62979 4541 62980
rect 7843 62979 7901 62980
rect 9955 62979 10013 62980
rect 5923 62936 5981 62937
rect 10915 62936 10973 62937
rect 11212 62936 11252 63064
rect 11299 63020 11357 63021
rect 13228 63020 13268 63064
rect 21283 63063 21341 63064
rect 21424 63044 21504 63064
rect 11299 62980 11308 63020
rect 11348 62980 13268 63020
rect 19555 63020 19613 63021
rect 19555 62980 19564 63020
rect 19604 62980 19948 63020
rect 19988 62980 19997 63020
rect 11299 62979 11357 62980
rect 19555 62979 19613 62980
rect 0 62896 1612 62936
rect 1652 62896 1661 62936
rect 2659 62896 2668 62936
rect 2708 62896 2717 62936
rect 5923 62896 5932 62936
rect 5972 62896 6028 62936
rect 6068 62896 6077 62936
rect 10723 62896 10732 62936
rect 10772 62896 10924 62936
rect 10964 62896 10973 62936
rect 11203 62896 11212 62936
rect 11252 62896 11261 62936
rect 0 62876 80 62896
rect 1603 62895 1661 62896
rect 5923 62895 5981 62896
rect 10915 62895 10973 62896
rect 2371 62852 2429 62853
rect 6115 62852 6173 62853
rect 2371 62812 2380 62852
rect 2420 62812 6124 62852
rect 6164 62812 6173 62852
rect 2371 62811 2429 62812
rect 6115 62811 6173 62812
rect 7555 62852 7613 62853
rect 7555 62812 7564 62852
rect 7604 62812 7660 62852
rect 7700 62812 7709 62852
rect 11587 62812 11596 62852
rect 11636 62812 11788 62852
rect 11828 62812 11837 62852
rect 7555 62811 7613 62812
rect 2659 62768 2717 62769
rect 9187 62768 9245 62769
rect 2659 62728 2668 62768
rect 2708 62728 2764 62768
rect 2804 62728 2813 62768
rect 3043 62728 3052 62768
rect 3092 62728 3724 62768
rect 3764 62728 3773 62768
rect 4919 62728 4928 62768
rect 4968 62728 5010 62768
rect 5050 62728 5092 62768
rect 5132 62728 5174 62768
rect 5214 62728 5256 62768
rect 5296 62728 5305 62768
rect 9187 62728 9196 62768
rect 9236 62728 12460 62768
rect 12500 62728 12509 62768
rect 15235 62728 15244 62768
rect 15284 62728 16396 62768
rect 16436 62728 16445 62768
rect 20039 62728 20048 62768
rect 20088 62728 20130 62768
rect 20170 62728 20212 62768
rect 20252 62728 20294 62768
rect 20334 62728 20376 62768
rect 20416 62728 20425 62768
rect 2659 62727 2717 62728
rect 9187 62727 9245 62728
rect 4771 62684 4829 62685
rect 9667 62684 9725 62685
rect 2467 62644 2476 62684
rect 2516 62644 4300 62684
rect 4340 62644 4780 62684
rect 4820 62644 5452 62684
rect 5492 62644 7084 62684
rect 7124 62644 7133 62684
rect 9667 62644 9676 62684
rect 9716 62644 21004 62684
rect 21044 62644 21053 62684
rect 4771 62643 4829 62644
rect 9667 62643 9725 62644
rect 0 62600 80 62620
rect 13507 62600 13565 62601
rect 0 62560 1996 62600
rect 2036 62560 2045 62600
rect 4483 62560 4492 62600
rect 4532 62560 4780 62600
rect 4820 62560 4829 62600
rect 6883 62560 6892 62600
rect 6932 62560 9196 62600
rect 9236 62560 9245 62600
rect 9379 62560 9388 62600
rect 9428 62560 9676 62600
rect 9716 62560 9725 62600
rect 9859 62560 9868 62600
rect 9908 62560 10348 62600
rect 10388 62560 10397 62600
rect 13507 62560 13516 62600
rect 13556 62560 13708 62600
rect 13748 62560 13757 62600
rect 15043 62560 15052 62600
rect 15092 62560 16588 62600
rect 16628 62560 16637 62600
rect 0 62540 80 62560
rect 13507 62559 13565 62560
rect 8323 62516 8381 62517
rect 8323 62476 8332 62516
rect 8372 62476 20524 62516
rect 20564 62476 20573 62516
rect 8323 62475 8381 62476
rect 1507 62432 1565 62433
rect 10627 62432 10685 62433
rect 21424 62432 21504 62452
rect 1507 62392 1516 62432
rect 1556 62392 1708 62432
rect 1748 62392 1757 62432
rect 4195 62392 4204 62432
rect 4244 62392 6316 62432
rect 6356 62392 6365 62432
rect 6883 62392 6892 62432
rect 6932 62392 7276 62432
rect 7316 62392 7468 62432
rect 7508 62392 7517 62432
rect 8995 62392 9004 62432
rect 9044 62392 9772 62432
rect 9812 62392 9821 62432
rect 10147 62392 10156 62432
rect 10196 62392 10636 62432
rect 10676 62392 10685 62432
rect 12451 62392 12460 62432
rect 12500 62392 15532 62432
rect 15572 62392 16012 62432
rect 16052 62392 16061 62432
rect 21283 62392 21292 62432
rect 21332 62392 21504 62432
rect 1507 62391 1565 62392
rect 10627 62391 10685 62392
rect 21424 62372 21504 62392
rect 9091 62308 9100 62348
rect 9140 62308 9676 62348
rect 9716 62308 9725 62348
rect 0 62264 80 62284
rect 7939 62264 7997 62265
rect 0 62224 7948 62264
rect 7988 62224 7997 62264
rect 0 62204 80 62224
rect 7939 62223 7997 62224
rect 10147 62264 10205 62265
rect 10147 62224 10156 62264
rect 10196 62224 10252 62264
rect 10292 62224 10301 62264
rect 11683 62224 11692 62264
rect 11732 62224 11980 62264
rect 12020 62224 12029 62264
rect 12547 62224 12556 62264
rect 12596 62224 14668 62264
rect 14708 62224 14717 62264
rect 15043 62224 15052 62264
rect 15092 62224 15340 62264
rect 15380 62224 15389 62264
rect 10147 62223 10205 62224
rect 3139 62180 3197 62181
rect 11683 62180 11741 62181
rect 12163 62180 12221 62181
rect 3054 62140 3148 62180
rect 3188 62140 3197 62180
rect 5827 62140 5836 62180
rect 5876 62140 11692 62180
rect 11732 62140 12172 62180
rect 12212 62140 12221 62180
rect 16003 62140 16012 62180
rect 16052 62140 16492 62180
rect 16532 62140 16541 62180
rect 3139 62139 3197 62140
rect 11683 62139 11741 62140
rect 12163 62139 12221 62140
rect 9763 62096 9821 62097
rect 17539 62096 17597 62097
rect 9763 62056 9772 62096
rect 9812 62056 17548 62096
rect 17588 62056 17597 62096
rect 9763 62055 9821 62056
rect 17539 62055 17597 62056
rect 3679 61972 3688 62012
rect 3728 61972 3770 62012
rect 3810 61972 3852 62012
rect 3892 61972 3934 62012
rect 3974 61972 4016 62012
rect 4056 61972 4065 62012
rect 18799 61972 18808 62012
rect 18848 61972 18890 62012
rect 18930 61972 18972 62012
rect 19012 61972 19054 62012
rect 19094 61972 19136 62012
rect 19176 61972 19185 62012
rect 0 61928 80 61948
rect 2659 61928 2717 61929
rect 0 61888 1612 61928
rect 1652 61888 1661 61928
rect 2659 61888 2668 61928
rect 2708 61888 5740 61928
rect 5780 61888 5789 61928
rect 7939 61888 7948 61928
rect 7988 61888 9580 61928
rect 9620 61888 9629 61928
rect 0 61868 80 61888
rect 2659 61887 2717 61888
rect 6403 61844 6461 61845
rect 7939 61844 7997 61845
rect 15523 61844 15581 61845
rect 3427 61804 3436 61844
rect 3476 61804 3724 61844
rect 3764 61804 3773 61844
rect 6403 61804 6412 61844
rect 6452 61804 7948 61844
rect 7988 61804 7997 61844
rect 8419 61804 8428 61844
rect 8468 61804 8840 61844
rect 15235 61804 15244 61844
rect 15284 61804 15532 61844
rect 15572 61804 15581 61844
rect 6403 61803 6461 61804
rect 7939 61803 7997 61804
rect 3907 61760 3965 61761
rect 3822 61720 3916 61760
rect 3956 61720 3965 61760
rect 3907 61719 3965 61720
rect 7747 61760 7805 61761
rect 8800 61760 8840 61804
rect 15523 61803 15581 61804
rect 21424 61760 21504 61780
rect 7747 61720 7756 61760
rect 7796 61720 7948 61760
rect 7988 61720 7997 61760
rect 8800 61720 9004 61760
rect 9044 61720 9053 61760
rect 15811 61720 15820 61760
rect 15860 61720 15869 61760
rect 17620 61720 20180 61760
rect 20707 61720 20716 61760
rect 20756 61720 21504 61760
rect 7747 61719 7805 61720
rect 2092 61636 2380 61676
rect 2420 61636 2429 61676
rect 3235 61636 3244 61676
rect 3284 61636 3820 61676
rect 3860 61636 4780 61676
rect 4820 61636 6988 61676
rect 7028 61636 7037 61676
rect 8707 61636 8716 61676
rect 8756 61636 10924 61676
rect 10964 61636 11360 61676
rect 13891 61636 13900 61676
rect 13940 61636 14956 61676
rect 14996 61636 15724 61676
rect 15764 61636 15773 61676
rect 0 61592 80 61612
rect 2092 61592 2132 61636
rect 11320 61592 11360 61636
rect 15820 61592 15860 61720
rect 15907 61676 15965 61677
rect 17620 61676 17660 61720
rect 15907 61636 15916 61676
rect 15956 61636 17660 61676
rect 15907 61635 15965 61636
rect 20140 61592 20180 61720
rect 21424 61700 21504 61720
rect 0 61552 2132 61592
rect 2179 61552 2188 61592
rect 2228 61552 2540 61592
rect 6499 61552 6508 61592
rect 6548 61552 6700 61592
rect 6740 61552 8332 61592
rect 8372 61552 8381 61592
rect 9667 61552 9676 61592
rect 9716 61552 11212 61592
rect 11252 61552 11261 61592
rect 11320 61552 11500 61592
rect 11540 61552 13420 61592
rect 13460 61552 13469 61592
rect 15811 61552 15820 61592
rect 15860 61552 15869 61592
rect 20140 61552 21388 61592
rect 21428 61552 21437 61592
rect 0 61532 80 61552
rect 2500 61508 2540 61552
rect 2500 61468 7564 61508
rect 7604 61468 7613 61508
rect 14371 61468 14380 61508
rect 14420 61468 15436 61508
rect 15476 61468 15485 61508
rect 14851 61384 14860 61424
rect 14900 61384 15724 61424
rect 15764 61384 15773 61424
rect 15916 61384 17452 61424
rect 17492 61384 17501 61424
rect 13027 61340 13085 61341
rect 15436 61340 15476 61384
rect 15916 61340 15956 61384
rect 6691 61300 6700 61340
rect 6740 61300 13036 61340
rect 13076 61300 13085 61340
rect 14947 61300 14956 61340
rect 14996 61300 15244 61340
rect 15284 61300 15293 61340
rect 15427 61300 15436 61340
rect 15476 61300 15485 61340
rect 15619 61300 15628 61340
rect 15668 61300 15956 61340
rect 16003 61340 16061 61341
rect 16003 61300 16012 61340
rect 16052 61300 17164 61340
rect 17204 61300 17213 61340
rect 13027 61299 13085 61300
rect 16003 61299 16061 61300
rect 0 61256 80 61276
rect 2179 61256 2237 61257
rect 0 61216 2188 61256
rect 2228 61216 3148 61256
rect 3188 61216 3197 61256
rect 4919 61216 4928 61256
rect 4968 61216 5010 61256
rect 5050 61216 5092 61256
rect 5132 61216 5174 61256
rect 5214 61216 5256 61256
rect 5296 61216 5305 61256
rect 14755 61216 14764 61256
rect 14804 61216 15916 61256
rect 15956 61216 15965 61256
rect 20039 61216 20048 61256
rect 20088 61216 20130 61256
rect 20170 61216 20212 61256
rect 20252 61216 20294 61256
rect 20334 61216 20376 61256
rect 20416 61216 20425 61256
rect 0 61196 80 61216
rect 2179 61215 2237 61216
rect 3331 61172 3389 61173
rect 15523 61172 15581 61173
rect 3331 61132 3340 61172
rect 3380 61132 6740 61172
rect 6787 61132 6796 61172
rect 6836 61132 7468 61172
rect 7508 61132 9484 61172
rect 9524 61132 9533 61172
rect 14179 61132 14188 61172
rect 14228 61132 14956 61172
rect 14996 61132 15005 61172
rect 15331 61132 15340 61172
rect 15380 61132 15532 61172
rect 15572 61132 15581 61172
rect 3331 61131 3389 61132
rect 4771 61088 4829 61089
rect 6700 61088 6740 61132
rect 15523 61131 15581 61132
rect 10819 61088 10877 61089
rect 11107 61088 11165 61089
rect 12259 61088 12317 61089
rect 13027 61088 13085 61089
rect 21424 61088 21504 61108
rect 2947 61048 2956 61088
rect 2996 61048 4780 61088
rect 4820 61048 4829 61088
rect 5635 61048 5644 61088
rect 5684 61048 6604 61088
rect 6644 61048 6653 61088
rect 6700 61048 9716 61088
rect 4771 61047 4829 61048
rect 4579 61004 4637 61005
rect 2755 60964 2764 61004
rect 2804 60964 3572 61004
rect 4494 60964 4588 61004
rect 4628 60964 4637 61004
rect 7843 60964 7852 61004
rect 7892 60964 8716 61004
rect 8756 60964 8765 61004
rect 8899 60964 8908 61004
rect 8948 60964 9100 61004
rect 9140 60964 9149 61004
rect 0 60920 80 60940
rect 3532 60920 3572 60964
rect 4579 60963 4637 60964
rect 5731 60920 5789 60921
rect 0 60860 116 60920
rect 2659 60880 2668 60920
rect 2708 60880 3436 60920
rect 3476 60880 3485 60920
rect 3532 60880 5068 60920
rect 5108 60880 5740 60920
rect 5780 60880 5789 60920
rect 6787 60880 6796 60920
rect 6836 60880 7180 60920
rect 7220 60880 8620 60920
rect 8660 60880 8669 60920
rect 5731 60879 5789 60880
rect 76 60836 116 60860
rect 76 60796 9292 60836
rect 9332 60796 9580 60836
rect 9620 60796 9629 60836
rect 4099 60712 4108 60752
rect 4148 60712 6700 60752
rect 6740 60712 6749 60752
rect 7843 60712 7852 60752
rect 7892 60712 8044 60752
rect 8084 60712 8093 60752
rect 9676 60668 9716 61048
rect 10819 61048 10828 61088
rect 10868 61048 10924 61088
rect 10964 61048 10973 61088
rect 11107 61048 11116 61088
rect 11156 61048 11250 61088
rect 12259 61048 12268 61088
rect 12308 61048 12364 61088
rect 12404 61048 12413 61088
rect 12739 61048 12748 61088
rect 12788 61048 13036 61088
rect 13076 61048 13085 61088
rect 14371 61048 14380 61088
rect 14420 61048 14429 61088
rect 14563 61048 14572 61088
rect 14612 61048 15628 61088
rect 15668 61048 15677 61088
rect 16003 61048 16012 61088
rect 16052 61048 16588 61088
rect 16628 61048 16637 61088
rect 21187 61048 21196 61088
rect 21236 61048 21504 61088
rect 10819 61047 10877 61048
rect 11107 61047 11165 61048
rect 12259 61047 12317 61048
rect 13027 61047 13085 61048
rect 12067 60964 12076 61004
rect 12116 60964 13996 61004
rect 14036 60964 14045 61004
rect 14380 60920 14420 61048
rect 21424 61028 21504 61048
rect 14467 60964 14476 61004
rect 14516 60964 15860 61004
rect 15820 60920 15860 60964
rect 12355 60880 12364 60920
rect 12404 60880 12413 60920
rect 12643 60880 12652 60920
rect 12692 60880 12844 60920
rect 12884 60880 12893 60920
rect 13027 60880 13036 60920
rect 13076 60880 13516 60920
rect 13556 60880 13565 60920
rect 14380 60880 14572 60920
rect 14612 60880 14621 60920
rect 15811 60880 15820 60920
rect 15860 60880 15869 60920
rect 16387 60880 16396 60920
rect 16436 60880 16684 60920
rect 16724 60880 16733 60920
rect 16963 60880 16972 60920
rect 17012 60880 17644 60920
rect 17684 60880 19468 60920
rect 19508 60880 19517 60920
rect 12364 60836 12404 60880
rect 13411 60836 13469 60837
rect 9763 60796 9772 60836
rect 9812 60796 11596 60836
rect 11636 60796 11884 60836
rect 11924 60796 11933 60836
rect 12364 60796 13420 60836
rect 13460 60796 13469 60836
rect 13411 60795 13469 60796
rect 10915 60712 10924 60752
rect 10964 60712 11212 60752
rect 11252 60712 11261 60752
rect 11971 60712 11980 60752
rect 12020 60712 18220 60752
rect 18260 60712 18269 60752
rect 15523 60668 15581 60669
rect 5155 60628 5164 60668
rect 5204 60628 8812 60668
rect 8852 60628 8861 60668
rect 9676 60628 12116 60668
rect 0 60584 80 60604
rect 12076 60584 12116 60628
rect 15523 60628 15532 60668
rect 15572 60628 15820 60668
rect 15860 60628 15869 60668
rect 17548 60628 17836 60668
rect 17876 60628 17885 60668
rect 15523 60627 15581 60628
rect 17548 60584 17588 60628
rect 0 60544 2284 60584
rect 2324 60544 3340 60584
rect 3380 60544 3389 60584
rect 5347 60544 5356 60584
rect 5396 60544 5836 60584
rect 5876 60544 5885 60584
rect 8515 60544 8524 60584
rect 8564 60544 8756 60584
rect 12076 60544 15628 60584
rect 15668 60544 15677 60584
rect 17539 60544 17548 60584
rect 17588 60544 17597 60584
rect 0 60524 80 60544
rect 6307 60500 6365 60501
rect 8611 60500 8669 60501
rect 3679 60460 3688 60500
rect 3728 60460 3770 60500
rect 3810 60460 3852 60500
rect 3892 60460 3934 60500
rect 3974 60460 4016 60500
rect 4056 60460 4065 60500
rect 5251 60460 5260 60500
rect 5300 60460 6316 60500
rect 6356 60460 8620 60500
rect 8660 60460 8669 60500
rect 6307 60459 6365 60460
rect 8611 60459 8669 60460
rect 8716 60500 8756 60544
rect 8716 60460 10444 60500
rect 10484 60460 14380 60500
rect 14420 60460 14429 60500
rect 17635 60460 17644 60500
rect 17684 60460 18124 60500
rect 18164 60460 18173 60500
rect 18799 60460 18808 60500
rect 18848 60460 18890 60500
rect 18930 60460 18972 60500
rect 19012 60460 19054 60500
rect 19094 60460 19136 60500
rect 19176 60460 19185 60500
rect 8716 60416 8756 60460
rect 11683 60416 11741 60417
rect 20995 60416 21053 60417
rect 21424 60416 21504 60436
rect 2500 60376 2956 60416
rect 2996 60376 4684 60416
rect 4724 60376 4733 60416
rect 5155 60376 5164 60416
rect 5204 60376 5548 60416
rect 5588 60376 5597 60416
rect 6403 60376 6412 60416
rect 6452 60376 7660 60416
rect 7700 60376 7709 60416
rect 8707 60376 8716 60416
rect 8756 60376 8765 60416
rect 8995 60376 9004 60416
rect 9044 60376 9868 60416
rect 9908 60376 9917 60416
rect 11598 60376 11692 60416
rect 11732 60376 11741 60416
rect 0 60248 80 60268
rect 2500 60248 2540 60376
rect 11683 60375 11741 60376
rect 12556 60376 13228 60416
rect 13268 60376 17740 60416
rect 17780 60376 18316 60416
rect 18356 60376 18365 60416
rect 20995 60376 21004 60416
rect 21044 60376 21504 60416
rect 2755 60332 2813 60333
rect 4675 60332 4733 60333
rect 5539 60332 5597 60333
rect 12556 60332 12596 60376
rect 20995 60375 21053 60376
rect 21424 60356 21504 60376
rect 13219 60332 13277 60333
rect 2755 60292 2764 60332
rect 2804 60292 3628 60332
rect 3668 60292 3677 60332
rect 4675 60292 4684 60332
rect 4724 60292 5548 60332
rect 5588 60292 5597 60332
rect 6595 60292 6604 60332
rect 6644 60292 12556 60332
rect 12596 60292 12605 60332
rect 13219 60292 13228 60332
rect 13268 60292 18604 60332
rect 18644 60292 18653 60332
rect 2755 60291 2813 60292
rect 4675 60291 4733 60292
rect 5539 60291 5597 60292
rect 13219 60291 13277 60292
rect 7459 60248 7517 60249
rect 0 60208 2540 60248
rect 5731 60208 5740 60248
rect 5780 60208 7468 60248
rect 7508 60208 7517 60248
rect 9283 60208 9292 60248
rect 9332 60208 16300 60248
rect 16340 60208 16349 60248
rect 0 60188 80 60208
rect 7459 60207 7517 60208
rect 8227 60164 8285 60165
rect 12259 60164 12317 60165
rect 2500 60124 6892 60164
rect 6932 60124 6941 60164
rect 7084 60124 7660 60164
rect 7700 60124 8236 60164
rect 8276 60124 8285 60164
rect 8899 60124 8908 60164
rect 8948 60124 8957 60164
rect 10915 60124 10924 60164
rect 10964 60124 11212 60164
rect 11252 60124 11261 60164
rect 12259 60124 12268 60164
rect 12308 60124 12460 60164
rect 12500 60124 12509 60164
rect 19075 60124 19084 60164
rect 19124 60124 19660 60164
rect 19700 60124 19709 60164
rect 2500 59996 2540 60124
rect 7084 60080 7124 60124
rect 8227 60123 8285 60124
rect 7075 60040 7084 60080
rect 7124 60040 7133 60080
rect 7267 60040 7276 60080
rect 7316 60040 8428 60080
rect 8468 60040 8477 60080
rect 1603 59956 1612 59996
rect 1652 59956 2540 59996
rect 2947 59956 2956 59996
rect 2996 59956 3340 59996
rect 3380 59956 3389 59996
rect 0 59912 80 59932
rect 8908 59912 8948 60124
rect 12259 60123 12317 60124
rect 12355 60080 12413 60081
rect 10723 60040 10732 60080
rect 10772 60040 10781 60080
rect 12355 60040 12364 60080
rect 12404 60040 12748 60080
rect 12788 60040 12797 60080
rect 14371 60040 14380 60080
rect 14420 60040 14764 60080
rect 14804 60040 14813 60080
rect 10732 59996 10772 60040
rect 12355 60039 12413 60040
rect 10732 59956 10828 59996
rect 10868 59956 10877 59996
rect 12835 59956 12844 59996
rect 12884 59956 13900 59996
rect 13940 59956 14668 59996
rect 14708 59956 14717 59996
rect 0 59872 212 59912
rect 2851 59872 2860 59912
rect 2900 59872 4780 59912
rect 4820 59872 4829 59912
rect 7267 59872 7276 59912
rect 7316 59872 8524 59912
rect 8564 59872 8573 59912
rect 8908 59872 9100 59912
rect 9140 59872 9149 59912
rect 10339 59872 10348 59912
rect 10388 59872 10924 59912
rect 10964 59872 10973 59912
rect 11683 59872 11692 59912
rect 11732 59872 15820 59912
rect 15860 59872 15869 59912
rect 18691 59872 18700 59912
rect 18740 59872 19276 59912
rect 19316 59872 19325 59912
rect 0 59852 80 59872
rect 172 59660 212 59872
rect 9571 59828 9629 59829
rect 2659 59788 2668 59828
rect 2708 59788 2956 59828
rect 2996 59788 3005 59828
rect 8995 59788 9004 59828
rect 9044 59788 9580 59828
rect 9620 59788 9629 59828
rect 10051 59788 10060 59828
rect 10100 59788 20812 59828
rect 20852 59788 20861 59828
rect 9571 59787 9629 59788
rect 21424 59744 21504 59764
rect 1507 59704 1516 59744
rect 1556 59704 4396 59744
rect 4436 59704 4445 59744
rect 4919 59704 4928 59744
rect 4968 59704 5010 59744
rect 5050 59704 5092 59744
rect 5132 59704 5174 59744
rect 5214 59704 5256 59744
rect 5296 59704 5305 59744
rect 20039 59704 20048 59744
rect 20088 59704 20130 59744
rect 20170 59704 20212 59744
rect 20252 59704 20294 59744
rect 20334 59704 20376 59744
rect 20416 59704 20425 59744
rect 20611 59704 20620 59744
rect 20660 59704 21504 59744
rect 21424 59684 21504 59704
rect 172 59620 9292 59660
rect 9332 59620 9341 59660
rect 0 59576 80 59596
rect 0 59536 2540 59576
rect 4387 59536 4396 59576
rect 4436 59536 6796 59576
rect 6836 59536 9868 59576
rect 9908 59536 9917 59576
rect 13795 59536 13804 59576
rect 13844 59536 14380 59576
rect 14420 59536 14429 59576
rect 0 59516 80 59536
rect 2500 59492 2540 59536
rect 16579 59492 16637 59493
rect 2500 59452 2668 59492
rect 2708 59452 12076 59492
rect 12116 59452 12364 59492
rect 12404 59452 12413 59492
rect 13027 59452 13036 59492
rect 13076 59452 13324 59492
rect 13364 59452 13373 59492
rect 16494 59452 16588 59492
rect 16628 59452 19276 59492
rect 19316 59452 19325 59492
rect 16579 59451 16637 59452
rect 9475 59408 9533 59409
rect 12643 59408 12701 59409
rect 13411 59408 13469 59409
rect 15619 59408 15677 59409
rect 2092 59368 5452 59408
rect 5492 59368 5501 59408
rect 6979 59368 6988 59408
rect 7028 59368 8913 59408
rect 8953 59368 8962 59408
rect 9390 59368 9484 59408
rect 9524 59368 9533 59408
rect 10435 59368 10444 59408
rect 10484 59368 10732 59408
rect 10772 59368 10781 59408
rect 12643 59368 12652 59408
rect 12692 59368 12940 59408
rect 12980 59368 12989 59408
rect 13411 59368 13420 59408
rect 13460 59368 14188 59408
rect 14228 59368 14237 59408
rect 15619 59368 15628 59408
rect 15668 59368 16300 59408
rect 16340 59368 16349 59408
rect 17251 59368 17260 59408
rect 17300 59368 17548 59408
rect 17588 59368 17597 59408
rect 2092 59324 2132 59368
rect 9475 59367 9533 59368
rect 12643 59367 12701 59368
rect 13411 59367 13469 59368
rect 15619 59367 15677 59368
rect 5635 59324 5693 59325
rect 2083 59284 2092 59324
rect 2132 59284 2141 59324
rect 5635 59284 5644 59324
rect 5684 59284 11308 59324
rect 11348 59284 14956 59324
rect 14996 59284 15005 59324
rect 17731 59284 17740 59324
rect 17780 59284 18124 59324
rect 18164 59284 18173 59324
rect 5635 59283 5693 59284
rect 0 59240 80 59260
rect 2659 59240 2717 59241
rect 6403 59240 6461 59241
rect 0 59200 500 59240
rect 0 59180 80 59200
rect 460 59156 500 59200
rect 2500 59200 2668 59240
rect 2708 59200 2717 59240
rect 5347 59200 5356 59240
rect 5396 59200 6412 59240
rect 6452 59200 6461 59240
rect 7747 59200 7756 59240
rect 7796 59200 8620 59240
rect 8660 59200 8669 59240
rect 10147 59200 10156 59240
rect 10196 59200 11788 59240
rect 11828 59200 11837 59240
rect 15235 59200 15244 59240
rect 15284 59200 16876 59240
rect 16916 59200 16925 59240
rect 17356 59200 17644 59240
rect 17684 59200 17693 59240
rect 18028 59200 18316 59240
rect 18356 59200 18365 59240
rect 2500 59156 2540 59200
rect 2659 59199 2717 59200
rect 6403 59199 6461 59200
rect 17356 59156 17396 59200
rect 17539 59156 17597 59157
rect 18028 59156 18068 59200
rect 460 59116 2540 59156
rect 17347 59116 17356 59156
rect 17396 59116 17405 59156
rect 17539 59116 17548 59156
rect 17588 59116 18028 59156
rect 18068 59116 18077 59156
rect 19075 59116 19084 59156
rect 19124 59116 19852 59156
rect 19892 59116 19901 59156
rect 17539 59115 17597 59116
rect 21424 59072 21504 59092
rect 4579 59032 4588 59072
rect 4628 59032 11596 59072
rect 11636 59032 11645 59072
rect 12355 59032 12364 59072
rect 12404 59032 12556 59072
rect 12596 59032 12605 59072
rect 20995 59032 21004 59072
rect 21044 59032 21504 59072
rect 21424 59012 21504 59032
rect 6403 58988 6461 58989
rect 3679 58948 3688 58988
rect 3728 58948 3770 58988
rect 3810 58948 3852 58988
rect 3892 58948 3934 58988
rect 3974 58948 4016 58988
rect 4056 58948 4065 58988
rect 6403 58948 6412 58988
rect 6452 58948 16012 58988
rect 16052 58948 16061 58988
rect 18799 58948 18808 58988
rect 18848 58948 18890 58988
rect 18930 58948 18972 58988
rect 19012 58948 19054 58988
rect 19094 58948 19136 58988
rect 19176 58948 19185 58988
rect 6403 58947 6461 58948
rect 0 58904 80 58924
rect 0 58864 1900 58904
rect 1940 58864 1949 58904
rect 3724 58864 11020 58904
rect 11060 58864 11069 58904
rect 11203 58864 11212 58904
rect 11252 58864 14092 58904
rect 14132 58864 14141 58904
rect 0 58844 80 58864
rect 3724 58820 3764 58864
rect 13411 58820 13469 58821
rect 3715 58780 3724 58820
rect 3764 58780 3773 58820
rect 6595 58780 6604 58820
rect 6644 58780 7180 58820
rect 7220 58780 7229 58820
rect 13411 58780 13420 58820
rect 13460 58780 13612 58820
rect 13652 58780 13661 58820
rect 16099 58780 16108 58820
rect 16148 58780 16588 58820
rect 16628 58780 16637 58820
rect 13411 58779 13469 58780
rect 4771 58736 4829 58737
rect 15331 58736 15389 58737
rect 2563 58696 2572 58736
rect 2612 58696 4780 58736
rect 4820 58696 4972 58736
rect 5012 58696 9964 58736
rect 10004 58696 11020 58736
rect 11060 58696 11069 58736
rect 11875 58696 11884 58736
rect 11924 58696 13652 58736
rect 4771 58695 4829 58696
rect 3331 58612 3340 58652
rect 3380 58612 5356 58652
rect 5396 58612 9004 58652
rect 9044 58612 9053 58652
rect 12547 58612 12556 58652
rect 12596 58612 12839 58652
rect 12879 58612 13516 58652
rect 13556 58612 13565 58652
rect 0 58568 80 58588
rect 13612 58568 13652 58696
rect 15331 58696 15340 58736
rect 15380 58696 15532 58736
rect 15572 58696 15581 58736
rect 15331 58695 15389 58696
rect 15427 58612 15436 58652
rect 15476 58612 16012 58652
rect 16052 58612 16340 58652
rect 16300 58568 16340 58612
rect 0 58528 11308 58568
rect 11348 58528 11357 58568
rect 11971 58528 11980 58568
rect 12020 58528 12940 58568
rect 12980 58528 12989 58568
rect 13603 58528 13612 58568
rect 13652 58528 13661 58568
rect 15139 58528 15148 58568
rect 15188 58528 16108 58568
rect 16148 58528 16157 58568
rect 16291 58528 16300 58568
rect 16340 58528 16349 58568
rect 0 58508 80 58528
rect 11299 58484 11357 58485
rect 6691 58444 6700 58484
rect 6740 58444 7084 58484
rect 7124 58444 7372 58484
rect 7412 58444 7421 58484
rect 8995 58444 9004 58484
rect 9044 58444 11308 58484
rect 11348 58444 11357 58484
rect 11299 58443 11357 58444
rect 12259 58484 12317 58485
rect 12259 58444 12268 58484
rect 12308 58444 20180 58484
rect 12259 58443 12317 58444
rect 20140 58400 20180 58444
rect 21424 58400 21504 58420
rect 5155 58360 5164 58400
rect 5204 58360 5548 58400
rect 5588 58360 5597 58400
rect 9955 58360 9964 58400
rect 10004 58360 10444 58400
rect 10484 58360 10493 58400
rect 11107 58360 11116 58400
rect 11156 58360 13036 58400
rect 13076 58360 13085 58400
rect 13219 58360 13228 58400
rect 13268 58360 13804 58400
rect 13844 58360 13853 58400
rect 20140 58360 21504 58400
rect 21424 58340 21504 58360
rect 1507 58276 1516 58316
rect 1556 58276 3724 58316
rect 3764 58276 3773 58316
rect 8800 58276 9772 58316
rect 9812 58276 18412 58316
rect 18452 58276 18461 58316
rect 0 58232 80 58252
rect 0 58192 4588 58232
rect 4628 58192 4637 58232
rect 4919 58192 4928 58232
rect 4968 58192 5010 58232
rect 5050 58192 5092 58232
rect 5132 58192 5174 58232
rect 5214 58192 5256 58232
rect 5296 58192 5305 58232
rect 0 58172 80 58192
rect 8800 58148 8840 58276
rect 10627 58192 10636 58232
rect 10676 58192 16780 58232
rect 16820 58192 16829 58232
rect 18211 58192 18220 58232
rect 18260 58192 18700 58232
rect 18740 58192 18749 58232
rect 20039 58192 20048 58232
rect 20088 58192 20130 58232
rect 20170 58192 20212 58232
rect 20252 58192 20294 58232
rect 20334 58192 20376 58232
rect 20416 58192 20425 58232
rect 6307 58108 6316 58148
rect 6356 58108 8840 58148
rect 10147 58108 10156 58148
rect 10196 58108 12556 58148
rect 12596 58108 12605 58148
rect 17827 58108 17836 58148
rect 17876 58108 18124 58148
rect 18164 58108 18173 58148
rect 4291 58024 4300 58064
rect 4340 58024 9620 58064
rect 9580 57981 9620 58024
rect 9571 57980 9629 57981
rect 5059 57940 5068 57980
rect 5108 57940 6124 57980
rect 6164 57940 6604 57980
rect 6644 57940 6653 57980
rect 9571 57940 9580 57980
rect 9620 57940 9629 57980
rect 11011 57940 11020 57980
rect 11060 57940 12940 57980
rect 12980 57940 12989 57980
rect 14083 57940 14092 57980
rect 14132 57940 19276 57980
rect 19316 57940 20044 57980
rect 20084 57940 20093 57980
rect 9571 57939 9629 57940
rect 0 57896 80 57916
rect 3139 57896 3197 57897
rect 6307 57896 6365 57897
rect 8515 57896 8573 57897
rect 0 57856 556 57896
rect 596 57856 605 57896
rect 3139 57856 3148 57896
rect 3188 57856 3628 57896
rect 3668 57856 3677 57896
rect 6222 57856 6316 57896
rect 6356 57856 6365 57896
rect 7555 57856 7564 57896
rect 7604 57856 8044 57896
rect 8084 57856 8180 57896
rect 8430 57856 8524 57896
rect 8564 57856 8573 57896
rect 9187 57856 9196 57896
rect 9236 57856 9580 57896
rect 9620 57856 9629 57896
rect 11683 57856 11692 57896
rect 11732 57856 11884 57896
rect 11924 57856 11933 57896
rect 16003 57856 16012 57896
rect 16052 57856 17644 57896
rect 17684 57856 17693 57896
rect 0 57836 80 57856
rect 3139 57855 3197 57856
rect 6307 57855 6365 57856
rect 8140 57812 8180 57856
rect 8515 57855 8573 57856
rect 9187 57812 9245 57813
rect 4099 57772 4108 57812
rect 4148 57772 4492 57812
rect 4532 57772 7852 57812
rect 7892 57772 7901 57812
rect 8140 57772 9196 57812
rect 9236 57772 10252 57812
rect 10292 57772 13516 57812
rect 13556 57772 14476 57812
rect 14516 57772 15340 57812
rect 15380 57772 15389 57812
rect 9187 57771 9245 57772
rect 17251 57728 17309 57729
rect 21424 57728 21504 57748
rect 8131 57688 8140 57728
rect 8180 57688 8812 57728
rect 8852 57688 8861 57728
rect 13315 57688 13324 57728
rect 13364 57688 13804 57728
rect 13844 57688 13853 57728
rect 17251 57688 17260 57728
rect 17300 57688 21504 57728
rect 17251 57687 17309 57688
rect 21424 57668 21504 57688
rect 6403 57644 6461 57645
rect 13027 57644 13085 57645
rect 6307 57604 6316 57644
rect 6356 57604 6412 57644
rect 6452 57604 6461 57644
rect 12163 57604 12172 57644
rect 12212 57604 13036 57644
rect 13076 57604 16396 57644
rect 16436 57604 17164 57644
rect 17204 57604 17213 57644
rect 6403 57603 6461 57604
rect 13027 57603 13085 57604
rect 0 57560 80 57580
rect 0 57520 1804 57560
rect 1844 57520 1853 57560
rect 9571 57520 9580 57560
rect 9620 57520 14764 57560
rect 14804 57520 15916 57560
rect 15956 57520 16876 57560
rect 16916 57520 19852 57560
rect 19892 57520 19901 57560
rect 0 57500 80 57520
rect 3679 57436 3688 57476
rect 3728 57436 3770 57476
rect 3810 57436 3852 57476
rect 3892 57436 3934 57476
rect 3974 57436 4016 57476
rect 4056 57436 4065 57476
rect 9859 57436 9868 57476
rect 9908 57436 10348 57476
rect 10388 57436 10397 57476
rect 11491 57436 11500 57476
rect 11540 57436 13324 57476
rect 13364 57436 13373 57476
rect 18799 57436 18808 57476
rect 18848 57436 18890 57476
rect 18930 57436 18972 57476
rect 19012 57436 19054 57476
rect 19094 57436 19136 57476
rect 19176 57436 19185 57476
rect 15331 57392 15389 57393
rect 15246 57352 15340 57392
rect 15380 57352 15389 57392
rect 15331 57351 15389 57352
rect 12931 57308 12989 57309
rect 16387 57308 16445 57309
rect 12931 57268 12940 57308
rect 12980 57268 14284 57308
rect 14324 57268 14333 57308
rect 16291 57268 16300 57308
rect 16340 57268 16396 57308
rect 16436 57268 16445 57308
rect 12931 57267 12989 57268
rect 16387 57267 16445 57268
rect 0 57224 80 57244
rect 0 57184 12364 57224
rect 12404 57184 12413 57224
rect 13891 57184 13900 57224
rect 13940 57184 13949 57224
rect 14371 57184 14380 57224
rect 14420 57184 14860 57224
rect 14900 57184 14909 57224
rect 18883 57184 18892 57224
rect 18932 57184 19564 57224
rect 19604 57184 19613 57224
rect 0 57164 80 57184
rect 7747 57100 7756 57140
rect 7796 57100 8044 57140
rect 8084 57100 8093 57140
rect 9667 57100 9676 57140
rect 9716 57100 10156 57140
rect 10196 57100 10205 57140
rect 11320 57100 12460 57140
rect 12500 57100 12509 57140
rect 6211 57056 6269 57057
rect 11320 57056 11360 57100
rect 13699 57056 13757 57057
rect 13900 57056 13940 57184
rect 14275 57100 14284 57140
rect 14324 57100 17836 57140
rect 17876 57100 18604 57140
rect 18644 57100 18653 57140
rect 21424 57056 21504 57076
rect 2947 57016 2956 57056
rect 2996 57016 3436 57056
rect 3476 57016 3485 57056
rect 3811 57016 3820 57056
rect 3860 57016 4396 57056
rect 4436 57016 4445 57056
rect 5443 57016 5452 57056
rect 5492 57016 5740 57056
rect 5780 57016 6220 57056
rect 6260 57016 6269 57056
rect 6691 57016 6700 57056
rect 6740 57016 6988 57056
rect 7028 57016 7037 57056
rect 7267 57016 7276 57056
rect 7316 57016 7564 57056
rect 7604 57016 7613 57056
rect 8227 57016 8236 57056
rect 8276 57016 8524 57056
rect 8564 57016 11360 57056
rect 11587 57016 11596 57056
rect 11636 57016 11645 57056
rect 13699 57016 13708 57056
rect 13748 57016 14860 57056
rect 14900 57016 14909 57056
rect 16867 57016 16876 57056
rect 16916 57016 17548 57056
rect 17588 57016 17597 57056
rect 19555 57016 19564 57056
rect 19604 57016 21504 57056
rect 6211 57015 6269 57016
rect 11596 56972 11636 57016
rect 13699 57015 13757 57016
rect 21424 56996 21504 57016
rect 4195 56932 4204 56972
rect 4244 56932 8908 56972
rect 8948 56932 9292 56972
rect 9332 56932 9341 56972
rect 11299 56932 11308 56972
rect 11348 56932 11636 56972
rect 13891 56932 13900 56972
rect 13940 56932 17260 56972
rect 17300 56932 17932 56972
rect 17972 56932 17981 56972
rect 0 56888 80 56908
rect 0 56848 748 56888
rect 788 56848 797 56888
rect 3235 56848 3244 56888
rect 3284 56848 3628 56888
rect 3668 56848 3677 56888
rect 6883 56848 6892 56888
rect 6932 56848 7508 56888
rect 17827 56848 17836 56888
rect 17876 56848 18028 56888
rect 18068 56848 18077 56888
rect 0 56828 80 56848
rect 7468 56804 7508 56848
rect 13411 56804 13469 56805
rect 7459 56764 7468 56804
rect 7508 56764 7517 56804
rect 11203 56764 11212 56804
rect 11252 56764 11596 56804
rect 11636 56764 11645 56804
rect 13315 56764 13324 56804
rect 13364 56764 13420 56804
rect 13460 56764 13469 56804
rect 13411 56763 13469 56764
rect 18691 56804 18749 56805
rect 18691 56764 18700 56804
rect 18740 56764 20908 56804
rect 20948 56764 20957 56804
rect 18691 56763 18749 56764
rect 4919 56680 4928 56720
rect 4968 56680 5010 56720
rect 5050 56680 5092 56720
rect 5132 56680 5174 56720
rect 5214 56680 5256 56720
rect 5296 56680 5305 56720
rect 7939 56680 7948 56720
rect 7988 56680 8428 56720
rect 8468 56680 8477 56720
rect 12259 56680 12268 56720
rect 12308 56680 13132 56720
rect 13172 56680 13804 56720
rect 13844 56680 13853 56720
rect 14659 56680 14668 56720
rect 14708 56680 17068 56720
rect 17108 56680 17117 56720
rect 20039 56680 20048 56720
rect 20088 56680 20130 56720
rect 20170 56680 20212 56720
rect 20252 56680 20294 56720
rect 20334 56680 20376 56720
rect 20416 56680 20425 56720
rect 11107 56596 11116 56636
rect 11156 56596 12076 56636
rect 12116 56596 14284 56636
rect 14324 56596 14572 56636
rect 14612 56596 14621 56636
rect 0 56552 80 56572
rect 9475 56552 9533 56553
rect 16867 56552 16925 56553
rect 0 56512 1612 56552
rect 1652 56512 1661 56552
rect 2851 56512 2860 56552
rect 2900 56512 3340 56552
rect 3380 56512 3389 56552
rect 3715 56512 3724 56552
rect 3764 56512 4684 56552
rect 4724 56512 4733 56552
rect 5731 56512 5740 56552
rect 5780 56512 9484 56552
rect 9524 56512 9533 56552
rect 16782 56512 16876 56552
rect 16916 56512 16925 56552
rect 0 56492 80 56512
rect 5740 56468 5780 56512
rect 9475 56511 9533 56512
rect 16867 56511 16925 56512
rect 16003 56468 16061 56469
rect 4387 56428 4396 56468
rect 4436 56428 5780 56468
rect 7171 56428 7180 56468
rect 7220 56428 9004 56468
rect 9044 56428 9053 56468
rect 15619 56428 15628 56468
rect 15668 56428 16012 56468
rect 16052 56428 19180 56468
rect 19220 56428 19229 56468
rect 16003 56427 16061 56428
rect 2755 56384 2813 56385
rect 17539 56384 17597 56385
rect 21424 56384 21504 56404
rect 2670 56344 2764 56384
rect 2804 56344 2813 56384
rect 7651 56344 7660 56384
rect 7700 56344 7948 56384
rect 7988 56344 7997 56384
rect 14467 56344 14476 56384
rect 14516 56344 16300 56384
rect 16340 56344 16349 56384
rect 16483 56344 16492 56384
rect 16532 56344 17548 56384
rect 17588 56344 17597 56384
rect 2755 56343 2813 56344
rect 17539 56343 17597 56344
rect 21388 56324 21504 56384
rect 3235 56300 3293 56301
rect 10819 56300 10877 56301
rect 3235 56260 3244 56300
rect 3284 56260 4300 56300
rect 4340 56260 5644 56300
rect 5684 56260 5693 56300
rect 9283 56260 9292 56300
rect 9332 56260 10100 56300
rect 3235 56259 3293 56260
rect 0 56216 80 56236
rect 10060 56217 10100 56260
rect 10819 56260 10828 56300
rect 10868 56260 11020 56300
rect 11060 56260 11980 56300
rect 12020 56260 12029 56300
rect 15043 56260 15052 56300
rect 15092 56260 15532 56300
rect 15572 56260 15581 56300
rect 15907 56260 15916 56300
rect 15956 56260 17356 56300
rect 17396 56260 17740 56300
rect 17780 56260 18028 56300
rect 18068 56260 18077 56300
rect 10819 56259 10877 56260
rect 10051 56216 10109 56217
rect 21388 56216 21428 56324
rect 0 56176 9484 56216
rect 9524 56176 9533 56216
rect 10051 56176 10060 56216
rect 10100 56176 15244 56216
rect 15284 56176 15293 56216
rect 18115 56176 18124 56216
rect 18164 56176 18604 56216
rect 18644 56176 18653 56216
rect 21388 56176 21484 56216
rect 0 56156 80 56176
rect 10051 56175 10109 56176
rect 21444 56132 21484 56176
rect 5731 56092 5740 56132
rect 5780 56092 6220 56132
rect 6260 56092 9196 56132
rect 9236 56092 9245 56132
rect 10531 56092 10540 56132
rect 10580 56092 21484 56132
rect 2659 56008 2668 56048
rect 2708 56008 2956 56048
rect 2996 56008 3005 56048
rect 9571 56008 9580 56048
rect 9620 56008 11884 56048
rect 11924 56008 11933 56048
rect 3679 55924 3688 55964
rect 3728 55924 3770 55964
rect 3810 55924 3852 55964
rect 3892 55924 3934 55964
rect 3974 55924 4016 55964
rect 4056 55924 4065 55964
rect 10339 55924 10348 55964
rect 10388 55924 10636 55964
rect 10676 55924 10685 55964
rect 14371 55924 14380 55964
rect 14420 55924 14668 55964
rect 14708 55924 14717 55964
rect 16579 55924 16588 55964
rect 16628 55924 16972 55964
rect 17012 55924 17021 55964
rect 18799 55924 18808 55964
rect 18848 55924 18890 55964
rect 18930 55924 18972 55964
rect 19012 55924 19054 55964
rect 19094 55924 19136 55964
rect 19176 55924 19185 55964
rect 0 55880 80 55900
rect 0 55840 14860 55880
rect 14900 55840 14909 55880
rect 0 55820 80 55840
rect 11299 55796 11357 55797
rect 2500 55756 6892 55796
rect 6932 55756 6941 55796
rect 11299 55756 11308 55796
rect 11348 55756 19372 55796
rect 19412 55756 19421 55796
rect 2500 55712 2540 55756
rect 11299 55755 11357 55756
rect 21424 55712 21504 55732
rect 2083 55672 2092 55712
rect 2132 55672 2540 55712
rect 4675 55672 4684 55712
rect 4724 55672 5260 55712
rect 5300 55672 5309 55712
rect 9667 55672 9676 55712
rect 9716 55672 9964 55712
rect 10004 55672 10013 55712
rect 11299 55672 11308 55712
rect 11348 55672 14380 55712
rect 14420 55672 14429 55712
rect 19555 55672 19564 55712
rect 19604 55672 21504 55712
rect 21424 55652 21504 55672
rect 3331 55628 3389 55629
rect 3331 55588 3340 55628
rect 3380 55588 3436 55628
rect 3476 55588 3485 55628
rect 6892 55588 11360 55628
rect 16291 55588 16300 55628
rect 16340 55588 16876 55628
rect 16916 55588 16925 55628
rect 3331 55587 3389 55588
rect 0 55544 80 55564
rect 6892 55544 6932 55588
rect 10147 55544 10205 55545
rect 11320 55544 11360 55588
rect 0 55504 6932 55544
rect 9859 55504 9868 55544
rect 9908 55504 10156 55544
rect 10196 55504 10205 55544
rect 10723 55504 10732 55544
rect 10772 55504 11020 55544
rect 11060 55504 11069 55544
rect 11320 55504 15820 55544
rect 15860 55504 15869 55544
rect 16963 55504 16972 55544
rect 17012 55504 18124 55544
rect 18164 55504 18173 55544
rect 0 55484 80 55504
rect 10147 55503 10205 55504
rect 2563 55420 2572 55460
rect 2612 55420 4684 55460
rect 4724 55420 4733 55460
rect 15972 55420 16012 55460
rect 16052 55420 16061 55460
rect 2755 55376 2813 55377
rect 16012 55376 16052 55420
rect 2755 55336 2764 55376
rect 2804 55336 3916 55376
rect 3956 55336 3965 55376
rect 13699 55336 13708 55376
rect 13748 55336 14092 55376
rect 14132 55336 14141 55376
rect 16012 55336 16780 55376
rect 16820 55336 16829 55376
rect 2755 55335 2813 55336
rect 2500 55252 9868 55292
rect 9908 55252 9917 55292
rect 11683 55252 11692 55292
rect 11732 55252 12364 55292
rect 12404 55252 17452 55292
rect 17492 55252 17501 55292
rect 0 55208 80 55228
rect 2500 55208 2540 55252
rect 0 55168 2540 55208
rect 4919 55168 4928 55208
rect 4968 55168 5010 55208
rect 5050 55168 5092 55208
rect 5132 55168 5174 55208
rect 5214 55168 5256 55208
rect 5296 55168 5305 55208
rect 6595 55168 6604 55208
rect 6644 55168 8524 55208
rect 8564 55168 8573 55208
rect 16387 55168 16396 55208
rect 16436 55168 16588 55208
rect 16628 55168 16637 55208
rect 20039 55168 20048 55208
rect 20088 55168 20130 55208
rect 20170 55168 20212 55208
rect 20252 55168 20294 55208
rect 20334 55168 20376 55208
rect 20416 55168 20425 55208
rect 0 55148 80 55168
rect 1987 55084 1996 55124
rect 2036 55084 2045 55124
rect 2851 55084 2860 55124
rect 2900 55084 3340 55124
rect 3380 55084 6220 55124
rect 6260 55084 7756 55124
rect 7796 55084 7805 55124
rect 9859 55084 9868 55124
rect 9908 55084 10156 55124
rect 10196 55084 10205 55124
rect 13699 55084 13708 55124
rect 13748 55084 15052 55124
rect 15092 55084 17644 55124
rect 17684 55084 17693 55124
rect 1996 55040 2036 55084
rect 16579 55040 16637 55041
rect 21424 55040 21504 55060
rect 1996 55000 5068 55040
rect 5108 55000 5117 55040
rect 16291 55000 16300 55040
rect 16340 55000 16588 55040
rect 16628 55000 16637 55040
rect 20227 55000 20236 55040
rect 20276 55000 21504 55040
rect 16579 54999 16637 55000
rect 21424 54980 21504 55000
rect 2947 54956 3005 54957
rect 10819 54956 10877 54957
rect 2947 54916 2956 54956
rect 2996 54916 3340 54956
rect 3380 54916 4396 54956
rect 4436 54916 4445 54956
rect 10734 54916 10828 54956
rect 10868 54916 10877 54956
rect 2947 54915 3005 54916
rect 10819 54915 10877 54916
rect 12556 54916 14380 54956
rect 14420 54916 14429 54956
rect 14755 54916 14764 54956
rect 14804 54916 17260 54956
rect 17300 54916 17932 54956
rect 17972 54916 17981 54956
rect 0 54872 80 54892
rect 4099 54872 4157 54873
rect 9187 54872 9245 54873
rect 12556 54872 12596 54916
rect 14275 54872 14333 54873
rect 0 54832 3052 54872
rect 3092 54832 3101 54872
rect 3811 54832 3820 54872
rect 3860 54832 4108 54872
rect 4148 54832 5356 54872
rect 5396 54832 5405 54872
rect 7555 54832 7564 54872
rect 7604 54832 7948 54872
rect 7988 54832 7997 54872
rect 9102 54832 9196 54872
rect 9236 54832 9245 54872
rect 10435 54832 10444 54872
rect 10484 54832 11308 54872
rect 11348 54832 11357 54872
rect 12547 54832 12556 54872
rect 12596 54832 12605 54872
rect 14083 54832 14092 54872
rect 14132 54832 14284 54872
rect 14324 54832 15532 54872
rect 15572 54832 15581 54872
rect 16675 54832 16684 54872
rect 16724 54832 17356 54872
rect 17396 54832 17405 54872
rect 0 54812 80 54832
rect 4099 54831 4157 54832
rect 9187 54831 9245 54832
rect 14275 54831 14333 54832
rect 3427 54788 3485 54789
rect 1987 54748 1996 54788
rect 2036 54748 2540 54788
rect 3342 54748 3436 54788
rect 3476 54748 3485 54788
rect 13507 54748 13516 54788
rect 13556 54748 15148 54788
rect 15188 54748 15197 54788
rect 16099 54748 16108 54788
rect 16148 54748 18316 54788
rect 18356 54748 18365 54788
rect 19843 54748 19852 54788
rect 19892 54748 20044 54788
rect 20084 54748 20093 54788
rect 2500 54704 2540 54748
rect 3427 54747 3485 54748
rect 2500 54664 3052 54704
rect 3092 54664 3101 54704
rect 11395 54664 11404 54704
rect 11444 54664 12076 54704
rect 12116 54664 12125 54704
rect 2500 54580 19276 54620
rect 19316 54580 19325 54620
rect 0 54536 80 54556
rect 2500 54536 2540 54580
rect 0 54496 2540 54536
rect 10819 54496 10828 54536
rect 10868 54496 15052 54536
rect 15092 54496 15101 54536
rect 17635 54496 17644 54536
rect 17684 54496 18508 54536
rect 18548 54496 19660 54536
rect 19700 54496 19709 54536
rect 0 54476 80 54496
rect 3679 54412 3688 54452
rect 3728 54412 3770 54452
rect 3810 54412 3852 54452
rect 3892 54412 3934 54452
rect 3974 54412 4016 54452
rect 4056 54412 4065 54452
rect 11299 54412 11308 54452
rect 11348 54412 15532 54452
rect 15572 54412 15581 54452
rect 18799 54412 18808 54452
rect 18848 54412 18890 54452
rect 18930 54412 18972 54452
rect 19012 54412 19054 54452
rect 19094 54412 19136 54452
rect 19176 54412 19185 54452
rect 21424 54368 21504 54388
rect 2947 54328 2956 54368
rect 2996 54328 4780 54368
rect 4820 54328 4829 54368
rect 11779 54328 11788 54368
rect 11828 54328 12268 54368
rect 12308 54328 12317 54368
rect 12931 54328 12940 54368
rect 12980 54328 13420 54368
rect 13460 54328 13469 54368
rect 19843 54328 19852 54368
rect 19892 54328 21504 54368
rect 21424 54308 21504 54328
rect 2500 54244 16588 54284
rect 16628 54244 16637 54284
rect 18307 54244 18316 54284
rect 18356 54244 19180 54284
rect 19220 54244 19229 54284
rect 0 54200 80 54220
rect 2500 54200 2540 54244
rect 0 54160 2540 54200
rect 2947 54160 2956 54200
rect 2996 54160 3724 54200
rect 3764 54160 3773 54200
rect 4387 54160 4396 54200
rect 4436 54160 6220 54200
rect 6260 54160 6269 54200
rect 6691 54160 6700 54200
rect 6740 54160 6749 54200
rect 8332 54160 9964 54200
rect 10004 54160 10013 54200
rect 10339 54160 10348 54200
rect 10388 54160 11212 54200
rect 11252 54160 11261 54200
rect 15043 54160 15052 54200
rect 15092 54160 16780 54200
rect 16820 54160 16829 54200
rect 0 54140 80 54160
rect 6700 54032 6740 54160
rect 8332 54116 8372 54160
rect 7555 54076 7564 54116
rect 7604 54076 8332 54116
rect 8372 54076 8381 54116
rect 11395 54076 11404 54116
rect 11444 54076 17164 54116
rect 17204 54076 17213 54116
rect 17443 54076 17452 54116
rect 17492 54076 19852 54116
rect 19892 54076 19901 54116
rect 10147 54032 10205 54033
rect 3811 53992 3820 54032
rect 3860 53992 4492 54032
rect 4532 53992 4541 54032
rect 6700 53992 7084 54032
rect 7124 53992 7948 54032
rect 7988 53992 9620 54032
rect 10032 53992 10060 54032
rect 10100 53992 10156 54032
rect 10196 53992 10348 54032
rect 10388 53992 10397 54032
rect 11971 53992 11980 54032
rect 12020 53992 12748 54032
rect 12788 53992 12797 54032
rect 13411 53992 13420 54032
rect 13460 53992 13804 54032
rect 13844 53992 13853 54032
rect 15811 53992 15820 54032
rect 15860 53992 19084 54032
rect 19124 53992 19133 54032
rect 2275 53948 2333 53949
rect 9580 53948 9620 53992
rect 10147 53991 10205 53992
rect 1315 53908 1324 53948
rect 1364 53908 2284 53948
rect 2324 53908 2333 53948
rect 3619 53908 3628 53948
rect 3668 53908 3916 53948
rect 3956 53908 3965 53948
rect 5923 53908 5932 53948
rect 5972 53908 6700 53948
rect 6740 53908 6749 53948
rect 9571 53908 9580 53948
rect 9620 53908 12556 53948
rect 12596 53908 12605 53948
rect 13123 53908 13132 53948
rect 13172 53908 13612 53948
rect 13652 53908 13661 53948
rect 2275 53907 2333 53908
rect 0 53864 80 53884
rect 0 53824 1708 53864
rect 1748 53824 1757 53864
rect 5539 53824 5548 53864
rect 5588 53824 7564 53864
rect 7604 53824 7613 53864
rect 10147 53824 10156 53864
rect 10196 53824 11360 53864
rect 13987 53824 13996 53864
rect 14036 53824 14764 53864
rect 14804 53824 14813 53864
rect 16675 53824 16684 53864
rect 16724 53824 16972 53864
rect 17012 53824 17021 53864
rect 20035 53824 20044 53864
rect 20084 53824 21428 53864
rect 0 53804 80 53824
rect 11320 53780 11360 53824
rect 547 53740 556 53780
rect 596 53740 2572 53780
rect 2612 53740 2621 53780
rect 11320 53740 21332 53780
rect 15907 53696 15965 53697
rect 4919 53656 4928 53696
rect 4968 53656 5010 53696
rect 5050 53656 5092 53696
rect 5132 53656 5174 53696
rect 5214 53656 5256 53696
rect 5296 53656 5305 53696
rect 11779 53656 11788 53696
rect 11828 53656 15916 53696
rect 15956 53656 15965 53696
rect 20039 53656 20048 53696
rect 20088 53656 20130 53696
rect 20170 53656 20212 53696
rect 20252 53656 20294 53696
rect 20334 53656 20376 53696
rect 20416 53656 20425 53696
rect 15907 53655 15965 53656
rect 6307 53612 6365 53613
rect 6307 53572 6316 53612
rect 6356 53572 19468 53612
rect 19508 53572 19517 53612
rect 6307 53571 6365 53572
rect 0 53528 80 53548
rect 21292 53528 21332 53740
rect 21388 53716 21428 53824
rect 21388 53656 21504 53716
rect 21424 53636 21504 53656
rect 0 53488 1804 53528
rect 1844 53488 1853 53528
rect 3619 53488 3628 53528
rect 3668 53488 8716 53528
rect 8756 53488 9292 53528
rect 9332 53488 9341 53528
rect 12163 53488 12172 53528
rect 12212 53488 12364 53528
rect 12404 53488 12413 53528
rect 13987 53488 13996 53528
rect 14036 53488 14380 53528
rect 14420 53488 14429 53528
rect 16867 53488 16876 53528
rect 16916 53488 17356 53528
rect 17396 53488 17405 53528
rect 21292 53488 21484 53528
rect 0 53468 80 53488
rect 8803 53444 8861 53445
rect 8803 53404 8812 53444
rect 8852 53404 14572 53444
rect 14612 53404 14621 53444
rect 17251 53404 17260 53444
rect 17300 53404 18740 53444
rect 8803 53403 8861 53404
rect 1507 53360 1565 53361
rect 11116 53360 11156 53404
rect 18700 53360 18740 53404
rect 1422 53320 1516 53360
rect 1556 53320 1565 53360
rect 3427 53320 3436 53360
rect 3476 53320 4204 53360
rect 4244 53320 4780 53360
rect 4820 53320 4829 53360
rect 9091 53320 9100 53360
rect 9140 53320 9772 53360
rect 9812 53320 9821 53360
rect 11107 53320 11116 53360
rect 11156 53320 11196 53360
rect 15715 53320 15724 53360
rect 15764 53320 16300 53360
rect 16340 53320 16349 53360
rect 18691 53320 18700 53360
rect 18740 53320 19756 53360
rect 19796 53320 19805 53360
rect 1507 53319 1565 53320
rect 21444 53276 21484 53488
rect 2755 53236 2764 53276
rect 2804 53236 5068 53276
rect 5108 53236 6412 53276
rect 6452 53236 9196 53276
rect 9236 53236 9964 53276
rect 10004 53236 10732 53276
rect 10772 53236 11596 53276
rect 11636 53236 13844 53276
rect 15619 53236 15628 53276
rect 15668 53236 18220 53276
rect 18260 53236 18269 53276
rect 21388 53236 21484 53276
rect 0 53192 80 53212
rect 0 53152 11980 53192
rect 12020 53152 12029 53192
rect 0 53132 80 53152
rect 13804 53108 13844 53236
rect 14275 53192 14333 53193
rect 21388 53192 21428 53236
rect 13987 53152 13996 53192
rect 14036 53152 14284 53192
rect 14324 53152 14333 53192
rect 14275 53151 14333 53152
rect 21292 53152 21428 53192
rect 2755 53068 2764 53108
rect 2804 53068 3724 53108
rect 3764 53068 3773 53108
rect 3907 53068 3916 53108
rect 3956 53068 4300 53108
rect 4340 53068 8620 53108
rect 8660 53068 8669 53108
rect 10339 53068 10348 53108
rect 10388 53068 10924 53108
rect 10964 53068 10973 53108
rect 13804 53068 15820 53108
rect 15860 53068 15869 53108
rect 16579 53068 16588 53108
rect 16628 53068 17068 53108
rect 17108 53068 17117 53108
rect 6307 53024 6365 53025
rect 21292 53024 21332 53152
rect 21424 53024 21504 53044
rect 4771 52984 4780 53024
rect 4820 52984 5836 53024
rect 5876 52984 6316 53024
rect 6356 52984 6365 53024
rect 12739 52984 12748 53024
rect 12788 52984 15148 53024
rect 15188 52984 15197 53024
rect 21292 52984 21504 53024
rect 6307 52983 6365 52984
rect 21424 52964 21504 52984
rect 3235 52940 3293 52941
rect 5635 52940 5693 52941
rect 739 52900 748 52940
rect 788 52900 2956 52940
rect 2996 52900 3005 52940
rect 3235 52900 3244 52940
rect 3284 52900 3436 52940
rect 3476 52900 3485 52940
rect 3679 52900 3688 52940
rect 3728 52900 3770 52940
rect 3810 52900 3852 52940
rect 3892 52900 3934 52940
rect 3974 52900 4016 52940
rect 4056 52900 4065 52940
rect 5539 52900 5548 52940
rect 5588 52900 5644 52940
rect 5684 52900 5693 52940
rect 7363 52900 7372 52940
rect 7412 52900 8044 52940
rect 8084 52900 8093 52940
rect 11971 52900 11980 52940
rect 12020 52900 13228 52940
rect 13268 52900 17452 52940
rect 17492 52900 17501 52940
rect 18799 52900 18808 52940
rect 18848 52900 18890 52940
rect 18930 52900 18972 52940
rect 19012 52900 19054 52940
rect 19094 52900 19136 52940
rect 19176 52900 19185 52940
rect 3235 52899 3293 52900
rect 5635 52899 5693 52900
rect 0 52856 80 52876
rect 17539 52856 17597 52857
rect 0 52816 17548 52856
rect 17588 52816 17597 52856
rect 0 52796 80 52816
rect 17539 52815 17597 52816
rect 18307 52856 18365 52857
rect 20611 52856 20669 52857
rect 18307 52816 18316 52856
rect 18356 52816 20620 52856
rect 20660 52816 20669 52856
rect 18307 52815 18365 52816
rect 20611 52815 20669 52816
rect 2563 52772 2621 52773
rect 1891 52732 1900 52772
rect 1940 52732 2572 52772
rect 2612 52732 2621 52772
rect 2563 52731 2621 52732
rect 3427 52772 3485 52773
rect 3427 52732 3436 52772
rect 3476 52732 3724 52772
rect 3764 52732 4396 52772
rect 4436 52732 4445 52772
rect 7267 52732 7276 52772
rect 7316 52732 19756 52772
rect 19796 52732 19805 52772
rect 3427 52731 3485 52732
rect 1315 52648 1324 52688
rect 1364 52648 2188 52688
rect 2228 52648 2237 52688
rect 12643 52648 12652 52688
rect 12692 52648 13036 52688
rect 13076 52648 13085 52688
rect 13795 52648 13804 52688
rect 13844 52648 13996 52688
rect 14036 52648 14045 52688
rect 1411 52564 1420 52604
rect 1460 52564 1940 52604
rect 1987 52564 1996 52604
rect 2036 52564 6796 52604
rect 6836 52564 6845 52604
rect 8131 52564 8140 52604
rect 8180 52564 8189 52604
rect 11395 52564 11404 52604
rect 11444 52564 12364 52604
rect 12404 52564 16204 52604
rect 16244 52564 16253 52604
rect 0 52520 80 52540
rect 0 52480 1844 52520
rect 0 52460 80 52480
rect 1804 52436 1844 52480
rect 1900 52436 1940 52564
rect 3331 52520 3389 52521
rect 3331 52480 3340 52520
rect 3380 52480 3628 52520
rect 3668 52480 3677 52520
rect 3811 52480 3820 52520
rect 3860 52480 5548 52520
rect 5588 52480 5597 52520
rect 6979 52480 6988 52520
rect 7028 52480 7660 52520
rect 7700 52480 7852 52520
rect 7892 52480 7901 52520
rect 3331 52479 3389 52480
rect 6403 52436 6461 52437
rect 1795 52396 1804 52436
rect 1844 52396 1853 52436
rect 1900 52396 2420 52436
rect 2380 52352 2420 52396
rect 6403 52396 6412 52436
rect 6452 52396 7372 52436
rect 7412 52396 7421 52436
rect 6403 52395 6461 52396
rect 1699 52312 1708 52352
rect 1748 52312 2092 52352
rect 2132 52312 2141 52352
rect 2371 52312 2380 52352
rect 2420 52312 2429 52352
rect 2563 52312 2572 52352
rect 2612 52312 2860 52352
rect 2900 52312 2909 52352
rect 8140 52268 8180 52564
rect 19747 52396 19756 52436
rect 19796 52396 20044 52436
rect 20084 52396 20093 52436
rect 21424 52352 21504 52372
rect 13219 52312 13228 52352
rect 13268 52312 13804 52352
rect 13844 52312 13853 52352
rect 15715 52312 15724 52352
rect 15764 52312 16012 52352
rect 16052 52312 16061 52352
rect 19651 52312 19660 52352
rect 19700 52312 21504 52352
rect 21424 52292 21504 52312
rect 7084 52228 7180 52268
rect 7220 52228 7229 52268
rect 7459 52228 7468 52268
rect 7508 52228 8524 52268
rect 8564 52228 8573 52268
rect 13123 52228 13132 52268
rect 13172 52228 13516 52268
rect 13556 52228 13708 52268
rect 13748 52228 13757 52268
rect 0 52184 80 52204
rect 0 52144 1420 52184
rect 1460 52144 1469 52184
rect 2083 52144 2092 52184
rect 2132 52144 2572 52184
rect 2612 52144 2621 52184
rect 4919 52144 4928 52184
rect 4968 52144 5010 52184
rect 5050 52144 5092 52184
rect 5132 52144 5174 52184
rect 5214 52144 5256 52184
rect 5296 52144 5305 52184
rect 0 52124 80 52144
rect 7084 52100 7124 52228
rect 13027 52144 13036 52184
rect 13076 52144 19276 52184
rect 19316 52144 19325 52184
rect 20039 52144 20048 52184
rect 20088 52144 20130 52184
rect 20170 52144 20212 52184
rect 20252 52144 20294 52184
rect 20334 52144 20376 52184
rect 20416 52144 20425 52184
rect 2659 52060 2668 52100
rect 2708 52060 4108 52100
rect 4148 52060 4157 52100
rect 7075 52060 7084 52100
rect 7124 52060 7133 52100
rect 12259 52060 12268 52100
rect 12308 52060 16780 52100
rect 16820 52060 16829 52100
rect 17251 52060 17260 52100
rect 17300 52060 17452 52100
rect 17492 52060 17501 52100
rect 19363 52060 19372 52100
rect 19412 52060 19660 52100
rect 19700 52060 19709 52100
rect 6403 51976 6412 52016
rect 6452 51976 7180 52016
rect 7220 51976 7229 52016
rect 16003 51976 16012 52016
rect 16052 51976 16204 52016
rect 16244 51976 16253 52016
rect 16963 51976 16972 52016
rect 17012 51976 17548 52016
rect 17588 51976 17597 52016
rect 19555 51976 19564 52016
rect 19604 51976 20044 52016
rect 20084 51976 20093 52016
rect 2563 51932 2621 51933
rect 1411 51892 1420 51932
rect 1460 51892 2572 51932
rect 2612 51892 7276 51932
rect 7316 51892 7325 51932
rect 11320 51892 12364 51932
rect 12404 51892 12413 51932
rect 13315 51892 13324 51932
rect 13364 51892 13612 51932
rect 13652 51892 13661 51932
rect 18307 51892 18316 51932
rect 18356 51892 18796 51932
rect 18836 51892 18845 51932
rect 2563 51891 2621 51892
rect 0 51848 80 51868
rect 11320 51848 11360 51892
rect 0 51808 11360 51848
rect 12643 51808 12652 51848
rect 12692 51808 13132 51848
rect 13172 51808 14188 51848
rect 14228 51808 14764 51848
rect 14804 51808 14813 51848
rect 15235 51808 15244 51848
rect 15284 51808 15820 51848
rect 15860 51808 17740 51848
rect 17780 51808 18412 51848
rect 18452 51808 18461 51848
rect 0 51788 80 51808
rect 2755 51764 2813 51765
rect 8131 51764 8189 51765
rect 15244 51764 15284 51808
rect 1891 51724 1900 51764
rect 1940 51724 2380 51764
rect 2420 51724 2429 51764
rect 2755 51724 2764 51764
rect 2804 51724 3628 51764
rect 3668 51724 3677 51764
rect 8035 51724 8044 51764
rect 8084 51724 8140 51764
rect 8180 51724 8189 51764
rect 9379 51724 9388 51764
rect 9428 51724 15284 51764
rect 15619 51724 15628 51764
rect 15668 51724 16204 51764
rect 16244 51724 18796 51764
rect 18836 51724 18845 51764
rect 2755 51723 2813 51724
rect 8131 51723 8189 51724
rect 6499 51680 6557 51681
rect 21424 51680 21504 51700
rect 2755 51640 2764 51680
rect 2804 51640 3148 51680
rect 3188 51640 3197 51680
rect 6499 51640 6508 51680
rect 6548 51640 8332 51680
rect 8372 51640 8381 51680
rect 8611 51640 8620 51680
rect 8660 51640 9292 51680
rect 9332 51640 9580 51680
rect 9620 51640 9629 51680
rect 10243 51640 10252 51680
rect 10292 51640 11212 51680
rect 11252 51640 11261 51680
rect 11320 51640 11500 51680
rect 11540 51640 11549 51680
rect 19939 51640 19948 51680
rect 19988 51640 21504 51680
rect 6499 51639 6557 51640
rect 11320 51596 11360 51640
rect 21424 51620 21504 51640
rect 6883 51556 6892 51596
rect 6932 51556 7372 51596
rect 7412 51556 7421 51596
rect 9859 51556 9868 51596
rect 9908 51556 11360 51596
rect 0 51512 80 51532
rect 6595 51512 6653 51513
rect 0 51472 6604 51512
rect 6644 51472 6653 51512
rect 0 51452 80 51472
rect 6595 51471 6653 51472
rect 3679 51388 3688 51428
rect 3728 51388 3770 51428
rect 3810 51388 3852 51428
rect 3892 51388 3934 51428
rect 3974 51388 4016 51428
rect 4056 51388 4065 51428
rect 4579 51388 4588 51428
rect 4628 51388 4972 51428
rect 5012 51388 5021 51428
rect 18799 51388 18808 51428
rect 18848 51388 18890 51428
rect 18930 51388 18972 51428
rect 19012 51388 19054 51428
rect 19094 51388 19136 51428
rect 19176 51388 19185 51428
rect 1219 51304 1228 51344
rect 1268 51304 9196 51344
rect 9236 51304 19948 51344
rect 19988 51304 19997 51344
rect 12643 51260 12701 51261
rect 13507 51260 13565 51261
rect 4291 51220 4300 51260
rect 4340 51220 4588 51260
rect 4628 51220 6124 51260
rect 6164 51220 6173 51260
rect 7747 51220 7756 51260
rect 7796 51220 8620 51260
rect 8660 51220 8669 51260
rect 11320 51220 12652 51260
rect 12692 51220 13516 51260
rect 13556 51220 13565 51260
rect 17251 51220 17260 51260
rect 17300 51220 17644 51260
rect 17684 51220 17693 51260
rect 0 51176 80 51196
rect 0 51136 2764 51176
rect 2804 51136 2813 51176
rect 0 51116 80 51136
rect 3043 51052 3052 51092
rect 3092 51052 9292 51092
rect 9332 51052 9341 51092
rect 3331 50968 3340 51008
rect 3380 50968 4012 51008
rect 4052 50968 4780 51008
rect 4820 50968 4829 51008
rect 5923 50968 5932 51008
rect 5972 50968 8140 51008
rect 8180 50968 8189 51008
rect 10051 50968 10060 51008
rect 10100 50968 10444 51008
rect 10484 50968 10493 51008
rect 1507 50924 1565 50925
rect 11320 50924 11360 51220
rect 12643 51219 12701 51220
rect 13507 51219 13565 51220
rect 11683 51052 11692 51092
rect 11732 51052 12172 51092
rect 12212 51052 12221 51092
rect 15139 51052 15148 51092
rect 15188 51052 15820 51092
rect 15860 51052 16204 51092
rect 16244 51052 16253 51092
rect 17059 51052 17068 51092
rect 17108 51052 19180 51092
rect 19220 51052 19229 51092
rect 21424 51008 21504 51028
rect 11491 50968 11500 51008
rect 11540 50968 11788 51008
rect 11828 50968 11837 51008
rect 12739 50968 12748 51008
rect 12788 50968 13324 51008
rect 13364 50968 13373 51008
rect 13987 50968 13996 51008
rect 14036 50968 14284 51008
rect 14324 50968 14333 51008
rect 15235 50968 15244 51008
rect 15284 50968 15916 51008
rect 15956 50968 16780 51008
rect 16820 50968 17452 51008
rect 17492 50968 17501 51008
rect 20131 50968 20140 51008
rect 20180 50968 21504 51008
rect 21424 50948 21504 50968
rect 1507 50884 1516 50924
rect 1556 50884 11360 50924
rect 1507 50883 1565 50884
rect 0 50840 80 50860
rect 0 50800 1516 50840
rect 1556 50800 1565 50840
rect 2659 50800 2668 50840
rect 2708 50800 4108 50840
rect 4148 50800 4157 50840
rect 4771 50800 4780 50840
rect 4820 50800 6412 50840
rect 6452 50800 6461 50840
rect 11011 50800 11020 50840
rect 11060 50800 14476 50840
rect 14516 50800 14956 50840
rect 14996 50800 15005 50840
rect 19171 50800 19180 50840
rect 19220 50800 19372 50840
rect 19412 50800 19421 50840
rect 19555 50800 19564 50840
rect 19604 50800 19613 50840
rect 0 50780 80 50800
rect 19564 50756 19604 50800
rect 2947 50716 2956 50756
rect 2996 50716 19604 50756
rect 4919 50632 4928 50672
rect 4968 50632 5010 50672
rect 5050 50632 5092 50672
rect 5132 50632 5174 50672
rect 5214 50632 5256 50672
rect 5296 50632 5305 50672
rect 6220 50632 7660 50672
rect 7700 50632 7709 50672
rect 16195 50632 16204 50672
rect 16244 50632 19948 50672
rect 19988 50632 19997 50672
rect 20039 50632 20048 50672
rect 20088 50632 20130 50672
rect 20170 50632 20212 50672
rect 20252 50632 20294 50672
rect 20334 50632 20376 50672
rect 20416 50632 20425 50672
rect 2563 50588 2621 50589
rect 6220 50588 6260 50632
rect 2083 50548 2092 50588
rect 2132 50548 2572 50588
rect 2612 50548 2621 50588
rect 5443 50548 5452 50588
rect 5492 50548 6220 50588
rect 6260 50548 6269 50588
rect 7267 50548 7276 50588
rect 7316 50548 7564 50588
rect 7604 50548 7613 50588
rect 10531 50548 10540 50588
rect 10580 50548 12268 50588
rect 12308 50548 12317 50588
rect 13996 50548 17932 50588
rect 17972 50548 17981 50588
rect 2563 50547 2621 50548
rect 0 50504 80 50524
rect 0 50464 13228 50504
rect 13268 50464 13277 50504
rect 0 50444 80 50464
rect 1507 50420 1565 50421
rect 1422 50380 1516 50420
rect 1556 50380 1565 50420
rect 1507 50379 1565 50380
rect 2563 50420 2621 50421
rect 13123 50420 13181 50421
rect 13996 50420 14036 50548
rect 18307 50504 18365 50505
rect 17251 50464 17260 50504
rect 17300 50464 17548 50504
rect 17588 50464 17597 50504
rect 18307 50464 18316 50504
rect 18356 50464 18604 50504
rect 18644 50464 18653 50504
rect 19267 50464 19276 50504
rect 19316 50464 19756 50504
rect 19796 50464 19805 50504
rect 18307 50463 18365 50464
rect 17923 50420 17981 50421
rect 2563 50380 2572 50420
rect 2612 50380 4684 50420
rect 4724 50380 4733 50420
rect 13123 50380 13132 50420
rect 13172 50380 13996 50420
rect 14036 50380 14045 50420
rect 15427 50380 15436 50420
rect 15476 50380 16684 50420
rect 16724 50380 16733 50420
rect 17059 50380 17068 50420
rect 17108 50380 17452 50420
rect 17492 50380 17501 50420
rect 17923 50380 17932 50420
rect 17972 50380 19852 50420
rect 19892 50380 19901 50420
rect 2563 50379 2621 50380
rect 13123 50379 13181 50380
rect 17923 50379 17981 50380
rect 21424 50336 21504 50356
rect 2659 50296 2668 50336
rect 2708 50296 4300 50336
rect 4340 50296 4349 50336
rect 6499 50296 6508 50336
rect 6548 50296 6796 50336
rect 6836 50296 7564 50336
rect 7604 50296 7613 50336
rect 10243 50296 10252 50336
rect 10292 50296 11596 50336
rect 11636 50296 11645 50336
rect 12835 50296 12844 50336
rect 12884 50296 14476 50336
rect 14516 50296 14525 50336
rect 15340 50296 19660 50336
rect 19700 50296 19709 50336
rect 20035 50296 20044 50336
rect 20084 50296 21504 50336
rect 5827 50212 5836 50252
rect 5876 50212 8716 50252
rect 8756 50212 8765 50252
rect 10435 50212 10444 50252
rect 10484 50212 10636 50252
rect 10676 50212 11404 50252
rect 11444 50212 11453 50252
rect 0 50168 80 50188
rect 15340 50168 15380 50296
rect 21424 50276 21504 50296
rect 16003 50212 16012 50252
rect 16052 50212 17068 50252
rect 17108 50212 17117 50252
rect 0 50128 15380 50168
rect 16963 50128 16972 50168
rect 17012 50128 17164 50168
rect 17204 50128 17213 50168
rect 17827 50128 17836 50168
rect 17876 50128 18220 50168
rect 18260 50128 19852 50168
rect 19892 50128 19901 50168
rect 0 50108 80 50128
rect 6595 50084 6653 50085
rect 2467 50044 2476 50084
rect 2516 50044 2860 50084
rect 2900 50044 2909 50084
rect 4003 50044 4012 50084
rect 4052 50044 4300 50084
rect 4340 50044 4349 50084
rect 4483 50044 4492 50084
rect 4532 50044 4876 50084
rect 4916 50044 4925 50084
rect 6595 50044 6604 50084
rect 6644 50044 15820 50084
rect 15860 50044 15869 50084
rect 16579 50044 16588 50084
rect 16628 50044 17548 50084
rect 17588 50044 19468 50084
rect 19508 50044 19517 50084
rect 6595 50043 6653 50044
rect 5635 50000 5693 50001
rect 3043 49960 3052 50000
rect 3092 49960 5644 50000
rect 5684 49960 6028 50000
rect 6068 49960 6077 50000
rect 7075 49960 7084 50000
rect 7124 49960 8812 50000
rect 8852 49960 8861 50000
rect 5635 49959 5693 49960
rect 1891 49876 1900 49916
rect 1940 49876 1949 49916
rect 3679 49876 3688 49916
rect 3728 49876 3770 49916
rect 3810 49876 3852 49916
rect 3892 49876 3934 49916
rect 3974 49876 4016 49916
rect 4056 49876 4065 49916
rect 18799 49876 18808 49916
rect 18848 49876 18890 49916
rect 18930 49876 18972 49916
rect 19012 49876 19054 49916
rect 19094 49876 19136 49916
rect 19176 49876 19185 49916
rect 0 49832 80 49852
rect 1900 49832 1940 49876
rect 0 49792 1940 49832
rect 12067 49792 12076 49832
rect 12116 49792 17932 49832
rect 17972 49792 17981 49832
rect 18115 49792 18124 49832
rect 18164 49792 18508 49832
rect 18548 49792 18557 49832
rect 0 49772 80 49792
rect 17539 49748 17597 49749
rect 12739 49708 12748 49748
rect 12788 49708 14764 49748
rect 14804 49708 16396 49748
rect 16436 49708 16445 49748
rect 16579 49708 16588 49748
rect 16628 49708 16876 49748
rect 16916 49708 16925 49748
rect 17539 49708 17548 49748
rect 17588 49708 18988 49748
rect 19028 49708 19037 49748
rect 17539 49707 17597 49708
rect 21424 49664 21504 49684
rect 11299 49624 11308 49664
rect 11348 49624 11596 49664
rect 11636 49624 11645 49664
rect 13507 49624 13516 49664
rect 13556 49624 13996 49664
rect 14036 49624 14045 49664
rect 14563 49624 14572 49664
rect 14612 49624 19372 49664
rect 19412 49624 19421 49664
rect 19651 49624 19660 49664
rect 19700 49624 21504 49664
rect 21424 49604 21504 49624
rect 13699 49580 13757 49581
rect 8707 49540 8716 49580
rect 8756 49540 10348 49580
rect 10388 49540 10397 49580
rect 12163 49540 12172 49580
rect 12212 49540 13708 49580
rect 13748 49540 15052 49580
rect 15092 49540 15101 49580
rect 15523 49540 15532 49580
rect 15572 49540 15916 49580
rect 15956 49540 18028 49580
rect 18068 49540 18077 49580
rect 13699 49539 13757 49540
rect 0 49496 80 49516
rect 0 49456 1516 49496
rect 1556 49456 1565 49496
rect 2947 49456 2956 49496
rect 2996 49456 5356 49496
rect 5396 49456 5405 49496
rect 5827 49456 5836 49496
rect 5876 49456 6700 49496
rect 6740 49456 6749 49496
rect 8611 49456 8620 49496
rect 8660 49456 8908 49496
rect 8948 49456 9868 49496
rect 9908 49456 9917 49496
rect 11107 49456 11116 49496
rect 11156 49456 11360 49496
rect 12931 49456 12940 49496
rect 12980 49456 13516 49496
rect 13556 49456 13565 49496
rect 15715 49456 15724 49496
rect 15764 49456 16396 49496
rect 16436 49456 16588 49496
rect 16628 49456 16637 49496
rect 18691 49456 18700 49496
rect 18740 49456 18749 49496
rect 0 49436 80 49456
rect 5356 49412 5396 49456
rect 11320 49412 11360 49456
rect 1699 49372 1708 49412
rect 1748 49372 2284 49412
rect 2324 49372 2333 49412
rect 3907 49372 3916 49412
rect 3956 49372 4204 49412
rect 4244 49372 4492 49412
rect 4532 49372 4541 49412
rect 5356 49372 8428 49412
rect 8468 49372 8477 49412
rect 11320 49372 12844 49412
rect 12884 49372 12893 49412
rect 13516 49328 13556 49456
rect 15139 49372 15148 49412
rect 15188 49372 15436 49412
rect 15476 49372 17644 49412
rect 17684 49372 18124 49412
rect 18164 49372 18173 49412
rect 18700 49328 18740 49456
rect 4579 49288 4588 49328
rect 4628 49288 6316 49328
rect 6356 49288 7084 49328
rect 7124 49288 7133 49328
rect 13516 49288 18740 49328
rect 556 49204 12844 49244
rect 12884 49204 12893 49244
rect 0 49160 80 49180
rect 556 49160 596 49204
rect 15628 49160 15668 49288
rect 0 49120 596 49160
rect 4919 49120 4928 49160
rect 4968 49120 5010 49160
rect 5050 49120 5092 49160
rect 5132 49120 5174 49160
rect 5214 49120 5256 49160
rect 5296 49120 5305 49160
rect 6787 49120 6796 49160
rect 6836 49120 7276 49160
rect 7316 49120 7325 49160
rect 13507 49120 13516 49160
rect 13556 49120 14572 49160
rect 14612 49120 14621 49160
rect 15427 49120 15436 49160
rect 15476 49120 15628 49160
rect 15668 49120 15677 49160
rect 15811 49120 15820 49160
rect 15860 49120 17356 49160
rect 17396 49120 17405 49160
rect 20039 49120 20048 49160
rect 20088 49120 20130 49160
rect 20170 49120 20212 49160
rect 20252 49120 20294 49160
rect 20334 49120 20376 49160
rect 20416 49120 20425 49160
rect 0 49100 80 49120
rect 3427 49036 3436 49076
rect 3476 49036 4396 49076
rect 4436 49036 4445 49076
rect 5347 49036 5356 49076
rect 5396 49036 5836 49076
rect 5876 49036 7372 49076
rect 7412 49036 7948 49076
rect 7988 49036 7997 49076
rect 21424 48992 21504 49012
rect 2500 48952 7756 48992
rect 7796 48952 7805 48992
rect 19171 48952 19180 48992
rect 19220 48952 19756 48992
rect 19796 48952 19805 48992
rect 19939 48952 19948 48992
rect 19988 48952 21504 48992
rect 2500 48908 2540 48952
rect 21424 48932 21504 48952
rect 2371 48868 2380 48908
rect 2420 48868 2540 48908
rect 4204 48868 16204 48908
rect 16244 48868 16253 48908
rect 18403 48868 18412 48908
rect 18452 48868 18461 48908
rect 0 48824 80 48844
rect 4204 48824 4244 48868
rect 6211 48824 6269 48825
rect 8899 48824 8957 48825
rect 9379 48824 9437 48825
rect 13123 48824 13181 48825
rect 0 48784 4244 48824
rect 5059 48784 5068 48824
rect 5108 48784 6220 48824
rect 6260 48784 6269 48824
rect 8814 48784 8908 48824
rect 8948 48784 9100 48824
rect 9140 48784 9149 48824
rect 9294 48784 9388 48824
rect 9428 48784 9437 48824
rect 11491 48784 11500 48824
rect 11540 48784 13132 48824
rect 13172 48784 13420 48824
rect 13460 48784 13469 48824
rect 13987 48784 13996 48824
rect 14036 48784 17644 48824
rect 17684 48784 18316 48824
rect 18356 48784 18365 48824
rect 0 48764 80 48784
rect 6211 48783 6269 48784
rect 8899 48783 8957 48784
rect 9379 48783 9437 48784
rect 13123 48783 13181 48784
rect 3043 48700 3052 48740
rect 3092 48700 5260 48740
rect 5300 48700 5309 48740
rect 13123 48700 13132 48740
rect 13172 48700 13804 48740
rect 13844 48700 13853 48740
rect 13699 48656 13757 48657
rect 1219 48616 1228 48656
rect 1268 48616 1996 48656
rect 2036 48616 11884 48656
rect 11924 48616 11933 48656
rect 13614 48616 13708 48656
rect 13748 48616 13757 48656
rect 18412 48656 18452 48868
rect 18412 48616 18604 48656
rect 18644 48616 18653 48656
rect 13699 48615 13757 48616
rect 2275 48532 2284 48572
rect 2324 48532 2668 48572
rect 2708 48532 2717 48572
rect 3148 48532 5932 48572
rect 5972 48532 5981 48572
rect 13219 48532 13228 48572
rect 13268 48532 13612 48572
rect 13652 48532 13661 48572
rect 14563 48532 14572 48572
rect 14612 48532 20716 48572
rect 20756 48532 20765 48572
rect 0 48488 80 48508
rect 0 48448 1516 48488
rect 1556 48448 1565 48488
rect 0 48428 80 48448
rect 3148 48320 3188 48532
rect 6211 48488 6269 48489
rect 5539 48448 5548 48488
rect 5588 48448 5597 48488
rect 5731 48448 5740 48488
rect 5780 48448 6220 48488
rect 6260 48448 19948 48488
rect 19988 48448 19997 48488
rect 5548 48404 5588 48448
rect 6211 48447 6269 48448
rect 6115 48404 6173 48405
rect 3679 48364 3688 48404
rect 3728 48364 3770 48404
rect 3810 48364 3852 48404
rect 3892 48364 3934 48404
rect 3974 48364 4016 48404
rect 4056 48364 4065 48404
rect 5548 48364 6124 48404
rect 6164 48364 6173 48404
rect 18799 48364 18808 48404
rect 18848 48364 18890 48404
rect 18930 48364 18972 48404
rect 19012 48364 19054 48404
rect 19094 48364 19136 48404
rect 19176 48364 19185 48404
rect 6115 48363 6173 48364
rect 21424 48320 21504 48340
rect 3139 48280 3148 48320
rect 3188 48280 3197 48320
rect 4867 48280 4876 48320
rect 4916 48280 5356 48320
rect 5396 48280 5405 48320
rect 5539 48280 5548 48320
rect 5588 48280 8140 48320
rect 8180 48280 8189 48320
rect 19843 48280 19852 48320
rect 19892 48280 21504 48320
rect 21424 48260 21504 48280
rect 2851 48196 2860 48236
rect 2900 48196 5932 48236
rect 5972 48196 6124 48236
rect 6164 48196 6173 48236
rect 6307 48196 6316 48236
rect 6356 48196 6508 48236
rect 6548 48196 9004 48236
rect 9044 48196 15820 48236
rect 15860 48196 15869 48236
rect 0 48152 80 48172
rect 0 48112 1708 48152
rect 1748 48112 1757 48152
rect 2467 48112 2476 48152
rect 2516 48112 3244 48152
rect 3284 48112 3293 48152
rect 3619 48112 3628 48152
rect 3668 48112 5068 48152
rect 5108 48112 5117 48152
rect 5347 48112 5356 48152
rect 5396 48112 6932 48152
rect 8131 48112 8140 48152
rect 8180 48112 8908 48152
rect 8948 48112 8957 48152
rect 0 48092 80 48112
rect 6892 48068 6932 48112
rect 1795 48028 1804 48068
rect 1844 48028 6700 48068
rect 6740 48028 6749 48068
rect 6883 48028 6892 48068
rect 6932 48028 9388 48068
rect 9428 48028 9868 48068
rect 9908 48028 9917 48068
rect 11320 48028 19852 48068
rect 19892 48028 19901 48068
rect 5923 47984 5981 47985
rect 1411 47944 1420 47984
rect 1460 47944 1996 47984
rect 2036 47944 2045 47984
rect 2563 47944 2572 47984
rect 2612 47944 3628 47984
rect 3668 47944 3677 47984
rect 5443 47944 5452 47984
rect 5492 47944 5932 47984
rect 5972 47944 5981 47984
rect 5923 47943 5981 47944
rect 6115 47984 6173 47985
rect 6115 47944 6124 47984
rect 6164 47944 7124 47984
rect 8227 47944 8236 47984
rect 8276 47944 9484 47984
rect 9524 47944 9533 47984
rect 6115 47943 6173 47944
rect 2755 47900 2813 47901
rect 7084 47900 7124 47944
rect 11320 47900 11360 48028
rect 14467 47944 14476 47984
rect 14516 47944 14860 47984
rect 14900 47944 14909 47984
rect 16867 47944 16876 47984
rect 16916 47944 17836 47984
rect 17876 47944 19468 47984
rect 19508 47944 19517 47984
rect 2670 47860 2764 47900
rect 2804 47860 2813 47900
rect 5059 47860 5068 47900
rect 5108 47860 6988 47900
rect 7028 47860 7037 47900
rect 7084 47860 11360 47900
rect 13411 47860 13420 47900
rect 13460 47860 18356 47900
rect 2755 47859 2813 47860
rect 0 47816 80 47836
rect 18316 47816 18356 47860
rect 0 47776 2540 47816
rect 3427 47776 3436 47816
rect 3476 47776 3820 47816
rect 3860 47776 3869 47816
rect 8995 47776 9004 47816
rect 9044 47776 9292 47816
rect 9332 47776 9341 47816
rect 14179 47776 14188 47816
rect 14228 47776 14476 47816
rect 14516 47776 14525 47816
rect 17731 47776 17740 47816
rect 17780 47776 18028 47816
rect 18068 47776 18077 47816
rect 18307 47776 18316 47816
rect 18356 47776 18365 47816
rect 20131 47776 20140 47816
rect 20180 47776 21332 47816
rect 0 47756 80 47776
rect 2500 47732 2540 47776
rect 2500 47692 10636 47732
rect 10676 47692 10685 47732
rect 6115 47648 6173 47649
rect 21292 47648 21332 47776
rect 21424 47648 21504 47668
rect 4919 47608 4928 47648
rect 4968 47608 5010 47648
rect 5050 47608 5092 47648
rect 5132 47608 5174 47648
rect 5214 47608 5256 47648
rect 5296 47608 5305 47648
rect 5635 47608 5644 47648
rect 5684 47608 6124 47648
rect 6164 47608 6173 47648
rect 20039 47608 20048 47648
rect 20088 47608 20130 47648
rect 20170 47608 20212 47648
rect 20252 47608 20294 47648
rect 20334 47608 20376 47648
rect 20416 47608 20425 47648
rect 21292 47608 21504 47648
rect 6115 47607 6173 47608
rect 21424 47588 21504 47608
rect 19267 47524 19276 47564
rect 19316 47524 19468 47564
rect 19508 47524 19517 47564
rect 0 47480 80 47500
rect 0 47440 15284 47480
rect 16387 47440 16396 47480
rect 16436 47440 16780 47480
rect 16820 47440 16829 47480
rect 0 47420 80 47440
rect 4099 47396 4157 47397
rect 13027 47396 13085 47397
rect 2380 47356 4108 47396
rect 4148 47356 13036 47396
rect 13076 47356 13085 47396
rect 15244 47396 15284 47440
rect 15244 47356 19276 47396
rect 19316 47356 19325 47396
rect 2380 47312 2420 47356
rect 4099 47355 4157 47356
rect 13027 47355 13085 47356
rect 2371 47272 2380 47312
rect 2420 47272 2429 47312
rect 3043 47272 3052 47312
rect 3092 47272 3340 47312
rect 3380 47272 3389 47312
rect 5443 47272 5452 47312
rect 5492 47272 6412 47312
rect 6452 47272 6461 47312
rect 12739 47272 12748 47312
rect 12788 47272 13516 47312
rect 13556 47272 13565 47312
rect 16963 47272 16972 47312
rect 17012 47272 17260 47312
rect 17300 47272 17309 47312
rect 17059 47228 17117 47229
rect 1987 47188 1996 47228
rect 2036 47188 4012 47228
rect 4052 47188 4061 47228
rect 11491 47188 11500 47228
rect 11540 47188 12364 47228
rect 12404 47188 13996 47228
rect 14036 47188 17068 47228
rect 17108 47188 18220 47228
rect 18260 47188 19852 47228
rect 19892 47188 19901 47228
rect 17059 47187 17117 47188
rect 0 47144 80 47164
rect 0 47104 1900 47144
rect 1940 47104 1949 47144
rect 0 47084 80 47104
rect 11779 47020 11788 47060
rect 11828 47020 12364 47060
rect 12404 47020 12413 47060
rect 17923 47020 17932 47060
rect 17972 47020 18412 47060
rect 18452 47020 18461 47060
rect 21424 46976 21504 46996
rect 19939 46936 19948 46976
rect 19988 46936 21504 46976
rect 21424 46916 21504 46936
rect 13507 46892 13565 46893
rect 3679 46852 3688 46892
rect 3728 46852 3770 46892
rect 3810 46852 3852 46892
rect 3892 46852 3934 46892
rect 3974 46852 4016 46892
rect 4056 46852 4065 46892
rect 13507 46852 13516 46892
rect 13556 46852 16148 46892
rect 18307 46852 18316 46892
rect 18356 46852 18700 46892
rect 18740 46852 18749 46892
rect 18799 46852 18808 46892
rect 18848 46852 18890 46892
rect 18930 46852 18972 46892
rect 19012 46852 19054 46892
rect 19094 46852 19136 46892
rect 19176 46852 19185 46892
rect 13507 46851 13565 46852
rect 0 46808 80 46828
rect 16108 46808 16148 46852
rect 0 46768 1516 46808
rect 1556 46768 1565 46808
rect 11107 46768 11116 46808
rect 11156 46768 15244 46808
rect 15284 46768 16012 46808
rect 16052 46768 16061 46808
rect 16108 46768 19892 46808
rect 0 46748 80 46768
rect 18307 46724 18365 46725
rect 9964 46684 11404 46724
rect 11444 46684 11453 46724
rect 12355 46684 12364 46724
rect 12404 46684 18316 46724
rect 18356 46684 18365 46724
rect 18979 46684 18988 46724
rect 19028 46684 19468 46724
rect 19508 46684 19517 46724
rect 5923 46640 5981 46641
rect 5838 46600 5932 46640
rect 5972 46600 5981 46640
rect 7075 46600 7084 46640
rect 7124 46600 7133 46640
rect 5923 46599 5981 46600
rect 7084 46556 7124 46600
rect 7084 46516 7468 46556
rect 7508 46516 7517 46556
rect 0 46472 80 46492
rect 9964 46472 10004 46684
rect 18307 46683 18365 46684
rect 19852 46556 19892 46768
rect 10339 46516 10348 46556
rect 10388 46516 10732 46556
rect 10772 46516 10781 46556
rect 12259 46516 12268 46556
rect 12308 46516 13612 46556
rect 13652 46516 13661 46556
rect 19843 46516 19852 46556
rect 19892 46516 19901 46556
rect 13027 46472 13085 46473
rect 0 46432 2540 46472
rect 8131 46432 8140 46472
rect 8180 46432 8620 46472
rect 8660 46432 8669 46472
rect 9475 46432 9484 46472
rect 9524 46432 9964 46472
rect 10004 46432 10013 46472
rect 10531 46432 10540 46472
rect 10580 46432 10924 46472
rect 10964 46432 10973 46472
rect 12942 46432 13036 46472
rect 13076 46432 13085 46472
rect 0 46412 80 46432
rect 2500 46388 2540 46432
rect 13027 46431 13085 46432
rect 18307 46472 18365 46473
rect 18307 46432 18316 46472
rect 18356 46432 18508 46472
rect 18548 46432 18557 46472
rect 18307 46431 18365 46432
rect 2500 46348 13708 46388
rect 13748 46348 13757 46388
rect 2275 46304 2333 46305
rect 21424 46304 21504 46324
rect 1219 46264 1228 46304
rect 1268 46264 2284 46304
rect 2324 46264 2333 46304
rect 2659 46264 2668 46304
rect 2708 46264 4012 46304
rect 4052 46264 4061 46304
rect 7075 46264 7084 46304
rect 7124 46264 7564 46304
rect 7604 46264 7613 46304
rect 9571 46264 9580 46304
rect 9620 46264 9868 46304
rect 9908 46264 9917 46304
rect 10051 46264 10060 46304
rect 10100 46264 10109 46304
rect 12643 46264 12652 46304
rect 12692 46264 13324 46304
rect 13364 46264 13373 46304
rect 14659 46264 14668 46304
rect 14708 46264 14860 46304
rect 14900 46264 14909 46304
rect 20035 46264 20044 46304
rect 20084 46264 21504 46304
rect 2275 46263 2333 46264
rect 10060 46220 10100 46264
rect 21424 46244 21504 46264
rect 7363 46180 7372 46220
rect 7412 46180 8908 46220
rect 8948 46180 9388 46220
rect 9428 46180 9437 46220
rect 9667 46180 9676 46220
rect 9716 46180 10100 46220
rect 10915 46180 10924 46220
rect 10964 46180 16108 46220
rect 16148 46180 16157 46220
rect 0 46136 80 46156
rect 0 46096 2540 46136
rect 4919 46096 4928 46136
rect 4968 46096 5010 46136
rect 5050 46096 5092 46136
rect 5132 46096 5174 46136
rect 5214 46096 5256 46136
rect 5296 46096 5305 46136
rect 10051 46096 10060 46136
rect 10100 46096 10444 46136
rect 10484 46096 15724 46136
rect 15764 46096 15773 46136
rect 20039 46096 20048 46136
rect 20088 46096 20130 46136
rect 20170 46096 20212 46136
rect 20252 46096 20294 46136
rect 20334 46096 20376 46136
rect 20416 46096 20425 46136
rect 0 46076 80 46096
rect 2500 46052 2540 46096
rect 2500 46012 8812 46052
rect 8852 46012 8861 46052
rect 12067 46012 12076 46052
rect 12116 46012 21484 46052
rect 6307 45928 6316 45968
rect 6356 45928 6700 45968
rect 6740 45928 9196 45968
rect 9236 45928 18892 45968
rect 18932 45928 18941 45968
rect 4099 45844 4108 45884
rect 4148 45844 7276 45884
rect 7316 45844 7325 45884
rect 9667 45844 9676 45884
rect 9716 45844 19564 45884
rect 19604 45844 19613 45884
rect 0 45800 80 45820
rect 21444 45800 21484 46012
rect 0 45760 1228 45800
rect 1268 45760 1277 45800
rect 2275 45760 2284 45800
rect 2324 45760 2476 45800
rect 2516 45760 2668 45800
rect 2708 45760 5356 45800
rect 5396 45760 7564 45800
rect 7604 45760 7613 45800
rect 15235 45760 15244 45800
rect 15284 45760 16780 45800
rect 16820 45760 16829 45800
rect 18883 45760 18892 45800
rect 18932 45760 19276 45800
rect 19316 45760 19325 45800
rect 21388 45760 21484 45800
rect 0 45740 80 45760
rect 10051 45716 10109 45717
rect 1699 45676 1708 45716
rect 1748 45676 2380 45716
rect 2420 45676 2429 45716
rect 9955 45676 9964 45716
rect 10004 45676 10060 45716
rect 10100 45676 10348 45716
rect 10388 45676 10397 45716
rect 18211 45676 18220 45716
rect 18260 45676 18700 45716
rect 18740 45676 18749 45716
rect 18979 45676 18988 45716
rect 19028 45676 19660 45716
rect 19700 45676 19709 45716
rect 10051 45675 10109 45676
rect 21388 45652 21428 45760
rect 3331 45632 3389 45633
rect 3331 45592 3340 45632
rect 3380 45592 3916 45632
rect 3956 45592 16012 45632
rect 16052 45592 16061 45632
rect 21388 45592 21504 45652
rect 3331 45591 3389 45592
rect 21424 45572 21504 45592
rect 16387 45548 16445 45549
rect 7171 45508 7180 45548
rect 7220 45508 7756 45548
rect 7796 45508 7805 45548
rect 16387 45508 16396 45548
rect 16436 45508 18796 45548
rect 18836 45508 18845 45548
rect 19075 45508 19084 45548
rect 19124 45508 19133 45548
rect 19363 45508 19372 45548
rect 19412 45508 19660 45548
rect 19700 45508 19709 45548
rect 16387 45507 16445 45508
rect 0 45464 80 45484
rect 19084 45464 19124 45508
rect 0 45424 1516 45464
rect 1556 45424 1565 45464
rect 6211 45424 6220 45464
rect 6260 45424 6269 45464
rect 19084 45424 19316 45464
rect 0 45404 80 45424
rect 2275 45380 2333 45381
rect 6220 45380 6260 45424
rect 2275 45340 2284 45380
rect 2324 45340 3572 45380
rect 3679 45340 3688 45380
rect 3728 45340 3770 45380
rect 3810 45340 3852 45380
rect 3892 45340 3934 45380
rect 3974 45340 4016 45380
rect 4056 45340 4065 45380
rect 5635 45340 5644 45380
rect 5684 45340 6260 45380
rect 6979 45340 6988 45380
rect 7028 45340 7276 45380
rect 7316 45340 7325 45380
rect 11875 45340 11884 45380
rect 11924 45340 12268 45380
rect 12308 45340 12317 45380
rect 13315 45340 13324 45380
rect 13364 45340 15532 45380
rect 15572 45340 15581 45380
rect 17059 45340 17068 45380
rect 17108 45340 17836 45380
rect 17876 45340 17885 45380
rect 18799 45340 18808 45380
rect 18848 45340 18890 45380
rect 18930 45340 18972 45380
rect 19012 45340 19054 45380
rect 19094 45340 19136 45380
rect 19176 45340 19185 45380
rect 2275 45339 2333 45340
rect 3532 45296 3572 45340
rect 2083 45256 2092 45296
rect 2132 45256 2540 45296
rect 3532 45256 18932 45296
rect 2500 45212 2540 45256
rect 18892 45212 18932 45256
rect 2500 45172 7372 45212
rect 7412 45172 7421 45212
rect 8803 45172 8812 45212
rect 8852 45172 16876 45212
rect 16916 45172 16925 45212
rect 17923 45172 17932 45212
rect 17972 45172 18508 45212
rect 18548 45172 18557 45212
rect 18883 45172 18892 45212
rect 18932 45172 18941 45212
rect 0 45128 80 45148
rect 19276 45128 19316 45424
rect 0 45088 11404 45128
rect 11444 45088 11453 45128
rect 12067 45088 12076 45128
rect 12116 45088 14188 45128
rect 14228 45088 18124 45128
rect 18164 45088 18173 45128
rect 18979 45088 18988 45128
rect 19028 45088 19316 45128
rect 0 45068 80 45088
rect 2083 45004 2092 45044
rect 2132 45004 7276 45044
rect 7316 45004 7325 45044
rect 7939 45004 7948 45044
rect 7988 45004 9004 45044
rect 9044 45004 19852 45044
rect 19892 45004 19901 45044
rect 2851 44960 2909 44961
rect 21424 44960 21504 44980
rect 2851 44920 2860 44960
rect 2900 44920 3628 44960
rect 3668 44920 3677 44960
rect 4003 44920 4012 44960
rect 4052 44920 4588 44960
rect 4628 44920 4637 44960
rect 7555 44920 7564 44960
rect 7604 44920 9196 44960
rect 9236 44920 10828 44960
rect 10868 44920 11212 44960
rect 11252 44920 13324 44960
rect 13364 44920 13804 44960
rect 13844 44920 14668 44960
rect 14708 44920 14717 44960
rect 15235 44920 15244 44960
rect 15284 44920 15436 44960
rect 15476 44920 15485 44960
rect 17731 44920 17740 44960
rect 17780 44920 18988 44960
rect 19028 44920 19037 44960
rect 19747 44920 19756 44960
rect 19796 44920 21504 44960
rect 2851 44919 2909 44920
rect 14668 44876 14708 44920
rect 21424 44900 21504 44920
rect 3523 44836 3532 44876
rect 3572 44836 5932 44876
rect 5972 44836 6220 44876
rect 6260 44836 6269 44876
rect 14668 44836 16492 44876
rect 16532 44836 18316 44876
rect 18356 44836 18365 44876
rect 0 44792 80 44812
rect 0 44752 2540 44792
rect 3043 44752 3052 44792
rect 3092 44752 6700 44792
rect 6740 44752 6749 44792
rect 18883 44752 18892 44792
rect 18932 44752 19852 44792
rect 19892 44752 19901 44792
rect 0 44732 80 44752
rect 2500 44540 2540 44752
rect 3811 44668 3820 44708
rect 3860 44668 4300 44708
rect 4340 44668 4349 44708
rect 13516 44668 13900 44708
rect 13940 44668 13949 44708
rect 13516 44624 13556 44668
rect 4919 44584 4928 44624
rect 4968 44584 5010 44624
rect 5050 44584 5092 44624
rect 5132 44584 5174 44624
rect 5214 44584 5256 44624
rect 5296 44584 5305 44624
rect 13507 44584 13516 44624
rect 13556 44584 13565 44624
rect 13699 44584 13708 44624
rect 13748 44584 16108 44624
rect 16148 44584 17548 44624
rect 17588 44584 17597 44624
rect 20039 44584 20048 44624
rect 20088 44584 20130 44624
rect 20170 44584 20212 44624
rect 20252 44584 20294 44624
rect 20334 44584 20376 44624
rect 20416 44584 20425 44624
rect 16387 44540 16445 44541
rect 2500 44500 16396 44540
rect 16436 44500 16445 44540
rect 17635 44500 17644 44540
rect 17684 44500 18124 44540
rect 18164 44500 19756 44540
rect 19796 44500 19805 44540
rect 16387 44499 16445 44500
rect 0 44456 80 44476
rect 0 44416 1900 44456
rect 1940 44416 1949 44456
rect 3532 44416 9676 44456
rect 9716 44416 9725 44456
rect 11299 44416 11308 44456
rect 11348 44416 12460 44456
rect 12500 44416 12509 44456
rect 15427 44416 15436 44456
rect 15476 44416 15724 44456
rect 15764 44416 15773 44456
rect 0 44396 80 44416
rect 1987 44164 1996 44204
rect 2036 44164 2476 44204
rect 2516 44164 2525 44204
rect 0 44120 80 44140
rect 3532 44120 3572 44416
rect 16195 44372 16253 44373
rect 5635 44332 5644 44372
rect 5684 44332 16204 44372
rect 16244 44332 16253 44372
rect 16195 44331 16253 44332
rect 6211 44288 6269 44289
rect 17059 44288 17117 44289
rect 21424 44288 21504 44308
rect 3619 44248 3628 44288
rect 3668 44248 6220 44288
rect 6260 44248 6269 44288
rect 10051 44248 10060 44288
rect 10100 44248 13708 44288
rect 13748 44248 13757 44288
rect 13987 44248 13996 44288
rect 14036 44248 14188 44288
rect 14228 44248 14237 44288
rect 15235 44248 15244 44288
rect 15284 44248 17068 44288
rect 17108 44248 17117 44288
rect 18307 44248 18316 44288
rect 18356 44248 19372 44288
rect 19412 44248 19421 44288
rect 19939 44248 19948 44288
rect 19988 44248 21504 44288
rect 6211 44247 6269 44248
rect 17059 44247 17117 44248
rect 21424 44228 21504 44248
rect 5059 44164 5068 44204
rect 5108 44164 7468 44204
rect 7508 44164 7517 44204
rect 9859 44164 9868 44204
rect 9908 44164 10636 44204
rect 10676 44164 10685 44204
rect 15811 44164 15820 44204
rect 15860 44164 17164 44204
rect 17204 44164 18220 44204
rect 18260 44164 18269 44204
rect 6211 44120 6269 44121
rect 0 44080 3572 44120
rect 5251 44080 5260 44120
rect 5300 44080 5548 44120
rect 5588 44080 5597 44120
rect 6211 44080 6220 44120
rect 6260 44080 6269 44120
rect 12835 44080 12844 44120
rect 12884 44080 17740 44120
rect 17780 44080 17789 44120
rect 0 44060 80 44080
rect 6211 44079 6269 44080
rect 6220 44036 6260 44079
rect 9379 44036 9437 44037
rect 2179 43996 2188 44036
rect 2228 43996 2668 44036
rect 2708 43996 2717 44036
rect 4003 43996 4012 44036
rect 4052 43996 4061 44036
rect 6211 43996 6220 44036
rect 6260 43996 6271 44036
rect 9379 43996 9388 44036
rect 9428 43996 9484 44036
rect 9524 43996 9533 44036
rect 4012 43952 4052 43996
rect 9379 43995 9437 43996
rect 8899 43952 8957 43953
rect 4012 43912 8908 43952
rect 8948 43912 8957 43952
rect 9283 43912 9292 43952
rect 9332 43912 9868 43952
rect 9908 43912 9917 43952
rect 8899 43911 8957 43912
rect 3679 43828 3688 43868
rect 3728 43828 3770 43868
rect 3810 43828 3852 43868
rect 3892 43828 3934 43868
rect 3974 43828 4016 43868
rect 4056 43828 4065 43868
rect 9763 43828 9772 43868
rect 9812 43828 15052 43868
rect 15092 43828 15101 43868
rect 18799 43828 18808 43868
rect 18848 43828 18890 43868
rect 18930 43828 18972 43868
rect 19012 43828 19054 43868
rect 19094 43828 19136 43868
rect 19176 43828 19185 43868
rect 0 43784 80 43804
rect 0 43744 17452 43784
rect 17492 43744 17501 43784
rect 0 43724 80 43744
rect 21187 43700 21245 43701
rect 19171 43660 19180 43700
rect 19220 43660 21196 43700
rect 21236 43660 21245 43700
rect 21187 43659 21245 43660
rect 21424 43616 21504 43636
rect 3139 43576 3148 43616
rect 3188 43576 3724 43616
rect 3764 43576 3773 43616
rect 13315 43576 13324 43616
rect 13364 43576 13804 43616
rect 13844 43576 13853 43616
rect 19939 43576 19948 43616
rect 19988 43576 21504 43616
rect 21424 43556 21504 43576
rect 2851 43492 2860 43532
rect 2900 43492 3436 43532
rect 3476 43492 3628 43532
rect 3668 43492 3677 43532
rect 4099 43492 4108 43532
rect 4148 43492 4780 43532
rect 4820 43492 4829 43532
rect 7459 43492 7468 43532
rect 7508 43492 8812 43532
rect 8852 43492 9388 43532
rect 9428 43492 9437 43532
rect 17731 43492 17740 43532
rect 17780 43492 18988 43532
rect 19028 43492 19037 43532
rect 0 43448 80 43468
rect 0 43408 13900 43448
rect 13940 43408 13949 43448
rect 15811 43408 15820 43448
rect 15860 43408 16108 43448
rect 16148 43408 16157 43448
rect 0 43388 80 43408
rect 9379 43364 9437 43365
rect 12163 43364 12221 43365
rect 8419 43324 8428 43364
rect 8468 43324 9388 43364
rect 9428 43324 9437 43364
rect 12078 43324 12172 43364
rect 12212 43324 12221 43364
rect 9379 43323 9437 43324
rect 12163 43323 12221 43324
rect 8899 43280 8957 43281
rect 9859 43280 9917 43281
rect 8899 43240 8908 43280
rect 8948 43240 9004 43280
rect 9044 43240 9053 43280
rect 9859 43240 9868 43280
rect 9908 43240 19948 43280
rect 19988 43240 19997 43280
rect 8899 43239 8957 43240
rect 9859 43239 9917 43240
rect 2500 43156 8908 43196
rect 8948 43156 8957 43196
rect 15523 43156 15532 43196
rect 15572 43156 15820 43196
rect 15860 43156 15869 43196
rect 0 43112 80 43132
rect 2500 43112 2540 43156
rect 0 43072 2540 43112
rect 4919 43072 4928 43112
rect 4968 43072 5010 43112
rect 5050 43072 5092 43112
rect 5132 43072 5174 43112
rect 5214 43072 5256 43112
rect 5296 43072 5305 43112
rect 20039 43072 20048 43112
rect 20088 43072 20130 43112
rect 20170 43072 20212 43112
rect 20252 43072 20294 43112
rect 20334 43072 20376 43112
rect 20416 43072 20425 43112
rect 0 43052 80 43072
rect 21424 42944 21504 42964
rect 3235 42904 3244 42944
rect 3284 42904 3532 42944
rect 3572 42904 3581 42944
rect 18019 42904 18028 42944
rect 18068 42904 21504 42944
rect 21424 42884 21504 42904
rect 15715 42860 15773 42861
rect 16387 42860 16445 42861
rect 17635 42860 17693 42861
rect 2659 42820 2668 42860
rect 2708 42820 4204 42860
rect 4244 42820 4253 42860
rect 4300 42820 6700 42860
rect 6740 42820 6749 42860
rect 6979 42820 6988 42860
rect 7028 42820 11360 42860
rect 0 42776 80 42796
rect 4300 42776 4340 42820
rect 0 42736 1268 42776
rect 2947 42736 2956 42776
rect 2996 42736 4340 42776
rect 4387 42776 4445 42777
rect 6019 42776 6077 42777
rect 4387 42736 4396 42776
rect 4436 42736 5068 42776
rect 5108 42736 5117 42776
rect 5934 42736 6028 42776
rect 6068 42736 6077 42776
rect 8131 42736 8140 42776
rect 8180 42736 8189 42776
rect 0 42716 80 42736
rect 1228 42608 1268 42736
rect 4387 42735 4445 42736
rect 6019 42735 6077 42736
rect 6028 42692 6068 42735
rect 1315 42652 1324 42692
rect 1364 42652 4820 42692
rect 4867 42652 4876 42692
rect 4916 42652 6068 42692
rect 4780 42608 4820 42652
rect 8140 42608 8180 42736
rect 11320 42692 11360 42820
rect 15715 42820 15724 42860
rect 15764 42820 16396 42860
rect 16436 42820 16445 42860
rect 17539 42820 17548 42860
rect 17588 42820 17644 42860
rect 17684 42820 17693 42860
rect 15715 42819 15773 42820
rect 16387 42819 16445 42820
rect 17635 42819 17693 42820
rect 11320 42652 19756 42692
rect 19796 42652 19805 42692
rect 21379 42608 21437 42609
rect 1228 42568 2540 42608
rect 4780 42568 5260 42608
rect 5300 42568 8180 42608
rect 19171 42568 19180 42608
rect 19220 42568 21388 42608
rect 21428 42568 21437 42608
rect 2500 42524 2540 42568
rect 21379 42567 21437 42568
rect 10243 42524 10301 42525
rect 18787 42524 18845 42525
rect 2500 42484 5164 42524
rect 5204 42484 5213 42524
rect 5443 42484 5452 42524
rect 5492 42484 5740 42524
rect 5780 42484 10252 42524
rect 10292 42484 10301 42524
rect 18702 42484 18796 42524
rect 18836 42484 18845 42524
rect 18979 42484 18988 42524
rect 19028 42484 19037 42524
rect 10243 42483 10301 42484
rect 18787 42483 18845 42484
rect 0 42440 80 42460
rect 18988 42440 19028 42484
rect 0 42400 6604 42440
rect 6644 42400 6653 42440
rect 9187 42400 9196 42440
rect 9236 42400 16972 42440
rect 17012 42400 17021 42440
rect 18700 42400 19028 42440
rect 0 42380 80 42400
rect 3679 42316 3688 42356
rect 3728 42316 3770 42356
rect 3810 42316 3852 42356
rect 3892 42316 3934 42356
rect 3974 42316 4016 42356
rect 4056 42316 4065 42356
rect 5155 42316 5164 42356
rect 5204 42316 6028 42356
rect 6068 42316 14860 42356
rect 14900 42316 14909 42356
rect 18700 42272 18740 42400
rect 18799 42316 18808 42356
rect 18848 42316 18890 42356
rect 18930 42316 18972 42356
rect 19012 42316 19054 42356
rect 19094 42316 19136 42356
rect 19176 42316 19185 42356
rect 21424 42272 21504 42292
rect 2500 42232 17932 42272
rect 17972 42232 18740 42272
rect 19651 42232 19660 42272
rect 19700 42232 21504 42272
rect 0 42104 80 42124
rect 2500 42104 2540 42232
rect 21424 42212 21504 42232
rect 14947 42188 15005 42189
rect 18691 42188 18749 42189
rect 14947 42148 14956 42188
rect 14996 42148 17164 42188
rect 17204 42148 17213 42188
rect 18691 42148 18700 42188
rect 18740 42148 19276 42188
rect 19316 42148 19325 42188
rect 19843 42148 19852 42188
rect 19892 42148 19901 42188
rect 14947 42147 15005 42148
rect 18691 42147 18749 42148
rect 13795 42104 13853 42105
rect 0 42064 2540 42104
rect 8803 42064 8812 42104
rect 8852 42064 10444 42104
rect 10484 42064 11116 42104
rect 11156 42064 11165 42104
rect 13795 42064 13804 42104
rect 13844 42064 18892 42104
rect 18932 42064 18941 42104
rect 0 42044 80 42064
rect 13795 42063 13853 42064
rect 2500 41980 18028 42020
rect 18068 41980 18508 42020
rect 18548 41980 18557 42020
rect 0 41768 80 41788
rect 2500 41768 2540 41980
rect 2659 41896 2668 41936
rect 2708 41896 4012 41936
rect 4052 41896 4061 41936
rect 10819 41896 10828 41936
rect 10868 41896 10908 41936
rect 11107 41896 11116 41936
rect 11156 41896 12076 41936
rect 12116 41896 12940 41936
rect 12980 41896 12989 41936
rect 2947 41852 3005 41853
rect 8611 41852 8669 41853
rect 10828 41852 10868 41896
rect 19852 41852 19892 42148
rect 2947 41812 2956 41852
rect 2996 41812 3532 41852
rect 3572 41812 3581 41852
rect 3907 41812 3916 41852
rect 3956 41812 4108 41852
rect 4148 41812 8620 41852
rect 8660 41812 8669 41852
rect 10051 41812 10060 41852
rect 10100 41812 18700 41852
rect 18740 41812 18749 41852
rect 19843 41812 19852 41852
rect 19892 41812 19901 41852
rect 2947 41811 3005 41812
rect 8611 41811 8669 41812
rect 19651 41768 19709 41769
rect 0 41728 2540 41768
rect 8995 41728 9004 41768
rect 9044 41728 9388 41768
rect 9428 41728 9437 41768
rect 12547 41728 12556 41768
rect 12596 41728 18508 41768
rect 18548 41728 18557 41768
rect 19566 41728 19660 41768
rect 19700 41728 19709 41768
rect 0 41708 80 41728
rect 19651 41727 19709 41728
rect 7555 41684 7613 41685
rect 11299 41684 11357 41685
rect 7470 41644 7564 41684
rect 7604 41644 11308 41684
rect 11348 41644 11357 41684
rect 19939 41644 19948 41684
rect 19988 41644 21044 41684
rect 7555 41643 7613 41644
rect 11299 41643 11357 41644
rect 4387 41600 4445 41601
rect 10723 41600 10781 41601
rect 3523 41560 3532 41600
rect 3572 41560 4396 41600
rect 4436 41560 4445 41600
rect 4919 41560 4928 41600
rect 4968 41560 5010 41600
rect 5050 41560 5092 41600
rect 5132 41560 5174 41600
rect 5214 41560 5256 41600
rect 5296 41560 5305 41600
rect 8803 41560 8812 41600
rect 8852 41560 9004 41600
rect 9044 41560 9053 41600
rect 9283 41560 9292 41600
rect 9332 41560 9484 41600
rect 9524 41560 10732 41600
rect 10772 41560 10781 41600
rect 4387 41559 4445 41560
rect 10723 41559 10781 41560
rect 11587 41600 11645 41601
rect 21004 41600 21044 41644
rect 21424 41600 21504 41620
rect 11587 41560 11596 41600
rect 11636 41560 19372 41600
rect 19412 41560 19421 41600
rect 20039 41560 20048 41600
rect 20088 41560 20130 41600
rect 20170 41560 20212 41600
rect 20252 41560 20294 41600
rect 20334 41560 20376 41600
rect 20416 41560 20425 41600
rect 21004 41560 21504 41600
rect 11587 41559 11645 41560
rect 21424 41540 21504 41560
rect 11875 41516 11933 41517
rect 2467 41476 2476 41516
rect 2516 41476 3340 41516
rect 3380 41476 3389 41516
rect 10531 41476 10540 41516
rect 10580 41476 11596 41516
rect 11636 41476 11884 41516
rect 11924 41476 11933 41516
rect 11875 41475 11933 41476
rect 12844 41476 15956 41516
rect 16003 41476 16012 41516
rect 16052 41476 19660 41516
rect 19700 41476 19709 41516
rect 0 41432 80 41452
rect 12844 41432 12884 41476
rect 13219 41432 13277 41433
rect 0 41392 12884 41432
rect 12931 41392 12940 41432
rect 12980 41392 13228 41432
rect 13268 41392 13277 41432
rect 15916 41432 15956 41476
rect 19843 41432 19901 41433
rect 15916 41392 18892 41432
rect 18932 41392 18941 41432
rect 19075 41392 19084 41432
rect 19124 41392 19852 41432
rect 19892 41392 19901 41432
rect 0 41372 80 41392
rect 13219 41391 13277 41392
rect 19843 41391 19901 41392
rect 9091 41308 9100 41348
rect 9140 41308 10444 41348
rect 10484 41308 10493 41348
rect 11320 41308 19372 41348
rect 19412 41308 19421 41348
rect 5443 41264 5501 41265
rect 6787 41264 6845 41265
rect 11320 41264 11360 41308
rect 11491 41264 11549 41265
rect 1891 41224 1900 41264
rect 1940 41224 4300 41264
rect 4340 41224 4349 41264
rect 4483 41224 4492 41264
rect 4532 41224 4876 41264
rect 4916 41224 4925 41264
rect 5358 41224 5452 41264
rect 5492 41224 5501 41264
rect 6403 41224 6412 41264
rect 6452 41224 6796 41264
rect 6836 41224 6845 41264
rect 5443 41223 5501 41224
rect 6787 41223 6845 41224
rect 6892 41224 11360 41264
rect 11406 41224 11500 41264
rect 11540 41224 11549 41264
rect 12355 41224 12364 41264
rect 12404 41224 20044 41264
rect 20084 41224 20093 41264
rect 5731 41180 5789 41181
rect 1411 41140 1420 41180
rect 1460 41140 2540 41180
rect 0 41096 80 41116
rect 2500 41096 2540 41140
rect 5731 41140 5740 41180
rect 5780 41140 5836 41180
rect 5876 41140 5885 41180
rect 5731 41139 5789 41140
rect 6892 41096 6932 41224
rect 11491 41223 11549 41224
rect 10915 41180 10973 41181
rect 10830 41140 10924 41180
rect 10964 41140 10973 41180
rect 10915 41139 10973 41140
rect 11320 41140 19276 41180
rect 19316 41140 19325 41180
rect 11320 41096 11360 41140
rect 19747 41096 19805 41097
rect 0 41056 212 41096
rect 2500 41056 6932 41096
rect 7267 41056 7276 41096
rect 7316 41056 11360 41096
rect 18979 41056 18988 41096
rect 19028 41056 19756 41096
rect 19796 41056 19805 41096
rect 0 41036 80 41056
rect 172 40928 212 41056
rect 7276 41012 7316 41056
rect 19747 41055 19805 41056
rect 19459 41012 19517 41013
rect 2947 40972 2956 41012
rect 2996 40972 3628 41012
rect 3668 40972 7316 41012
rect 8236 40972 18316 41012
rect 18356 40972 18365 41012
rect 18883 40972 18892 41012
rect 18932 40972 18941 41012
rect 19374 40972 19468 41012
rect 19508 40972 19517 41012
rect 19843 40972 19852 41012
rect 19892 40972 20180 41012
rect 4483 40928 4541 40929
rect 5923 40928 5981 40929
rect 8131 40928 8189 40929
rect 172 40888 4492 40928
rect 4532 40888 5780 40928
rect 5838 40888 5932 40928
rect 5972 40888 8140 40928
rect 8180 40888 8189 40928
rect 4483 40887 4541 40888
rect 5740 40844 5780 40888
rect 5923 40887 5981 40888
rect 8131 40887 8189 40888
rect 8236 40844 8276 40972
rect 18892 40928 18932 40972
rect 19459 40971 19517 40972
rect 3679 40804 3688 40844
rect 3728 40804 3770 40844
rect 3810 40804 3852 40844
rect 3892 40804 3934 40844
rect 3974 40804 4016 40844
rect 4056 40804 4065 40844
rect 5740 40804 8276 40844
rect 11320 40888 18932 40928
rect 20140 40928 20180 40972
rect 21424 40928 21504 40948
rect 20140 40888 21504 40928
rect 0 40760 80 40780
rect 0 40720 2324 40760
rect 4867 40720 4876 40760
rect 4916 40720 5164 40760
rect 5204 40720 6508 40760
rect 6548 40720 7180 40760
rect 7220 40720 7229 40760
rect 8995 40720 9004 40760
rect 9044 40720 10636 40760
rect 10676 40720 10685 40760
rect 0 40700 80 40720
rect 2284 40677 2324 40720
rect 2275 40676 2333 40677
rect 11320 40676 11360 40888
rect 21424 40868 21504 40888
rect 18799 40804 18808 40844
rect 18848 40804 18890 40844
rect 18930 40804 18972 40844
rect 19012 40804 19054 40844
rect 19094 40804 19136 40844
rect 19176 40804 19185 40844
rect 17155 40676 17213 40677
rect 19459 40676 19517 40677
rect 2275 40636 2284 40676
rect 2324 40636 11360 40676
rect 13219 40636 13228 40676
rect 13268 40636 14572 40676
rect 14612 40636 14621 40676
rect 17155 40636 17164 40676
rect 17204 40636 19084 40676
rect 19124 40636 19133 40676
rect 19374 40636 19468 40676
rect 19508 40636 19517 40676
rect 2275 40635 2333 40636
rect 17155 40635 17213 40636
rect 19459 40635 19517 40636
rect 2851 40552 2860 40592
rect 2900 40552 5932 40592
rect 5972 40552 7660 40592
rect 7700 40552 19564 40592
rect 19604 40552 19613 40592
rect 9571 40508 9629 40509
rect 1228 40468 1420 40508
rect 1460 40468 1708 40508
rect 1748 40468 1757 40508
rect 3907 40468 3916 40508
rect 3956 40468 4396 40508
rect 4436 40468 5684 40508
rect 6595 40468 6604 40508
rect 6644 40468 6988 40508
rect 7028 40468 9004 40508
rect 9044 40468 9053 40508
rect 9571 40468 9580 40508
rect 9620 40468 9964 40508
rect 10004 40468 10013 40508
rect 11491 40468 11500 40508
rect 11540 40468 13036 40508
rect 13076 40468 13085 40508
rect 19651 40468 19660 40508
rect 19700 40468 19948 40508
rect 19988 40468 19997 40508
rect 0 40424 80 40444
rect 1228 40424 1268 40468
rect 4771 40424 4829 40425
rect 0 40384 1268 40424
rect 1315 40384 1324 40424
rect 1364 40384 2572 40424
rect 2612 40384 2621 40424
rect 4771 40384 4780 40424
rect 4820 40384 5164 40424
rect 5204 40384 5213 40424
rect 5539 40384 5548 40424
rect 5588 40384 5597 40424
rect 0 40364 80 40384
rect 4771 40383 4829 40384
rect 5548 40340 5588 40384
rect 2371 40300 2380 40340
rect 2420 40300 2668 40340
rect 2708 40300 3148 40340
rect 3188 40300 3197 40340
rect 4099 40300 4108 40340
rect 4148 40300 5588 40340
rect 5644 40340 5684 40468
rect 9571 40467 9629 40468
rect 8419 40424 8477 40425
rect 9859 40424 9917 40425
rect 10435 40424 10493 40425
rect 7171 40384 7180 40424
rect 7220 40384 7756 40424
rect 7796 40384 8428 40424
rect 8468 40384 8908 40424
rect 8948 40384 8957 40424
rect 9774 40384 9868 40424
rect 9908 40384 9917 40424
rect 10350 40384 10444 40424
rect 10484 40384 10493 40424
rect 10627 40384 10636 40424
rect 10676 40384 17740 40424
rect 17780 40384 17789 40424
rect 8419 40383 8477 40384
rect 9859 40383 9917 40384
rect 10435 40383 10493 40384
rect 5644 40300 12748 40340
rect 12788 40300 12797 40340
rect 16867 40256 16925 40257
rect 21424 40256 21504 40276
rect 11011 40216 11020 40256
rect 11060 40216 16876 40256
rect 16916 40216 16925 40256
rect 19843 40216 19852 40256
rect 19892 40216 21504 40256
rect 16867 40215 16925 40216
rect 21424 40196 21504 40216
rect 6787 40132 6796 40172
rect 6836 40132 7180 40172
rect 7220 40132 7229 40172
rect 9763 40132 9772 40172
rect 9812 40132 18988 40172
rect 19028 40132 19037 40172
rect 0 40088 80 40108
rect 0 40048 2860 40088
rect 2900 40048 2909 40088
rect 4919 40048 4928 40088
rect 4968 40048 5010 40088
rect 5050 40048 5092 40088
rect 5132 40048 5174 40088
rect 5214 40048 5256 40088
rect 5296 40048 5305 40088
rect 5347 40048 5356 40088
rect 5396 40048 5740 40088
rect 5780 40048 5789 40088
rect 9955 40048 9964 40088
rect 10004 40048 11360 40088
rect 20039 40048 20048 40088
rect 20088 40048 20130 40088
rect 20170 40048 20212 40088
rect 20252 40048 20294 40088
rect 20334 40048 20376 40088
rect 20416 40048 20425 40088
rect 0 40028 80 40048
rect 11320 40004 11360 40048
rect 16579 40004 16637 40005
rect 20995 40004 21053 40005
rect 2500 39964 10060 40004
rect 10100 39964 10109 40004
rect 11320 39964 16588 40004
rect 16628 39964 16637 40004
rect 19555 39964 19564 40004
rect 19604 39964 21004 40004
rect 21044 39964 21053 40004
rect 2500 39920 2540 39964
rect 16579 39963 16637 39964
rect 20995 39963 21053 39964
rect 1507 39880 1516 39920
rect 1556 39880 2540 39920
rect 3043 39880 3052 39920
rect 3092 39880 5740 39920
rect 5780 39880 5789 39920
rect 5836 39880 11360 39920
rect 19939 39880 19948 39920
rect 19988 39880 21196 39920
rect 21236 39880 21245 39920
rect 5836 39836 5876 39880
rect 2563 39796 2572 39836
rect 2612 39796 5876 39836
rect 11320 39836 11360 39880
rect 11320 39796 19604 39836
rect 0 39752 80 39772
rect 19564 39752 19604 39796
rect 0 39712 1420 39752
rect 1460 39712 2956 39752
rect 2996 39712 3005 39752
rect 3427 39712 3436 39752
rect 3476 39712 4012 39752
rect 4052 39712 4061 39752
rect 6211 39712 6220 39752
rect 6260 39712 6700 39752
rect 6740 39712 6749 39752
rect 6796 39712 6897 39752
rect 6937 39712 7564 39752
rect 7604 39712 7613 39752
rect 8131 39712 8140 39752
rect 8180 39712 8908 39752
rect 8948 39712 10636 39752
rect 10676 39712 10685 39752
rect 11875 39712 11884 39752
rect 11924 39712 15724 39752
rect 15764 39712 19372 39752
rect 19412 39712 19421 39752
rect 19555 39712 19564 39752
rect 19604 39712 19613 39752
rect 0 39692 80 39712
rect 643 39668 701 39669
rect 6796 39668 6836 39712
rect 643 39628 652 39668
rect 692 39628 4588 39668
rect 4628 39628 4637 39668
rect 6115 39628 6124 39668
rect 6164 39628 6836 39668
rect 16291 39628 16300 39668
rect 16340 39628 19756 39668
rect 19796 39628 19805 39668
rect 643 39627 701 39628
rect 9283 39584 9341 39585
rect 13603 39584 13661 39585
rect 21424 39584 21504 39604
rect 76 39544 1516 39584
rect 1556 39544 1804 39584
rect 1844 39544 1853 39584
rect 2755 39544 2764 39584
rect 2804 39544 3340 39584
rect 3380 39544 3389 39584
rect 6499 39544 6508 39584
rect 6548 39544 7468 39584
rect 7508 39544 7517 39584
rect 9198 39544 9292 39584
rect 9332 39544 9341 39584
rect 12835 39544 12844 39584
rect 12884 39544 13228 39584
rect 13268 39544 13277 39584
rect 13603 39544 13612 39584
rect 13652 39544 14572 39584
rect 14612 39544 14621 39584
rect 20515 39544 20524 39584
rect 20564 39544 21504 39584
rect 76 39436 116 39544
rect 9283 39543 9341 39544
rect 13603 39543 13661 39544
rect 21424 39524 21504 39544
rect 931 39460 940 39500
rect 980 39460 4108 39500
rect 4148 39460 4157 39500
rect 15139 39460 15148 39500
rect 15188 39460 19372 39500
rect 19412 39460 19421 39500
rect 0 39376 116 39436
rect 163 39416 221 39417
rect 163 39376 172 39416
rect 212 39376 4492 39416
rect 4532 39376 4541 39416
rect 7939 39376 7948 39416
rect 7988 39376 19660 39416
rect 19700 39376 19709 39416
rect 0 39356 80 39376
rect 163 39375 221 39376
rect 355 39332 413 39333
rect 643 39332 701 39333
rect 355 39292 364 39332
rect 404 39292 652 39332
rect 692 39292 701 39332
rect 3679 39292 3688 39332
rect 3728 39292 3770 39332
rect 3810 39292 3852 39332
rect 3892 39292 3934 39332
rect 3974 39292 4016 39332
rect 4056 39292 4065 39332
rect 355 39291 413 39292
rect 643 39291 701 39292
rect 3331 39248 3389 39249
rect 7948 39248 7988 39376
rect 18799 39292 18808 39332
rect 18848 39292 18890 39332
rect 18930 39292 18972 39332
rect 19012 39292 19054 39332
rect 19094 39292 19136 39332
rect 19176 39292 19185 39332
rect 76 39208 3340 39248
rect 3380 39208 7988 39248
rect 10627 39208 10636 39248
rect 10676 39208 12748 39248
rect 12788 39208 14476 39248
rect 14516 39208 14860 39248
rect 14900 39208 14909 39248
rect 76 39100 116 39208
rect 3331 39207 3389 39208
rect 11683 39124 11692 39164
rect 11732 39124 16300 39164
rect 16340 39124 16349 39164
rect 0 39040 116 39100
rect 18403 39080 18461 39081
rect 20707 39080 20765 39081
rect 1987 39040 1996 39080
rect 2036 39040 2668 39080
rect 2708 39040 2717 39080
rect 6787 39040 6796 39080
rect 6836 39040 8044 39080
rect 8084 39040 8093 39080
rect 9091 39040 9100 39080
rect 9140 39040 10156 39080
rect 10196 39040 10205 39080
rect 14371 39040 14380 39080
rect 14420 39040 15244 39080
rect 15284 39040 15293 39080
rect 18403 39040 18412 39080
rect 18452 39040 20716 39080
rect 20756 39040 20765 39080
rect 0 39020 80 39040
rect 18403 39039 18461 39040
rect 20707 39039 20765 39040
rect 5251 38956 5260 38996
rect 5300 38956 6028 38996
rect 6068 38956 6077 38996
rect 6883 38956 6892 38996
rect 6932 38956 7276 38996
rect 7316 38956 7325 38996
rect 7651 38956 7660 38996
rect 7700 38956 8332 38996
rect 8372 38956 9196 38996
rect 9236 38956 9245 38996
rect 12931 38956 12940 38996
rect 12980 38956 13132 38996
rect 13172 38956 13181 38996
rect 3235 38912 3293 38913
rect 11683 38912 11741 38913
rect 13411 38912 13469 38913
rect 21424 38912 21504 38932
rect 1315 38872 1324 38912
rect 1364 38872 1996 38912
rect 2036 38872 2045 38912
rect 3150 38872 3244 38912
rect 3284 38872 3293 38912
rect 5923 38872 5932 38912
rect 5972 38872 8716 38912
rect 8756 38872 8765 38912
rect 11683 38872 11692 38912
rect 11732 38872 13420 38912
rect 13460 38872 13469 38912
rect 19267 38872 19276 38912
rect 19316 38872 21504 38912
rect 3235 38871 3293 38872
rect 11683 38871 11741 38872
rect 13411 38871 13469 38872
rect 3244 38828 3284 38871
rect 21424 38852 21504 38872
rect 4771 38828 4829 38829
rect 3244 38788 4780 38828
rect 4820 38788 6508 38828
rect 6548 38788 6557 38828
rect 20140 38788 21292 38828
rect 21332 38788 21341 38828
rect 4771 38787 4829 38788
rect 0 38744 80 38764
rect 2467 38744 2525 38745
rect 10435 38744 10493 38745
rect 20140 38744 20180 38788
rect 0 38704 2476 38744
rect 2516 38704 2525 38744
rect 10339 38704 10348 38744
rect 10388 38704 10444 38744
rect 10484 38704 10493 38744
rect 14659 38704 14668 38744
rect 14708 38704 20180 38744
rect 0 38684 80 38704
rect 2467 38703 2525 38704
rect 10435 38703 10493 38704
rect 7075 38660 7133 38661
rect 14083 38660 14141 38661
rect 1987 38620 1996 38660
rect 2036 38620 7084 38660
rect 7124 38620 7133 38660
rect 9667 38620 9676 38660
rect 9716 38620 14092 38660
rect 14132 38620 14141 38660
rect 7075 38619 7133 38620
rect 14083 38619 14141 38620
rect 4919 38536 4928 38576
rect 4968 38536 5010 38576
rect 5050 38536 5092 38576
rect 5132 38536 5174 38576
rect 5214 38536 5256 38576
rect 5296 38536 5305 38576
rect 7171 38536 7180 38576
rect 7220 38536 8812 38576
rect 8852 38536 8861 38576
rect 20039 38536 20048 38576
rect 20088 38536 20130 38576
rect 20170 38536 20212 38576
rect 20252 38536 20294 38576
rect 20334 38536 20376 38576
rect 20416 38536 20425 38576
rect 7075 38492 7133 38493
rect 4291 38452 4300 38492
rect 4340 38452 6644 38492
rect 0 38408 80 38428
rect 1411 38408 1469 38409
rect 0 38368 1420 38408
rect 1460 38368 1469 38408
rect 6604 38408 6644 38452
rect 7075 38452 7084 38492
rect 7124 38452 18700 38492
rect 18740 38452 18749 38492
rect 7075 38451 7133 38452
rect 6604 38368 19276 38408
rect 19316 38368 19325 38408
rect 0 38348 80 38368
rect 1411 38367 1469 38368
rect 1603 38284 1612 38324
rect 1652 38284 4396 38324
rect 4436 38284 4445 38324
rect 5155 38284 5164 38324
rect 5204 38284 6988 38324
rect 7028 38284 7037 38324
rect 21424 38240 21504 38260
rect 2275 38200 2284 38240
rect 2324 38200 2860 38240
rect 2900 38200 2909 38240
rect 3139 38200 3148 38240
rect 3188 38200 3724 38240
rect 3764 38200 3773 38240
rect 5539 38200 5548 38240
rect 5588 38200 6124 38240
rect 6164 38200 6173 38240
rect 8515 38200 8524 38240
rect 8564 38200 8908 38240
rect 8948 38200 8957 38240
rect 11491 38200 11500 38240
rect 11540 38200 11692 38240
rect 11732 38200 11741 38240
rect 13027 38200 13036 38240
rect 13076 38200 13516 38240
rect 13556 38200 13565 38240
rect 13891 38200 13900 38240
rect 13940 38200 14092 38240
rect 14132 38200 14141 38240
rect 19555 38200 19564 38240
rect 19604 38200 21504 38240
rect 2860 38156 2900 38200
rect 21424 38180 21504 38200
rect 5827 38156 5885 38157
rect 2860 38116 4780 38156
rect 4820 38116 4972 38156
rect 5012 38116 5021 38156
rect 5827 38116 5836 38156
rect 5876 38116 6028 38156
rect 6068 38116 6077 38156
rect 5827 38115 5885 38116
rect 0 38072 80 38092
rect 8707 38072 8765 38073
rect 0 38032 1612 38072
rect 1652 38032 1661 38072
rect 6979 38032 6988 38072
rect 7028 38032 7276 38072
rect 7316 38032 7325 38072
rect 8707 38032 8716 38072
rect 8756 38032 19564 38072
rect 19604 38032 19613 38072
rect 0 38012 80 38032
rect 8707 38031 8765 38032
rect 12739 37948 12748 37988
rect 12788 37948 12940 37988
rect 12980 37948 12989 37988
rect 14179 37948 14188 37988
rect 14228 37948 15052 37988
rect 15092 37948 15101 37988
rect 2563 37864 2572 37904
rect 2612 37864 6700 37904
rect 6740 37864 7948 37904
rect 7988 37864 7997 37904
rect 10243 37864 10252 37904
rect 10292 37864 10301 37904
rect 11404 37864 13132 37904
rect 13172 37864 13324 37904
rect 13364 37864 13373 37904
rect 13507 37864 13516 37904
rect 13556 37864 13900 37904
rect 13940 37864 13949 37904
rect 15427 37864 15436 37904
rect 15476 37864 15820 37904
rect 15860 37864 15869 37904
rect 3139 37780 3148 37820
rect 3188 37780 3284 37820
rect 3679 37780 3688 37820
rect 3728 37780 3770 37820
rect 3810 37780 3852 37820
rect 3892 37780 3934 37820
rect 3974 37780 4016 37820
rect 4056 37780 4065 37820
rect 0 37736 80 37756
rect 3244 37736 3284 37780
rect 10252 37736 10292 37864
rect 11404 37820 11444 37864
rect 11587 37820 11645 37821
rect 10444 37780 11404 37820
rect 11444 37780 11453 37820
rect 11502 37780 11596 37820
rect 11636 37780 11645 37820
rect 10444 37736 10484 37780
rect 11587 37779 11645 37780
rect 14284 37780 14476 37820
rect 14516 37780 14525 37820
rect 18799 37780 18808 37820
rect 18848 37780 18890 37820
rect 18930 37780 18972 37820
rect 19012 37780 19054 37820
rect 19094 37780 19136 37820
rect 19176 37780 19185 37820
rect 13603 37736 13661 37737
rect 0 37696 1324 37736
rect 1364 37696 1373 37736
rect 3244 37696 3380 37736
rect 9763 37696 9772 37736
rect 9812 37696 10292 37736
rect 10339 37696 10348 37736
rect 10388 37696 10444 37736
rect 10484 37696 10493 37736
rect 11020 37696 11308 37736
rect 11348 37696 11357 37736
rect 12643 37696 12652 37736
rect 12692 37696 13612 37736
rect 13652 37696 13661 37736
rect 0 37676 80 37696
rect 3340 37652 3380 37696
rect 11020 37652 11060 37696
rect 13603 37695 13661 37696
rect 3340 37612 9676 37652
rect 9716 37612 11060 37652
rect 11107 37652 11165 37653
rect 14284 37652 14324 37780
rect 11107 37612 11116 37652
rect 11156 37612 13612 37652
rect 13652 37612 14324 37652
rect 16099 37652 16157 37653
rect 16099 37612 16108 37652
rect 16148 37612 19948 37652
rect 19988 37612 19997 37652
rect 11107 37611 11165 37612
rect 16099 37611 16157 37612
rect 21424 37568 21504 37588
rect 3523 37528 3532 37568
rect 3572 37528 7276 37568
rect 7316 37528 7325 37568
rect 7843 37528 7852 37568
rect 7892 37528 14380 37568
rect 14420 37528 14429 37568
rect 18691 37528 18700 37568
rect 18740 37528 21504 37568
rect 21424 37508 21504 37528
rect 12067 37484 12125 37485
rect 19555 37484 19613 37485
rect 1411 37444 1420 37484
rect 1460 37444 1900 37484
rect 1940 37444 1949 37484
rect 5443 37444 5452 37484
rect 5492 37444 5836 37484
rect 5876 37444 6644 37484
rect 6691 37444 6700 37484
rect 6740 37444 7083 37484
rect 7123 37444 7132 37484
rect 9955 37444 9964 37484
rect 10004 37444 10444 37484
rect 10484 37444 10493 37484
rect 12067 37444 12076 37484
rect 12116 37444 12172 37484
rect 12212 37444 12221 37484
rect 19470 37444 19564 37484
rect 19604 37444 19613 37484
rect 0 37400 80 37420
rect 3043 37400 3101 37401
rect 6604 37400 6644 37444
rect 12067 37443 12125 37444
rect 19555 37443 19613 37444
rect 0 37360 2572 37400
rect 2612 37360 2621 37400
rect 2851 37360 2860 37400
rect 2900 37360 3052 37400
rect 3092 37360 3101 37400
rect 3619 37360 3628 37400
rect 3668 37360 4436 37400
rect 6595 37360 6604 37400
rect 6644 37360 9772 37400
rect 9812 37360 9821 37400
rect 11587 37360 11596 37400
rect 11636 37360 12556 37400
rect 12596 37360 12605 37400
rect 0 37340 80 37360
rect 3043 37359 3101 37360
rect 1315 37316 1373 37317
rect 4396 37316 4436 37360
rect 11596 37316 11636 37360
rect 1315 37276 1324 37316
rect 1364 37276 4300 37316
rect 4340 37276 4349 37316
rect 4396 37276 9044 37316
rect 10915 37276 10924 37316
rect 10964 37276 11636 37316
rect 12163 37276 12172 37316
rect 12212 37276 13036 37316
rect 13076 37276 13085 37316
rect 18979 37276 18988 37316
rect 19028 37276 19660 37316
rect 19700 37276 19709 37316
rect 1315 37275 1373 37276
rect 835 37232 893 37233
rect 8035 37232 8093 37233
rect 9004 37232 9044 37276
rect 11107 37232 11165 37233
rect 11587 37232 11645 37233
rect 835 37192 844 37232
rect 884 37192 4108 37232
rect 4148 37192 4157 37232
rect 7747 37192 7756 37232
rect 7796 37192 8044 37232
rect 8084 37192 8093 37232
rect 8995 37192 9004 37232
rect 9044 37192 11116 37232
rect 11156 37192 11165 37232
rect 835 37191 893 37192
rect 8035 37191 8093 37192
rect 11107 37191 11165 37192
rect 11320 37192 11596 37232
rect 11636 37192 11732 37232
rect 11779 37192 11788 37232
rect 11828 37192 12844 37232
rect 12884 37192 12893 37232
rect 18883 37192 18892 37232
rect 18932 37192 19468 37232
rect 19508 37192 19517 37232
rect 7459 37148 7517 37149
rect 11320 37148 11360 37192
rect 11587 37191 11645 37192
rect 4291 37108 4300 37148
rect 4340 37108 7468 37148
rect 7508 37108 7852 37148
rect 7892 37108 7901 37148
rect 7948 37108 11360 37148
rect 11692 37148 11732 37192
rect 11692 37108 19756 37148
rect 19796 37108 19805 37148
rect 7459 37107 7517 37108
rect 0 37064 80 37084
rect 0 37024 1420 37064
rect 1460 37024 1469 37064
rect 4919 37024 4928 37064
rect 4968 37024 5010 37064
rect 5050 37024 5092 37064
rect 5132 37024 5174 37064
rect 5214 37024 5256 37064
rect 5296 37024 5305 37064
rect 7171 37024 7180 37064
rect 7220 37024 7468 37064
rect 7508 37024 7517 37064
rect 0 37004 80 37024
rect 6883 36980 6941 36981
rect 7948 36980 7988 37108
rect 11203 37024 11212 37064
rect 11252 37024 12652 37064
rect 12692 37024 12701 37064
rect 13315 37024 13324 37064
rect 13364 37024 13804 37064
rect 13844 37024 13853 37064
rect 20039 37024 20048 37064
rect 20088 37024 20130 37064
rect 20170 37024 20212 37064
rect 20252 37024 20294 37064
rect 20334 37024 20376 37064
rect 20416 37024 20425 37064
rect 2467 36940 2476 36980
rect 2516 36940 6740 36980
rect 1603 36856 1612 36896
rect 1652 36856 2956 36896
rect 2996 36856 3005 36896
rect 5347 36812 5405 36813
rect 5155 36772 5164 36812
rect 5204 36772 5356 36812
rect 5396 36772 5405 36812
rect 6700 36812 6740 36940
rect 6883 36940 6892 36980
rect 6932 36940 7988 36980
rect 10147 36940 10156 36980
rect 10196 36940 10732 36980
rect 10772 36940 10781 36980
rect 10828 36940 12076 36980
rect 12116 36940 12125 36980
rect 6883 36939 6941 36940
rect 8419 36896 8477 36897
rect 10828 36896 10868 36940
rect 13219 36896 13277 36897
rect 21424 36896 21504 36916
rect 8419 36856 8428 36896
rect 8468 36856 8716 36896
rect 8756 36856 10060 36896
rect 10100 36856 10109 36896
rect 10819 36856 10828 36896
rect 10868 36856 10877 36896
rect 12259 36856 12268 36896
rect 12308 36856 13036 36896
rect 13076 36856 13085 36896
rect 13219 36856 13228 36896
rect 13268 36856 13362 36896
rect 19171 36856 19180 36896
rect 19220 36856 21504 36896
rect 8419 36855 8477 36856
rect 13219 36855 13277 36856
rect 21424 36836 21504 36856
rect 10243 36812 10301 36813
rect 17443 36812 17501 36813
rect 6700 36772 10252 36812
rect 10292 36772 10388 36812
rect 12835 36772 12844 36812
rect 12884 36772 14036 36812
rect 5347 36771 5405 36772
rect 10243 36771 10301 36772
rect 0 36728 80 36748
rect 6883 36728 6941 36729
rect 10348 36728 10388 36772
rect 12931 36728 12989 36729
rect 13996 36728 14036 36772
rect 17443 36772 17452 36812
rect 17492 36772 19564 36812
rect 19604 36772 19613 36812
rect 17443 36771 17501 36772
rect 0 36688 6892 36728
rect 6932 36688 6941 36728
rect 7459 36688 7468 36728
rect 7508 36688 9676 36728
rect 9716 36688 9725 36728
rect 10339 36688 10348 36728
rect 10388 36688 10397 36728
rect 11011 36688 11020 36728
rect 11060 36688 11788 36728
rect 11828 36688 11837 36728
rect 12846 36688 12940 36728
rect 12980 36688 12989 36728
rect 13987 36688 13996 36728
rect 14036 36688 14045 36728
rect 0 36668 80 36688
rect 6883 36687 6941 36688
rect 12931 36687 12989 36688
rect 11683 36644 11741 36645
rect 11971 36644 12029 36645
rect 2275 36604 2284 36644
rect 2324 36604 2476 36644
rect 2516 36604 4108 36644
rect 4148 36604 4157 36644
rect 5539 36604 5548 36644
rect 5588 36604 7084 36644
rect 7124 36604 7133 36644
rect 7267 36604 7276 36644
rect 7316 36604 7564 36644
rect 7604 36604 7613 36644
rect 10051 36604 10060 36644
rect 10100 36604 10828 36644
rect 10868 36604 10877 36644
rect 11587 36604 11596 36644
rect 11636 36604 11692 36644
rect 11732 36604 11980 36644
rect 12020 36604 12029 36644
rect 12739 36604 12748 36644
rect 12788 36604 13900 36644
rect 13940 36604 13949 36644
rect 19363 36604 19372 36644
rect 19412 36604 19660 36644
rect 19700 36604 19709 36644
rect 11683 36603 11741 36604
rect 11971 36603 12029 36604
rect 18595 36560 18653 36561
rect 20515 36560 20573 36561
rect 2947 36520 2956 36560
rect 2996 36520 3628 36560
rect 3668 36520 3677 36560
rect 6211 36520 6220 36560
rect 6260 36520 8716 36560
rect 8756 36520 8765 36560
rect 10531 36520 10540 36560
rect 10580 36520 12460 36560
rect 12500 36520 12509 36560
rect 18595 36520 18604 36560
rect 18644 36520 20524 36560
rect 20564 36520 20573 36560
rect 18595 36519 18653 36520
rect 20515 36519 20573 36520
rect 13603 36476 13661 36477
rect 7555 36436 7564 36476
rect 7604 36436 11308 36476
rect 11348 36436 11357 36476
rect 11980 36436 13612 36476
rect 13652 36436 13661 36476
rect 18883 36436 18892 36476
rect 18932 36436 18941 36476
rect 0 36392 80 36412
rect 1603 36392 1661 36393
rect 7843 36392 7901 36393
rect 10435 36392 10493 36393
rect 0 36352 1612 36392
rect 1652 36352 1661 36392
rect 2083 36352 2092 36392
rect 2132 36352 7852 36392
rect 7892 36352 10060 36392
rect 10100 36352 10109 36392
rect 10339 36352 10348 36392
rect 10388 36352 10444 36392
rect 10484 36352 10493 36392
rect 0 36332 80 36352
rect 1603 36351 1661 36352
rect 7843 36351 7901 36352
rect 10435 36351 10493 36352
rect 11980 36308 12020 36436
rect 13603 36435 13661 36436
rect 18892 36392 18932 36436
rect 3679 36268 3688 36308
rect 3728 36268 3770 36308
rect 3810 36268 3852 36308
rect 3892 36268 3934 36308
rect 3974 36268 4016 36308
rect 4056 36268 4065 36308
rect 6892 36268 12020 36308
rect 12076 36352 18932 36392
rect 2371 36184 2380 36224
rect 2420 36184 2668 36224
rect 2708 36184 2717 36224
rect 2083 36140 2141 36141
rect 6892 36140 6932 36268
rect 12076 36224 12116 36352
rect 13315 36268 13324 36308
rect 13364 36268 13708 36308
rect 13748 36268 13757 36308
rect 18799 36268 18808 36308
rect 18848 36268 18890 36308
rect 18930 36268 18972 36308
rect 19012 36268 19054 36308
rect 19094 36268 19136 36308
rect 19176 36268 19185 36308
rect 19555 36268 19564 36308
rect 19604 36268 21100 36308
rect 21140 36268 21149 36308
rect 21424 36224 21504 36244
rect 9571 36184 9580 36224
rect 9620 36184 11252 36224
rect 11299 36184 11308 36224
rect 11348 36184 12116 36224
rect 12172 36184 15340 36224
rect 15380 36184 15389 36224
rect 19267 36184 19276 36224
rect 19316 36184 21504 36224
rect 10819 36140 10877 36141
rect 2083 36100 2092 36140
rect 2132 36100 2188 36140
rect 2228 36100 6932 36140
rect 7084 36100 10828 36140
rect 10868 36100 10877 36140
rect 11212 36140 11252 36184
rect 12172 36140 12212 36184
rect 21424 36164 21504 36184
rect 11212 36100 12212 36140
rect 12259 36100 12268 36140
rect 12308 36100 12844 36140
rect 12884 36100 12893 36140
rect 2083 36099 2141 36100
rect 0 36056 80 36076
rect 7084 36056 7124 36100
rect 10819 36099 10877 36100
rect 0 36016 2540 36056
rect 3235 36016 3244 36056
rect 3284 36016 7124 36056
rect 10243 36016 10252 36056
rect 10292 36016 10540 36056
rect 10580 36016 10589 36056
rect 10723 36016 10732 36056
rect 10772 36016 10924 36056
rect 10964 36016 10973 36056
rect 12643 36016 12652 36056
rect 12692 36016 13228 36056
rect 13268 36016 13277 36056
rect 19171 36016 19180 36056
rect 19220 36016 20620 36056
rect 20660 36016 20669 36056
rect 0 35996 80 36016
rect 2500 35972 2540 36016
rect 10540 35972 10580 36016
rect 2500 35932 5836 35972
rect 5876 35932 9580 35972
rect 9620 35932 9629 35972
rect 10540 35932 11020 35972
rect 11060 35932 11069 35972
rect 12931 35932 12940 35972
rect 12980 35932 14476 35972
rect 14516 35932 14525 35972
rect 3235 35888 3293 35889
rect 1315 35848 1324 35888
rect 1364 35848 1900 35888
rect 1940 35848 1949 35888
rect 2659 35848 2668 35888
rect 2708 35848 3244 35888
rect 3284 35848 4108 35888
rect 4148 35848 4157 35888
rect 4675 35848 4684 35888
rect 4724 35848 4972 35888
rect 5012 35848 5021 35888
rect 6595 35848 6604 35888
rect 6644 35848 6892 35888
rect 6932 35848 6941 35888
rect 10051 35848 10060 35888
rect 10100 35848 10580 35888
rect 10627 35848 10636 35888
rect 10676 35848 11788 35888
rect 11828 35848 11837 35888
rect 12067 35848 12076 35888
rect 12116 35848 12556 35888
rect 12596 35848 12605 35888
rect 13411 35848 13420 35888
rect 13460 35848 13469 35888
rect 14179 35848 14188 35888
rect 14228 35848 14860 35888
rect 14900 35848 14909 35888
rect 3235 35847 3293 35848
rect 10540 35804 10580 35848
rect 13420 35804 13460 35848
rect 2563 35764 2572 35804
rect 2612 35764 2860 35804
rect 2900 35764 7564 35804
rect 7604 35764 7613 35804
rect 10540 35764 10732 35804
rect 10772 35764 10781 35804
rect 10924 35764 11596 35804
rect 11636 35764 11645 35804
rect 13420 35764 21388 35804
rect 21428 35764 21437 35804
rect 0 35720 80 35740
rect 1315 35720 1373 35721
rect 10924 35720 10964 35764
rect 13507 35720 13565 35721
rect 0 35680 1324 35720
rect 1364 35680 1373 35720
rect 10531 35680 10540 35720
rect 10580 35680 10964 35720
rect 11011 35680 11020 35720
rect 11060 35680 11308 35720
rect 11348 35680 11357 35720
rect 11491 35680 11500 35720
rect 11540 35680 11828 35720
rect 12739 35680 12748 35720
rect 12788 35680 13228 35720
rect 13268 35680 13516 35720
rect 13556 35680 13565 35720
rect 0 35660 80 35680
rect 1315 35679 1373 35680
rect 3139 35636 3197 35637
rect 11491 35636 11549 35637
rect 11788 35636 11828 35680
rect 13507 35679 13565 35680
rect 12259 35636 12317 35637
rect 3139 35596 3148 35636
rect 3188 35596 4588 35636
rect 4628 35596 11500 35636
rect 11540 35596 11549 35636
rect 11779 35596 11788 35636
rect 11828 35596 11837 35636
rect 12259 35596 12268 35636
rect 12308 35596 19948 35636
rect 19988 35596 19997 35636
rect 3139 35595 3197 35596
rect 11491 35595 11549 35596
rect 12259 35595 12317 35596
rect 18019 35552 18077 35553
rect 21424 35552 21504 35572
rect 4919 35512 4928 35552
rect 4968 35512 5010 35552
rect 5050 35512 5092 35552
rect 5132 35512 5174 35552
rect 5214 35512 5256 35552
rect 5296 35512 5305 35552
rect 7747 35512 7756 35552
rect 7796 35512 8140 35552
rect 8180 35512 8189 35552
rect 9379 35512 9388 35552
rect 9428 35512 9676 35552
rect 9716 35512 9725 35552
rect 10819 35512 10828 35552
rect 10868 35512 11308 35552
rect 11348 35512 11357 35552
rect 11404 35512 18028 35552
rect 18068 35512 18077 35552
rect 20039 35512 20048 35552
rect 20088 35512 20130 35552
rect 20170 35512 20212 35552
rect 20252 35512 20294 35552
rect 20334 35512 20376 35552
rect 20416 35512 20425 35552
rect 21379 35512 21388 35552
rect 21428 35512 21504 35552
rect 10819 35468 10877 35469
rect 11404 35468 11444 35512
rect 18019 35511 18077 35512
rect 21424 35492 21504 35512
rect 10819 35428 10828 35468
rect 10868 35428 11444 35468
rect 13219 35428 13228 35468
rect 13268 35428 13804 35468
rect 13844 35428 13853 35468
rect 10819 35427 10877 35428
rect 0 35384 80 35404
rect 1315 35384 1373 35385
rect 0 35344 1324 35384
rect 1364 35344 1373 35384
rect 4483 35344 4492 35384
rect 4532 35344 4541 35384
rect 5155 35344 5164 35384
rect 5204 35344 5452 35384
rect 5492 35344 5501 35384
rect 6499 35344 6508 35384
rect 6548 35344 6557 35384
rect 6883 35344 6892 35384
rect 6932 35344 8044 35384
rect 8084 35344 8093 35384
rect 12652 35344 13324 35384
rect 13364 35344 13516 35384
rect 13556 35344 13565 35384
rect 0 35324 80 35344
rect 1315 35343 1373 35344
rect 4492 35300 4532 35344
rect 5827 35300 5885 35301
rect 6508 35300 6548 35344
rect 7651 35300 7709 35301
rect 12652 35300 12692 35344
rect 13411 35300 13469 35301
rect 2851 35260 2860 35300
rect 2900 35260 4108 35300
rect 4148 35260 4532 35300
rect 5742 35260 5836 35300
rect 5876 35260 5885 35300
rect 6019 35260 6028 35300
rect 6068 35260 6548 35300
rect 6595 35260 6604 35300
rect 6644 35260 7660 35300
rect 7700 35260 7709 35300
rect 5827 35259 5885 35260
rect 7651 35259 7709 35260
rect 10540 35260 11360 35300
rect 3043 35176 3052 35216
rect 3092 35176 4300 35216
rect 4340 35176 4349 35216
rect 5443 35176 5452 35216
rect 5492 35176 5740 35216
rect 5780 35176 6220 35216
rect 6260 35176 6269 35216
rect 6979 35176 6988 35216
rect 7028 35176 7037 35216
rect 5539 35132 5597 35133
rect 6787 35132 6845 35133
rect 3811 35092 3820 35132
rect 3860 35092 5548 35132
rect 5588 35092 5597 35132
rect 6702 35092 6796 35132
rect 6836 35092 6845 35132
rect 0 35048 80 35068
rect 3811 35048 3869 35049
rect 4492 35048 4532 35092
rect 5539 35091 5597 35092
rect 6787 35091 6845 35092
rect 6988 35048 7028 35176
rect 10540 35132 10580 35260
rect 11320 35216 11360 35260
rect 11404 35260 11884 35300
rect 11924 35260 12692 35300
rect 12739 35260 12748 35300
rect 12788 35260 13420 35300
rect 13460 35260 13469 35300
rect 19171 35260 19180 35300
rect 19220 35260 21004 35300
rect 21044 35260 21053 35300
rect 11404 35216 11444 35260
rect 13411 35259 13469 35260
rect 11779 35216 11837 35217
rect 11107 35176 11116 35216
rect 11156 35176 11165 35216
rect 11320 35176 11404 35216
rect 11444 35176 11453 35216
rect 11694 35176 11788 35216
rect 11828 35176 11837 35216
rect 12067 35176 12076 35216
rect 12116 35176 13036 35216
rect 13076 35176 13085 35216
rect 14275 35176 14284 35216
rect 14324 35176 14764 35216
rect 14804 35176 14813 35216
rect 15523 35176 15532 35216
rect 15572 35176 19756 35216
rect 19796 35176 19805 35216
rect 11116 35132 11156 35176
rect 11779 35175 11837 35176
rect 13795 35132 13853 35133
rect 10531 35092 10540 35132
rect 10580 35092 10589 35132
rect 11116 35092 11444 35132
rect 11491 35092 11500 35132
rect 11540 35092 12172 35132
rect 12212 35092 12221 35132
rect 12547 35092 12556 35132
rect 12596 35092 13132 35132
rect 13172 35092 13181 35132
rect 13795 35092 13804 35132
rect 13844 35092 19372 35132
rect 19412 35092 19421 35132
rect 11107 35048 11165 35049
rect 11404 35048 11444 35092
rect 13795 35091 13853 35092
rect 21283 35048 21341 35049
rect 0 35008 1996 35048
rect 2036 35008 2045 35048
rect 3715 35008 3724 35048
rect 3764 35008 3820 35048
rect 3860 35008 4436 35048
rect 4483 35008 4492 35048
rect 4532 35008 4572 35048
rect 4771 35008 4780 35048
rect 4820 35008 7028 35048
rect 10051 35008 10060 35048
rect 10100 35008 10444 35048
rect 10484 35008 10493 35048
rect 10819 35008 10828 35048
rect 10868 35008 11116 35048
rect 11156 35008 11165 35048
rect 11395 35008 11404 35048
rect 11444 35008 11453 35048
rect 12643 35008 12652 35048
rect 12692 35008 12940 35048
rect 12980 35008 13516 35048
rect 13556 35008 14092 35048
rect 14132 35008 14476 35048
rect 14516 35008 14525 35048
rect 18307 35008 18316 35048
rect 18356 35008 18978 35048
rect 19018 35008 19027 35048
rect 19555 35008 19564 35048
rect 19604 35008 21292 35048
rect 21332 35008 21341 35048
rect 0 34988 80 35008
rect 3811 35007 3869 35008
rect 4396 34964 4436 35008
rect 11107 35007 11165 35008
rect 21283 35007 21341 35008
rect 172 34924 2956 34964
rect 2996 34924 3005 34964
rect 3235 34924 3244 34964
rect 3284 34924 3532 34964
rect 3572 34924 4108 34964
rect 4148 34924 4157 34964
rect 4396 34924 10252 34964
rect 10292 34924 10636 34964
rect 10676 34924 10685 34964
rect 11107 34924 11116 34964
rect 11156 34924 11500 34964
rect 11540 34924 11549 34964
rect 13411 34924 13420 34964
rect 13460 34924 14188 34964
rect 14228 34924 14237 34964
rect 16579 34924 16588 34964
rect 16628 34924 20180 34964
rect 172 34880 212 34924
rect 9571 34880 9629 34881
rect 20140 34880 20180 34924
rect 21424 34880 21504 34900
rect 67 34840 76 34880
rect 116 34840 212 34880
rect 2371 34840 2380 34880
rect 2420 34840 4588 34880
rect 4628 34840 9580 34880
rect 9620 34840 9629 34880
rect 13315 34840 13324 34880
rect 13364 34840 13708 34880
rect 13748 34840 13757 34880
rect 15340 34840 19468 34880
rect 19508 34840 19517 34880
rect 20140 34840 21504 34880
rect 9571 34839 9629 34840
rect 8419 34796 8477 34797
rect 15340 34796 15380 34840
rect 21424 34820 21504 34840
rect 1219 34756 1228 34796
rect 1268 34756 1420 34796
rect 1460 34756 2612 34796
rect 3679 34756 3688 34796
rect 3728 34756 3770 34796
rect 3810 34756 3852 34796
rect 3892 34756 3934 34796
rect 3974 34756 4016 34796
rect 4056 34756 4065 34796
rect 4108 34756 6892 34796
rect 6932 34756 8428 34796
rect 8468 34756 15380 34796
rect 18799 34756 18808 34796
rect 18848 34756 18890 34796
rect 18930 34756 18972 34796
rect 19012 34756 19054 34796
rect 19094 34756 19136 34796
rect 19176 34756 19185 34796
rect 0 34712 80 34732
rect 2572 34712 2612 34756
rect 4108 34712 4148 34756
rect 8419 34755 8477 34756
rect 9571 34712 9629 34713
rect 0 34672 76 34712
rect 116 34672 125 34712
rect 2572 34672 4148 34712
rect 5251 34672 5260 34712
rect 5300 34672 5932 34712
rect 5972 34672 5981 34712
rect 6691 34672 6700 34712
rect 6740 34672 7948 34712
rect 7988 34672 7997 34712
rect 9571 34672 9580 34712
rect 9620 34672 15532 34712
rect 15572 34672 15581 34712
rect 0 34652 80 34672
rect 9571 34671 9629 34672
rect 10243 34628 10301 34629
rect 13123 34628 13181 34629
rect 13795 34628 13853 34629
rect 17251 34628 17309 34629
rect 6403 34588 6412 34628
rect 6452 34588 7468 34628
rect 7508 34588 7517 34628
rect 10243 34588 10252 34628
rect 10292 34588 11116 34628
rect 11156 34588 11165 34628
rect 11320 34588 13132 34628
rect 13172 34588 13804 34628
rect 13844 34588 13853 34628
rect 14371 34588 14380 34628
rect 14420 34588 14429 34628
rect 17251 34588 17260 34628
rect 17300 34588 19564 34628
rect 19604 34588 19613 34628
rect 10243 34587 10301 34588
rect 2659 34504 2668 34544
rect 2708 34504 10924 34544
rect 10964 34504 10973 34544
rect 11320 34460 11360 34588
rect 13123 34587 13181 34588
rect 13795 34587 13853 34588
rect 14380 34544 14420 34588
rect 17251 34587 17309 34588
rect 11587 34504 11596 34544
rect 11636 34504 11980 34544
rect 12020 34504 12940 34544
rect 12980 34504 12989 34544
rect 13036 34504 13228 34544
rect 13268 34504 13277 34544
rect 13795 34504 13804 34544
rect 13844 34504 14188 34544
rect 14228 34504 14237 34544
rect 14380 34504 19756 34544
rect 19796 34504 19805 34544
rect 13036 34460 13076 34504
rect 1987 34420 1996 34460
rect 2036 34420 2540 34460
rect 0 34376 80 34396
rect 2179 34376 2237 34377
rect 0 34336 1652 34376
rect 2094 34336 2188 34376
rect 2228 34336 2237 34376
rect 2500 34376 2540 34420
rect 2668 34420 11360 34460
rect 12067 34420 12076 34460
rect 12116 34420 12556 34460
rect 12596 34420 12605 34460
rect 13027 34420 13036 34460
rect 13076 34420 13085 34460
rect 14563 34420 14572 34460
rect 14612 34420 14621 34460
rect 2668 34376 2708 34420
rect 6019 34376 6077 34377
rect 8323 34376 8381 34377
rect 9091 34376 9149 34377
rect 2500 34336 2708 34376
rect 3811 34336 3820 34376
rect 3860 34336 4204 34376
rect 4244 34336 4396 34376
rect 4436 34336 4445 34376
rect 5059 34336 5068 34376
rect 5108 34336 5548 34376
rect 5588 34336 5597 34376
rect 6019 34336 6028 34376
rect 6068 34336 6124 34376
rect 6164 34336 6173 34376
rect 6307 34336 6316 34376
rect 6356 34336 7756 34376
rect 7796 34336 8140 34376
rect 8180 34336 8189 34376
rect 8323 34336 8332 34376
rect 8372 34336 8524 34376
rect 8564 34336 8573 34376
rect 8995 34336 9004 34376
rect 9044 34336 9100 34376
rect 9140 34336 9149 34376
rect 10051 34336 10060 34376
rect 10100 34336 10732 34376
rect 10772 34336 11596 34376
rect 11636 34336 11645 34376
rect 12451 34336 12460 34376
rect 12500 34336 13708 34376
rect 13748 34336 13757 34376
rect 0 34316 80 34336
rect 1612 34292 1652 34336
rect 2179 34335 2237 34336
rect 6019 34335 6077 34336
rect 8323 34335 8381 34336
rect 9091 34335 9149 34336
rect 3907 34292 3965 34293
rect 14572 34292 14612 34420
rect 1612 34252 2956 34292
rect 2996 34252 3005 34292
rect 3822 34252 3916 34292
rect 3956 34252 3965 34292
rect 6019 34252 6028 34292
rect 6068 34252 6796 34292
rect 6836 34252 6845 34292
rect 7267 34252 7276 34292
rect 7316 34252 7948 34292
rect 7988 34252 7997 34292
rect 14380 34252 14612 34292
rect 3907 34251 3965 34252
rect 4387 34208 4445 34209
rect 12643 34208 12701 34209
rect 14380 34208 14420 34252
rect 21424 34208 21504 34228
rect 2500 34168 2668 34208
rect 2708 34168 3244 34208
rect 3284 34168 3293 34208
rect 4302 34168 4396 34208
rect 4436 34168 4445 34208
rect 5059 34168 5068 34208
rect 5108 34168 6316 34208
rect 6356 34168 6365 34208
rect 6595 34168 6604 34208
rect 6644 34168 10156 34208
rect 10196 34168 10205 34208
rect 12643 34168 12652 34208
rect 12692 34168 12844 34208
rect 12884 34168 12893 34208
rect 13507 34168 13516 34208
rect 13556 34168 13804 34208
rect 13844 34168 13853 34208
rect 14371 34168 14380 34208
rect 14420 34168 14429 34208
rect 14563 34168 14572 34208
rect 14612 34168 14621 34208
rect 19843 34168 19852 34208
rect 19892 34168 21504 34208
rect 2500 34124 2540 34168
rect 4387 34167 4445 34168
rect 12643 34167 12701 34168
rect 14572 34124 14612 34168
rect 21424 34148 21504 34168
rect 259 34084 268 34124
rect 308 34084 2540 34124
rect 8803 34084 8812 34124
rect 8852 34084 9580 34124
rect 9620 34084 9629 34124
rect 10915 34084 10924 34124
rect 10964 34084 11692 34124
rect 11732 34084 11741 34124
rect 11875 34084 11884 34124
rect 11924 34084 12940 34124
rect 12980 34084 14612 34124
rect 0 34040 80 34060
rect 13603 34040 13661 34041
rect 13900 34040 13940 34084
rect 19363 34040 19421 34041
rect 0 34000 1132 34040
rect 1172 34000 1181 34040
rect 4919 34000 4928 34040
rect 4968 34000 5010 34040
rect 5050 34000 5092 34040
rect 5132 34000 5174 34040
rect 5214 34000 5256 34040
rect 5296 34000 5305 34040
rect 6211 34000 6220 34040
rect 6260 34000 6269 34040
rect 6499 34000 6508 34040
rect 6548 34000 7756 34040
rect 7796 34000 7805 34040
rect 12259 34000 12268 34040
rect 12308 34000 12748 34040
rect 12788 34000 12797 34040
rect 13603 34000 13612 34040
rect 13652 34000 13708 34040
rect 13748 34000 13757 34040
rect 13891 34000 13900 34040
rect 13940 34000 13949 34040
rect 13994 34000 14003 34040
rect 14043 34000 14052 34040
rect 14755 34000 14764 34040
rect 14804 34000 14956 34040
rect 14996 34000 15005 34040
rect 19278 34000 19372 34040
rect 19412 34000 19421 34040
rect 20039 34000 20048 34040
rect 20088 34000 20130 34040
rect 20170 34000 20212 34040
rect 20252 34000 20294 34040
rect 20334 34000 20376 34040
rect 20416 34000 20425 34040
rect 0 33980 80 34000
rect 6220 33956 6260 34000
rect 13603 33999 13661 34000
rect 7747 33956 7805 33957
rect 13996 33956 14036 34000
rect 19363 33999 19421 34000
rect 3139 33916 3148 33956
rect 3188 33916 3724 33956
rect 3764 33916 3773 33956
rect 5635 33916 5644 33956
rect 5684 33916 5932 33956
rect 5972 33916 6260 33956
rect 7075 33916 7084 33956
rect 7124 33916 7276 33956
rect 7316 33916 7325 33956
rect 7555 33916 7564 33956
rect 7604 33916 7756 33956
rect 7796 33916 8332 33956
rect 8372 33916 8381 33956
rect 11683 33916 11692 33956
rect 11732 33916 14036 33956
rect 7747 33915 7805 33916
rect 2851 33832 2860 33872
rect 2900 33832 3476 33872
rect 6211 33832 6220 33872
rect 6260 33832 7468 33872
rect 7508 33832 7517 33872
rect 9763 33832 9772 33872
rect 9812 33832 9964 33872
rect 10004 33832 10013 33872
rect 11203 33832 11212 33872
rect 11252 33832 11788 33872
rect 11828 33832 11837 33872
rect 12739 33832 12748 33872
rect 12788 33832 13420 33872
rect 13460 33832 13469 33872
rect 3436 33788 3476 33832
rect 1708 33748 2572 33788
rect 2612 33748 2621 33788
rect 3427 33748 3436 33788
rect 3476 33748 3485 33788
rect 5635 33748 5644 33788
rect 5684 33748 7508 33788
rect 0 33704 80 33724
rect 1708 33704 1748 33748
rect 7468 33704 7508 33748
rect 0 33664 1652 33704
rect 1699 33664 1708 33704
rect 1748 33664 1757 33704
rect 2467 33664 2476 33704
rect 2516 33664 2956 33704
rect 2996 33664 3340 33704
rect 3380 33664 3389 33704
rect 6115 33664 6124 33704
rect 6164 33664 6604 33704
rect 6644 33664 7276 33704
rect 7316 33664 7325 33704
rect 7459 33664 7468 33704
rect 7508 33664 7517 33704
rect 8227 33664 8236 33704
rect 8276 33664 8716 33704
rect 8756 33664 9580 33704
rect 9620 33664 11212 33704
rect 11252 33664 11261 33704
rect 11395 33664 11404 33704
rect 11444 33664 11884 33704
rect 11924 33664 12076 33704
rect 12116 33664 12125 33704
rect 13411 33664 13420 33704
rect 13460 33664 13612 33704
rect 13652 33664 13661 33704
rect 14467 33664 14476 33704
rect 14516 33664 14668 33704
rect 14708 33664 14717 33704
rect 15715 33664 15724 33704
rect 15764 33664 16204 33704
rect 16244 33664 16253 33704
rect 0 33644 80 33664
rect 1612 33620 1652 33664
rect 4387 33620 4445 33621
rect 10531 33620 10589 33621
rect 1612 33580 2188 33620
rect 2228 33580 2237 33620
rect 4387 33580 4396 33620
rect 4436 33580 6028 33620
rect 6068 33580 6077 33620
rect 6883 33580 6892 33620
rect 6932 33580 10348 33620
rect 10388 33580 10397 33620
rect 10531 33580 10540 33620
rect 10580 33580 20180 33620
rect 4387 33579 4445 33580
rect 10531 33579 10589 33580
rect 20140 33536 20180 33580
rect 21424 33536 21504 33556
rect 4195 33496 4204 33536
rect 4244 33496 16012 33536
rect 16052 33496 16492 33536
rect 16532 33496 18316 33536
rect 18356 33496 18365 33536
rect 20140 33496 21504 33536
rect 21424 33476 21504 33496
rect 7267 33412 7276 33452
rect 7316 33412 7564 33452
rect 7604 33412 7613 33452
rect 12163 33412 12172 33452
rect 12212 33412 12556 33452
rect 12596 33412 12605 33452
rect 13507 33412 13516 33452
rect 13556 33412 13900 33452
rect 13940 33412 14092 33452
rect 14132 33412 14141 33452
rect 0 33368 80 33388
rect 0 33328 4684 33368
rect 4724 33328 11692 33368
rect 11732 33328 16108 33368
rect 16148 33328 18220 33368
rect 18260 33328 18700 33368
rect 18740 33328 18749 33368
rect 0 33308 80 33328
rect 8227 33284 8285 33285
rect 3679 33244 3688 33284
rect 3728 33244 3770 33284
rect 3810 33244 3852 33284
rect 3892 33244 3934 33284
rect 3974 33244 4016 33284
rect 4056 33244 4065 33284
rect 7363 33244 7372 33284
rect 7412 33244 8236 33284
rect 8276 33244 8285 33284
rect 8227 33243 8285 33244
rect 12067 33284 12125 33285
rect 12067 33244 12076 33284
rect 12116 33244 12172 33284
rect 12212 33244 12221 33284
rect 13507 33244 13516 33284
rect 13556 33244 13996 33284
rect 14036 33244 14045 33284
rect 18799 33244 18808 33284
rect 18848 33244 18890 33284
rect 18930 33244 18972 33284
rect 19012 33244 19054 33284
rect 19094 33244 19136 33284
rect 19176 33244 19185 33284
rect 12067 33243 12125 33244
rect 1411 33200 1469 33201
rect 7555 33200 7613 33201
rect 1325 33160 1420 33200
rect 1460 33160 6124 33200
rect 6164 33160 7564 33200
rect 7604 33160 7613 33200
rect 7939 33160 7948 33200
rect 7988 33160 8332 33200
rect 8372 33160 8381 33200
rect 9955 33160 9964 33200
rect 10004 33160 11360 33200
rect 1411 33159 1469 33160
rect 7555 33159 7613 33160
rect 11320 33116 11360 33160
rect 2179 33076 2188 33116
rect 2228 33076 4724 33116
rect 7075 33076 7084 33116
rect 7124 33076 8524 33116
rect 8564 33076 10444 33116
rect 10484 33076 10493 33116
rect 11320 33076 13996 33116
rect 14036 33076 14045 33116
rect 0 33032 80 33052
rect 4684 33032 4724 33076
rect 0 32992 4204 33032
rect 4244 32992 4253 33032
rect 4684 32992 13364 33032
rect 13411 32992 13420 33032
rect 13460 32992 14188 33032
rect 14228 32992 14237 33032
rect 0 32972 80 32992
rect 13324 32948 13364 32992
rect 7171 32908 7180 32948
rect 7220 32908 7660 32948
rect 7700 32908 7709 32948
rect 8035 32908 8044 32948
rect 8084 32908 8428 32948
rect 8468 32908 8477 32948
rect 13324 32908 16204 32948
rect 16244 32908 16253 32948
rect 19363 32864 19421 32865
rect 163 32824 172 32864
rect 212 32824 2092 32864
rect 2132 32824 2764 32864
rect 2804 32824 2813 32864
rect 2956 32824 3340 32864
rect 3380 32824 3389 32864
rect 6691 32824 6700 32864
rect 6740 32824 7988 32864
rect 12067 32824 12076 32864
rect 12116 32824 13228 32864
rect 13268 32824 13277 32864
rect 13987 32824 13996 32864
rect 14036 32824 19372 32864
rect 19412 32824 19421 32864
rect 2956 32780 2996 32824
rect 3235 32780 3293 32781
rect 5347 32780 5405 32781
rect 7948 32780 7988 32824
rect 19363 32823 19421 32824
rect 19939 32864 19997 32865
rect 21424 32864 21504 32884
rect 19939 32824 19948 32864
rect 19988 32824 21504 32864
rect 19939 32823 19997 32824
rect 21424 32804 21504 32824
rect 2851 32740 2860 32780
rect 2900 32740 2996 32780
rect 3043 32740 3052 32780
rect 3092 32740 3244 32780
rect 3284 32740 3532 32780
rect 3572 32740 3724 32780
rect 3764 32740 3773 32780
rect 4387 32740 4396 32780
rect 4436 32740 5356 32780
rect 5396 32740 5405 32780
rect 7940 32740 7949 32780
rect 7989 32740 7998 32780
rect 12268 32740 13132 32780
rect 13172 32740 13181 32780
rect 3235 32739 3293 32740
rect 5347 32739 5405 32740
rect 0 32696 80 32716
rect 7651 32696 7709 32697
rect 12268 32696 12308 32740
rect 13219 32696 13277 32697
rect 0 32656 2284 32696
rect 2324 32656 2333 32696
rect 3235 32656 3244 32696
rect 3284 32656 6796 32696
rect 6836 32656 6845 32696
rect 7555 32656 7564 32696
rect 7604 32656 7660 32696
rect 7700 32656 7756 32696
rect 7796 32656 7824 32696
rect 12259 32656 12268 32696
rect 12308 32656 12317 32696
rect 13219 32656 13228 32696
rect 13268 32656 14764 32696
rect 14804 32656 16588 32696
rect 16628 32656 17452 32696
rect 17492 32656 17501 32696
rect 0 32636 80 32656
rect 7651 32655 7709 32656
rect 13219 32655 13277 32656
rect 6211 32572 6220 32612
rect 6260 32572 7852 32612
rect 7892 32572 7901 32612
rect 7747 32528 7805 32529
rect 4919 32488 4928 32528
rect 4968 32488 5010 32528
rect 5050 32488 5092 32528
rect 5132 32488 5174 32528
rect 5214 32488 5256 32528
rect 5296 32488 5305 32528
rect 7662 32488 7756 32528
rect 7796 32488 7805 32528
rect 20039 32488 20048 32528
rect 20088 32488 20130 32528
rect 20170 32488 20212 32528
rect 20252 32488 20294 32528
rect 20334 32488 20376 32528
rect 20416 32488 20425 32528
rect 7747 32487 7805 32488
rect 5539 32404 5548 32444
rect 5588 32404 5836 32444
rect 5876 32404 6508 32444
rect 6548 32404 8236 32444
rect 8276 32404 8285 32444
rect 0 32360 80 32380
rect 15715 32360 15773 32361
rect 0 32320 4396 32360
rect 4436 32320 9964 32360
rect 10004 32320 10013 32360
rect 11203 32320 11212 32360
rect 11252 32320 12076 32360
rect 12116 32320 12460 32360
rect 12500 32320 12509 32360
rect 15331 32320 15340 32360
rect 15380 32320 15724 32360
rect 15764 32320 16300 32360
rect 16340 32320 16349 32360
rect 0 32300 80 32320
rect 15715 32319 15773 32320
rect 6019 32276 6077 32277
rect 5923 32236 5932 32276
rect 5972 32236 6028 32276
rect 6068 32236 6077 32276
rect 7555 32236 7564 32276
rect 7604 32236 8332 32276
rect 8372 32236 8381 32276
rect 12643 32236 12652 32276
rect 12692 32236 13516 32276
rect 13556 32236 19660 32276
rect 19700 32236 19709 32276
rect 6019 32235 6077 32236
rect 7459 32192 7517 32193
rect 16963 32192 17021 32193
rect 21424 32192 21504 32212
rect 7459 32152 7468 32192
rect 7508 32152 7660 32192
rect 7700 32152 7709 32192
rect 7843 32152 7852 32192
rect 7892 32152 8716 32192
rect 8756 32152 8765 32192
rect 12355 32152 12364 32192
rect 12404 32152 12844 32192
rect 12884 32152 12893 32192
rect 13027 32152 13036 32192
rect 13076 32152 13085 32192
rect 13411 32152 13420 32192
rect 13460 32152 14380 32192
rect 14420 32152 14429 32192
rect 14659 32152 14668 32192
rect 14708 32152 14717 32192
rect 15139 32152 15148 32192
rect 15188 32152 15436 32192
rect 15476 32152 15820 32192
rect 15860 32152 15869 32192
rect 16963 32152 16972 32192
rect 17012 32152 21504 32192
rect 7459 32151 7517 32152
rect 6787 32108 6845 32109
rect 6403 32068 6412 32108
rect 6452 32068 6796 32108
rect 6836 32068 6845 32108
rect 6787 32067 6845 32068
rect 0 32024 80 32044
rect 7651 32024 7709 32025
rect 13036 32024 13076 32152
rect 14668 32108 14708 32152
rect 16963 32151 17021 32152
rect 21424 32132 21504 32152
rect 14668 32068 15916 32108
rect 15956 32068 15965 32108
rect 0 31984 3244 32024
rect 3284 31984 3293 32024
rect 4195 31984 4204 32024
rect 4244 31984 4492 32024
rect 4532 31984 4541 32024
rect 7363 31984 7372 32024
rect 7412 31984 7660 32024
rect 7700 31984 7709 32024
rect 11011 31984 11020 32024
rect 11060 31984 13076 32024
rect 14659 31984 14668 32024
rect 14708 31984 14860 32024
rect 14900 31984 14909 32024
rect 0 31964 80 31984
rect 7651 31983 7709 31984
rect 4099 31940 4157 31941
rect 3715 31900 3724 31940
rect 3764 31900 4108 31940
rect 4148 31900 4157 31940
rect 16099 31900 16108 31940
rect 16148 31900 16780 31940
rect 16820 31900 16829 31940
rect 4099 31899 4157 31900
rect 2467 31856 2525 31857
rect 2381 31816 2476 31856
rect 2516 31816 6892 31856
rect 6932 31816 6941 31856
rect 14563 31816 14572 31856
rect 14612 31816 14860 31856
rect 14900 31816 14909 31856
rect 2467 31815 2525 31816
rect 3679 31732 3688 31772
rect 3728 31732 3770 31772
rect 3810 31732 3852 31772
rect 3892 31732 3934 31772
rect 3974 31732 4016 31772
rect 4056 31732 4065 31772
rect 4291 31732 4300 31772
rect 4340 31732 5932 31772
rect 5972 31732 5981 31772
rect 6892 31732 14188 31772
rect 14228 31732 14237 31772
rect 18799 31732 18808 31772
rect 18848 31732 18890 31772
rect 18930 31732 18972 31772
rect 19012 31732 19054 31772
rect 19094 31732 19136 31772
rect 19176 31732 19185 31772
rect 0 31688 80 31708
rect 6892 31688 6932 31732
rect 0 31648 6932 31688
rect 10339 31688 10397 31689
rect 10339 31648 10348 31688
rect 10388 31648 21332 31688
rect 0 31628 80 31648
rect 10339 31647 10397 31648
rect 8995 31604 9053 31605
rect 11587 31604 11645 31605
rect 739 31564 748 31604
rect 788 31564 6316 31604
rect 6356 31564 6365 31604
rect 6883 31564 6892 31604
rect 6932 31564 9004 31604
rect 9044 31564 9196 31604
rect 9236 31564 9245 31604
rect 11491 31564 11500 31604
rect 11540 31564 11596 31604
rect 11636 31564 11884 31604
rect 11924 31564 11933 31604
rect 12931 31564 12940 31604
rect 12980 31564 13228 31604
rect 13268 31564 13277 31604
rect 14371 31564 14380 31604
rect 14420 31564 19276 31604
rect 19316 31564 19325 31604
rect 8995 31563 9053 31564
rect 11587 31563 11645 31564
rect 2179 31520 2237 31521
rect 15331 31520 15389 31521
rect 2179 31480 2188 31520
rect 2228 31480 2668 31520
rect 2708 31480 2717 31520
rect 2851 31480 2860 31520
rect 2900 31480 2909 31520
rect 3043 31480 3052 31520
rect 3092 31480 3436 31520
rect 3476 31480 5068 31520
rect 5108 31480 5117 31520
rect 5347 31480 5356 31520
rect 5396 31480 5405 31520
rect 11395 31480 11404 31520
rect 11444 31480 12748 31520
rect 12788 31480 12797 31520
rect 14467 31480 14476 31520
rect 14516 31480 14956 31520
rect 14996 31480 15005 31520
rect 15235 31480 15244 31520
rect 15284 31480 15340 31520
rect 15380 31480 15389 31520
rect 21292 31520 21332 31648
rect 21424 31520 21504 31540
rect 21292 31480 21504 31520
rect 2179 31479 2237 31480
rect 2860 31436 2900 31480
rect 5356 31436 5396 31480
rect 15331 31479 15389 31480
rect 21424 31460 21504 31480
rect 14371 31436 14429 31437
rect 16675 31436 16733 31437
rect 2371 31396 2380 31436
rect 2420 31396 2900 31436
rect 3715 31396 3724 31436
rect 3764 31396 4780 31436
rect 4820 31396 4829 31436
rect 5356 31396 7276 31436
rect 7316 31396 8140 31436
rect 8180 31396 8189 31436
rect 8323 31396 8332 31436
rect 8372 31396 9292 31436
rect 9332 31396 10636 31436
rect 10676 31396 10685 31436
rect 10732 31396 13556 31436
rect 0 31352 80 31372
rect 10732 31352 10772 31396
rect 11395 31352 11453 31353
rect 12259 31352 12317 31353
rect 13516 31352 13556 31396
rect 14371 31396 14380 31436
rect 14420 31396 16684 31436
rect 16724 31396 16733 31436
rect 14371 31395 14429 31396
rect 16675 31395 16733 31396
rect 0 31312 1268 31352
rect 1987 31312 1996 31352
rect 2036 31312 2860 31352
rect 2900 31312 2909 31352
rect 3043 31312 3052 31352
rect 3092 31312 5356 31352
rect 5396 31312 5548 31352
rect 5588 31312 5597 31352
rect 6691 31312 6700 31352
rect 6740 31312 8236 31352
rect 8276 31312 9868 31352
rect 9908 31312 9917 31352
rect 10444 31312 10772 31352
rect 11203 31312 11212 31352
rect 11252 31312 11404 31352
rect 11444 31312 12268 31352
rect 12308 31312 12317 31352
rect 13507 31312 13516 31352
rect 13556 31312 13565 31352
rect 17731 31312 17740 31352
rect 17780 31312 19468 31352
rect 19508 31312 19517 31352
rect 0 31292 80 31312
rect 1228 31268 1268 31312
rect 9955 31268 10013 31269
rect 1228 31228 9964 31268
rect 10004 31228 10013 31268
rect 9955 31227 10013 31228
rect 10444 31184 10484 31312
rect 11395 31311 11453 31312
rect 12259 31311 12317 31312
rect 15427 31268 15485 31269
rect 10627 31228 10636 31268
rect 10676 31228 10685 31268
rect 15331 31228 15340 31268
rect 15380 31228 15436 31268
rect 15476 31228 15485 31268
rect 17827 31228 17836 31268
rect 17876 31228 18412 31268
rect 18452 31228 18461 31268
rect 2947 31144 2956 31184
rect 2996 31144 3916 31184
rect 3956 31144 3965 31184
rect 4675 31144 4684 31184
rect 4724 31144 4972 31184
rect 5012 31144 5021 31184
rect 7075 31144 7084 31184
rect 7124 31144 7276 31184
rect 7316 31144 7325 31184
rect 8035 31144 8044 31184
rect 8084 31144 10484 31184
rect 10636 31184 10676 31228
rect 15427 31227 15485 31228
rect 19939 31184 19997 31185
rect 10636 31144 11308 31184
rect 11348 31144 11357 31184
rect 12931 31144 12940 31184
rect 12980 31144 13228 31184
rect 13268 31144 13277 31184
rect 15235 31144 15244 31184
rect 15284 31144 16108 31184
rect 16148 31144 16157 31184
rect 19939 31144 19948 31184
rect 19988 31144 20044 31184
rect 20084 31144 20093 31184
rect 19939 31143 19997 31144
rect 9475 31100 9533 31101
rect 2467 31060 2476 31100
rect 2516 31060 3628 31100
rect 3668 31060 3677 31100
rect 9379 31060 9388 31100
rect 9428 31060 9484 31100
rect 9524 31060 9533 31100
rect 12739 31060 12748 31100
rect 12788 31060 13324 31100
rect 13364 31060 13373 31100
rect 14563 31060 14572 31100
rect 14612 31060 16204 31100
rect 16244 31060 16253 31100
rect 9475 31059 9533 31060
rect 0 31016 80 31036
rect 8803 31016 8861 31017
rect 11107 31016 11165 31017
rect 18691 31016 18749 31017
rect 0 30976 1556 31016
rect 3331 30976 3340 31016
rect 3380 30976 3724 31016
rect 3764 30976 3773 31016
rect 4919 30976 4928 31016
rect 4968 30976 5010 31016
rect 5050 30976 5092 31016
rect 5132 30976 5174 31016
rect 5214 30976 5256 31016
rect 5296 30976 5305 31016
rect 8718 30976 8812 31016
rect 8852 30976 8861 31016
rect 9187 30976 9196 31016
rect 9236 30976 9964 31016
rect 10004 30976 10013 31016
rect 10531 30976 10540 31016
rect 10580 30976 11116 31016
rect 11156 30976 11165 31016
rect 16579 30976 16588 31016
rect 16628 30976 18700 31016
rect 18740 30976 18749 31016
rect 19267 30976 19276 31016
rect 19316 30976 19948 31016
rect 19988 30976 19997 31016
rect 20039 30976 20048 31016
rect 20088 30976 20130 31016
rect 20170 30976 20212 31016
rect 20252 30976 20294 31016
rect 20334 30976 20376 31016
rect 20416 30976 20425 31016
rect 0 30956 80 30976
rect 0 30680 80 30700
rect 0 30640 1420 30680
rect 1460 30640 1469 30680
rect 0 30620 80 30640
rect 1516 30428 1556 30976
rect 8803 30975 8861 30976
rect 11107 30975 11165 30976
rect 18691 30975 18749 30976
rect 1699 30892 1708 30932
rect 1748 30892 3244 30932
rect 3284 30892 3293 30932
rect 5827 30892 5836 30932
rect 5876 30892 9676 30932
rect 9716 30892 9725 30932
rect 10339 30892 10348 30932
rect 10388 30892 11212 30932
rect 11252 30892 11261 30932
rect 12163 30892 12172 30932
rect 12212 30892 18796 30932
rect 18836 30892 18845 30932
rect 2179 30848 2237 30849
rect 5836 30848 5876 30892
rect 1891 30808 1900 30848
rect 1940 30808 2036 30848
rect 2083 30808 2092 30848
rect 2132 30808 2188 30848
rect 2228 30808 2237 30848
rect 3811 30808 3820 30848
rect 3860 30808 4492 30848
rect 4532 30808 4541 30848
rect 5059 30808 5068 30848
rect 5108 30808 5876 30848
rect 6979 30848 7037 30849
rect 21424 30848 21504 30868
rect 6979 30808 6988 30848
rect 7028 30808 21504 30848
rect 1996 30596 2036 30808
rect 2179 30807 2237 30808
rect 6979 30807 7037 30808
rect 21424 30788 21504 30808
rect 5827 30764 5885 30765
rect 11779 30764 11837 30765
rect 2500 30724 2764 30764
rect 2804 30724 3148 30764
rect 3188 30724 3197 30764
rect 4579 30724 4588 30764
rect 4628 30724 4637 30764
rect 5742 30724 5836 30764
rect 5876 30724 5885 30764
rect 9379 30724 9388 30764
rect 9428 30724 9676 30764
rect 9716 30724 9725 30764
rect 10435 30724 10444 30764
rect 10484 30724 11212 30764
rect 11252 30724 11261 30764
rect 11779 30724 11788 30764
rect 11828 30724 11980 30764
rect 12020 30724 12460 30764
rect 12500 30724 12509 30764
rect 13219 30724 13228 30764
rect 13268 30724 13420 30764
rect 13460 30724 13469 30764
rect 14668 30724 17740 30764
rect 17780 30724 17789 30764
rect 2500 30680 2540 30724
rect 4588 30680 4628 30724
rect 5827 30723 5885 30724
rect 11779 30723 11837 30724
rect 12355 30680 12413 30681
rect 2179 30640 2188 30680
rect 2228 30640 2540 30680
rect 3043 30640 3052 30680
rect 3092 30640 4204 30680
rect 4244 30640 4628 30680
rect 6115 30640 6124 30680
rect 6164 30640 7220 30680
rect 8515 30640 8524 30680
rect 8564 30640 8812 30680
rect 8852 30640 9484 30680
rect 9524 30640 10828 30680
rect 10868 30640 10877 30680
rect 12270 30640 12364 30680
rect 12404 30640 12413 30680
rect 13795 30640 13804 30680
rect 13844 30640 14572 30680
rect 14612 30640 14621 30680
rect 1987 30556 1996 30596
rect 2036 30556 2045 30596
rect 2947 30556 2956 30596
rect 2996 30556 7084 30596
rect 7124 30556 7133 30596
rect 2083 30472 2092 30512
rect 2132 30472 2476 30512
rect 2516 30472 3340 30512
rect 3380 30472 3389 30512
rect 3619 30472 3628 30512
rect 3668 30472 5836 30512
rect 5876 30472 5885 30512
rect 7084 30428 7124 30556
rect 7180 30512 7220 30640
rect 12355 30639 12413 30640
rect 14668 30596 14708 30724
rect 14755 30640 14764 30680
rect 14804 30640 15148 30680
rect 15188 30640 18604 30680
rect 18644 30640 18653 30680
rect 19939 30640 19948 30680
rect 19988 30640 20236 30680
rect 20276 30640 20285 30680
rect 10339 30556 10348 30596
rect 10388 30556 10732 30596
rect 10772 30556 10781 30596
rect 11299 30556 11308 30596
rect 11348 30556 14708 30596
rect 15235 30556 15244 30596
rect 15284 30556 15628 30596
rect 15668 30556 15677 30596
rect 7180 30472 8620 30512
rect 8660 30472 8812 30512
rect 8852 30472 8861 30512
rect 10915 30472 10924 30512
rect 10964 30472 11500 30512
rect 11540 30472 11549 30512
rect 12739 30472 12748 30512
rect 12788 30472 13132 30512
rect 13172 30472 13181 30512
rect 15043 30472 15052 30512
rect 15092 30472 15724 30512
rect 15764 30472 16588 30512
rect 16628 30472 16637 30512
rect 18019 30472 18028 30512
rect 18068 30472 18700 30512
rect 18740 30472 18749 30512
rect 19267 30472 19276 30512
rect 19316 30472 20620 30512
rect 20660 30472 20669 30512
rect 15715 30428 15773 30429
rect 1516 30388 2860 30428
rect 2900 30388 4588 30428
rect 4628 30388 4637 30428
rect 7084 30388 15724 30428
rect 15764 30388 15773 30428
rect 19075 30388 19084 30428
rect 19124 30388 20524 30428
rect 20564 30388 20573 30428
rect 15715 30387 15773 30388
rect 0 30344 80 30364
rect 3139 30344 3197 30345
rect 8803 30344 8861 30345
rect 9475 30344 9533 30345
rect 0 30304 3148 30344
rect 3188 30304 3197 30344
rect 0 30284 80 30304
rect 3139 30303 3197 30304
rect 3532 30304 5068 30344
rect 5108 30304 5117 30344
rect 8803 30304 8812 30344
rect 8852 30304 8908 30344
rect 8948 30304 8957 30344
rect 9379 30304 9388 30344
rect 9428 30304 9484 30344
rect 9524 30304 9533 30344
rect 17923 30304 17932 30344
rect 17972 30304 17981 30344
rect 3532 30260 3572 30304
rect 8803 30303 8861 30304
rect 9475 30303 9533 30304
rect 17932 30260 17972 30304
rect 19939 30260 19997 30261
rect 1411 30220 1420 30260
rect 1460 30220 1708 30260
rect 1748 30220 3572 30260
rect 3679 30220 3688 30260
rect 3728 30220 3770 30260
rect 3810 30220 3852 30260
rect 3892 30220 3934 30260
rect 3974 30220 4016 30260
rect 4056 30220 4065 30260
rect 5443 30220 5452 30260
rect 5492 30220 6412 30260
rect 6452 30220 6461 30260
rect 6979 30220 6988 30260
rect 7028 30220 9004 30260
rect 9044 30220 9053 30260
rect 14659 30220 14668 30260
rect 14708 30220 15820 30260
rect 15860 30220 15869 30260
rect 16195 30220 16204 30260
rect 16244 30220 17644 30260
rect 17684 30220 17693 30260
rect 17932 30220 18412 30260
rect 18452 30220 18461 30260
rect 18799 30220 18808 30260
rect 18848 30220 18890 30260
rect 18930 30220 18972 30260
rect 19012 30220 19054 30260
rect 19094 30220 19136 30260
rect 19176 30220 19185 30260
rect 19651 30220 19660 30260
rect 19700 30220 19948 30260
rect 19988 30220 19997 30260
rect 19939 30219 19997 30220
rect 2179 30176 2237 30177
rect 21424 30176 21504 30196
rect 2094 30136 2188 30176
rect 2228 30136 2237 30176
rect 2179 30135 2237 30136
rect 2500 30136 10924 30176
rect 10964 30136 10973 30176
rect 11320 30136 21504 30176
rect 1603 30092 1661 30093
rect 1987 30092 2045 30093
rect 2500 30092 2540 30136
rect 9763 30092 9821 30093
rect 11320 30092 11360 30136
rect 21424 30116 21504 30136
rect 15331 30092 15389 30093
rect 1603 30052 1612 30092
rect 1652 30052 1996 30092
rect 2036 30052 2540 30092
rect 4387 30052 4396 30092
rect 4436 30052 5644 30092
rect 5684 30052 5693 30092
rect 9763 30052 9772 30092
rect 9812 30052 11360 30092
rect 13699 30052 13708 30092
rect 13748 30052 14668 30092
rect 14708 30052 14717 30092
rect 15331 30052 15340 30092
rect 15380 30052 15724 30092
rect 15764 30052 15773 30092
rect 17347 30052 17356 30092
rect 17396 30052 20180 30092
rect 1603 30051 1661 30052
rect 1987 30051 2045 30052
rect 9763 30051 9821 30052
rect 15331 30051 15389 30052
rect 0 30008 80 30028
rect 20140 30008 20180 30052
rect 0 29968 2540 30008
rect 9187 29968 9196 30008
rect 9236 29968 10444 30008
rect 10484 29968 10493 30008
rect 11107 29968 11116 30008
rect 11156 29968 11596 30008
rect 11636 29968 11645 30008
rect 15235 29968 15244 30008
rect 15284 29968 19468 30008
rect 19508 29968 19852 30008
rect 19892 29968 19901 30008
rect 20140 29968 21388 30008
rect 21428 29968 21437 30008
rect 0 29948 80 29968
rect 2500 29924 2540 29968
rect 2500 29884 12460 29924
rect 12500 29884 12509 29924
rect 16675 29884 16684 29924
rect 16724 29884 18124 29924
rect 18164 29884 18316 29924
rect 18356 29884 18365 29924
rect 4099 29840 4157 29841
rect 1123 29800 1132 29840
rect 1172 29800 2956 29840
rect 2996 29800 3005 29840
rect 3619 29800 3628 29840
rect 3668 29800 4108 29840
rect 4148 29800 4204 29840
rect 4244 29800 5548 29840
rect 5588 29800 6124 29840
rect 6164 29800 6173 29840
rect 6403 29800 6412 29840
rect 6452 29800 8332 29840
rect 8372 29800 8381 29840
rect 9187 29800 9196 29840
rect 9236 29800 10540 29840
rect 10580 29800 10589 29840
rect 10915 29800 10924 29840
rect 10964 29800 13900 29840
rect 13940 29800 13949 29840
rect 14467 29800 14476 29840
rect 14516 29800 14764 29840
rect 14804 29800 14813 29840
rect 15619 29800 15628 29840
rect 15668 29800 15916 29840
rect 15956 29800 15965 29840
rect 17539 29800 17548 29840
rect 17588 29800 18412 29840
rect 18452 29800 19564 29840
rect 19604 29800 19613 29840
rect 4099 29799 4157 29800
rect 11299 29756 11357 29757
rect 14476 29756 14516 29800
rect 2083 29716 2092 29756
rect 2132 29716 5356 29756
rect 5396 29716 5405 29756
rect 8707 29716 8716 29756
rect 8756 29716 11308 29756
rect 11348 29716 11357 29756
rect 13123 29716 13132 29756
rect 13172 29716 14516 29756
rect 15331 29716 15340 29756
rect 15380 29716 19948 29756
rect 19988 29716 19997 29756
rect 11299 29715 11357 29716
rect 0 29672 80 29692
rect 8227 29672 8285 29673
rect 10243 29672 10301 29673
rect 13123 29672 13181 29673
rect 15820 29672 15860 29716
rect 0 29632 3436 29672
rect 3476 29632 3485 29672
rect 8227 29632 8236 29672
rect 8276 29632 9484 29672
rect 9524 29632 9868 29672
rect 9908 29632 9917 29672
rect 10243 29632 10252 29672
rect 10292 29632 10540 29672
rect 10580 29632 10589 29672
rect 11875 29632 11884 29672
rect 11924 29632 12364 29672
rect 12404 29632 12413 29672
rect 13027 29632 13036 29672
rect 13076 29632 13132 29672
rect 13172 29632 13181 29672
rect 15811 29632 15820 29672
rect 15860 29632 15900 29672
rect 18115 29632 18124 29672
rect 18164 29632 18173 29672
rect 19075 29632 19084 29672
rect 19124 29632 20044 29672
rect 20084 29632 20093 29672
rect 0 29612 80 29632
rect 8227 29631 8285 29632
rect 10243 29631 10301 29632
rect 13123 29631 13181 29632
rect 18124 29588 18164 29632
rect 2947 29548 2956 29588
rect 2996 29548 14380 29588
rect 14420 29548 14429 29588
rect 15235 29548 15244 29588
rect 15284 29548 16300 29588
rect 16340 29548 18164 29588
rect 4919 29464 4928 29504
rect 4968 29464 5010 29504
rect 5050 29464 5092 29504
rect 5132 29464 5174 29504
rect 5214 29464 5256 29504
rect 5296 29464 5305 29504
rect 5827 29464 5836 29504
rect 5876 29464 8812 29504
rect 8852 29464 11116 29504
rect 11156 29464 11165 29504
rect 11587 29464 11596 29504
rect 11636 29464 12172 29504
rect 12212 29464 13132 29504
rect 13172 29464 13181 29504
rect 17731 29464 17740 29504
rect 17780 29464 18604 29504
rect 18644 29464 19564 29504
rect 19604 29464 19613 29504
rect 4588 29380 6316 29420
rect 6356 29380 6365 29420
rect 10243 29380 10252 29420
rect 10292 29380 10540 29420
rect 10580 29380 10589 29420
rect 16483 29380 16492 29420
rect 16532 29380 17644 29420
rect 17684 29380 17693 29420
rect 0 29336 80 29356
rect 4588 29336 4628 29380
rect 15235 29336 15293 29337
rect 17059 29336 17117 29337
rect 19948 29336 19988 29632
rect 20803 29504 20861 29505
rect 21424 29504 21504 29524
rect 20039 29464 20048 29504
rect 20088 29464 20130 29504
rect 20170 29464 20212 29504
rect 20252 29464 20294 29504
rect 20334 29464 20376 29504
rect 20416 29464 20425 29504
rect 20803 29464 20812 29504
rect 20852 29464 21504 29504
rect 20803 29463 20861 29464
rect 21424 29444 21504 29464
rect 0 29296 4628 29336
rect 4675 29296 4684 29336
rect 4724 29296 7948 29336
rect 7988 29296 7997 29336
rect 9955 29296 9964 29336
rect 10004 29296 10636 29336
rect 10676 29296 10685 29336
rect 11971 29296 11980 29336
rect 12020 29296 12172 29336
rect 12212 29296 12221 29336
rect 13603 29296 13612 29336
rect 13652 29296 15244 29336
rect 15284 29296 15293 29336
rect 16291 29296 16300 29336
rect 16340 29296 16684 29336
rect 16724 29296 16733 29336
rect 17059 29296 17068 29336
rect 17108 29296 17164 29336
rect 17204 29296 17213 29336
rect 19948 29296 20140 29336
rect 20180 29296 20189 29336
rect 0 29276 80 29296
rect 15235 29295 15293 29296
rect 17059 29295 17117 29296
rect 10723 29252 10781 29253
rect 2083 29212 2092 29252
rect 2132 29212 8620 29252
rect 8660 29212 8669 29252
rect 10723 29212 10732 29252
rect 10772 29212 11020 29252
rect 11060 29212 11069 29252
rect 16483 29212 16492 29252
rect 16532 29212 16972 29252
rect 17012 29212 17021 29252
rect 18115 29212 18124 29252
rect 18164 29212 19660 29252
rect 19700 29212 19709 29252
rect 10723 29211 10781 29212
rect 4195 29168 4253 29169
rect 5539 29168 5597 29169
rect 67 29128 76 29168
rect 116 29128 1900 29168
rect 1940 29128 1949 29168
rect 2659 29128 2668 29168
rect 2708 29128 3628 29168
rect 3668 29128 3677 29168
rect 4110 29128 4204 29168
rect 4244 29128 4253 29168
rect 5347 29128 5356 29168
rect 5396 29128 5548 29168
rect 5588 29128 5597 29168
rect 4195 29127 4253 29128
rect 5539 29127 5597 29128
rect 6883 29168 6941 29169
rect 6883 29128 6892 29168
rect 6932 29128 6988 29168
rect 7028 29128 7037 29168
rect 7363 29128 7372 29168
rect 7412 29128 9580 29168
rect 9620 29128 9629 29168
rect 10147 29128 10156 29168
rect 10196 29128 10924 29168
rect 10964 29128 10973 29168
rect 11683 29128 11692 29168
rect 11732 29128 12020 29168
rect 12067 29128 12076 29168
rect 12116 29128 12125 29168
rect 16771 29128 16780 29168
rect 16820 29128 17740 29168
rect 17780 29128 17789 29168
rect 18019 29128 18028 29168
rect 18068 29128 19948 29168
rect 19988 29128 19997 29168
rect 6883 29127 6941 29128
rect 1315 29084 1373 29085
rect 4771 29084 4829 29085
rect 460 29044 1036 29084
rect 1076 29044 1085 29084
rect 1315 29044 1324 29084
rect 1364 29044 2956 29084
rect 2996 29044 3005 29084
rect 3427 29044 3436 29084
rect 3476 29044 4780 29084
rect 4820 29044 4829 29084
rect 0 29000 80 29020
rect 460 29000 500 29044
rect 1315 29043 1373 29044
rect 4771 29043 4829 29044
rect 10828 29044 11308 29084
rect 11348 29044 11357 29084
rect 0 28960 500 29000
rect 1987 29000 2045 29001
rect 2947 29000 3005 29001
rect 10828 29000 10868 29044
rect 1987 28960 1996 29000
rect 2036 28960 2284 29000
rect 2324 28960 2333 29000
rect 2467 28960 2476 29000
rect 2516 28960 2668 29000
rect 2708 28960 2717 29000
rect 2947 28960 2956 29000
rect 2996 28960 3005 29000
rect 6403 28960 6412 29000
rect 6452 28960 6604 29000
rect 6644 28960 6653 29000
rect 10788 28960 10828 29000
rect 10868 28960 10877 29000
rect 0 28940 80 28960
rect 1987 28959 2045 28960
rect 2947 28959 3005 28960
rect 2755 28916 2813 28917
rect 2956 28916 2996 28959
rect 10723 28916 10781 28917
rect 11980 28916 12020 29128
rect 12076 29084 12116 29128
rect 17443 29084 17501 29085
rect 12076 29044 12308 29084
rect 16387 29044 16396 29084
rect 16436 29044 17220 29084
rect 17260 29044 17269 29084
rect 17443 29044 17452 29084
rect 17492 29044 17548 29084
rect 17588 29044 17597 29084
rect 12268 29000 12308 29044
rect 17443 29043 17501 29044
rect 12228 28960 12268 29000
rect 12308 28960 12317 29000
rect 17059 28916 17117 28917
rect 2755 28876 2764 28916
rect 2804 28876 2996 28916
rect 3139 28876 3148 28916
rect 3188 28876 4012 28916
rect 4052 28876 4061 28916
rect 10627 28876 10636 28916
rect 10676 28876 10732 28916
rect 10772 28876 10781 28916
rect 11971 28876 11980 28916
rect 12020 28876 12029 28916
rect 15523 28876 15532 28916
rect 15572 28876 16684 28916
rect 16724 28876 17068 28916
rect 17108 28876 17117 28916
rect 2755 28875 2813 28876
rect 10723 28875 10781 28876
rect 17059 28875 17117 28876
rect 7267 28832 7325 28833
rect 21424 28832 21504 28852
rect 7267 28792 7276 28832
rect 7316 28792 21504 28832
rect 7267 28791 7325 28792
rect 21424 28772 21504 28792
rect 3679 28708 3688 28748
rect 3728 28708 3770 28748
rect 3810 28708 3852 28748
rect 3892 28708 3934 28748
rect 3974 28708 4016 28748
rect 4056 28708 4065 28748
rect 4771 28708 4780 28748
rect 4820 28708 6412 28748
rect 6452 28708 6461 28748
rect 18799 28708 18808 28748
rect 18848 28708 18890 28748
rect 18930 28708 18972 28748
rect 19012 28708 19054 28748
rect 19094 28708 19136 28748
rect 19176 28708 19185 28748
rect 0 28664 80 28684
rect 0 28624 1940 28664
rect 1987 28624 1996 28664
rect 2036 28624 5932 28664
rect 5972 28624 5981 28664
rect 11491 28624 11500 28664
rect 11540 28624 12076 28664
rect 12116 28624 12125 28664
rect 0 28604 80 28624
rect 1900 28580 1940 28624
rect 1900 28540 5452 28580
rect 5492 28540 5501 28580
rect 10339 28540 10348 28580
rect 10388 28540 11212 28580
rect 11252 28540 11261 28580
rect 11875 28540 11884 28580
rect 11924 28540 12172 28580
rect 12212 28540 12221 28580
rect 12739 28540 12748 28580
rect 12788 28540 13228 28580
rect 13268 28540 13277 28580
rect 13315 28496 13373 28497
rect 3619 28456 3628 28496
rect 3668 28456 4108 28496
rect 4148 28456 4157 28496
rect 5539 28456 5548 28496
rect 5588 28456 5836 28496
rect 5876 28456 5885 28496
rect 6883 28456 6892 28496
rect 6932 28456 13324 28496
rect 13364 28456 13373 28496
rect 13315 28455 13373 28456
rect 19555 28496 19613 28497
rect 19555 28456 19564 28496
rect 19604 28456 20044 28496
rect 20084 28456 20093 28496
rect 19555 28455 19613 28456
rect 547 28412 605 28413
rect 547 28372 556 28412
rect 596 28372 3244 28412
rect 3284 28372 7988 28412
rect 8995 28372 9004 28412
rect 9044 28372 12652 28412
rect 12692 28372 17836 28412
rect 17876 28372 17885 28412
rect 547 28371 605 28372
rect 0 28328 80 28348
rect 0 28288 1708 28328
rect 1748 28288 1757 28328
rect 4099 28288 4108 28328
rect 4148 28288 4157 28328
rect 6307 28288 6316 28328
rect 6356 28288 6700 28328
rect 6740 28288 6749 28328
rect 0 28268 80 28288
rect 3139 28244 3197 28245
rect 4108 28244 4148 28288
rect 7948 28244 7988 28372
rect 19939 28328 19997 28329
rect 8323 28288 8332 28328
rect 8372 28288 9868 28328
rect 9908 28288 12748 28328
rect 12788 28288 12797 28328
rect 14179 28288 14188 28328
rect 14228 28288 14956 28328
rect 14996 28288 15005 28328
rect 19854 28288 19948 28328
rect 19988 28288 19997 28328
rect 19939 28287 19997 28288
rect 10819 28244 10877 28245
rect 13507 28244 13565 28245
rect 1315 28204 1324 28244
rect 1364 28204 3148 28244
rect 3188 28204 4148 28244
rect 5347 28204 5356 28244
rect 5396 28204 7084 28244
rect 7124 28204 7852 28244
rect 7892 28204 7901 28244
rect 7948 28204 10828 28244
rect 10868 28204 13516 28244
rect 13556 28204 13565 28244
rect 3139 28203 3197 28204
rect 10819 28203 10877 28204
rect 13507 28203 13565 28204
rect 4291 28160 4349 28161
rect 21424 28160 21504 28180
rect 3427 28120 3436 28160
rect 3476 28120 3724 28160
rect 3764 28120 3773 28160
rect 4206 28120 4300 28160
rect 4340 28120 4349 28160
rect 6787 28120 6796 28160
rect 6836 28120 8140 28160
rect 8180 28120 9292 28160
rect 9332 28120 10156 28160
rect 10196 28120 11116 28160
rect 11156 28120 11360 28160
rect 11779 28120 11788 28160
rect 11828 28120 21504 28160
rect 4291 28119 4349 28120
rect 4099 28036 4108 28076
rect 4148 28036 4684 28076
rect 4724 28036 4733 28076
rect 5923 28036 5932 28076
rect 5972 28036 6316 28076
rect 6356 28036 6365 28076
rect 0 27992 80 28012
rect 2275 27992 2333 27993
rect 11320 27992 11360 28120
rect 21424 28100 21504 28120
rect 18691 27992 18749 27993
rect 0 27932 116 27992
rect 2275 27952 2284 27992
rect 2324 27952 4244 27992
rect 4919 27952 4928 27992
rect 4968 27952 5010 27992
rect 5050 27952 5092 27992
rect 5132 27952 5174 27992
rect 5214 27952 5256 27992
rect 5296 27952 5305 27992
rect 7555 27952 7564 27992
rect 7604 27952 8044 27992
rect 8084 27952 8093 27992
rect 11320 27952 15436 27992
rect 15476 27952 15485 27992
rect 18307 27952 18316 27992
rect 18356 27952 18700 27992
rect 18740 27952 19756 27992
rect 19796 27952 19805 27992
rect 20039 27952 20048 27992
rect 20088 27952 20130 27992
rect 20170 27952 20212 27992
rect 20252 27952 20294 27992
rect 20334 27952 20376 27992
rect 20416 27952 20425 27992
rect 2275 27951 2333 27952
rect 76 27908 116 27932
rect 4204 27908 4244 27952
rect 18691 27951 18749 27952
rect 12451 27908 12509 27909
rect 76 27868 4148 27908
rect 4204 27868 5932 27908
rect 5972 27868 5981 27908
rect 9283 27868 9292 27908
rect 9332 27868 11884 27908
rect 11924 27868 11933 27908
rect 12366 27868 12460 27908
rect 12500 27868 12509 27908
rect 4108 27824 4148 27868
rect 12451 27867 12509 27868
rect 19276 27868 19468 27908
rect 19508 27868 19517 27908
rect 6979 27824 7037 27825
rect 2563 27784 2572 27824
rect 2612 27784 2860 27824
rect 2900 27784 2909 27824
rect 4108 27784 6932 27824
rect 2275 27740 2333 27741
rect 6892 27740 6932 27784
rect 6979 27784 6988 27824
rect 7028 27784 17836 27824
rect 17876 27784 18124 27824
rect 18164 27784 18173 27824
rect 6979 27783 7037 27784
rect 11107 27740 11165 27741
rect 1315 27700 1324 27740
rect 1364 27700 2284 27740
rect 2324 27700 2333 27740
rect 3811 27700 3820 27740
rect 3860 27700 4012 27740
rect 4052 27700 5644 27740
rect 5684 27700 5693 27740
rect 6892 27700 9100 27740
rect 9140 27700 9149 27740
rect 11011 27700 11020 27740
rect 11060 27700 11116 27740
rect 11156 27700 11165 27740
rect 2275 27699 2333 27700
rect 11107 27699 11165 27700
rect 16003 27740 16061 27741
rect 19276 27740 19316 27868
rect 19843 27784 19852 27824
rect 19892 27784 20180 27824
rect 20140 27740 20180 27784
rect 16003 27700 16012 27740
rect 16052 27700 16204 27740
rect 16244 27700 16253 27740
rect 17731 27700 17740 27740
rect 17780 27700 19316 27740
rect 20131 27700 20140 27740
rect 20180 27700 20189 27740
rect 16003 27699 16061 27700
rect 0 27656 80 27676
rect 0 27616 4052 27656
rect 4771 27616 4780 27656
rect 4820 27616 5260 27656
rect 5300 27616 5309 27656
rect 5443 27616 5452 27656
rect 5492 27616 5501 27656
rect 8611 27616 8620 27656
rect 8660 27616 9484 27656
rect 9524 27616 10540 27656
rect 10580 27616 10589 27656
rect 12163 27616 12172 27656
rect 12212 27616 13228 27656
rect 13268 27616 14284 27656
rect 14324 27616 14764 27656
rect 14804 27616 15532 27656
rect 15572 27616 15581 27656
rect 15715 27616 15724 27656
rect 15764 27616 17068 27656
rect 17108 27616 17117 27656
rect 0 27596 80 27616
rect 1795 27448 1804 27488
rect 1844 27448 2860 27488
rect 2900 27448 2909 27488
rect 4012 27404 4052 27616
rect 5452 27572 5492 27616
rect 4108 27532 5492 27572
rect 7075 27572 7133 27573
rect 15811 27572 15869 27573
rect 7075 27532 7084 27572
rect 7124 27532 10924 27572
rect 10964 27532 10973 27572
rect 14659 27532 14668 27572
rect 14708 27532 15628 27572
rect 15668 27532 15677 27572
rect 15811 27532 15820 27572
rect 15860 27532 15916 27572
rect 15956 27532 18220 27572
rect 18260 27532 18700 27572
rect 18740 27532 18749 27572
rect 4108 27488 4148 27532
rect 7075 27531 7133 27532
rect 15811 27531 15869 27532
rect 4291 27488 4349 27489
rect 21424 27488 21504 27508
rect 4099 27448 4108 27488
rect 4148 27448 4157 27488
rect 4291 27448 4300 27488
rect 4340 27448 4434 27488
rect 10147 27448 10156 27488
rect 10196 27448 10732 27488
rect 10772 27448 10781 27488
rect 11683 27448 11692 27488
rect 11732 27448 12268 27488
rect 12308 27448 12317 27488
rect 13411 27448 13420 27488
rect 13460 27448 14476 27488
rect 14516 27448 16588 27488
rect 16628 27448 17164 27488
rect 17204 27448 17213 27488
rect 19939 27448 19948 27488
rect 19988 27448 21504 27488
rect 4291 27447 4349 27448
rect 21424 27428 21504 27448
rect 6979 27404 7037 27405
rect 2467 27364 2476 27404
rect 2516 27364 2764 27404
rect 2804 27364 3956 27404
rect 4012 27364 6988 27404
rect 7028 27364 7037 27404
rect 11779 27364 11788 27404
rect 11828 27364 12364 27404
rect 12404 27364 12413 27404
rect 20035 27364 20044 27404
rect 20084 27364 20093 27404
rect 0 27320 80 27340
rect 3916 27320 3956 27364
rect 6979 27363 7037 27364
rect 20044 27320 20084 27364
rect 0 27280 2540 27320
rect 3916 27280 4204 27320
rect 4244 27280 4253 27320
rect 4771 27280 4780 27320
rect 4820 27280 6796 27320
rect 6836 27280 6845 27320
rect 10915 27280 10924 27320
rect 10964 27280 17260 27320
rect 17300 27280 17309 27320
rect 19459 27280 19468 27320
rect 19508 27280 20084 27320
rect 0 27260 80 27280
rect 2500 27152 2540 27280
rect 13795 27236 13853 27237
rect 3679 27196 3688 27236
rect 3728 27196 3770 27236
rect 3810 27196 3852 27236
rect 3892 27196 3934 27236
rect 3974 27196 4016 27236
rect 4056 27196 4065 27236
rect 10243 27196 10252 27236
rect 10292 27196 11308 27236
rect 11348 27196 11357 27236
rect 13795 27196 13804 27236
rect 13844 27196 18028 27236
rect 18068 27196 18077 27236
rect 18799 27196 18808 27236
rect 18848 27196 18890 27236
rect 18930 27196 18972 27236
rect 19012 27196 19054 27236
rect 19094 27196 19136 27236
rect 19176 27196 19185 27236
rect 19267 27196 19276 27236
rect 19316 27196 19660 27236
rect 19700 27196 19852 27236
rect 19892 27196 19901 27236
rect 13795 27195 13853 27196
rect 4195 27152 4253 27153
rect 2500 27112 4204 27152
rect 4244 27112 4253 27152
rect 4195 27111 4253 27112
rect 7660 27112 9964 27152
rect 10004 27112 18412 27152
rect 18452 27112 18461 27152
rect 3427 27068 3485 27069
rect 7660 27068 7700 27112
rect 9475 27068 9533 27069
rect 3427 27028 3436 27068
rect 3476 27028 7700 27068
rect 7747 27028 7756 27068
rect 7796 27028 9484 27068
rect 9524 27028 14188 27068
rect 14228 27028 14237 27068
rect 3427 27027 3485 27028
rect 9475 27027 9533 27028
rect 0 26984 80 27004
rect 2467 26984 2525 26985
rect 11587 26984 11645 26985
rect 12451 26984 12509 26985
rect 0 26944 2476 26984
rect 2516 26944 2525 26984
rect 4195 26944 4204 26984
rect 4244 26944 5740 26984
rect 5780 26944 8332 26984
rect 8372 26944 11360 26984
rect 11491 26944 11500 26984
rect 11540 26944 11596 26984
rect 11636 26944 11645 26984
rect 11971 26944 11980 26984
rect 12020 26944 12172 26984
rect 12212 26944 12221 26984
rect 12366 26944 12460 26984
rect 12500 26944 12509 26984
rect 13411 26944 13420 26984
rect 13460 26944 13469 26984
rect 16099 26944 16108 26984
rect 16148 26944 16588 26984
rect 16628 26944 16637 26984
rect 0 26924 80 26944
rect 2467 26943 2525 26944
rect 2179 26900 2237 26901
rect 11320 26900 11360 26944
rect 11587 26943 11645 26944
rect 12451 26943 12509 26944
rect 13420 26900 13460 26944
rect 2179 26860 2188 26900
rect 2228 26860 3572 26900
rect 6403 26860 6412 26900
rect 6452 26860 6796 26900
rect 6836 26860 6845 26900
rect 9763 26860 9772 26900
rect 9812 26860 9821 26900
rect 10051 26860 10060 26900
rect 10100 26860 11116 26900
rect 11156 26860 11165 26900
rect 11320 26860 13460 26900
rect 2179 26859 2237 26860
rect 3532 26817 3572 26860
rect 2563 26816 2621 26817
rect 3523 26816 3581 26817
rect 6595 26816 6653 26817
rect 8803 26816 8861 26817
rect 9571 26816 9629 26817
rect 2467 26776 2476 26816
rect 2516 26776 2572 26816
rect 2612 26776 3284 26816
rect 2563 26775 2621 26776
rect 739 26732 797 26733
rect 3244 26732 3284 26776
rect 3523 26776 3532 26816
rect 3572 26776 3724 26816
rect 3764 26776 3773 26816
rect 4483 26776 4492 26816
rect 4532 26776 4684 26816
rect 4724 26776 6604 26816
rect 6644 26776 6653 26816
rect 6883 26776 6892 26816
rect 6932 26776 7276 26816
rect 7316 26776 7325 26816
rect 8803 26776 8812 26816
rect 8852 26776 9580 26816
rect 9620 26776 9629 26816
rect 3523 26775 3581 26776
rect 6595 26775 6653 26776
rect 8803 26775 8861 26776
rect 9571 26775 9629 26776
rect 739 26692 748 26732
rect 788 26692 3148 26732
rect 3188 26692 3197 26732
rect 3244 26692 5260 26732
rect 5300 26692 5309 26732
rect 5923 26692 5932 26732
rect 5972 26692 6220 26732
rect 6260 26692 6269 26732
rect 7747 26692 7756 26732
rect 7796 26692 8140 26732
rect 8180 26692 8189 26732
rect 739 26691 797 26692
rect 0 26648 80 26668
rect 4579 26648 4637 26649
rect 7075 26648 7133 26649
rect 0 26608 748 26648
rect 788 26608 797 26648
rect 1123 26608 1132 26648
rect 1172 26608 3724 26648
rect 3764 26608 3773 26648
rect 4579 26608 4588 26648
rect 4628 26608 7084 26648
rect 7124 26608 7133 26648
rect 0 26588 80 26608
rect 4579 26607 4637 26608
rect 7075 26607 7133 26608
rect 9772 26564 9812 26860
rect 12451 26816 12509 26817
rect 21424 26816 21504 26836
rect 10627 26776 10636 26816
rect 10676 26776 10828 26816
rect 10868 26776 10877 26816
rect 11212 26776 11596 26816
rect 11636 26776 11645 26816
rect 12451 26776 12460 26816
rect 12500 26776 17932 26816
rect 17972 26776 17981 26816
rect 18691 26776 18700 26816
rect 18740 26776 19372 26816
rect 19412 26776 19421 26816
rect 19747 26776 19756 26816
rect 19796 26776 19805 26816
rect 20716 26776 21504 26816
rect 11212 26732 11252 26776
rect 12451 26775 12509 26776
rect 11587 26732 11645 26733
rect 19756 26732 19796 26776
rect 20716 26732 20756 26776
rect 21424 26756 21504 26776
rect 10339 26692 10348 26732
rect 10388 26692 11252 26732
rect 11320 26692 11596 26732
rect 11636 26692 11645 26732
rect 17347 26692 17356 26732
rect 17396 26692 17644 26732
rect 17684 26692 19796 26732
rect 19939 26692 19948 26732
rect 19988 26692 20756 26732
rect 11320 26648 11360 26692
rect 11587 26691 11645 26692
rect 10819 26608 10828 26648
rect 10868 26608 11360 26648
rect 12931 26648 12989 26649
rect 19939 26648 19997 26649
rect 12931 26608 12940 26648
rect 12980 26608 13516 26648
rect 13556 26608 13565 26648
rect 15907 26608 15916 26648
rect 15956 26608 17068 26648
rect 17108 26608 17117 26648
rect 19555 26608 19564 26648
rect 19604 26608 19948 26648
rect 19988 26608 19997 26648
rect 12931 26607 12989 26608
rect 19939 26607 19997 26608
rect 19843 26564 19901 26565
rect 5548 26524 6932 26564
rect 9772 26524 10252 26564
rect 10292 26524 11020 26564
rect 11060 26524 11069 26564
rect 11395 26524 11404 26564
rect 11444 26524 14572 26564
rect 14612 26524 17452 26564
rect 17492 26524 17501 26564
rect 19084 26524 19852 26564
rect 19892 26524 19901 26564
rect 4387 26480 4445 26481
rect 5548 26480 5588 26524
rect 6892 26480 6932 26524
rect 19084 26480 19124 26524
rect 19843 26523 19901 26524
rect 19555 26480 19613 26481
rect 2947 26440 2956 26480
rect 2996 26440 3436 26480
rect 3476 26440 3485 26480
rect 4302 26440 4396 26480
rect 4436 26440 4445 26480
rect 4919 26440 4928 26480
rect 4968 26440 5010 26480
rect 5050 26440 5092 26480
rect 5132 26440 5174 26480
rect 5214 26440 5256 26480
rect 5296 26440 5305 26480
rect 5539 26440 5548 26480
rect 5588 26440 5597 26480
rect 6892 26440 12268 26480
rect 12308 26440 12317 26480
rect 19075 26440 19084 26480
rect 19124 26440 19133 26480
rect 19267 26440 19276 26480
rect 19316 26440 19564 26480
rect 19604 26440 19613 26480
rect 20039 26440 20048 26480
rect 20088 26440 20130 26480
rect 20170 26440 20212 26480
rect 20252 26440 20294 26480
rect 20334 26440 20376 26480
rect 20416 26440 20425 26480
rect 4387 26439 4445 26440
rect 19555 26439 19613 26440
rect 0 26312 80 26332
rect 4675 26312 4733 26313
rect 7459 26312 7517 26313
rect 0 26272 4684 26312
rect 4724 26272 4733 26312
rect 5059 26272 5068 26312
rect 5108 26272 5452 26312
rect 5492 26272 5501 26312
rect 7374 26272 7468 26312
rect 7508 26272 7517 26312
rect 0 26252 80 26272
rect 4675 26271 4733 26272
rect 7459 26271 7517 26272
rect 9667 26312 9725 26313
rect 11203 26312 11261 26313
rect 9667 26272 9676 26312
rect 9716 26272 9964 26312
rect 10004 26272 10013 26312
rect 11118 26272 11212 26312
rect 11252 26272 11261 26312
rect 9667 26271 9725 26272
rect 11203 26271 11261 26272
rect 2467 26228 2525 26229
rect 2467 26188 2476 26228
rect 2516 26188 3148 26228
rect 3188 26188 3197 26228
rect 7756 26188 11500 26228
rect 11540 26188 11549 26228
rect 12355 26188 12364 26228
rect 12404 26188 14956 26228
rect 14996 26188 15188 26228
rect 15811 26188 15820 26228
rect 15860 26188 16972 26228
rect 17012 26188 17021 26228
rect 2467 26187 2525 26188
rect 3523 26144 3581 26145
rect 6115 26144 6173 26145
rect 7555 26144 7613 26145
rect 7756 26144 7796 26188
rect 15148 26144 15188 26188
rect 17635 26144 17693 26145
rect 21424 26144 21504 26164
rect 1507 26104 1516 26144
rect 1556 26104 2188 26144
rect 2228 26104 2237 26144
rect 2851 26104 2860 26144
rect 2900 26104 3244 26144
rect 3284 26104 3293 26144
rect 3438 26104 3532 26144
rect 3572 26104 3581 26144
rect 4483 26104 4492 26144
rect 4532 26104 5260 26144
rect 5300 26104 5309 26144
rect 6115 26104 6124 26144
rect 6164 26104 7084 26144
rect 7124 26104 7372 26144
rect 7412 26104 7421 26144
rect 7555 26104 7564 26144
rect 7604 26104 7756 26144
rect 7796 26104 7805 26144
rect 8803 26104 8812 26144
rect 8852 26104 9004 26144
rect 9044 26104 9053 26144
rect 10060 26104 14668 26144
rect 14708 26104 14717 26144
rect 15139 26104 15148 26144
rect 15188 26104 15197 26144
rect 15427 26104 15436 26144
rect 15476 26104 16204 26144
rect 16244 26104 16253 26144
rect 17635 26104 17644 26144
rect 17684 26104 21504 26144
rect 3523 26103 3581 26104
rect 6115 26103 6173 26104
rect 7555 26103 7613 26104
rect 10060 26060 10100 26104
rect 17635 26103 17693 26104
rect 21424 26084 21504 26104
rect 14563 26060 14621 26061
rect 1027 26020 1036 26060
rect 1076 26020 10060 26060
rect 10100 26020 10109 26060
rect 14478 26020 14572 26060
rect 14612 26020 14621 26060
rect 14563 26019 14621 26020
rect 0 25976 80 25996
rect 2851 25976 2909 25977
rect 0 25936 2860 25976
rect 2900 25936 2909 25976
rect 0 25916 80 25936
rect 2851 25935 2909 25936
rect 3331 25976 3389 25977
rect 3331 25936 3340 25976
rect 3380 25936 4780 25976
rect 4820 25936 4829 25976
rect 7468 25936 11980 25976
rect 12020 25936 12029 25976
rect 3331 25935 3389 25936
rect 5923 25892 5981 25893
rect 7468 25892 7508 25936
rect 8419 25892 8477 25893
rect 2179 25852 2188 25892
rect 2228 25852 3532 25892
rect 3572 25852 3581 25892
rect 5923 25852 5932 25892
rect 5972 25852 6028 25892
rect 6068 25852 7508 25892
rect 7555 25852 7564 25892
rect 7604 25852 7756 25892
rect 7796 25852 7805 25892
rect 8419 25852 8428 25892
rect 8468 25852 13132 25892
rect 13172 25852 13181 25892
rect 16003 25852 16012 25892
rect 16052 25852 16684 25892
rect 16724 25852 16733 25892
rect 5923 25851 5981 25852
rect 8419 25851 8477 25852
rect 2659 25808 2717 25809
rect 2371 25768 2380 25808
rect 2420 25768 2429 25808
rect 2659 25768 2668 25808
rect 2708 25768 9100 25808
rect 9140 25768 9149 25808
rect 9955 25768 9964 25808
rect 10004 25768 10252 25808
rect 10292 25768 10301 25808
rect 2380 25724 2420 25768
rect 2659 25767 2717 25768
rect 4771 25724 4829 25725
rect 1507 25684 1516 25724
rect 1556 25684 2420 25724
rect 3679 25684 3688 25724
rect 3728 25684 3770 25724
rect 3810 25684 3852 25724
rect 3892 25684 3934 25724
rect 3974 25684 4016 25724
rect 4056 25684 4065 25724
rect 4195 25684 4204 25724
rect 4244 25684 4780 25724
rect 4820 25684 6604 25724
rect 6644 25684 6653 25724
rect 9187 25684 9196 25724
rect 9236 25684 9484 25724
rect 9524 25684 9533 25724
rect 18799 25684 18808 25724
rect 18848 25684 18890 25724
rect 18930 25684 18972 25724
rect 19012 25684 19054 25724
rect 19094 25684 19136 25724
rect 19176 25684 19185 25724
rect 4771 25683 4829 25684
rect 0 25640 80 25660
rect 4963 25640 5021 25641
rect 0 25600 1996 25640
rect 2036 25600 2045 25640
rect 4963 25600 4972 25640
rect 5012 25600 5780 25640
rect 14659 25600 14668 25640
rect 14708 25600 15244 25640
rect 15284 25600 15293 25640
rect 0 25580 80 25600
rect 4963 25599 5021 25600
rect 2467 25516 2476 25556
rect 2516 25516 2764 25556
rect 2804 25516 2813 25556
rect 3139 25516 3148 25556
rect 3188 25516 5164 25556
rect 5204 25516 5213 25556
rect 2179 25432 2188 25472
rect 2228 25432 4684 25472
rect 4724 25432 4733 25472
rect 5251 25432 5260 25472
rect 5300 25432 5644 25472
rect 5684 25432 5693 25472
rect 2659 25388 2717 25389
rect 3427 25388 3485 25389
rect 5740 25388 5780 25600
rect 5827 25516 5836 25556
rect 5876 25516 7660 25556
rect 7700 25516 7709 25556
rect 14083 25516 14092 25556
rect 14132 25516 14572 25556
rect 14612 25516 14956 25556
rect 14996 25516 15005 25556
rect 15139 25516 15148 25556
rect 15188 25516 16108 25556
rect 16148 25516 16157 25556
rect 11107 25472 11165 25473
rect 21424 25472 21504 25492
rect 11107 25432 11116 25472
rect 11156 25432 11404 25472
rect 11444 25432 11453 25472
rect 16291 25432 16300 25472
rect 16340 25432 17164 25472
rect 17204 25432 17213 25472
rect 20908 25432 21504 25472
rect 11107 25431 11165 25432
rect 11299 25388 11357 25389
rect 20908 25388 20948 25432
rect 21424 25412 21504 25432
rect 2284 25348 2668 25388
rect 2708 25348 2717 25388
rect 2851 25348 2860 25388
rect 2900 25348 3436 25388
rect 3476 25348 3485 25388
rect 0 25304 80 25324
rect 2284 25304 2324 25348
rect 2659 25347 2717 25348
rect 3427 25347 3485 25348
rect 4780 25348 5164 25388
rect 5204 25348 5213 25388
rect 5740 25348 5836 25388
rect 5876 25348 5885 25388
rect 11299 25348 11308 25388
rect 11348 25348 20948 25388
rect 4780 25304 4820 25348
rect 0 25264 2324 25304
rect 2371 25264 2380 25304
rect 2420 25264 3148 25304
rect 3188 25264 3197 25304
rect 3811 25264 3820 25304
rect 3860 25264 4204 25304
rect 4244 25264 4253 25304
rect 4771 25264 4780 25304
rect 4820 25264 4829 25304
rect 0 25244 80 25264
rect 4771 25220 4829 25221
rect 4291 25180 4300 25220
rect 4340 25180 4780 25220
rect 4820 25180 4829 25220
rect 4771 25179 4829 25180
rect 5059 25220 5117 25221
rect 5740 25220 5780 25348
rect 11299 25347 11357 25348
rect 7075 25304 7133 25305
rect 8995 25304 9053 25305
rect 6403 25264 6412 25304
rect 6452 25264 6700 25304
rect 6740 25264 6749 25304
rect 7075 25264 7084 25304
rect 7124 25264 7276 25304
rect 7316 25264 7325 25304
rect 8995 25264 9004 25304
rect 9044 25264 9772 25304
rect 9812 25264 9821 25304
rect 10243 25264 10252 25304
rect 10292 25264 10924 25304
rect 10964 25264 10973 25304
rect 14947 25264 14956 25304
rect 14996 25264 15340 25304
rect 15380 25264 15389 25304
rect 7075 25263 7133 25264
rect 8995 25263 9053 25264
rect 5059 25180 5068 25220
rect 5108 25180 5119 25220
rect 5443 25180 5452 25220
rect 5492 25180 5780 25220
rect 6307 25220 6365 25221
rect 6307 25180 6316 25220
rect 6356 25180 6796 25220
rect 6836 25180 6845 25220
rect 6979 25180 6988 25220
rect 7028 25180 7948 25220
rect 7988 25180 7997 25220
rect 14371 25180 14380 25220
rect 14420 25180 15436 25220
rect 15476 25180 16492 25220
rect 16532 25180 17836 25220
rect 17876 25180 18220 25220
rect 18260 25180 18269 25220
rect 5059 25179 5117 25180
rect 6307 25179 6365 25180
rect 5068 25136 5108 25179
rect 5251 25136 5309 25137
rect 12451 25136 12509 25137
rect 5059 25096 5068 25136
rect 5108 25096 5117 25136
rect 5251 25096 5260 25136
rect 5300 25096 12460 25136
rect 12500 25096 12509 25136
rect 5251 25095 5309 25096
rect 12451 25095 12509 25096
rect 4387 25052 4445 25053
rect 2467 25012 2476 25052
rect 2516 25012 2668 25052
rect 2708 25012 2717 25052
rect 4387 25012 4396 25052
rect 4436 25012 5972 25052
rect 6307 25012 6316 25052
rect 6356 25012 6892 25052
rect 6932 25012 6941 25052
rect 8419 25012 8428 25052
rect 8468 25012 8716 25052
rect 8756 25012 8765 25052
rect 4387 25011 4445 25012
rect 0 24968 80 24988
rect 835 24968 893 24969
rect 5932 24968 5972 25012
rect 0 24928 844 24968
rect 884 24928 893 24968
rect 1315 24928 1324 24968
rect 1364 24928 1804 24968
rect 1844 24928 1853 24968
rect 4919 24928 4928 24968
rect 4968 24928 5010 24968
rect 5050 24928 5092 24968
rect 5132 24928 5174 24968
rect 5214 24928 5256 24968
rect 5296 24928 5305 24968
rect 5731 24928 5740 24968
rect 5780 24928 5876 24968
rect 5932 24928 11884 24968
rect 11924 24928 11933 24968
rect 20039 24928 20048 24968
rect 20088 24928 20130 24968
rect 20170 24928 20212 24968
rect 20252 24928 20294 24968
rect 20334 24928 20376 24968
rect 20416 24928 20425 24968
rect 0 24908 80 24928
rect 835 24927 893 24928
rect 5731 24884 5789 24885
rect 4195 24844 4204 24884
rect 4244 24844 5740 24884
rect 5780 24844 5789 24884
rect 5836 24884 5876 24928
rect 5836 24844 14092 24884
rect 14132 24844 14141 24884
rect 5731 24843 5789 24844
rect 4579 24800 4637 24801
rect 5635 24800 5693 24801
rect 8707 24800 8765 24801
rect 1795 24760 1804 24800
rect 1844 24760 4340 24800
rect 2275 24716 2333 24717
rect 4300 24716 4340 24760
rect 4579 24760 4588 24800
rect 4628 24760 4876 24800
rect 4916 24760 4925 24800
rect 5347 24760 5356 24800
rect 5396 24760 5644 24800
rect 5684 24760 6983 24800
rect 7023 24760 7032 24800
rect 7075 24760 7084 24800
rect 7124 24760 8716 24800
rect 8756 24760 8765 24800
rect 4579 24759 4637 24760
rect 5635 24759 5693 24760
rect 8707 24759 8765 24760
rect 9187 24800 9245 24801
rect 9763 24800 9821 24801
rect 15139 24800 15197 24801
rect 21424 24800 21504 24820
rect 9187 24760 9196 24800
rect 9236 24760 9292 24800
rect 9332 24760 9341 24800
rect 9763 24760 9772 24800
rect 9812 24760 9868 24800
rect 9908 24760 9917 24800
rect 11107 24760 11116 24800
rect 11156 24760 15148 24800
rect 15188 24760 15197 24800
rect 16099 24760 16108 24800
rect 16148 24760 16780 24800
rect 16820 24760 16972 24800
rect 17012 24760 17021 24800
rect 17347 24760 17356 24800
rect 17396 24760 21504 24800
rect 9187 24759 9245 24760
rect 9763 24759 9821 24760
rect 15139 24759 15197 24760
rect 21424 24740 21504 24760
rect 2275 24676 2284 24716
rect 2324 24676 4204 24716
rect 4244 24676 4253 24716
rect 4300 24676 11596 24716
rect 11636 24676 15380 24716
rect 2275 24675 2333 24676
rect 0 24632 80 24652
rect 9667 24632 9725 24633
rect 10435 24632 10493 24633
rect 11203 24632 11261 24633
rect 15340 24632 15380 24676
rect 15427 24632 15485 24633
rect 16963 24632 17021 24633
rect 0 24592 8372 24632
rect 0 24572 80 24592
rect 1315 24548 1373 24549
rect 3331 24548 3389 24549
rect 5539 24548 5597 24549
rect 7747 24548 7805 24549
rect 1230 24508 1324 24548
rect 1364 24508 1373 24548
rect 3139 24508 3148 24548
rect 3188 24508 3340 24548
rect 3380 24508 3389 24548
rect 4387 24508 4396 24548
rect 4436 24508 5548 24548
rect 5588 24508 5597 24548
rect 5923 24508 5932 24548
rect 5972 24508 7756 24548
rect 7796 24508 7852 24548
rect 7892 24508 7920 24548
rect 1315 24507 1373 24508
rect 3331 24507 3389 24508
rect 5539 24507 5597 24508
rect 7747 24507 7805 24508
rect 3340 24464 3380 24507
rect 6115 24464 6173 24465
rect 8332 24464 8372 24592
rect 9667 24592 9676 24632
rect 9716 24592 9868 24632
rect 9908 24592 9917 24632
rect 10435 24592 10444 24632
rect 10484 24592 11212 24632
rect 11252 24592 12652 24632
rect 12692 24592 12701 24632
rect 14371 24592 14380 24632
rect 14420 24592 14956 24632
rect 14996 24592 15005 24632
rect 15331 24592 15340 24632
rect 15380 24592 15436 24632
rect 15476 24592 15485 24632
rect 16867 24592 16876 24632
rect 16916 24592 16972 24632
rect 17012 24592 17021 24632
rect 9667 24591 9725 24592
rect 10435 24591 10493 24592
rect 11203 24591 11261 24592
rect 15427 24591 15485 24592
rect 16963 24591 17021 24592
rect 8611 24548 8669 24549
rect 8611 24508 8620 24548
rect 8660 24508 21292 24548
rect 21332 24508 21341 24548
rect 8611 24507 8669 24508
rect 2467 24424 2476 24464
rect 2516 24424 3052 24464
rect 3092 24424 3101 24464
rect 3340 24424 5356 24464
rect 5396 24424 5405 24464
rect 6030 24424 6124 24464
rect 6164 24424 6173 24464
rect 7363 24424 7372 24464
rect 7412 24424 8236 24464
rect 8276 24424 8285 24464
rect 8332 24424 16492 24464
rect 16532 24424 16541 24464
rect 6115 24423 6173 24424
rect 6499 24380 6557 24381
rect 7459 24380 7517 24381
rect 3235 24340 3244 24380
rect 3284 24340 6220 24380
rect 6260 24340 6269 24380
rect 6499 24340 6508 24380
rect 6548 24340 7084 24380
rect 7124 24340 7468 24380
rect 7508 24340 7517 24380
rect 6499 24339 6557 24340
rect 7459 24339 7517 24340
rect 9187 24380 9245 24381
rect 12355 24380 12413 24381
rect 9187 24340 9196 24380
rect 9236 24340 9388 24380
rect 9428 24340 9437 24380
rect 10531 24340 10540 24380
rect 10580 24340 11116 24380
rect 11156 24340 11165 24380
rect 12270 24340 12364 24380
rect 12404 24340 12413 24380
rect 9187 24339 9245 24340
rect 12355 24339 12413 24340
rect 0 24296 80 24316
rect 6019 24296 6077 24297
rect 0 24256 3340 24296
rect 3380 24256 3389 24296
rect 3532 24256 6028 24296
rect 6068 24256 6077 24296
rect 0 24236 80 24256
rect 3532 24212 3572 24256
rect 6019 24255 6077 24256
rect 6787 24296 6845 24297
rect 6787 24256 6796 24296
rect 6836 24256 7180 24296
rect 7220 24256 7229 24296
rect 8803 24256 8812 24296
rect 8852 24256 11308 24296
rect 11348 24256 11357 24296
rect 15139 24256 15148 24296
rect 15188 24256 15532 24296
rect 15572 24256 15581 24296
rect 6787 24255 6845 24256
rect 10435 24212 10493 24213
rect 11875 24212 11933 24213
rect 460 24172 3572 24212
rect 3679 24172 3688 24212
rect 3728 24172 3770 24212
rect 3810 24172 3852 24212
rect 3892 24172 3934 24212
rect 3974 24172 4016 24212
rect 4056 24172 4065 24212
rect 5635 24172 5644 24212
rect 5684 24172 10444 24212
rect 10484 24172 10493 24212
rect 11683 24172 11692 24212
rect 11732 24172 11884 24212
rect 11924 24172 11933 24212
rect 18799 24172 18808 24212
rect 18848 24172 18890 24212
rect 18930 24172 18972 24212
rect 19012 24172 19054 24212
rect 19094 24172 19136 24212
rect 19176 24172 19185 24212
rect 0 23960 80 23980
rect 460 23960 500 24172
rect 10435 24171 10493 24172
rect 11875 24171 11933 24172
rect 12451 24128 12509 24129
rect 21424 24128 21504 24148
rect 1699 24088 1708 24128
rect 1748 24088 2132 24128
rect 4387 24088 4396 24128
rect 4436 24088 4588 24128
rect 4628 24088 4637 24128
rect 5251 24088 5260 24128
rect 5300 24088 6028 24128
rect 6068 24088 6077 24128
rect 12366 24088 12460 24128
rect 12500 24088 12509 24128
rect 13699 24088 13708 24128
rect 13748 24088 14188 24128
rect 14228 24088 14237 24128
rect 15532 24088 15764 24128
rect 17251 24088 17260 24128
rect 17300 24088 21504 24128
rect 0 23920 500 23960
rect 0 23900 80 23920
rect 2092 23876 2132 24088
rect 12451 24087 12509 24088
rect 15532 24044 15572 24088
rect 15724 24044 15764 24088
rect 21424 24068 21504 24088
rect 3811 24004 3820 24044
rect 3860 24004 15572 24044
rect 15619 24004 15628 24044
rect 15668 24004 15677 24044
rect 15724 24004 20620 24044
rect 20660 24004 20669 24044
rect 7747 23960 7805 23961
rect 12643 23960 12701 23961
rect 15628 23960 15668 24004
rect 2659 23920 2668 23960
rect 2708 23920 3532 23960
rect 3572 23920 3581 23960
rect 4291 23920 4300 23960
rect 4340 23920 7564 23960
rect 7604 23920 7613 23960
rect 7747 23920 7756 23960
rect 7796 23920 8044 23960
rect 8084 23920 8093 23960
rect 11683 23920 11692 23960
rect 11732 23920 12404 23960
rect 7747 23919 7805 23920
rect 3427 23876 3485 23877
rect 7267 23876 7325 23877
rect 12364 23876 12404 23920
rect 12643 23920 12652 23960
rect 12692 23920 12748 23960
rect 12788 23920 12797 23960
rect 13123 23920 13132 23960
rect 13172 23920 13181 23960
rect 13987 23920 13996 23960
rect 14036 23920 14380 23960
rect 14420 23920 14429 23960
rect 14563 23920 14572 23960
rect 14612 23920 14621 23960
rect 15628 23920 17068 23960
rect 17108 23920 17117 23960
rect 17827 23920 17836 23960
rect 17876 23920 19372 23960
rect 19412 23920 19421 23960
rect 12643 23919 12701 23920
rect 2092 23836 2572 23876
rect 2612 23836 2621 23876
rect 3427 23836 3436 23876
rect 3476 23836 5836 23876
rect 5876 23836 5885 23876
rect 6307 23836 6316 23876
rect 6356 23836 6604 23876
rect 6644 23836 6653 23876
rect 7182 23836 7276 23876
rect 7316 23836 8140 23876
rect 8180 23836 8189 23876
rect 12355 23836 12364 23876
rect 12404 23836 12413 23876
rect 3427 23835 3485 23836
rect 7267 23835 7325 23836
rect 1411 23752 1420 23792
rect 1460 23752 2284 23792
rect 2324 23752 2476 23792
rect 2516 23752 2525 23792
rect 2851 23752 2860 23792
rect 2900 23752 3148 23792
rect 3188 23752 3197 23792
rect 5443 23752 5452 23792
rect 5492 23752 5740 23792
rect 5780 23752 6700 23792
rect 6740 23752 7756 23792
rect 7796 23752 7805 23792
rect 8323 23752 8332 23792
rect 8372 23752 8620 23792
rect 8660 23752 8669 23792
rect 8803 23752 8812 23792
rect 8852 23752 9484 23792
rect 9524 23752 9533 23792
rect 11203 23752 11212 23792
rect 11252 23752 11500 23792
rect 11540 23752 11884 23792
rect 11924 23752 11933 23792
rect 12067 23752 12076 23792
rect 12116 23752 12652 23792
rect 12692 23752 12701 23792
rect 1315 23668 1324 23708
rect 1364 23668 2188 23708
rect 2228 23668 2237 23708
rect 3523 23668 3532 23708
rect 3572 23668 6124 23708
rect 6164 23668 6173 23708
rect 7459 23668 7468 23708
rect 7508 23668 9100 23708
rect 9140 23668 9149 23708
rect 10723 23668 10732 23708
rect 10772 23668 11308 23708
rect 11348 23668 11357 23708
rect 0 23624 80 23644
rect 12355 23624 12413 23625
rect 13132 23624 13172 23920
rect 14572 23876 14612 23920
rect 13507 23836 13516 23876
rect 13556 23836 15724 23876
rect 15764 23836 15773 23876
rect 15907 23836 15916 23876
rect 15956 23836 18028 23876
rect 18068 23836 19180 23876
rect 19220 23836 19229 23876
rect 14083 23792 14141 23793
rect 13987 23752 13996 23792
rect 14036 23752 14092 23792
rect 14132 23752 14141 23792
rect 14275 23752 14284 23792
rect 14324 23752 14572 23792
rect 14612 23752 14621 23792
rect 15043 23752 15052 23792
rect 15092 23752 15820 23792
rect 15860 23752 15869 23792
rect 15916 23752 18124 23792
rect 18164 23752 18173 23792
rect 14083 23751 14141 23752
rect 15235 23668 15244 23708
rect 15284 23668 15532 23708
rect 15572 23668 15581 23708
rect 15916 23624 15956 23752
rect 17635 23668 17644 23708
rect 17684 23668 19852 23708
rect 19892 23668 19901 23708
rect 0 23584 8428 23624
rect 8468 23584 8477 23624
rect 8803 23584 8812 23624
rect 8852 23584 12364 23624
rect 12404 23584 12413 23624
rect 13123 23584 13132 23624
rect 13172 23584 13181 23624
rect 13507 23584 13516 23624
rect 13556 23584 15956 23624
rect 16099 23584 16108 23624
rect 16148 23584 16300 23624
rect 16340 23584 16349 23624
rect 19267 23584 19276 23624
rect 19316 23584 19564 23624
rect 19604 23584 19613 23624
rect 20035 23584 20044 23624
rect 20084 23584 20093 23624
rect 0 23564 80 23584
rect 12355 23583 12413 23584
rect 6499 23540 6557 23541
rect 8707 23540 8765 23541
rect 20044 23540 20084 23584
rect 1699 23500 1708 23540
rect 1748 23500 6508 23540
rect 6548 23500 6557 23540
rect 7651 23500 7660 23540
rect 7700 23500 8140 23540
rect 8180 23500 8189 23540
rect 8707 23500 8716 23540
rect 8756 23500 16780 23540
rect 16820 23500 16829 23540
rect 17827 23500 17836 23540
rect 17876 23500 18028 23540
rect 18068 23500 18077 23540
rect 19843 23500 19852 23540
rect 19892 23500 20084 23540
rect 6499 23499 6557 23500
rect 8707 23499 8765 23500
rect 21424 23456 21504 23476
rect 1027 23416 1036 23456
rect 1076 23416 4108 23456
rect 4148 23416 4157 23456
rect 4919 23416 4928 23456
rect 4968 23416 5010 23456
rect 5050 23416 5092 23456
rect 5132 23416 5174 23456
rect 5214 23416 5256 23456
rect 5296 23416 5305 23456
rect 6892 23416 12556 23456
rect 12596 23416 12605 23456
rect 14947 23416 14956 23456
rect 14996 23416 15244 23456
rect 15284 23416 15293 23456
rect 15523 23416 15532 23456
rect 15572 23416 16108 23456
rect 16148 23416 16684 23456
rect 16724 23416 16733 23456
rect 20039 23416 20048 23456
rect 20088 23416 20130 23456
rect 20170 23416 20212 23456
rect 20252 23416 20294 23456
rect 20334 23416 20376 23456
rect 20416 23416 20425 23456
rect 20611 23416 20620 23456
rect 20660 23416 21504 23456
rect 1987 23332 1996 23372
rect 2036 23332 2476 23372
rect 2516 23332 2525 23372
rect 0 23288 80 23308
rect 6892 23288 6932 23416
rect 21424 23396 21504 23416
rect 7564 23332 16396 23372
rect 16436 23332 16445 23372
rect 17827 23332 17836 23372
rect 17876 23332 18604 23372
rect 18644 23332 18653 23372
rect 7267 23288 7325 23289
rect 0 23248 6932 23288
rect 7075 23248 7084 23288
rect 7124 23248 7276 23288
rect 7316 23248 7325 23288
rect 0 23228 80 23248
rect 7267 23247 7325 23248
rect 4195 23204 4253 23205
rect 7564 23204 7604 23332
rect 7651 23288 7709 23289
rect 8707 23288 8765 23289
rect 7651 23248 7660 23288
rect 7700 23248 8716 23288
rect 8756 23248 8765 23288
rect 7651 23247 7709 23248
rect 8707 23247 8765 23248
rect 11320 23248 12076 23288
rect 12116 23248 12125 23288
rect 12547 23248 12556 23288
rect 12596 23248 12844 23288
rect 12884 23248 13612 23288
rect 13652 23248 13661 23288
rect 15427 23248 15436 23288
rect 15476 23248 15820 23288
rect 15860 23248 15869 23288
rect 4195 23164 4204 23204
rect 4244 23164 7604 23204
rect 9475 23164 9484 23204
rect 9524 23164 10444 23204
rect 10484 23164 10493 23204
rect 4195 23163 4253 23164
rect 11320 23120 11360 23248
rect 11491 23164 11500 23204
rect 11540 23164 13420 23204
rect 13460 23164 13469 23204
rect 15235 23164 15244 23204
rect 15284 23164 15668 23204
rect 11692 23120 11732 23164
rect 4003 23080 4012 23120
rect 4052 23080 10060 23120
rect 10100 23080 11360 23120
rect 11683 23080 11692 23120
rect 11732 23080 11772 23120
rect 12355 23080 12364 23120
rect 12404 23080 13612 23120
rect 13652 23080 15532 23120
rect 15572 23080 15581 23120
rect 4195 23036 4253 23037
rect 15427 23036 15485 23037
rect 2659 22996 2668 23036
rect 2708 22996 3916 23036
rect 3956 22996 4204 23036
rect 4244 22996 4253 23036
rect 6019 22996 6028 23036
rect 6068 22996 6892 23036
rect 6932 22996 8524 23036
rect 8564 22996 8573 23036
rect 11596 22996 12940 23036
rect 12980 22996 14284 23036
rect 14324 22996 14333 23036
rect 15342 22996 15436 23036
rect 15476 22996 15485 23036
rect 4195 22995 4253 22996
rect 0 22952 80 22972
rect 8524 22952 8564 22996
rect 9955 22952 10013 22953
rect 11596 22952 11636 22996
rect 15427 22995 15485 22996
rect 15628 22952 15668 23164
rect 0 22912 2092 22952
rect 2132 22912 2141 22952
rect 2275 22912 2284 22952
rect 2324 22912 3436 22952
rect 3476 22912 3485 22952
rect 8524 22912 8716 22952
rect 8756 22912 8765 22952
rect 9840 22912 9868 22952
rect 9908 22912 9964 22952
rect 10004 22912 11636 22952
rect 12067 22912 12076 22952
rect 12116 22912 15476 22952
rect 15523 22912 15532 22952
rect 15572 22912 15668 22952
rect 0 22892 80 22912
rect 9955 22911 10013 22912
rect 15436 22868 15476 22912
rect 15811 22868 15869 22869
rect 16108 22868 16148 23332
rect 17443 23248 17452 23288
rect 17492 23248 18220 23288
rect 18260 23248 18412 23288
rect 18452 23248 18461 23288
rect 18691 23080 18700 23120
rect 18740 23080 19756 23120
rect 19796 23080 19805 23120
rect 20131 22868 20189 22869
rect 1411 22828 1420 22868
rect 1460 22828 1996 22868
rect 2036 22828 5356 22868
rect 5396 22828 6604 22868
rect 6644 22828 6653 22868
rect 7075 22828 7084 22868
rect 7124 22828 8140 22868
rect 8180 22828 8189 22868
rect 8419 22828 8428 22868
rect 8468 22828 13708 22868
rect 13748 22828 13757 22868
rect 15436 22828 15820 22868
rect 15860 22828 15869 22868
rect 16099 22828 16108 22868
rect 16148 22828 16157 22868
rect 20131 22828 20140 22868
rect 20180 22828 20189 22868
rect 15811 22827 15869 22828
rect 20131 22827 20189 22828
rect 2563 22784 2621 22785
rect 20140 22784 20180 22827
rect 21424 22784 21504 22804
rect 2563 22744 2572 22784
rect 2612 22744 2706 22784
rect 15619 22744 15628 22784
rect 15668 22744 15916 22784
rect 15956 22744 15965 22784
rect 20140 22744 21504 22784
rect 2563 22743 2621 22744
rect 21424 22724 21504 22744
rect 3679 22660 3688 22700
rect 3728 22660 3770 22700
rect 3810 22660 3852 22700
rect 3892 22660 3934 22700
rect 3974 22660 4016 22700
rect 4056 22660 4065 22700
rect 10435 22660 10444 22700
rect 10484 22660 11980 22700
rect 12020 22660 13132 22700
rect 13172 22660 13181 22700
rect 16195 22660 16204 22700
rect 16244 22660 16972 22700
rect 17012 22660 17021 22700
rect 18799 22660 18808 22700
rect 18848 22660 18890 22700
rect 18930 22660 18972 22700
rect 19012 22660 19054 22700
rect 19094 22660 19136 22700
rect 19176 22660 19185 22700
rect 0 22616 80 22636
rect 0 22576 1900 22616
rect 1940 22576 1949 22616
rect 8515 22576 8524 22616
rect 8564 22576 14380 22616
rect 14420 22576 14429 22616
rect 16387 22576 16396 22616
rect 16436 22576 17356 22616
rect 17396 22576 17405 22616
rect 0 22556 80 22576
rect 11779 22492 11788 22532
rect 11828 22492 13996 22532
rect 14036 22492 17452 22532
rect 17492 22492 17501 22532
rect 2380 22408 9772 22448
rect 9812 22408 9821 22448
rect 12163 22408 12172 22448
rect 12212 22408 13132 22448
rect 13172 22408 13181 22448
rect 0 22280 80 22300
rect 2380 22280 2420 22408
rect 12451 22364 12509 22365
rect 3523 22324 3532 22364
rect 3572 22324 6412 22364
rect 6452 22324 6461 22364
rect 11875 22324 11884 22364
rect 11924 22324 12076 22364
rect 12116 22324 12125 22364
rect 12451 22324 12460 22364
rect 12500 22324 14092 22364
rect 14132 22324 14141 22364
rect 12451 22323 12509 22324
rect 3331 22280 3389 22281
rect 4483 22280 4541 22281
rect 13315 22280 13373 22281
rect 0 22240 2420 22280
rect 2467 22240 2476 22280
rect 2516 22240 3052 22280
rect 3092 22240 3340 22280
rect 3380 22240 3389 22280
rect 4398 22240 4492 22280
rect 4532 22240 4541 22280
rect 5443 22240 5452 22280
rect 5492 22240 5740 22280
rect 5780 22240 5789 22280
rect 6115 22240 6124 22280
rect 6164 22240 6173 22280
rect 6787 22240 6796 22280
rect 6836 22240 7660 22280
rect 7700 22240 7709 22280
rect 8323 22240 8332 22280
rect 8372 22240 8908 22280
rect 8948 22240 8957 22280
rect 11587 22240 11596 22280
rect 11636 22240 13036 22280
rect 13076 22240 13085 22280
rect 13230 22240 13324 22280
rect 13364 22240 13373 22280
rect 13699 22240 13708 22280
rect 13748 22240 16396 22280
rect 16436 22240 16445 22280
rect 0 22220 80 22240
rect 3331 22239 3389 22240
rect 4483 22239 4541 22240
rect 6124 22196 6164 22240
rect 1699 22156 1708 22196
rect 1748 22156 6164 22196
rect 6211 22156 6220 22196
rect 6260 22156 6700 22196
rect 6740 22156 6749 22196
rect 6796 22112 6836 22240
rect 13315 22239 13373 22240
rect 12163 22156 12172 22196
rect 12212 22156 12844 22196
rect 12884 22156 13228 22196
rect 13268 22156 13277 22196
rect 21424 22112 21504 22132
rect 4675 22072 4684 22112
rect 4724 22072 6836 22112
rect 8899 22072 8908 22112
rect 8948 22072 9388 22112
rect 9428 22072 9437 22112
rect 12547 22072 12556 22112
rect 12596 22072 16012 22112
rect 16052 22072 16061 22112
rect 17731 22072 17740 22112
rect 17780 22072 18604 22112
rect 18644 22072 18653 22112
rect 20140 22072 21504 22112
rect 12163 22028 12221 22029
rect 20140 22028 20180 22072
rect 21424 22052 21504 22072
rect 4771 21988 4780 22028
rect 4820 21988 6988 22028
rect 7028 21988 7037 22028
rect 12163 21988 12172 22028
rect 12212 21988 20180 22028
rect 12163 21987 12221 21988
rect 0 21944 80 21964
rect 7747 21944 7805 21945
rect 0 21904 2540 21944
rect 2947 21904 2956 21944
rect 2996 21904 4108 21944
rect 4148 21904 4157 21944
rect 4919 21904 4928 21944
rect 4968 21904 5010 21944
rect 5050 21904 5092 21944
rect 5132 21904 5174 21944
rect 5214 21904 5256 21944
rect 5296 21904 5305 21944
rect 6787 21904 6796 21944
rect 6836 21904 7756 21944
rect 7796 21904 7805 21944
rect 13123 21904 13132 21944
rect 13172 21904 13516 21944
rect 13556 21904 13565 21944
rect 20039 21904 20048 21944
rect 20088 21904 20130 21944
rect 20170 21904 20212 21944
rect 20252 21904 20294 21944
rect 20334 21904 20376 21944
rect 20416 21904 20425 21944
rect 0 21884 80 21904
rect 2500 21860 2540 21904
rect 7747 21903 7805 21904
rect 2500 21820 5548 21860
rect 5588 21820 5597 21860
rect 5923 21820 5932 21860
rect 5972 21820 6508 21860
rect 6548 21820 7372 21860
rect 7412 21820 7421 21860
rect 7555 21820 7564 21860
rect 7604 21820 7613 21860
rect 14083 21820 14092 21860
rect 14132 21820 16204 21860
rect 16244 21820 16253 21860
rect 16579 21820 16588 21860
rect 16628 21820 21484 21860
rect 3139 21736 3148 21776
rect 3188 21736 3532 21776
rect 3572 21736 3581 21776
rect 5155 21736 5164 21776
rect 5204 21736 6700 21776
rect 6740 21736 6749 21776
rect 3427 21692 3485 21693
rect 2755 21652 2764 21692
rect 2804 21652 3436 21692
rect 3476 21652 3724 21692
rect 3764 21652 3773 21692
rect 5347 21652 5356 21692
rect 5396 21652 7180 21692
rect 7220 21652 7229 21692
rect 3427 21651 3485 21652
rect 0 21608 80 21628
rect 1315 21608 1373 21609
rect 0 21568 268 21608
rect 308 21568 317 21608
rect 1315 21568 1324 21608
rect 1364 21568 1708 21608
rect 1748 21568 1757 21608
rect 2083 21568 2092 21608
rect 2132 21568 4204 21608
rect 4244 21568 4253 21608
rect 5155 21568 5164 21608
rect 5204 21568 5548 21608
rect 5588 21568 5597 21608
rect 5731 21568 5740 21608
rect 5780 21568 6316 21608
rect 6356 21568 6365 21608
rect 0 21548 80 21568
rect 1315 21567 1373 21568
rect 451 21524 509 21525
rect 451 21484 460 21524
rect 500 21484 5932 21524
rect 5972 21484 5981 21524
rect 451 21483 509 21484
rect 7564 21440 7604 21820
rect 12451 21736 12460 21776
rect 12500 21736 16492 21776
rect 16532 21736 18508 21776
rect 18548 21736 18557 21776
rect 8419 21692 8477 21693
rect 7651 21652 7660 21692
rect 7700 21652 7948 21692
rect 7988 21652 8428 21692
rect 8468 21652 8477 21692
rect 10435 21652 10444 21692
rect 10484 21652 11308 21692
rect 11348 21652 12652 21692
rect 12692 21652 14956 21692
rect 14996 21652 15005 21692
rect 15820 21652 19276 21692
rect 19316 21652 19325 21692
rect 8419 21651 8477 21652
rect 9187 21608 9245 21609
rect 9187 21568 9196 21608
rect 9236 21568 9388 21608
rect 9428 21568 9437 21608
rect 12739 21568 12748 21608
rect 12788 21568 13228 21608
rect 13268 21568 13277 21608
rect 13411 21568 13420 21608
rect 13460 21568 13612 21608
rect 13652 21568 15724 21608
rect 15764 21568 15773 21608
rect 9187 21567 9245 21568
rect 10147 21524 10205 21525
rect 15820 21524 15860 21652
rect 19363 21608 19421 21609
rect 21444 21608 21484 21820
rect 18979 21568 18988 21608
rect 19028 21568 19372 21608
rect 19412 21568 19421 21608
rect 19363 21567 19421 21568
rect 21292 21568 21484 21608
rect 9187 21484 9196 21524
rect 9236 21484 10156 21524
rect 10196 21484 10205 21524
rect 11395 21484 11404 21524
rect 11444 21484 12076 21524
rect 12116 21484 15860 21524
rect 16003 21484 16012 21524
rect 16052 21484 16588 21524
rect 16628 21484 16637 21524
rect 10147 21483 10205 21484
rect 21292 21440 21332 21568
rect 21424 21440 21504 21460
rect 2083 21400 2092 21440
rect 2132 21400 2860 21440
rect 2900 21400 2909 21440
rect 6019 21400 6028 21440
rect 6068 21400 7180 21440
rect 7220 21400 7229 21440
rect 7555 21400 7564 21440
rect 7604 21400 7613 21440
rect 12547 21400 12556 21440
rect 12596 21400 12844 21440
rect 12884 21400 12893 21440
rect 13411 21400 13420 21440
rect 13460 21400 13708 21440
rect 13748 21400 13757 21440
rect 16099 21400 16108 21440
rect 16148 21400 16396 21440
rect 16436 21400 16445 21440
rect 17155 21400 17164 21440
rect 17204 21400 17548 21440
rect 17588 21400 18028 21440
rect 18068 21400 18077 21440
rect 21292 21400 21504 21440
rect 21424 21380 21504 21400
rect 6595 21356 6653 21357
rect 9763 21356 9821 21357
rect 6595 21316 6604 21356
rect 6644 21316 6700 21356
rect 6740 21316 6749 21356
rect 9763 21316 9772 21356
rect 9812 21316 9868 21356
rect 9908 21316 9917 21356
rect 15427 21316 15436 21356
rect 15476 21316 16012 21356
rect 16052 21316 16061 21356
rect 6595 21315 6653 21316
rect 9763 21315 9821 21316
rect 0 21272 80 21292
rect 2083 21272 2141 21273
rect 0 21232 2092 21272
rect 2132 21232 7756 21272
rect 7796 21232 7805 21272
rect 8803 21232 8812 21272
rect 8852 21232 10828 21272
rect 10868 21232 10877 21272
rect 0 21212 80 21232
rect 2083 21231 2141 21232
rect 3679 21148 3688 21188
rect 3728 21148 3770 21188
rect 3810 21148 3852 21188
rect 3892 21148 3934 21188
rect 3974 21148 4016 21188
rect 4056 21148 4065 21188
rect 5347 21148 5356 21188
rect 5396 21148 10348 21188
rect 10388 21148 10397 21188
rect 18799 21148 18808 21188
rect 18848 21148 18890 21188
rect 18930 21148 18972 21188
rect 19012 21148 19054 21188
rect 19094 21148 19136 21188
rect 19176 21148 19185 21188
rect 18403 21104 18461 21105
rect 2755 21064 2764 21104
rect 2804 21064 7372 21104
rect 7412 21064 7421 21104
rect 10627 21064 10636 21104
rect 10676 21064 11308 21104
rect 11348 21064 11357 21104
rect 18115 21064 18124 21104
rect 18164 21064 18412 21104
rect 18452 21064 18461 21104
rect 18403 21063 18461 21064
rect 12643 21020 12701 21021
rect 3331 20980 3340 21020
rect 3380 20980 12652 21020
rect 12692 20980 14380 21020
rect 14420 20980 14429 21020
rect 12643 20979 12701 20980
rect 0 20936 80 20956
rect 0 20896 2956 20936
rect 2996 20896 3005 20936
rect 3427 20896 3436 20936
rect 3476 20896 3724 20936
rect 3764 20896 4684 20936
rect 4724 20896 5356 20936
rect 5396 20896 5405 20936
rect 6019 20896 6028 20936
rect 6068 20896 7084 20936
rect 7124 20896 7133 20936
rect 11320 20896 20180 20936
rect 0 20876 80 20896
rect 7843 20852 7901 20853
rect 3523 20812 3532 20852
rect 3572 20812 3916 20852
rect 3956 20812 5068 20852
rect 5108 20812 6988 20852
rect 7028 20812 7037 20852
rect 7758 20812 7852 20852
rect 7892 20812 7901 20852
rect 7843 20811 7901 20812
rect 3139 20768 3197 20769
rect 3427 20768 3485 20769
rect 1507 20728 1516 20768
rect 1556 20728 2668 20768
rect 2708 20728 2717 20768
rect 3139 20728 3148 20768
rect 3188 20728 3436 20768
rect 3476 20728 3485 20768
rect 3139 20727 3197 20728
rect 3427 20727 3485 20728
rect 4771 20768 4829 20769
rect 9475 20768 9533 20769
rect 4771 20728 4780 20768
rect 4820 20728 5164 20768
rect 5204 20728 5213 20768
rect 5347 20728 5356 20768
rect 5396 20728 5836 20768
rect 5876 20728 5885 20768
rect 9475 20728 9484 20768
rect 9524 20728 9580 20768
rect 9620 20728 9629 20768
rect 4771 20727 4829 20728
rect 9475 20727 9533 20728
rect 2755 20684 2813 20685
rect 11320 20684 11360 20896
rect 16204 20812 17164 20852
rect 17204 20812 17213 20852
rect 17347 20812 17356 20852
rect 17396 20812 18508 20852
rect 18548 20812 18557 20852
rect 12163 20768 12221 20769
rect 16204 20768 16244 20812
rect 20140 20768 20180 20896
rect 21424 20768 21504 20788
rect 12163 20728 12172 20768
rect 12212 20728 12268 20768
rect 12308 20728 12317 20768
rect 12643 20728 12652 20768
rect 12692 20728 13516 20768
rect 13556 20728 13565 20768
rect 13987 20728 13996 20768
rect 14036 20728 14764 20768
rect 14804 20728 14956 20768
rect 14996 20728 15628 20768
rect 15668 20728 15677 20768
rect 15811 20728 15820 20768
rect 15860 20728 16204 20768
rect 16244 20728 16253 20768
rect 16867 20728 16876 20768
rect 16916 20728 18124 20768
rect 18164 20728 18173 20768
rect 20140 20728 21504 20768
rect 12163 20727 12221 20728
rect 21424 20708 21504 20728
rect 748 20644 2540 20684
rect 0 20600 80 20620
rect 748 20600 788 20644
rect 0 20560 788 20600
rect 2500 20600 2540 20644
rect 2755 20644 2764 20684
rect 2804 20644 11360 20684
rect 16771 20644 16780 20684
rect 16820 20644 17548 20684
rect 17588 20644 17597 20684
rect 17827 20644 17836 20684
rect 17876 20644 18028 20684
rect 18068 20644 18077 20684
rect 2755 20643 2813 20644
rect 2500 20560 5780 20600
rect 6979 20560 6988 20600
rect 7028 20560 7276 20600
rect 7316 20560 7325 20600
rect 9571 20560 9580 20600
rect 9620 20560 9964 20600
rect 10004 20560 10013 20600
rect 10819 20560 10828 20600
rect 10868 20560 13996 20600
rect 14036 20560 14045 20600
rect 14467 20560 14476 20600
rect 14516 20560 14764 20600
rect 14804 20560 14813 20600
rect 16963 20560 16972 20600
rect 17012 20560 18700 20600
rect 18740 20560 18749 20600
rect 0 20540 80 20560
rect 5740 20516 5780 20560
rect 1315 20476 1324 20516
rect 1364 20476 5644 20516
rect 5684 20476 5693 20516
rect 5740 20476 10636 20516
rect 10676 20476 10685 20516
rect 16291 20476 16300 20516
rect 16340 20476 17164 20516
rect 17204 20476 17213 20516
rect 17731 20476 17740 20516
rect 17780 20476 18124 20516
rect 18164 20476 18173 20516
rect 6499 20432 6557 20433
rect 18403 20432 18461 20433
rect 4919 20392 4928 20432
rect 4968 20392 5010 20432
rect 5050 20392 5092 20432
rect 5132 20392 5174 20432
rect 5214 20392 5256 20432
rect 5296 20392 5305 20432
rect 5347 20392 5356 20432
rect 5396 20392 6508 20432
rect 6548 20392 6557 20432
rect 6787 20392 6796 20432
rect 6836 20392 8716 20432
rect 8756 20392 8765 20432
rect 18318 20392 18412 20432
rect 18452 20392 18461 20432
rect 20039 20392 20048 20432
rect 20088 20392 20130 20432
rect 20170 20392 20212 20432
rect 20252 20392 20294 20432
rect 20334 20392 20376 20432
rect 20416 20392 20425 20432
rect 6499 20391 6557 20392
rect 18403 20391 18461 20392
rect 2947 20308 2956 20348
rect 2996 20308 9868 20348
rect 9908 20308 9917 20348
rect 17347 20308 17356 20348
rect 17396 20308 18316 20348
rect 18356 20308 18365 20348
rect 0 20264 80 20284
rect 3043 20264 3101 20265
rect 0 20224 3052 20264
rect 3092 20224 3101 20264
rect 0 20204 80 20224
rect 3043 20223 3101 20224
rect 4396 20224 5684 20264
rect 18019 20224 18028 20264
rect 18068 20224 18356 20264
rect 3523 20096 3581 20097
rect 4396 20096 4436 20224
rect 4771 20180 4829 20181
rect 4771 20140 4780 20180
rect 4820 20140 4876 20180
rect 4916 20140 4925 20180
rect 4771 20139 4829 20140
rect 5644 20096 5684 20224
rect 18316 20180 18356 20224
rect 12259 20140 12268 20180
rect 12308 20140 12652 20180
rect 12692 20140 12701 20180
rect 14148 20140 14188 20180
rect 14228 20140 14237 20180
rect 18307 20140 18316 20180
rect 18356 20140 18365 20180
rect 10147 20096 10205 20097
rect 14188 20096 14228 20140
rect 18019 20096 18077 20097
rect 21424 20096 21504 20116
rect 3523 20056 3532 20096
rect 3572 20056 4436 20096
rect 4483 20056 4492 20096
rect 4532 20056 5548 20096
rect 5588 20056 5597 20096
rect 5644 20056 7468 20096
rect 7508 20056 9100 20096
rect 9140 20056 10156 20096
rect 10196 20056 10205 20096
rect 11395 20056 11404 20096
rect 11444 20056 14380 20096
rect 14420 20056 14429 20096
rect 17059 20056 17068 20096
rect 17108 20056 17740 20096
rect 17780 20056 17789 20096
rect 18019 20056 18028 20096
rect 18068 20056 21504 20096
rect 3523 20055 3581 20056
rect 10147 20055 10205 20056
rect 18019 20055 18077 20056
rect 21424 20036 21504 20056
rect 5635 20012 5693 20013
rect 8707 20012 8765 20013
rect 11875 20012 11933 20013
rect 3427 19972 3436 20012
rect 3476 19972 4396 20012
rect 4436 19972 4445 20012
rect 5251 19972 5260 20012
rect 5300 19972 5644 20012
rect 5684 19972 5693 20012
rect 7555 19972 7564 20012
rect 7604 19972 8428 20012
rect 8468 19972 8477 20012
rect 8622 19972 8716 20012
rect 8756 19972 8765 20012
rect 11790 19972 11884 20012
rect 11924 19972 11933 20012
rect 5635 19971 5693 19972
rect 8707 19971 8765 19972
rect 11875 19971 11933 19972
rect 12163 20012 12221 20013
rect 12163 19972 12172 20012
rect 12212 19972 12268 20012
rect 12308 19972 12317 20012
rect 14083 19972 14092 20012
rect 14132 19972 14141 20012
rect 16867 19972 16876 20012
rect 16916 19972 17836 20012
rect 17876 19972 17885 20012
rect 12163 19971 12221 19972
rect 0 19928 80 19948
rect 14092 19928 14132 19972
rect 0 19888 1612 19928
rect 1652 19888 1661 19928
rect 4675 19888 4684 19928
rect 4724 19888 6220 19928
rect 6260 19888 6269 19928
rect 12163 19888 12172 19928
rect 12212 19888 12364 19928
rect 12404 19888 12413 19928
rect 13987 19888 13996 19928
rect 14036 19888 14132 19928
rect 0 19868 80 19888
rect 12547 19844 12605 19845
rect 1699 19804 1708 19844
rect 1748 19804 1940 19844
rect 2467 19804 2476 19844
rect 2516 19804 6796 19844
rect 6836 19804 6845 19844
rect 10147 19804 10156 19844
rect 10196 19804 10636 19844
rect 10676 19804 10685 19844
rect 12462 19804 12556 19844
rect 12596 19804 12605 19844
rect 14467 19804 14476 19844
rect 14516 19804 15820 19844
rect 15860 19804 15869 19844
rect 17347 19804 17356 19844
rect 17396 19804 18604 19844
rect 18644 19804 18653 19844
rect 1900 19760 1940 19804
rect 12547 19803 12605 19804
rect 6115 19760 6173 19761
rect 1315 19720 1324 19760
rect 1364 19720 1804 19760
rect 1844 19720 1853 19760
rect 1900 19720 4148 19760
rect 5443 19720 5452 19760
rect 5492 19720 6124 19760
rect 6164 19720 7084 19760
rect 7124 19720 16876 19760
rect 16916 19720 16925 19760
rect 4108 19676 4148 19720
rect 6115 19719 6173 19720
rect 8803 19676 8861 19677
rect 9187 19676 9245 19677
rect 3679 19636 3688 19676
rect 3728 19636 3770 19676
rect 3810 19636 3852 19676
rect 3892 19636 3934 19676
rect 3974 19636 4016 19676
rect 4056 19636 4065 19676
rect 4108 19636 5740 19676
rect 5780 19636 5789 19676
rect 6595 19636 6604 19676
rect 6644 19636 6796 19676
rect 6836 19636 6845 19676
rect 8803 19636 8812 19676
rect 8852 19636 9196 19676
rect 9236 19636 9524 19676
rect 10243 19636 10252 19676
rect 10292 19636 14380 19676
rect 14420 19636 14429 19676
rect 18799 19636 18808 19676
rect 18848 19636 18890 19676
rect 18930 19636 18972 19676
rect 19012 19636 19054 19676
rect 19094 19636 19136 19676
rect 19176 19636 19185 19676
rect 8803 19635 8861 19636
rect 9187 19635 9245 19636
rect 0 19592 80 19612
rect 9484 19592 9524 19636
rect 0 19552 9388 19592
rect 9428 19552 9437 19592
rect 9484 19552 15628 19592
rect 15668 19552 15677 19592
rect 0 19532 80 19552
rect 2755 19468 2764 19508
rect 2804 19468 3052 19508
rect 3092 19468 3101 19508
rect 5635 19468 5644 19508
rect 5684 19468 11212 19508
rect 11252 19468 11261 19508
rect 3139 19424 3197 19425
rect 10051 19424 10109 19425
rect 21424 19424 21504 19444
rect 2563 19384 2572 19424
rect 2612 19384 2956 19424
rect 2996 19384 3005 19424
rect 3139 19384 3148 19424
rect 3188 19384 9100 19424
rect 9140 19384 9149 19424
rect 10051 19384 10060 19424
rect 10100 19384 21504 19424
rect 3139 19383 3197 19384
rect 10051 19383 10109 19384
rect 21424 19364 21504 19384
rect 4195 19340 4253 19341
rect 6307 19340 6365 19341
rect 6499 19340 6557 19341
rect 4110 19300 4204 19340
rect 4244 19300 6260 19340
rect 4195 19299 4253 19300
rect 0 19256 80 19276
rect 4387 19256 4445 19257
rect 6220 19256 6260 19300
rect 6307 19300 6316 19340
rect 6356 19300 6508 19340
rect 6548 19300 6557 19340
rect 6691 19300 6700 19340
rect 6740 19300 7372 19340
rect 7412 19300 7421 19340
rect 13315 19300 13324 19340
rect 13364 19300 13612 19340
rect 13652 19300 13661 19340
rect 13987 19300 13996 19340
rect 14036 19300 14284 19340
rect 14324 19300 14333 19340
rect 16867 19300 16876 19340
rect 16916 19300 18700 19340
rect 18740 19300 18749 19340
rect 6307 19299 6365 19300
rect 6499 19299 6557 19300
rect 6979 19256 7037 19257
rect 0 19216 4396 19256
rect 4436 19216 4445 19256
rect 5251 19216 5260 19256
rect 5300 19216 6124 19256
rect 6164 19216 6173 19256
rect 6220 19216 6316 19256
rect 6356 19216 6365 19256
rect 6595 19216 6604 19256
rect 6644 19216 6988 19256
rect 7028 19216 7037 19256
rect 7651 19216 7660 19256
rect 7700 19216 8332 19256
rect 8372 19216 8381 19256
rect 13507 19216 13516 19256
rect 13556 19216 14188 19256
rect 14228 19216 14237 19256
rect 17443 19216 17452 19256
rect 17492 19216 17501 19256
rect 0 19196 80 19216
rect 4387 19215 4445 19216
rect 6979 19215 7037 19216
rect 17452 19172 17492 19216
rect 6019 19132 6028 19172
rect 6068 19132 6700 19172
rect 6740 19132 6749 19172
rect 11203 19132 11212 19172
rect 11252 19132 12556 19172
rect 12596 19132 17492 19172
rect 10339 19088 10397 19089
rect 14755 19088 14813 19089
rect 5635 19048 5644 19088
rect 5684 19048 5932 19088
rect 5972 19048 5981 19088
rect 10254 19048 10348 19088
rect 10388 19048 10397 19088
rect 13891 19048 13900 19088
rect 13940 19048 14764 19088
rect 14804 19048 14813 19088
rect 10339 19047 10397 19048
rect 14755 19047 14813 19048
rect 14860 19048 17356 19088
rect 17396 19048 17405 19088
rect 18595 19048 18604 19088
rect 18644 19048 18892 19088
rect 18932 19048 18941 19088
rect 5347 19004 5405 19005
rect 8803 19004 8861 19005
rect 14860 19004 14900 19048
rect 5347 18964 5356 19004
rect 5396 18964 8812 19004
rect 8852 18964 8861 19004
rect 12451 18964 12460 19004
rect 12500 18964 13708 19004
rect 13748 18964 14900 19004
rect 15715 18964 15724 19004
rect 15764 18964 16300 19004
rect 16340 18964 16349 19004
rect 5347 18963 5405 18964
rect 8803 18963 8861 18964
rect 0 18920 80 18940
rect 3043 18920 3101 18921
rect 5923 18920 5981 18921
rect 8035 18920 8093 18921
rect 0 18880 172 18920
rect 212 18880 221 18920
rect 3043 18880 3052 18920
rect 3092 18880 3148 18920
rect 3188 18880 3197 18920
rect 4919 18880 4928 18920
rect 4968 18880 5010 18920
rect 5050 18880 5092 18920
rect 5132 18880 5174 18920
rect 5214 18880 5256 18920
rect 5296 18880 5305 18920
rect 5635 18880 5644 18920
rect 5684 18880 5932 18920
rect 5972 18880 5981 18920
rect 0 18860 80 18880
rect 3043 18879 3101 18880
rect 5923 18879 5981 18880
rect 6508 18880 7180 18920
rect 7220 18880 7229 18920
rect 8035 18880 8044 18920
rect 8084 18880 9196 18920
rect 9236 18880 9245 18920
rect 9292 18880 12748 18920
rect 12788 18880 12797 18920
rect 14563 18880 14572 18920
rect 14612 18880 15628 18920
rect 15668 18880 15677 18920
rect 20039 18880 20048 18920
rect 20088 18880 20130 18920
rect 20170 18880 20212 18920
rect 20252 18880 20294 18920
rect 20334 18880 20376 18920
rect 20416 18880 20425 18920
rect 6508 18836 6548 18880
rect 8035 18879 8093 18880
rect 6787 18836 6845 18837
rect 9292 18836 9332 18880
rect 11107 18836 11165 18837
rect 13795 18836 13853 18837
rect 15427 18836 15485 18837
rect 4771 18796 4780 18836
rect 4820 18796 6548 18836
rect 6595 18796 6604 18836
rect 6644 18796 6796 18836
rect 6836 18796 6845 18836
rect 8803 18796 8812 18836
rect 8852 18796 9332 18836
rect 10540 18796 10924 18836
rect 10964 18796 10973 18836
rect 11107 18796 11116 18836
rect 11156 18796 11250 18836
rect 12643 18796 12652 18836
rect 12692 18796 13804 18836
rect 13844 18796 13853 18836
rect 15342 18796 15436 18836
rect 15476 18796 15485 18836
rect 6787 18795 6845 18796
rect 2563 18712 2572 18752
rect 2612 18712 3340 18752
rect 3380 18712 3389 18752
rect 5539 18712 5548 18752
rect 5588 18712 6796 18752
rect 6836 18712 6845 18752
rect 7843 18668 7901 18669
rect 460 18628 7852 18668
rect 7892 18628 7901 18668
rect 0 18584 80 18604
rect 460 18584 500 18628
rect 7843 18627 7901 18628
rect 4579 18584 4637 18585
rect 0 18544 500 18584
rect 1795 18544 1804 18584
rect 1844 18544 4300 18584
rect 4340 18544 4588 18584
rect 4628 18544 4637 18584
rect 5347 18544 5356 18584
rect 5396 18544 5548 18584
rect 5588 18544 5597 18584
rect 6115 18544 6124 18584
rect 6164 18544 6412 18584
rect 6452 18544 6796 18584
rect 6836 18544 6845 18584
rect 7075 18544 7084 18584
rect 7124 18544 9580 18584
rect 9620 18544 9629 18584
rect 0 18524 80 18544
rect 4579 18543 4637 18544
rect 10540 18500 10580 18796
rect 11107 18795 11165 18796
rect 13795 18795 13853 18796
rect 15427 18795 15485 18796
rect 21424 18752 21504 18772
rect 11011 18712 11020 18752
rect 11060 18712 11069 18752
rect 13027 18712 13036 18752
rect 13076 18712 13804 18752
rect 13844 18712 13853 18752
rect 15907 18712 15916 18752
rect 15956 18712 16204 18752
rect 16244 18712 16253 18752
rect 18499 18712 18508 18752
rect 18548 18712 21504 18752
rect 11020 18668 11060 18712
rect 21424 18692 21504 18712
rect 12163 18668 12221 18669
rect 17443 18668 17501 18669
rect 11020 18628 11212 18668
rect 11252 18628 11261 18668
rect 12163 18628 12172 18668
rect 12212 18628 12748 18668
rect 12788 18628 12797 18668
rect 17443 18628 17452 18668
rect 17492 18628 17548 18668
rect 17588 18628 17597 18668
rect 12163 18627 12221 18628
rect 17443 18627 17501 18628
rect 16963 18584 17021 18585
rect 10627 18544 10636 18584
rect 10676 18544 13804 18584
rect 13844 18544 13853 18584
rect 16963 18544 16972 18584
rect 17012 18544 20620 18584
rect 20660 18544 20669 18584
rect 16963 18543 17021 18544
rect 5740 18460 6028 18500
rect 6068 18460 6077 18500
rect 10051 18460 10060 18500
rect 10100 18460 11596 18500
rect 11636 18460 11645 18500
rect 5740 18416 5780 18460
rect 5731 18376 5740 18416
rect 5780 18376 5789 18416
rect 5923 18376 5932 18416
rect 5972 18376 8812 18416
rect 8852 18376 8861 18416
rect 4099 18292 4108 18332
rect 4148 18292 7084 18332
rect 7124 18292 7133 18332
rect 14851 18292 14860 18332
rect 14900 18292 15244 18332
rect 15284 18292 15293 18332
rect 0 18248 80 18268
rect 10147 18248 10205 18249
rect 0 18208 9484 18248
rect 9524 18208 9964 18248
rect 10004 18208 10013 18248
rect 10147 18208 10156 18248
rect 10196 18208 10732 18248
rect 10772 18208 15628 18248
rect 15668 18208 15677 18248
rect 0 18188 80 18208
rect 10147 18207 10205 18208
rect 16675 18164 16733 18165
rect 3331 18124 3340 18164
rect 3380 18124 3532 18164
rect 3572 18124 3581 18164
rect 3679 18124 3688 18164
rect 3728 18124 3770 18164
rect 3810 18124 3852 18164
rect 3892 18124 3934 18164
rect 3974 18124 4016 18164
rect 4056 18124 4065 18164
rect 7267 18124 7276 18164
rect 7316 18124 11596 18164
rect 11636 18124 11645 18164
rect 12739 18124 12748 18164
rect 12788 18124 14956 18164
rect 14996 18124 16684 18164
rect 16724 18124 16733 18164
rect 18799 18124 18808 18164
rect 18848 18124 18890 18164
rect 18930 18124 18972 18164
rect 19012 18124 19054 18164
rect 19094 18124 19136 18164
rect 19176 18124 19185 18164
rect 16675 18123 16733 18124
rect 7459 18080 7517 18081
rect 10051 18080 10109 18081
rect 21424 18080 21504 18100
rect 2947 18040 2956 18080
rect 2996 18040 4684 18080
rect 4724 18040 7468 18080
rect 7508 18040 9676 18080
rect 9716 18040 9725 18080
rect 10051 18040 10060 18080
rect 10100 18040 12652 18080
rect 12692 18040 12701 18080
rect 21379 18040 21388 18080
rect 21428 18040 21504 18080
rect 7459 18039 7517 18040
rect 10051 18039 10109 18040
rect 21424 18020 21504 18040
rect 1315 17956 1324 17996
rect 1364 17956 3628 17996
rect 3668 17956 6892 17996
rect 6932 17956 6941 17996
rect 7075 17956 7084 17996
rect 7124 17956 7564 17996
rect 7604 17956 7613 17996
rect 8131 17956 8140 17996
rect 8180 17956 8524 17996
rect 8564 17956 8573 17996
rect 10147 17956 10156 17996
rect 10196 17956 10292 17996
rect 12547 17956 12556 17996
rect 12596 17956 12940 17996
rect 12980 17956 12989 17996
rect 14947 17956 14956 17996
rect 14996 17956 15724 17996
rect 15764 17956 15773 17996
rect 0 17912 80 17932
rect 0 17872 10060 17912
rect 10100 17872 10109 17912
rect 0 17852 80 17872
rect 3139 17828 3197 17829
rect 4483 17828 4541 17829
rect 10051 17828 10109 17829
rect 10252 17828 10292 17956
rect 15235 17872 15244 17912
rect 15284 17872 15820 17912
rect 15860 17872 15869 17912
rect 3139 17788 3148 17828
rect 3188 17788 3244 17828
rect 3284 17788 3293 17828
rect 4483 17788 4492 17828
rect 4532 17788 8908 17828
rect 8948 17788 10060 17828
rect 10100 17788 10109 17828
rect 10243 17788 10252 17828
rect 10292 17788 10301 17828
rect 10531 17788 10540 17828
rect 10580 17788 11404 17828
rect 11444 17788 12748 17828
rect 12788 17788 12797 17828
rect 15427 17788 15436 17828
rect 15476 17788 15485 17828
rect 3139 17787 3197 17788
rect 4483 17787 4541 17788
rect 10051 17787 10109 17788
rect 8707 17744 8765 17745
rect 10540 17744 10580 17788
rect 1507 17704 1516 17744
rect 1556 17704 2540 17744
rect 3715 17704 3724 17744
rect 3764 17704 5644 17744
rect 5684 17704 5693 17744
rect 8515 17704 8524 17744
rect 8564 17704 8716 17744
rect 8756 17704 8765 17744
rect 2500 17660 2540 17704
rect 8707 17703 8765 17704
rect 8812 17704 10156 17744
rect 10196 17704 10580 17744
rect 11587 17704 11596 17744
rect 11636 17704 12172 17744
rect 12212 17704 13516 17744
rect 13556 17704 13565 17744
rect 3043 17660 3101 17661
rect 8716 17660 8756 17703
rect 8812 17660 8852 17704
rect 15436 17660 15476 17788
rect 16003 17704 16012 17744
rect 16052 17704 17644 17744
rect 17684 17704 17693 17744
rect 2500 17620 2668 17660
rect 2708 17620 2860 17660
rect 2900 17620 2909 17660
rect 3043 17620 3052 17660
rect 3092 17620 3186 17660
rect 8716 17620 8812 17660
rect 8852 17620 8880 17660
rect 9283 17620 9292 17660
rect 9332 17620 9676 17660
rect 9716 17620 11360 17660
rect 14659 17620 14668 17660
rect 14708 17620 15476 17660
rect 18499 17620 18508 17660
rect 18548 17620 19084 17660
rect 19124 17620 19133 17660
rect 3043 17619 3101 17620
rect 0 17576 80 17596
rect 4387 17576 4445 17577
rect 0 17536 4396 17576
rect 4436 17536 4445 17576
rect 0 17516 80 17536
rect 4387 17535 4445 17536
rect 4579 17576 4637 17577
rect 5731 17576 5789 17577
rect 11320 17576 11360 17620
rect 4579 17536 4588 17576
rect 4628 17536 5260 17576
rect 5300 17536 5309 17576
rect 5731 17536 5740 17576
rect 5780 17536 9100 17576
rect 9140 17536 9149 17576
rect 11320 17536 13132 17576
rect 13172 17536 13181 17576
rect 15139 17536 15148 17576
rect 15188 17536 15916 17576
rect 15956 17536 15965 17576
rect 16483 17536 16492 17576
rect 16532 17536 16876 17576
rect 16916 17536 18892 17576
rect 18932 17536 19276 17576
rect 19316 17536 19325 17576
rect 4579 17535 4637 17536
rect 5731 17535 5789 17536
rect 2947 17492 3005 17493
rect 1795 17452 1804 17492
rect 1844 17452 2540 17492
rect 2862 17452 2956 17492
rect 2996 17452 3005 17492
rect 2500 17408 2540 17452
rect 2947 17451 3005 17452
rect 5347 17492 5405 17493
rect 5347 17452 5356 17492
rect 5396 17452 5490 17492
rect 11491 17452 11500 17492
rect 11540 17452 19372 17492
rect 19412 17452 19421 17492
rect 5347 17451 5405 17452
rect 3427 17408 3485 17409
rect 16483 17408 16541 17409
rect 21424 17408 21504 17428
rect 2500 17368 3436 17408
rect 3476 17368 3485 17408
rect 4919 17368 4928 17408
rect 4968 17368 5010 17408
rect 5050 17368 5092 17408
rect 5132 17368 5174 17408
rect 5214 17368 5256 17408
rect 5296 17368 5305 17408
rect 10531 17368 10540 17408
rect 10580 17368 11212 17408
rect 11252 17368 16492 17408
rect 16532 17368 16684 17408
rect 16724 17368 16733 17408
rect 20039 17368 20048 17408
rect 20088 17368 20130 17408
rect 20170 17368 20212 17408
rect 20252 17368 20294 17408
rect 20334 17368 20376 17408
rect 20416 17368 20425 17408
rect 20524 17368 21504 17408
rect 3427 17367 3485 17368
rect 16483 17367 16541 17368
rect 3436 17324 3476 17367
rect 8899 17324 8957 17325
rect 20524 17324 20564 17368
rect 21424 17348 21504 17368
rect 2851 17284 2860 17324
rect 2900 17284 3244 17324
rect 3284 17284 3293 17324
rect 3436 17284 6028 17324
rect 6068 17284 6077 17324
rect 8899 17284 8908 17324
rect 8948 17284 20564 17324
rect 8899 17283 8957 17284
rect 0 17240 80 17260
rect 15427 17240 15485 17241
rect 0 17200 8716 17240
rect 8756 17200 8765 17240
rect 8812 17200 11500 17240
rect 11540 17200 11549 17240
rect 15342 17200 15436 17240
rect 15476 17200 15485 17240
rect 0 17180 80 17200
rect 8812 17156 8852 17200
rect 15427 17199 15485 17200
rect 1603 17116 1612 17156
rect 1652 17116 2572 17156
rect 2612 17116 2956 17156
rect 2996 17116 3005 17156
rect 4771 17116 4780 17156
rect 4820 17116 5164 17156
rect 5204 17116 5213 17156
rect 8419 17116 8428 17156
rect 8468 17116 8852 17156
rect 9091 17116 9100 17156
rect 9140 17116 9388 17156
rect 9428 17116 9437 17156
rect 10915 17116 10924 17156
rect 10964 17116 11308 17156
rect 11348 17116 11357 17156
rect 15907 17116 15916 17156
rect 15956 17116 16204 17156
rect 16244 17116 18700 17156
rect 18740 17116 18749 17156
rect 3043 17072 3101 17073
rect 4099 17072 4157 17073
rect 5347 17072 5405 17073
rect 7651 17072 7709 17073
rect 7843 17072 7901 17073
rect 14755 17072 14813 17073
rect 1411 17032 1420 17072
rect 1460 17032 2860 17072
rect 2900 17032 2909 17072
rect 3043 17032 3052 17072
rect 3092 17032 4108 17072
rect 4148 17032 4972 17072
rect 5012 17032 5021 17072
rect 5262 17032 5356 17072
rect 5396 17032 6892 17072
rect 6932 17032 7276 17072
rect 7316 17032 7325 17072
rect 7566 17032 7660 17072
rect 7700 17032 7852 17072
rect 7892 17032 7901 17072
rect 9475 17032 9484 17072
rect 9524 17032 13516 17072
rect 13556 17032 13565 17072
rect 14755 17032 14764 17072
rect 14804 17032 15244 17072
rect 15284 17032 15293 17072
rect 17059 17032 17068 17072
rect 17108 17032 17117 17072
rect 3043 17031 3101 17032
rect 4099 17031 4157 17032
rect 5347 17031 5405 17032
rect 7651 17031 7709 17032
rect 7843 17031 7901 17032
rect 14755 17031 14813 17032
rect 6787 16988 6845 16989
rect 17068 16988 17108 17032
rect 5827 16948 5836 16988
rect 5876 16948 6796 16988
rect 6836 16948 6845 16988
rect 14563 16948 14572 16988
rect 14612 16948 14956 16988
rect 14996 16948 15005 16988
rect 16771 16948 16780 16988
rect 16820 16948 17108 16988
rect 6787 16947 6845 16948
rect 0 16904 80 16924
rect 16675 16904 16733 16905
rect 0 16864 11020 16904
rect 11060 16864 11069 16904
rect 14179 16864 14188 16904
rect 14228 16864 14860 16904
rect 14900 16864 16204 16904
rect 16244 16864 16253 16904
rect 16675 16864 16684 16904
rect 16724 16864 16876 16904
rect 16916 16864 16925 16904
rect 17827 16864 17836 16904
rect 17876 16864 18508 16904
rect 18548 16864 18557 16904
rect 0 16844 80 16864
rect 16675 16863 16733 16864
rect 6307 16820 6365 16821
rect 1219 16780 1228 16820
rect 1268 16780 3724 16820
rect 3764 16780 3773 16820
rect 4003 16780 4012 16820
rect 4052 16780 4300 16820
rect 4340 16780 4349 16820
rect 6222 16780 6316 16820
rect 6356 16780 6365 16820
rect 6307 16779 6365 16780
rect 6595 16820 6653 16821
rect 6595 16780 6604 16820
rect 6644 16780 6892 16820
rect 6932 16780 6941 16820
rect 12355 16780 12364 16820
rect 12404 16780 14228 16820
rect 14563 16780 14572 16820
rect 14612 16780 15052 16820
rect 15092 16780 15101 16820
rect 6595 16779 6653 16780
rect 5539 16736 5597 16737
rect 14188 16736 14228 16780
rect 21424 16736 21504 16756
rect 5539 16696 5548 16736
rect 5588 16696 12748 16736
rect 12788 16696 12797 16736
rect 14188 16696 21504 16736
rect 5539 16695 5597 16696
rect 21424 16676 21504 16696
rect 8035 16652 8093 16653
rect 3679 16612 3688 16652
rect 3728 16612 3770 16652
rect 3810 16612 3852 16652
rect 3892 16612 3934 16652
rect 3974 16612 4016 16652
rect 4056 16612 4065 16652
rect 4579 16612 4588 16652
rect 4628 16612 5548 16652
rect 5588 16612 5597 16652
rect 6019 16612 6028 16652
rect 6068 16612 8044 16652
rect 8084 16612 8428 16652
rect 8468 16612 8477 16652
rect 18799 16612 18808 16652
rect 18848 16612 18890 16652
rect 18930 16612 18972 16652
rect 19012 16612 19054 16652
rect 19094 16612 19136 16652
rect 19176 16612 19185 16652
rect 8035 16611 8093 16612
rect 0 16568 80 16588
rect 0 16528 9484 16568
rect 9524 16528 9533 16568
rect 0 16508 80 16528
rect 1891 16444 1900 16484
rect 1940 16444 2284 16484
rect 2324 16444 4108 16484
rect 4148 16444 9676 16484
rect 9716 16444 9725 16484
rect 15139 16444 15148 16484
rect 15188 16444 16300 16484
rect 16340 16444 16349 16484
rect 2467 16400 2525 16401
rect 3331 16400 3389 16401
rect 2467 16360 2476 16400
rect 2516 16360 2860 16400
rect 2900 16360 2909 16400
rect 3246 16360 3340 16400
rect 3380 16360 3389 16400
rect 4771 16360 4780 16400
rect 4820 16360 8044 16400
rect 8084 16360 8093 16400
rect 16195 16360 16204 16400
rect 16244 16360 17836 16400
rect 17876 16360 17885 16400
rect 2467 16359 2525 16360
rect 3331 16359 3389 16360
rect 6499 16276 6508 16316
rect 6548 16276 9868 16316
rect 9908 16276 9917 16316
rect 16387 16276 16396 16316
rect 16436 16276 16684 16316
rect 16724 16276 16733 16316
rect 0 16232 80 16252
rect 12835 16232 12893 16233
rect 0 16192 2764 16232
rect 2804 16192 2813 16232
rect 3139 16192 3148 16232
rect 3188 16192 3340 16232
rect 3380 16192 3389 16232
rect 3523 16192 3532 16232
rect 3572 16192 4300 16232
rect 4340 16192 4349 16232
rect 5923 16192 5932 16232
rect 5972 16192 9772 16232
rect 9812 16192 9821 16232
rect 10051 16192 10060 16232
rect 10100 16192 10348 16232
rect 10388 16192 10397 16232
rect 12835 16192 12844 16232
rect 12884 16192 17740 16232
rect 17780 16192 18028 16232
rect 18068 16192 18077 16232
rect 0 16172 80 16192
rect 12835 16191 12893 16192
rect 8899 16148 8957 16149
rect 6307 16108 6316 16148
rect 6356 16108 6508 16148
rect 6548 16108 6557 16148
rect 7075 16108 7084 16148
rect 7124 16108 8908 16148
rect 8948 16108 9388 16148
rect 9428 16108 9437 16148
rect 17251 16108 17260 16148
rect 17300 16108 17548 16148
rect 17588 16108 17597 16148
rect 8899 16107 8957 16108
rect 10147 16064 10205 16065
rect 21424 16064 21504 16084
rect 10147 16024 10156 16064
rect 10196 16024 11020 16064
rect 11060 16024 11069 16064
rect 20611 16024 20620 16064
rect 20660 16024 21504 16064
rect 10147 16023 10205 16024
rect 21424 16004 21504 16024
rect 6403 15940 6412 15980
rect 6452 15940 7468 15980
rect 7508 15940 8908 15980
rect 8948 15940 10156 15980
rect 10196 15940 10205 15980
rect 0 15896 80 15916
rect 0 15856 1516 15896
rect 1556 15856 1565 15896
rect 4919 15856 4928 15896
rect 4968 15856 5010 15896
rect 5050 15856 5092 15896
rect 5132 15856 5174 15896
rect 5214 15856 5256 15896
rect 5296 15856 5305 15896
rect 7363 15856 7372 15896
rect 7412 15856 8044 15896
rect 8084 15856 8236 15896
rect 8276 15856 8285 15896
rect 13123 15856 13132 15896
rect 13172 15856 13420 15896
rect 13460 15856 13469 15896
rect 20039 15856 20048 15896
rect 20088 15856 20130 15896
rect 20170 15856 20212 15896
rect 20252 15856 20294 15896
rect 20334 15856 20376 15896
rect 20416 15856 20425 15896
rect 0 15836 80 15856
rect 4291 15772 4300 15812
rect 4340 15772 5932 15812
rect 5972 15772 5981 15812
rect 12259 15772 12268 15812
rect 12308 15772 13996 15812
rect 14036 15772 14045 15812
rect 4291 15728 4349 15729
rect 2467 15688 2476 15728
rect 2516 15688 2764 15728
rect 2804 15688 3052 15728
rect 3092 15688 3101 15728
rect 3966 15688 3975 15728
rect 4015 15688 4300 15728
rect 4340 15688 4396 15728
rect 4436 15688 4445 15728
rect 11320 15688 14092 15728
rect 14132 15688 14141 15728
rect 4291 15687 4349 15688
rect 1603 15604 1612 15644
rect 1652 15604 7564 15644
rect 7604 15604 7613 15644
rect 0 15560 80 15580
rect 11320 15560 11360 15688
rect 15715 15560 15773 15561
rect 0 15520 1708 15560
rect 1748 15520 1757 15560
rect 3139 15520 3148 15560
rect 3188 15520 3820 15560
rect 3860 15520 3869 15560
rect 3916 15520 11360 15560
rect 11875 15520 11884 15560
rect 11924 15520 12748 15560
rect 12788 15520 13708 15560
rect 13748 15520 13757 15560
rect 15715 15520 15724 15560
rect 15764 15520 16588 15560
rect 16628 15520 16637 15560
rect 0 15500 80 15520
rect 3331 15436 3340 15476
rect 3380 15436 3532 15476
rect 3572 15436 3581 15476
rect 3916 15392 3956 15520
rect 15715 15519 15773 15520
rect 12835 15476 12893 15477
rect 4387 15436 4396 15476
rect 4436 15436 11360 15476
rect 11683 15436 11692 15476
rect 11732 15436 12076 15476
rect 12116 15436 12125 15476
rect 12750 15436 12844 15476
rect 12884 15436 12893 15476
rect 11320 15392 11360 15436
rect 12835 15435 12893 15436
rect 21424 15392 21504 15412
rect 2500 15352 3956 15392
rect 6691 15352 6700 15392
rect 6740 15352 6988 15392
rect 7028 15352 7037 15392
rect 11320 15352 15244 15392
rect 15284 15352 15293 15392
rect 21283 15352 21292 15392
rect 21332 15352 21504 15392
rect 2500 15308 2540 15352
rect 21424 15332 21504 15352
rect 3427 15308 3485 15309
rect 9187 15308 9245 15309
rect 1891 15268 1900 15308
rect 1940 15268 2540 15308
rect 3342 15268 3436 15308
rect 3476 15268 3485 15308
rect 5251 15268 5260 15308
rect 5300 15268 8428 15308
rect 8468 15268 9196 15308
rect 9236 15268 9245 15308
rect 12643 15268 12652 15308
rect 12692 15268 13612 15308
rect 13652 15268 14284 15308
rect 14324 15268 14333 15308
rect 15043 15268 15052 15308
rect 15092 15268 15724 15308
rect 15764 15268 15773 15308
rect 16579 15268 16588 15308
rect 16628 15268 17068 15308
rect 17108 15268 17117 15308
rect 3427 15267 3485 15268
rect 9187 15267 9245 15268
rect 0 15224 80 15244
rect 0 15184 1324 15224
rect 1364 15184 1373 15224
rect 1603 15184 1612 15224
rect 1652 15184 6796 15224
rect 6836 15184 6845 15224
rect 7651 15184 7660 15224
rect 7700 15184 9964 15224
rect 10004 15184 10013 15224
rect 0 15164 80 15184
rect 6499 15140 6557 15141
rect 3679 15100 3688 15140
rect 3728 15100 3770 15140
rect 3810 15100 3852 15140
rect 3892 15100 3934 15140
rect 3974 15100 4016 15140
rect 4056 15100 4065 15140
rect 6499 15100 6508 15140
rect 6548 15100 7564 15140
rect 7604 15100 7613 15140
rect 18799 15100 18808 15140
rect 18848 15100 18890 15140
rect 18930 15100 18972 15140
rect 19012 15100 19054 15140
rect 19094 15100 19136 15140
rect 19176 15100 19185 15140
rect 6499 15099 6557 15100
rect 8035 15056 8093 15057
rect 7950 15016 8044 15056
rect 8084 15016 8093 15056
rect 8035 15015 8093 15016
rect 3235 14972 3293 14973
rect 3235 14932 3244 14972
rect 3284 14932 5164 14972
rect 5204 14932 10060 14972
rect 10100 14932 10444 14972
rect 10484 14932 10493 14972
rect 3235 14931 3293 14932
rect 0 14888 80 14908
rect 0 14848 7660 14888
rect 7700 14848 7709 14888
rect 8131 14848 8140 14888
rect 8180 14848 8428 14888
rect 8468 14848 8477 14888
rect 12835 14848 12844 14888
rect 12884 14848 13228 14888
rect 13268 14848 13277 14888
rect 13987 14848 13996 14888
rect 14036 14848 15436 14888
rect 15476 14848 16492 14888
rect 16532 14848 16541 14888
rect 0 14828 80 14848
rect 4675 14764 4684 14804
rect 4724 14764 6220 14804
rect 6260 14764 6269 14804
rect 7843 14764 7852 14804
rect 7892 14764 8716 14804
rect 8756 14764 8765 14804
rect 12163 14764 12172 14804
rect 12212 14764 17260 14804
rect 17300 14764 17548 14804
rect 17588 14764 17597 14804
rect 4195 14720 4253 14721
rect 21424 14720 21504 14740
rect 2500 14680 4204 14720
rect 4244 14680 4253 14720
rect 9283 14680 9292 14720
rect 9332 14680 11020 14720
rect 11060 14680 11069 14720
rect 12739 14680 12748 14720
rect 12788 14680 13036 14720
rect 13076 14680 15532 14720
rect 15572 14680 15581 14720
rect 16771 14680 16780 14720
rect 16820 14680 17164 14720
rect 17204 14680 17213 14720
rect 17635 14680 17644 14720
rect 17684 14680 18220 14720
rect 18260 14680 18269 14720
rect 2500 14636 2540 14680
rect 4195 14679 4253 14680
rect 21388 14660 21504 14720
rect 13027 14636 13085 14637
rect 21388 14636 21428 14660
rect 2083 14596 2092 14636
rect 2132 14596 2540 14636
rect 2947 14596 2956 14636
rect 2996 14596 5836 14636
rect 5876 14596 5885 14636
rect 13027 14596 13036 14636
rect 13076 14596 21428 14636
rect 13027 14595 13085 14596
rect 0 14552 80 14572
rect 3331 14552 3389 14553
rect 0 14512 2860 14552
rect 2900 14512 2909 14552
rect 3246 14512 3340 14552
rect 3380 14512 3389 14552
rect 3523 14512 3532 14552
rect 3572 14512 6700 14552
rect 6740 14512 7372 14552
rect 7412 14512 7421 14552
rect 11683 14512 11692 14552
rect 11732 14512 12940 14552
rect 12980 14512 12989 14552
rect 14563 14512 14572 14552
rect 14612 14512 14956 14552
rect 14996 14512 15005 14552
rect 16483 14512 16492 14552
rect 16532 14512 18796 14552
rect 18836 14512 18845 14552
rect 0 14492 80 14512
rect 3331 14511 3389 14512
rect 9475 14468 9533 14469
rect 1987 14428 1996 14468
rect 2036 14428 9484 14468
rect 9524 14428 9533 14468
rect 13315 14428 13324 14468
rect 13364 14428 13516 14468
rect 13556 14428 13565 14468
rect 9475 14427 9533 14428
rect 3811 14344 3820 14384
rect 3860 14344 4300 14384
rect 4340 14344 4349 14384
rect 4919 14344 4928 14384
rect 4968 14344 5010 14384
rect 5050 14344 5092 14384
rect 5132 14344 5174 14384
rect 5214 14344 5256 14384
rect 5296 14344 5305 14384
rect 20039 14344 20048 14384
rect 20088 14344 20130 14384
rect 20170 14344 20212 14384
rect 20252 14344 20294 14384
rect 20334 14344 20376 14384
rect 20416 14344 20425 14384
rect 1507 14260 1516 14300
rect 1556 14260 17356 14300
rect 17396 14260 17405 14300
rect 0 14216 80 14236
rect 16483 14216 16541 14217
rect 0 14176 1804 14216
rect 1844 14176 1853 14216
rect 5827 14176 5836 14216
rect 5876 14176 9292 14216
rect 9332 14176 9341 14216
rect 16483 14176 16492 14216
rect 16532 14176 16684 14216
rect 16724 14176 16733 14216
rect 18595 14176 18604 14216
rect 18644 14176 19180 14216
rect 19220 14176 19229 14216
rect 0 14156 80 14176
rect 16483 14175 16541 14176
rect 4195 14132 4253 14133
rect 8899 14132 8957 14133
rect 4195 14092 4204 14132
rect 4244 14092 4972 14132
rect 5012 14092 5021 14132
rect 8800 14092 8908 14132
rect 8948 14092 9484 14132
rect 9524 14092 9533 14132
rect 14179 14092 14188 14132
rect 14228 14092 16108 14132
rect 16148 14092 18700 14132
rect 18740 14092 19276 14132
rect 19316 14092 19325 14132
rect 4195 14091 4253 14092
rect 2275 14008 2284 14048
rect 2324 14008 2668 14048
rect 2708 14008 3244 14048
rect 3284 14008 3293 14048
rect 3427 14008 3436 14048
rect 3476 14008 3820 14048
rect 3860 14008 5452 14048
rect 5492 14008 5501 14048
rect 6499 14008 6508 14048
rect 6548 14008 8620 14048
rect 8660 14008 8669 14048
rect 8800 13964 8840 14092
rect 8899 14091 8957 14092
rect 9379 14048 9437 14049
rect 21424 14048 21504 14068
rect 9379 14008 9388 14048
rect 9428 14008 21504 14048
rect 9379 14007 9437 14008
rect 21424 13988 21504 14008
rect 8707 13924 8716 13964
rect 8756 13924 8840 13964
rect 11203 13964 11261 13965
rect 11203 13924 11212 13964
rect 11252 13924 17644 13964
rect 17684 13924 17693 13964
rect 11203 13923 11261 13924
rect 0 13880 80 13900
rect 7459 13880 7517 13881
rect 10339 13880 10397 13881
rect 13123 13880 13181 13881
rect 0 13840 2228 13880
rect 0 13820 80 13840
rect 2188 13712 2228 13840
rect 2380 13840 3724 13880
rect 3764 13840 3773 13880
rect 7075 13840 7084 13880
rect 7124 13840 7468 13880
rect 7508 13840 7517 13880
rect 9571 13840 9580 13880
rect 9620 13840 10348 13880
rect 10388 13840 10397 13880
rect 13038 13840 13132 13880
rect 13172 13840 13181 13880
rect 15331 13840 15340 13880
rect 15380 13840 16012 13880
rect 16052 13840 16061 13880
rect 17155 13840 17164 13880
rect 17204 13840 18988 13880
rect 19028 13840 19037 13880
rect 2380 13712 2420 13840
rect 7459 13839 7517 13840
rect 10339 13839 10397 13840
rect 13123 13839 13181 13840
rect 9379 13756 9388 13796
rect 9428 13756 10252 13796
rect 10292 13756 10301 13796
rect 14659 13756 14668 13796
rect 14708 13756 15436 13796
rect 15476 13756 15485 13796
rect 2188 13672 2420 13712
rect 13795 13672 13804 13712
rect 13844 13672 15916 13712
rect 15956 13672 16204 13712
rect 16244 13672 16253 13712
rect 3679 13588 3688 13628
rect 3728 13588 3770 13628
rect 3810 13588 3852 13628
rect 3892 13588 3934 13628
rect 3974 13588 4016 13628
rect 4056 13588 4065 13628
rect 18799 13588 18808 13628
rect 18848 13588 18890 13628
rect 18930 13588 18972 13628
rect 19012 13588 19054 13628
rect 19094 13588 19136 13628
rect 19176 13588 19185 13628
rect 0 13544 80 13564
rect 0 13504 1228 13544
rect 1268 13504 1277 13544
rect 2563 13504 2572 13544
rect 2612 13504 2860 13544
rect 2900 13504 2909 13544
rect 0 13484 80 13504
rect 4579 13420 4588 13460
rect 4628 13420 5068 13460
rect 5108 13420 5117 13460
rect 17059 13420 17068 13460
rect 17108 13420 17356 13460
rect 17396 13420 17405 13460
rect 6211 13376 6269 13377
rect 21424 13376 21504 13396
rect 4675 13336 4684 13376
rect 4724 13336 6220 13376
rect 6260 13336 8428 13376
rect 8468 13336 8477 13376
rect 12259 13336 12268 13376
rect 12308 13336 13420 13376
rect 13460 13336 14188 13376
rect 14228 13336 14380 13376
rect 14420 13336 14429 13376
rect 15139 13336 15148 13376
rect 15188 13336 15628 13376
rect 15668 13336 15677 13376
rect 18307 13336 18316 13376
rect 18356 13336 21504 13376
rect 6211 13335 6269 13336
rect 21424 13316 21504 13336
rect 5635 13292 5693 13293
rect 15811 13292 15869 13293
rect 1219 13252 1228 13292
rect 1268 13252 4492 13292
rect 4532 13252 4541 13292
rect 5550 13252 5644 13292
rect 5684 13252 5693 13292
rect 6211 13252 6220 13292
rect 6260 13252 6508 13292
rect 6548 13252 8044 13292
rect 8084 13252 8093 13292
rect 13603 13252 13612 13292
rect 13652 13252 13900 13292
rect 13940 13252 13949 13292
rect 15811 13252 15820 13292
rect 15860 13252 15916 13292
rect 15956 13252 15965 13292
rect 16387 13252 16396 13292
rect 16436 13252 17068 13292
rect 17108 13252 17117 13292
rect 5635 13251 5693 13252
rect 15811 13251 15869 13252
rect 0 13208 80 13228
rect 4099 13208 4157 13209
rect 0 13168 76 13208
rect 116 13168 125 13208
rect 2467 13168 2476 13208
rect 2516 13168 2764 13208
rect 2804 13168 2813 13208
rect 4014 13168 4108 13208
rect 4148 13168 5836 13208
rect 5876 13168 5885 13208
rect 7267 13168 7276 13208
rect 7316 13168 8524 13208
rect 8564 13168 8573 13208
rect 11011 13168 11020 13217
rect 11060 13177 11146 13217
rect 11060 13168 11069 13177
rect 13123 13168 13132 13208
rect 13172 13168 13420 13208
rect 13460 13168 15532 13208
rect 15572 13168 15724 13208
rect 15764 13168 15773 13208
rect 0 13148 80 13168
rect 4099 13167 4157 13168
rect 11011 13167 11069 13168
rect 6787 13124 6845 13125
rect 4291 13084 4300 13124
rect 4340 13084 4588 13124
rect 4628 13084 4637 13124
rect 6787 13084 6796 13124
rect 6836 13084 9772 13124
rect 9812 13084 9821 13124
rect 6787 13083 6845 13084
rect 1603 13000 1612 13040
rect 1652 13000 15052 13040
rect 15092 13000 15101 13040
rect 6307 12956 6365 12957
rect 6307 12916 6316 12956
rect 6356 12916 7852 12956
rect 7892 12916 7901 12956
rect 6307 12915 6365 12916
rect 0 12872 80 12892
rect 0 12832 1708 12872
rect 1748 12832 1757 12872
rect 4919 12832 4928 12872
rect 4968 12832 5010 12872
rect 5050 12832 5092 12872
rect 5132 12832 5174 12872
rect 5214 12832 5256 12872
rect 5296 12832 5305 12872
rect 6019 12832 6028 12872
rect 6068 12832 6220 12872
rect 6260 12832 6269 12872
rect 8323 12832 8332 12872
rect 8372 12832 13420 12872
rect 13460 12832 13708 12872
rect 13748 12832 13757 12872
rect 20039 12832 20048 12872
rect 20088 12832 20130 12872
rect 20170 12832 20212 12872
rect 20252 12832 20294 12872
rect 20334 12832 20376 12872
rect 20416 12832 20425 12872
rect 0 12812 80 12832
rect 2083 12748 2092 12788
rect 2132 12748 6316 12788
rect 6356 12748 6365 12788
rect 16195 12704 16253 12705
rect 21424 12704 21504 12724
rect 2371 12664 2380 12704
rect 2420 12664 2668 12704
rect 2708 12664 2956 12704
rect 2996 12664 3005 12704
rect 16195 12664 16204 12704
rect 16244 12664 21504 12704
rect 16195 12663 16253 12664
rect 21424 12644 21504 12664
rect 11011 12620 11069 12621
rect 13123 12620 13181 12621
rect 15235 12620 15293 12621
rect 2179 12580 2188 12620
rect 2228 12580 2764 12620
rect 2804 12580 2813 12620
rect 3043 12580 3052 12620
rect 3092 12580 3101 12620
rect 3235 12580 3244 12620
rect 3284 12580 3628 12620
rect 3668 12580 3677 12620
rect 6979 12580 6988 12620
rect 7028 12580 7660 12620
rect 7700 12580 7709 12620
rect 9091 12580 9100 12620
rect 9140 12580 9964 12620
rect 10004 12580 10732 12620
rect 10772 12580 11020 12620
rect 11060 12580 13132 12620
rect 13172 12580 13181 12620
rect 15150 12580 15244 12620
rect 15284 12580 15293 12620
rect 15619 12580 15628 12620
rect 15668 12580 17260 12620
rect 17300 12580 17309 12620
rect 0 12536 80 12556
rect 3052 12536 3092 12580
rect 11011 12579 11069 12580
rect 13123 12579 13181 12580
rect 15235 12579 15293 12580
rect 7171 12536 7229 12537
rect 7747 12536 7805 12537
rect 15916 12536 15956 12580
rect 0 12496 212 12536
rect 1315 12496 1324 12536
rect 1364 12496 3092 12536
rect 3139 12496 3148 12536
rect 3188 12496 3916 12536
rect 3956 12496 3965 12536
rect 7171 12496 7180 12536
rect 7220 12496 7756 12536
rect 7796 12496 7805 12536
rect 15907 12496 15916 12536
rect 15956 12496 15996 12536
rect 16291 12496 16300 12536
rect 16340 12496 19564 12536
rect 19604 12496 19613 12536
rect 0 12476 80 12496
rect 172 12368 212 12496
rect 7171 12495 7229 12496
rect 7747 12495 7805 12496
rect 3043 12412 3052 12452
rect 3092 12412 3724 12452
rect 3764 12412 7084 12452
rect 7124 12412 7133 12452
rect 7459 12412 7468 12452
rect 7508 12412 7948 12452
rect 7988 12412 7997 12452
rect 172 12328 17644 12368
rect 17684 12328 17693 12368
rect 11011 12284 11069 12285
rect 11203 12284 11261 12285
rect 4387 12244 4396 12284
rect 4436 12244 8044 12284
rect 8084 12244 8093 12284
rect 9475 12244 9484 12284
rect 9524 12244 11020 12284
rect 11060 12244 11212 12284
rect 11252 12244 11261 12284
rect 12643 12244 12652 12284
rect 12692 12244 13036 12284
rect 13076 12244 13085 12284
rect 13603 12244 13612 12284
rect 13652 12244 14092 12284
rect 14132 12244 14141 12284
rect 11011 12243 11069 12244
rect 11203 12243 11261 12244
rect 0 12200 80 12220
rect 0 12160 7468 12200
rect 7508 12160 7517 12200
rect 0 12140 80 12160
rect 3679 12076 3688 12116
rect 3728 12076 3770 12116
rect 3810 12076 3852 12116
rect 3892 12076 3934 12116
rect 3974 12076 4016 12116
rect 4056 12076 4065 12116
rect 10915 12076 10924 12116
rect 10964 12076 11212 12116
rect 11252 12076 11261 12116
rect 18799 12076 18808 12116
rect 18848 12076 18890 12116
rect 18930 12076 18972 12116
rect 19012 12076 19054 12116
rect 19094 12076 19136 12116
rect 19176 12076 19185 12116
rect 21424 12032 21504 12052
rect 4483 11992 4492 12032
rect 4532 11992 5356 12032
rect 5396 11992 6316 12032
rect 6356 11992 21504 12032
rect 21424 11972 21504 11992
rect 1987 11908 1996 11948
rect 2036 11908 2188 11948
rect 2228 11908 2237 11948
rect 7075 11908 7084 11948
rect 7124 11908 7948 11948
rect 7988 11908 8620 11948
rect 8660 11908 16108 11948
rect 16148 11908 16157 11948
rect 0 11864 80 11884
rect 15811 11864 15869 11865
rect 0 11824 1708 11864
rect 1748 11824 1757 11864
rect 4963 11824 4972 11864
rect 5012 11824 5644 11864
rect 5684 11824 5693 11864
rect 8803 11824 8812 11864
rect 8852 11824 9868 11864
rect 9908 11824 9917 11864
rect 11203 11824 11212 11864
rect 11252 11824 15820 11864
rect 15860 11824 15869 11864
rect 0 11804 80 11824
rect 15811 11823 15869 11824
rect 16387 11780 16445 11781
rect 1987 11740 1996 11780
rect 2036 11740 12940 11780
rect 12980 11740 12989 11780
rect 16302 11740 16396 11780
rect 16436 11740 16445 11780
rect 16387 11739 16445 11740
rect 13123 11696 13181 11697
rect 7267 11656 7276 11696
rect 7316 11656 7852 11696
rect 7892 11656 7901 11696
rect 10531 11656 10540 11696
rect 10580 11656 10868 11696
rect 12451 11656 12460 11696
rect 12500 11656 13132 11696
rect 13172 11656 14956 11696
rect 14996 11656 15005 11696
rect 2500 11572 5644 11612
rect 5684 11572 5693 11612
rect 6979 11572 6988 11612
rect 7028 11572 9388 11612
rect 9428 11572 9437 11612
rect 0 11528 80 11548
rect 2500 11528 2540 11572
rect 4291 11528 4349 11529
rect 0 11488 1268 11528
rect 1891 11488 1900 11528
rect 1940 11488 2540 11528
rect 4099 11488 4108 11528
rect 4148 11488 4300 11528
rect 4340 11488 4349 11528
rect 5923 11488 5932 11528
rect 5972 11488 6220 11528
rect 6260 11488 6269 11528
rect 8131 11488 8140 11528
rect 8180 11488 8716 11528
rect 8756 11488 8765 11528
rect 10435 11488 10444 11528
rect 10484 11488 10493 11528
rect 0 11468 80 11488
rect 1228 11444 1268 11488
rect 4291 11487 4349 11488
rect 10444 11444 10484 11488
rect 10828 11444 10868 11656
rect 13123 11655 13181 11656
rect 13315 11572 13324 11612
rect 13364 11572 13804 11612
rect 13844 11572 13853 11612
rect 17443 11572 17452 11612
rect 17492 11572 17836 11612
rect 17876 11572 17885 11612
rect 14083 11488 14092 11528
rect 14132 11488 14860 11528
rect 14900 11488 14909 11528
rect 16963 11488 16972 11528
rect 17012 11488 17548 11528
rect 17588 11488 18412 11528
rect 18452 11488 18461 11528
rect 1228 11404 2380 11444
rect 2420 11404 2429 11444
rect 4684 11404 6028 11444
rect 6068 11404 10484 11444
rect 10819 11404 10828 11444
rect 10868 11404 10877 11444
rect 11299 11404 11308 11444
rect 11348 11404 20564 11444
rect 4684 11360 4724 11404
rect 20524 11360 20564 11404
rect 21424 11360 21504 11380
rect 4644 11320 4684 11360
rect 4724 11320 4733 11360
rect 4919 11320 4928 11360
rect 4968 11320 5010 11360
rect 5050 11320 5092 11360
rect 5132 11320 5174 11360
rect 5214 11320 5256 11360
rect 5296 11320 5305 11360
rect 9667 11320 9676 11360
rect 9716 11320 11212 11360
rect 11252 11320 11261 11360
rect 11683 11320 11692 11360
rect 11732 11320 11828 11360
rect 20039 11320 20048 11360
rect 20088 11320 20130 11360
rect 20170 11320 20212 11360
rect 20252 11320 20294 11360
rect 20334 11320 20376 11360
rect 20416 11320 20425 11360
rect 20524 11320 21504 11360
rect 4099 11276 4157 11277
rect 6211 11276 6269 11277
rect 3340 11236 4108 11276
rect 4148 11236 5356 11276
rect 5396 11236 5405 11276
rect 6115 11236 6124 11276
rect 6164 11236 6220 11276
rect 6260 11236 6269 11276
rect 6403 11236 6412 11276
rect 6452 11236 6700 11276
rect 6740 11236 7084 11276
rect 7124 11236 7133 11276
rect 11491 11236 11500 11276
rect 11540 11236 11732 11276
rect 0 11192 80 11212
rect 3340 11192 3380 11236
rect 4099 11235 4157 11236
rect 6124 11192 6164 11236
rect 6211 11235 6269 11236
rect 11692 11192 11732 11236
rect 0 11152 1420 11192
rect 1460 11152 1469 11192
rect 3043 11152 3052 11192
rect 3092 11152 3340 11192
rect 3380 11152 3389 11192
rect 4003 11152 4012 11192
rect 4052 11152 4780 11192
rect 4820 11152 6164 11192
rect 9859 11152 9868 11192
rect 9908 11152 10156 11192
rect 10196 11152 10205 11192
rect 11683 11152 11692 11192
rect 11732 11152 11741 11192
rect 0 11132 80 11152
rect 4579 11108 4637 11109
rect 11788 11108 11828 11320
rect 21424 11300 21504 11320
rect 14371 11192 14429 11193
rect 14286 11152 14380 11192
rect 14420 11152 14429 11192
rect 15907 11152 15916 11192
rect 15956 11152 16492 11192
rect 16532 11152 16541 11192
rect 14371 11151 14429 11152
rect 2179 11068 2188 11108
rect 2228 11068 4588 11108
rect 4628 11068 4637 11108
rect 10243 11068 10252 11108
rect 10292 11068 10636 11108
rect 10676 11068 10685 11108
rect 11491 11068 11500 11108
rect 11540 11068 11828 11108
rect 4579 11067 4637 11068
rect 10147 11024 10205 11025
rect 3427 10984 3436 11024
rect 3476 10984 5548 11024
rect 5588 10984 5597 11024
rect 10062 10984 10156 11024
rect 10196 10984 10205 11024
rect 10435 10984 10444 11024
rect 10484 10984 11404 11024
rect 11444 10984 11453 11024
rect 13027 10984 13036 11024
rect 13076 10984 13420 11024
rect 13460 10984 13469 11024
rect 14371 10984 14380 11024
rect 14420 10984 14956 11024
rect 14996 10984 16300 11024
rect 16340 10984 18028 11024
rect 18068 10984 18316 11024
rect 18356 10984 18508 11024
rect 18548 10984 18557 11024
rect 10147 10983 10205 10984
rect 1603 10900 1612 10940
rect 1652 10900 10060 10940
rect 10100 10900 10109 10940
rect 14179 10900 14188 10940
rect 14228 10900 15052 10940
rect 15092 10900 15101 10940
rect 0 10856 80 10876
rect 0 10816 10732 10856
rect 10772 10816 10781 10856
rect 12931 10816 12940 10856
rect 12980 10816 14668 10856
rect 14708 10816 14717 10856
rect 0 10796 80 10816
rect 6307 10732 6316 10772
rect 6356 10732 6604 10772
rect 6644 10732 6653 10772
rect 12067 10732 12076 10772
rect 12116 10732 12556 10772
rect 12596 10732 12605 10772
rect 21424 10688 21504 10708
rect 6115 10648 6124 10688
rect 6164 10648 7468 10688
rect 7508 10648 7517 10688
rect 11320 10648 11980 10688
rect 12020 10648 12029 10688
rect 18700 10648 21504 10688
rect 2563 10604 2621 10605
rect 11320 10604 11360 10648
rect 18700 10604 18740 10648
rect 21424 10628 21504 10648
rect 2467 10564 2476 10604
rect 2516 10564 2572 10604
rect 2612 10564 2621 10604
rect 3679 10564 3688 10604
rect 3728 10564 3770 10604
rect 3810 10564 3852 10604
rect 3892 10564 3934 10604
rect 3974 10564 4016 10604
rect 4056 10564 4065 10604
rect 6499 10564 6508 10604
rect 6548 10564 11360 10604
rect 11875 10564 11884 10604
rect 11924 10564 12076 10604
rect 12116 10564 12125 10604
rect 12739 10564 12748 10604
rect 12788 10564 13708 10604
rect 13748 10564 18028 10604
rect 18068 10564 18700 10604
rect 18740 10564 18749 10604
rect 18799 10564 18808 10604
rect 18848 10564 18890 10604
rect 18930 10564 18972 10604
rect 19012 10564 19054 10604
rect 19094 10564 19136 10604
rect 19176 10564 19185 10604
rect 2563 10563 2621 10564
rect 0 10520 80 10540
rect 0 10480 7948 10520
rect 7988 10480 7997 10520
rect 11971 10480 11980 10520
rect 12020 10480 14284 10520
rect 14324 10480 14333 10520
rect 0 10460 80 10480
rect 2467 10396 2476 10436
rect 2516 10396 10732 10436
rect 10772 10396 10781 10436
rect 11875 10396 11884 10436
rect 11924 10396 13748 10436
rect 15715 10396 15724 10436
rect 15764 10396 16012 10436
rect 16052 10396 16061 10436
rect 18691 10396 18700 10436
rect 18740 10396 19468 10436
rect 19508 10396 19517 10436
rect 13708 10352 13748 10396
rect 4387 10312 4396 10352
rect 4436 10312 5452 10352
rect 5492 10312 6412 10352
rect 6452 10312 6461 10352
rect 10531 10312 10540 10352
rect 10580 10312 12460 10352
rect 12500 10312 12509 10352
rect 13699 10312 13708 10352
rect 13748 10312 17068 10352
rect 17108 10312 17117 10352
rect 1603 10228 1612 10268
rect 1652 10228 14668 10268
rect 14708 10228 14717 10268
rect 0 10184 80 10204
rect 0 10144 2284 10184
rect 2324 10144 2333 10184
rect 3811 10144 3820 10184
rect 3860 10144 4204 10184
rect 4244 10144 4253 10184
rect 5539 10144 5548 10184
rect 5588 10144 5932 10184
rect 5972 10144 7660 10184
rect 7700 10144 8332 10184
rect 8372 10144 9964 10184
rect 10004 10144 10348 10184
rect 10388 10144 10540 10184
rect 10580 10144 10589 10184
rect 11107 10144 11116 10184
rect 11156 10144 11404 10184
rect 11444 10144 11453 10184
rect 11971 10144 11980 10184
rect 12020 10144 12029 10184
rect 12355 10144 12364 10184
rect 12404 10144 12652 10184
rect 12692 10144 13324 10184
rect 13364 10144 13373 10184
rect 14275 10144 14284 10184
rect 14324 10144 18412 10184
rect 18452 10144 18461 10184
rect 0 10124 80 10144
rect 11980 10100 12020 10144
rect 1891 10060 1900 10100
rect 1940 10060 4684 10100
rect 4724 10060 4733 10100
rect 7075 10060 7084 10100
rect 7124 10060 7372 10100
rect 7412 10060 7421 10100
rect 11299 10060 11308 10100
rect 11348 10060 12020 10100
rect 13987 10060 13996 10100
rect 14036 10060 17260 10100
rect 17300 10060 17309 10100
rect 2851 10016 2909 10017
rect 21424 10016 21504 10036
rect 2766 9976 2860 10016
rect 2900 9976 2909 10016
rect 3715 9976 3724 10016
rect 3764 9976 4492 10016
rect 4532 9976 4541 10016
rect 11320 9976 21504 10016
rect 2851 9975 2909 9976
rect 11320 9932 11360 9976
rect 21424 9956 21504 9976
rect 2083 9892 2092 9932
rect 2132 9892 6028 9932
rect 6068 9892 6316 9932
rect 6356 9892 6365 9932
rect 8803 9892 8812 9932
rect 8852 9892 11360 9932
rect 14371 9932 14429 9933
rect 14371 9892 14380 9932
rect 14420 9892 14668 9932
rect 14708 9892 14717 9932
rect 0 9848 80 9868
rect 2947 9848 3005 9849
rect 4675 9848 4733 9849
rect 0 9808 1900 9848
rect 1940 9808 1949 9848
rect 2862 9808 2956 9848
rect 2996 9808 3005 9848
rect 4579 9808 4588 9848
rect 4628 9808 4684 9848
rect 4724 9808 4733 9848
rect 4919 9808 4928 9848
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 5296 9808 5305 9848
rect 0 9788 80 9808
rect 2947 9807 3005 9808
rect 4675 9807 4733 9808
rect 7651 9764 7709 9765
rect 8812 9764 8852 9892
rect 14371 9891 14429 9892
rect 20039 9808 20048 9848
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20416 9808 20425 9848
rect 4099 9724 4108 9764
rect 4148 9724 7660 9764
rect 7700 9724 8852 9764
rect 16963 9724 16972 9764
rect 17012 9724 17260 9764
rect 17300 9724 17309 9764
rect 7651 9723 7709 9724
rect 6787 9680 6845 9681
rect 8611 9680 8669 9681
rect 3235 9640 3244 9680
rect 3284 9640 4780 9680
rect 4820 9640 4829 9680
rect 5827 9640 5836 9680
rect 5876 9640 6796 9680
rect 6836 9640 6845 9680
rect 8526 9640 8620 9680
rect 8660 9640 8669 9680
rect 10339 9640 10348 9680
rect 10388 9640 10828 9680
rect 10868 9640 10877 9680
rect 14179 9640 14188 9680
rect 14228 9640 17740 9680
rect 17780 9640 17789 9680
rect 6787 9639 6845 9640
rect 8611 9639 8669 9640
rect 15715 9596 15773 9597
rect 4003 9556 4012 9596
rect 4052 9556 5073 9596
rect 5113 9556 5122 9596
rect 9763 9556 9772 9596
rect 9812 9556 11788 9596
rect 11828 9556 15724 9596
rect 15764 9556 15773 9596
rect 15715 9555 15773 9556
rect 0 9512 80 9532
rect 0 9472 1324 9512
rect 1364 9472 1373 9512
rect 3043 9472 3052 9512
rect 3092 9472 3244 9512
rect 3284 9472 3293 9512
rect 3427 9472 3436 9512
rect 3476 9472 3820 9512
rect 3860 9472 3869 9512
rect 4291 9472 4300 9512
rect 4340 9472 4972 9512
rect 5012 9472 5260 9512
rect 5300 9472 5309 9512
rect 9091 9472 9100 9512
rect 9140 9472 9868 9512
rect 9908 9472 13612 9512
rect 13652 9472 14572 9512
rect 14612 9472 14621 9512
rect 14851 9472 14860 9512
rect 14900 9472 16012 9512
rect 16052 9472 16061 9512
rect 18307 9472 18316 9512
rect 18356 9472 19276 9512
rect 19316 9472 19325 9512
rect 0 9452 80 9472
rect 2083 9388 2092 9428
rect 2132 9388 17644 9428
rect 17684 9388 17693 9428
rect 21424 9344 21504 9364
rect 1315 9304 1324 9344
rect 1364 9304 2540 9344
rect 7363 9304 7372 9344
rect 7412 9304 13172 9344
rect 13219 9304 13228 9344
rect 13268 9304 14860 9344
rect 14900 9304 14909 9344
rect 20140 9304 21504 9344
rect 2500 9260 2540 9304
rect 7651 9260 7709 9261
rect 8611 9260 8669 9261
rect 1507 9220 1516 9260
rect 1556 9220 1565 9260
rect 2500 9220 7084 9260
rect 7124 9220 7133 9260
rect 7566 9220 7660 9260
rect 7700 9220 7709 9260
rect 8526 9220 8620 9260
rect 8660 9220 8669 9260
rect 13132 9260 13172 9304
rect 20140 9260 20180 9304
rect 21424 9284 21504 9304
rect 13132 9220 13708 9260
rect 13748 9220 20180 9260
rect 0 9176 80 9196
rect 1516 9176 1556 9220
rect 7651 9219 7709 9220
rect 8611 9219 8669 9220
rect 0 9136 1556 9176
rect 2659 9136 2668 9176
rect 2708 9136 4204 9176
rect 4244 9136 4253 9176
rect 8131 9136 8140 9176
rect 8180 9136 8428 9176
rect 8468 9136 10348 9176
rect 10388 9136 10397 9176
rect 0 9116 80 9136
rect 8899 9092 8957 9093
rect 2755 9052 2764 9092
rect 2804 9052 3052 9092
rect 3092 9052 3101 9092
rect 3679 9052 3688 9092
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 4056 9052 4065 9092
rect 8899 9052 8908 9092
rect 8948 9052 15820 9092
rect 15860 9052 18316 9092
rect 18356 9052 18365 9092
rect 18799 9052 18808 9092
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 19176 9052 19185 9092
rect 8899 9051 8957 9052
rect 2500 8968 12556 9008
rect 12596 8968 12605 9008
rect 2500 8924 2540 8968
rect 1411 8884 1420 8924
rect 1460 8884 2540 8924
rect 15331 8884 15340 8924
rect 15380 8884 15628 8924
rect 15668 8884 15677 8924
rect 17731 8884 17740 8924
rect 17780 8884 18124 8924
rect 18164 8884 18173 8924
rect 0 8840 80 8860
rect 0 8800 1228 8840
rect 1268 8800 1277 8840
rect 2371 8800 2380 8840
rect 2420 8800 3724 8840
rect 3764 8800 3773 8840
rect 4012 8800 7988 8840
rect 8323 8800 8332 8840
rect 8372 8800 10060 8840
rect 10100 8800 10109 8840
rect 11779 8800 11788 8840
rect 11828 8800 12460 8840
rect 12500 8800 14188 8840
rect 14228 8800 14237 8840
rect 17155 8800 17164 8840
rect 17204 8800 18700 8840
rect 18740 8800 18749 8840
rect 0 8780 80 8800
rect 4012 8756 4052 8800
rect 7843 8756 7901 8757
rect 1699 8716 1708 8756
rect 1748 8716 4052 8756
rect 4099 8716 4108 8756
rect 4148 8716 7852 8756
rect 7892 8716 7901 8756
rect 7948 8756 7988 8800
rect 7948 8716 10156 8756
rect 10196 8716 10205 8756
rect 10494 8716 10503 8756
rect 10543 8716 11212 8756
rect 11252 8716 12844 8756
rect 12884 8716 12893 8756
rect 15427 8716 15436 8756
rect 15476 8716 17068 8756
rect 17108 8716 17117 8756
rect 7843 8715 7901 8716
rect 13027 8672 13085 8673
rect 21424 8672 21504 8692
rect 2851 8632 2860 8672
rect 2900 8632 3340 8672
rect 3380 8632 3389 8672
rect 3459 8632 3468 8672
rect 3508 8632 4012 8672
rect 4052 8632 4061 8672
rect 5347 8632 5356 8672
rect 5396 8632 5492 8672
rect 6595 8632 6604 8672
rect 6644 8632 6892 8672
rect 6932 8632 6941 8672
rect 8227 8632 8236 8672
rect 8276 8632 9964 8672
rect 10004 8632 10013 8672
rect 12739 8632 12748 8672
rect 12788 8632 13036 8672
rect 13076 8632 13085 8672
rect 15523 8632 15532 8672
rect 15572 8632 16300 8672
rect 16340 8632 17548 8672
rect 17588 8632 17597 8672
rect 21379 8632 21388 8672
rect 21428 8632 21504 8672
rect 0 8504 80 8524
rect 5347 8504 5405 8505
rect 5452 8504 5492 8632
rect 13027 8631 13085 8632
rect 21424 8612 21504 8632
rect 5539 8548 5548 8588
rect 5588 8548 7468 8588
rect 7508 8548 7517 8588
rect 9571 8548 9580 8588
rect 9620 8548 10924 8588
rect 10964 8548 10973 8588
rect 0 8464 1900 8504
rect 1940 8464 1949 8504
rect 2467 8464 2476 8504
rect 2516 8464 3244 8504
rect 3284 8464 3293 8504
rect 5328 8464 5356 8504
rect 5396 8464 7180 8504
rect 7220 8464 8524 8504
rect 8564 8464 10060 8504
rect 10100 8464 10109 8504
rect 10339 8464 10348 8504
rect 10388 8464 11884 8504
rect 11924 8464 11933 8504
rect 0 8444 80 8464
rect 5347 8463 5405 8464
rect 2563 8420 2621 8421
rect 2563 8380 2572 8420
rect 2612 8380 2668 8420
rect 2708 8380 2717 8420
rect 3907 8380 3916 8420
rect 3956 8380 14572 8420
rect 14612 8380 14621 8420
rect 2563 8379 2621 8380
rect 11011 8336 11069 8337
rect 1795 8296 1804 8336
rect 1844 8296 2540 8336
rect 4919 8296 4928 8336
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 5296 8296 5305 8336
rect 6691 8296 6700 8336
rect 6740 8296 7084 8336
rect 7124 8296 7133 8336
rect 10915 8296 10924 8336
rect 10964 8296 11020 8336
rect 11060 8296 11069 8336
rect 20039 8296 20048 8336
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20416 8296 20425 8336
rect 2500 8252 2540 8296
rect 11011 8295 11069 8296
rect 2500 8212 8716 8252
rect 8756 8212 8765 8252
rect 10051 8212 10060 8252
rect 10100 8212 10444 8252
rect 10484 8212 12556 8252
rect 12596 8212 12940 8252
rect 12980 8212 12989 8252
rect 13603 8212 13612 8252
rect 13652 8212 15148 8252
rect 15188 8212 15197 8252
rect 16675 8212 16684 8252
rect 16724 8212 17260 8252
rect 17300 8212 17309 8252
rect 0 8168 80 8188
rect 7075 8168 7133 8169
rect 11011 8168 11069 8169
rect 0 8128 1516 8168
rect 1556 8128 1565 8168
rect 2851 8128 2860 8168
rect 2900 8128 3052 8168
rect 3092 8128 3101 8168
rect 5923 8128 5932 8168
rect 5972 8128 6700 8168
rect 6740 8128 6749 8168
rect 7075 8128 7084 8168
rect 7124 8128 8044 8168
rect 8084 8128 8093 8168
rect 11011 8128 11020 8168
rect 11060 8128 11154 8168
rect 11395 8128 11404 8168
rect 11444 8128 16780 8168
rect 16820 8128 16829 8168
rect 16963 8128 16972 8168
rect 17012 8128 17452 8168
rect 17492 8128 17501 8168
rect 21292 8128 21388 8168
rect 21428 8128 21437 8168
rect 0 8108 80 8128
rect 7075 8127 7133 8128
rect 11011 8127 11069 8128
rect 5347 8084 5405 8085
rect 21292 8084 21332 8128
rect 1516 8044 4108 8084
rect 4148 8044 4157 8084
rect 4867 8044 4876 8084
rect 4916 8044 5356 8084
rect 5396 8044 5405 8084
rect 11875 8044 11884 8084
rect 11924 8044 13900 8084
rect 13940 8044 14476 8084
rect 14516 8044 14525 8084
rect 14572 8044 21332 8084
rect 1516 8000 1556 8044
rect 5347 8043 5405 8044
rect 14572 8000 14612 8044
rect 16099 8000 16157 8001
rect 21424 8000 21504 8020
rect 1507 7960 1516 8000
rect 1556 7960 1565 8000
rect 3619 7960 3628 8000
rect 3668 7960 7276 8000
rect 7316 7960 7325 8000
rect 7459 7960 7468 8000
rect 7508 7960 7852 8000
rect 7892 7960 9580 8000
rect 9620 7960 12652 8000
rect 12692 7960 12940 8000
rect 12980 7960 14612 8000
rect 16014 7960 16108 8000
rect 16148 7960 16396 8000
rect 16436 7960 16445 8000
rect 17539 7960 17548 8000
rect 17588 7960 19372 8000
rect 19412 7960 21504 8000
rect 16099 7959 16157 7960
rect 21424 7940 21504 7960
rect 10819 7916 10877 7917
rect 1603 7876 1612 7916
rect 1652 7876 3380 7916
rect 3427 7876 3436 7916
rect 3476 7876 5740 7916
rect 5780 7876 5789 7916
rect 6595 7876 6604 7916
rect 6644 7876 8044 7916
rect 8084 7876 8093 7916
rect 8899 7876 8908 7916
rect 8948 7876 9196 7916
rect 9236 7876 9676 7916
rect 9716 7876 9725 7916
rect 10819 7876 10828 7916
rect 10868 7876 10924 7916
rect 10964 7876 10973 7916
rect 12259 7876 12268 7916
rect 12308 7876 12556 7916
rect 12596 7876 17164 7916
rect 17204 7876 17213 7916
rect 18787 7876 18796 7916
rect 18836 7876 19180 7916
rect 19220 7876 19229 7916
rect 0 7832 80 7852
rect 3340 7832 3380 7876
rect 10819 7875 10877 7876
rect 5539 7832 5597 7833
rect 0 7792 3244 7832
rect 3284 7792 3293 7832
rect 3340 7792 5260 7832
rect 5300 7792 5548 7832
rect 5588 7792 5597 7832
rect 6019 7792 6028 7832
rect 6068 7792 6508 7832
rect 6548 7792 7180 7832
rect 7220 7792 7229 7832
rect 13411 7792 13420 7832
rect 13460 7792 13804 7832
rect 13844 7792 16396 7832
rect 16436 7792 16445 7832
rect 0 7772 80 7792
rect 5539 7791 5597 7792
rect 2083 7708 2092 7748
rect 2132 7708 14092 7748
rect 14132 7708 14141 7748
rect 6211 7664 6269 7665
rect 1987 7624 1996 7664
rect 2036 7624 4588 7664
rect 4628 7624 4637 7664
rect 6211 7624 6220 7664
rect 6260 7624 7084 7664
rect 7124 7624 7133 7664
rect 6211 7623 6269 7624
rect 13027 7580 13085 7581
rect 3679 7540 3688 7580
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 4056 7540 4065 7580
rect 4771 7540 4780 7580
rect 4820 7540 5452 7580
rect 5492 7540 5501 7580
rect 8515 7540 8524 7580
rect 8564 7540 9004 7580
rect 9044 7540 9053 7580
rect 11107 7540 11116 7580
rect 11156 7540 13036 7580
rect 13076 7540 13085 7580
rect 18799 7540 18808 7580
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 19176 7540 19185 7580
rect 13027 7539 13085 7540
rect 0 7496 80 7516
rect 11395 7496 11453 7497
rect 0 7456 1324 7496
rect 1364 7456 1373 7496
rect 1699 7456 1708 7496
rect 1748 7456 2860 7496
rect 2900 7456 2909 7496
rect 10243 7456 10252 7496
rect 10292 7456 11020 7496
rect 11060 7456 11069 7496
rect 11280 7456 11297 7496
rect 11337 7456 11404 7496
rect 11444 7456 11453 7496
rect 12739 7456 12748 7496
rect 12788 7456 14380 7496
rect 14420 7456 14429 7496
rect 0 7436 80 7456
rect 11395 7455 11453 7456
rect 1603 7372 1612 7412
rect 1652 7372 14284 7412
rect 14324 7372 14333 7412
rect 14755 7328 14813 7329
rect 21424 7328 21504 7348
rect 3715 7288 3724 7328
rect 3764 7288 6604 7328
rect 6644 7288 6653 7328
rect 11203 7288 11212 7328
rect 11252 7288 11404 7328
rect 11444 7288 11453 7328
rect 11500 7288 14764 7328
rect 14804 7288 17164 7328
rect 17204 7288 17213 7328
rect 17635 7288 17644 7328
rect 17684 7288 21504 7328
rect 4771 7244 4829 7245
rect 11500 7244 11540 7288
rect 14755 7287 14813 7288
rect 21424 7268 21504 7288
rect 3331 7204 3340 7244
rect 3380 7204 4300 7244
rect 4340 7204 4349 7244
rect 4771 7204 4780 7244
rect 4820 7204 11500 7244
rect 11540 7204 11549 7244
rect 4771 7203 4829 7204
rect 0 7160 80 7180
rect 2371 7160 2429 7161
rect 0 7120 2380 7160
rect 2420 7120 2429 7160
rect 3523 7120 3532 7160
rect 3572 7120 5740 7160
rect 5780 7120 5789 7160
rect 9187 7120 9196 7160
rect 9236 7120 11360 7160
rect 13123 7120 13132 7160
rect 13172 7120 13612 7160
rect 13652 7120 13804 7160
rect 13844 7120 13853 7160
rect 14947 7120 14956 7160
rect 14996 7120 15436 7160
rect 15476 7120 16684 7160
rect 16724 7120 16733 7160
rect 0 7100 80 7120
rect 2371 7119 2429 7120
rect 11320 7076 11360 7120
rect 2755 7036 2764 7076
rect 2804 7036 5548 7076
rect 5588 7036 6124 7076
rect 6164 7036 6988 7076
rect 7028 7036 8236 7076
rect 8276 7036 8620 7076
rect 8660 7036 9388 7076
rect 9428 7036 9772 7076
rect 9812 7036 10444 7076
rect 10484 7036 10493 7076
rect 10915 7036 10924 7076
rect 10964 7036 11212 7076
rect 11252 7036 11261 7076
rect 11320 7036 11692 7076
rect 11732 7036 15476 7076
rect 11395 6992 11453 6993
rect 15436 6992 15476 7036
rect 2659 6952 2668 6992
rect 2708 6952 7412 6992
rect 7459 6952 7468 6992
rect 7508 6952 11404 6992
rect 11444 6952 13324 6992
rect 13364 6952 13373 6992
rect 15427 6952 15436 6992
rect 15476 6952 15485 6992
rect 0 6824 80 6844
rect 7372 6824 7412 6952
rect 11395 6951 11453 6952
rect 11203 6908 11261 6909
rect 8899 6868 8908 6908
rect 8948 6868 10252 6908
rect 10292 6868 11212 6908
rect 11252 6868 13612 6908
rect 13652 6868 13661 6908
rect 14371 6868 14380 6908
rect 14420 6868 16588 6908
rect 16628 6868 16637 6908
rect 11203 6867 11261 6868
rect 0 6784 1708 6824
rect 1748 6784 1757 6824
rect 2083 6784 2092 6824
rect 2132 6784 2668 6824
rect 2708 6784 2717 6824
rect 2851 6784 2860 6824
rect 2900 6784 3340 6824
rect 3380 6784 3389 6824
rect 4919 6784 4928 6824
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 5296 6784 5305 6824
rect 7372 6784 8332 6824
rect 8372 6784 17644 6824
rect 17684 6784 17693 6824
rect 20039 6784 20048 6824
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20416 6784 20425 6824
rect 0 6764 80 6784
rect 2275 6700 2284 6740
rect 2324 6700 2956 6740
rect 2996 6700 3005 6740
rect 3048 6700 3057 6740
rect 3097 6700 4593 6740
rect 4633 6700 4642 6740
rect 10627 6700 10636 6740
rect 10676 6700 13036 6740
rect 13076 6700 16204 6740
rect 16244 6700 16253 6740
rect 11587 6656 11645 6657
rect 1612 6616 3148 6656
rect 3188 6616 3197 6656
rect 8707 6616 8716 6656
rect 8756 6616 11116 6656
rect 11156 6616 11165 6656
rect 11587 6616 11596 6656
rect 11636 6616 11788 6656
rect 11828 6616 11837 6656
rect 12259 6616 12268 6656
rect 12308 6616 12556 6656
rect 12596 6616 12605 6656
rect 0 6488 80 6508
rect 1612 6488 1652 6616
rect 11587 6615 11645 6616
rect 2179 6532 2188 6572
rect 2228 6532 2540 6572
rect 3331 6532 3340 6572
rect 3380 6532 4876 6572
rect 4916 6532 4925 6572
rect 8995 6532 9004 6572
rect 9044 6532 9196 6572
rect 9236 6532 11212 6572
rect 11252 6532 11261 6572
rect 0 6448 1652 6488
rect 2500 6488 2540 6532
rect 4675 6488 4733 6489
rect 2500 6448 2572 6488
rect 2612 6448 2621 6488
rect 3235 6448 3244 6488
rect 3284 6448 3532 6488
rect 3572 6448 3581 6488
rect 3811 6448 3820 6488
rect 3860 6448 4492 6488
rect 4532 6448 4541 6488
rect 4675 6448 4684 6488
rect 4724 6448 6988 6488
rect 7028 6448 7037 6488
rect 10723 6448 10732 6488
rect 10772 6448 10924 6488
rect 10964 6448 10973 6488
rect 12163 6448 12172 6488
rect 12212 6448 12844 6488
rect 12884 6448 12893 6488
rect 13123 6448 13132 6488
rect 13172 6448 13516 6488
rect 13556 6448 16876 6488
rect 16916 6448 16925 6488
rect 0 6428 80 6448
rect 4675 6447 4733 6448
rect 2371 6364 2380 6404
rect 2420 6364 2668 6404
rect 2708 6364 2717 6404
rect 10732 6364 11356 6404
rect 11396 6364 11630 6404
rect 11670 6364 11679 6404
rect 13027 6364 13036 6404
rect 13076 6364 13324 6404
rect 13364 6364 13900 6404
rect 13940 6364 13949 6404
rect 10732 6320 10772 6364
rect 11011 6320 11069 6321
rect 11203 6320 11261 6321
rect 10723 6280 10732 6320
rect 10772 6280 10781 6320
rect 10926 6280 11020 6320
rect 11060 6280 11069 6320
rect 11118 6280 11212 6320
rect 11252 6280 11261 6320
rect 11011 6279 11069 6280
rect 11203 6279 11261 6280
rect 11320 6280 18508 6320
rect 18548 6280 18557 6320
rect 8035 6196 8044 6236
rect 8084 6196 8428 6236
rect 8468 6196 8477 6236
rect 0 6152 80 6172
rect 2371 6152 2429 6153
rect 11320 6152 11360 6280
rect 12163 6236 12221 6237
rect 11683 6196 11692 6236
rect 11732 6196 12172 6236
rect 12212 6196 12221 6236
rect 12163 6195 12221 6196
rect 11587 6152 11645 6153
rect 0 6112 1324 6152
rect 1364 6112 1373 6152
rect 2371 6112 2380 6152
rect 2420 6112 11360 6152
rect 11502 6112 11596 6152
rect 11636 6112 11645 6152
rect 0 6092 80 6112
rect 2371 6111 2429 6112
rect 11587 6111 11645 6112
rect 3679 6028 3688 6068
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 4056 6028 4065 6068
rect 4387 6028 4396 6068
rect 4436 6028 5356 6068
rect 5396 6028 5405 6068
rect 18799 6028 18808 6068
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 19176 6028 19185 6068
rect 8515 5944 8524 5984
rect 8564 5944 10540 5984
rect 10580 5944 11308 5984
rect 11348 5944 11357 5984
rect 2179 5860 2188 5900
rect 2228 5860 10156 5900
rect 10196 5860 10205 5900
rect 11320 5860 16300 5900
rect 16340 5860 16349 5900
rect 0 5816 80 5836
rect 11320 5816 11360 5860
rect 0 5776 2284 5816
rect 2324 5776 2333 5816
rect 6979 5776 6988 5816
rect 7028 5776 11360 5816
rect 0 5756 80 5776
rect 9091 5732 9149 5733
rect 4387 5692 4396 5732
rect 4436 5692 4588 5732
rect 4628 5692 6028 5732
rect 6068 5692 6077 5732
rect 6307 5692 6316 5732
rect 6356 5692 6508 5732
rect 6548 5692 6557 5732
rect 7075 5692 7084 5732
rect 7124 5692 9100 5732
rect 9140 5692 9149 5732
rect 9091 5691 9149 5692
rect 2851 5648 2909 5649
rect 4771 5648 4829 5649
rect 8323 5648 8381 5649
rect 2851 5608 2860 5648
rect 2900 5608 2956 5648
rect 2996 5608 3005 5648
rect 4686 5608 4780 5648
rect 4820 5608 4829 5648
rect 6595 5608 6604 5648
rect 6644 5608 8332 5648
rect 8372 5608 8381 5648
rect 9859 5608 9868 5648
rect 9908 5608 10252 5648
rect 10292 5608 10301 5648
rect 12451 5608 12460 5648
rect 12500 5608 12940 5648
rect 12980 5608 12989 5648
rect 2851 5607 2909 5608
rect 4771 5607 4829 5608
rect 2371 5564 2429 5565
rect 6604 5564 6644 5608
rect 8323 5607 8381 5608
rect 2371 5524 2380 5564
rect 2420 5524 6644 5564
rect 9955 5524 9964 5564
rect 10004 5524 10540 5564
rect 10580 5524 10589 5564
rect 12259 5524 12268 5564
rect 12308 5524 12556 5564
rect 12596 5524 14188 5564
rect 14228 5524 14237 5564
rect 15628 5524 17260 5564
rect 17300 5524 17309 5564
rect 2371 5523 2429 5524
rect 0 5480 80 5500
rect 15628 5480 15668 5524
rect 16099 5480 16157 5481
rect 0 5440 1900 5480
rect 1940 5440 1949 5480
rect 2500 5440 15668 5480
rect 15715 5440 15724 5480
rect 15764 5440 16108 5480
rect 16148 5440 16204 5480
rect 16244 5440 16253 5480
rect 0 5420 80 5440
rect 2500 5396 2540 5440
rect 16099 5439 16157 5440
rect 6979 5396 7037 5397
rect 1219 5356 1228 5396
rect 1268 5356 2540 5396
rect 6894 5356 6988 5396
rect 7028 5356 7037 5396
rect 10819 5356 10828 5396
rect 10868 5356 11980 5396
rect 12020 5356 12029 5396
rect 14755 5356 14764 5396
rect 14804 5356 15244 5396
rect 15284 5356 15293 5396
rect 16963 5356 16972 5396
rect 17012 5356 17260 5396
rect 17300 5356 17309 5396
rect 6979 5355 7037 5356
rect 2563 5272 2572 5312
rect 2612 5272 2860 5312
rect 2900 5272 2909 5312
rect 4919 5272 4928 5312
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 5296 5272 5305 5312
rect 6115 5272 6124 5312
rect 6164 5272 18892 5312
rect 18932 5272 18941 5312
rect 20039 5272 20048 5312
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20416 5272 20425 5312
rect 6019 5188 6028 5228
rect 6068 5188 6988 5228
rect 7028 5188 7037 5228
rect 8419 5188 8428 5228
rect 8468 5188 12460 5228
rect 12500 5188 12509 5228
rect 14179 5188 14188 5228
rect 14228 5188 16684 5228
rect 16724 5188 16733 5228
rect 0 5144 80 5164
rect 6979 5144 7037 5145
rect 0 5104 3052 5144
rect 3092 5104 3101 5144
rect 6691 5104 6700 5144
rect 6740 5104 6988 5144
rect 7028 5104 7037 5144
rect 9763 5104 9772 5144
rect 9812 5104 10156 5144
rect 10196 5104 10205 5144
rect 11875 5104 11884 5144
rect 11924 5104 12268 5144
rect 12308 5104 12317 5144
rect 13795 5104 13804 5144
rect 13844 5104 13853 5144
rect 0 5084 80 5104
rect 6979 5103 7037 5104
rect 13804 5060 13844 5104
rect 6211 5020 6220 5060
rect 6260 5020 6740 5060
rect 6787 5020 6796 5060
rect 6836 5020 7660 5060
rect 7700 5020 7709 5060
rect 11779 5020 11788 5060
rect 11828 5020 12556 5060
rect 12596 5020 12844 5060
rect 12884 5020 12893 5060
rect 13804 5020 15532 5060
rect 15572 5020 15581 5060
rect 15907 5020 15916 5060
rect 15956 5020 16492 5060
rect 16532 5020 16541 5060
rect 2947 4976 3005 4977
rect 6700 4976 6740 5020
rect 2947 4936 2956 4976
rect 2996 4936 5164 4976
rect 5204 4936 5213 4976
rect 6700 4936 7756 4976
rect 7796 4936 7805 4976
rect 2947 4935 3005 4936
rect 11980 4892 12020 5020
rect 13027 4976 13085 4977
rect 12067 4936 12076 4976
rect 12116 4936 12748 4976
rect 12788 4936 12797 4976
rect 12942 4936 13036 4976
rect 13076 4936 13085 4976
rect 13795 4936 13804 4976
rect 13844 4936 16108 4976
rect 16148 4936 16157 4976
rect 16771 4936 16780 4976
rect 16820 4936 16972 4976
rect 17012 4936 18412 4976
rect 18452 4936 18461 4976
rect 13027 4935 13085 4936
rect 2659 4852 2668 4892
rect 2708 4852 4588 4892
rect 4628 4852 4637 4892
rect 4867 4852 4876 4892
rect 4916 4852 5548 4892
rect 5588 4852 5597 4892
rect 6403 4852 6412 4892
rect 6452 4852 8812 4892
rect 8852 4852 8861 4892
rect 11980 4852 12172 4892
rect 12212 4852 12221 4892
rect 0 4808 80 4828
rect 4675 4808 4733 4809
rect 0 4768 1804 4808
rect 1844 4768 1853 4808
rect 3427 4768 3436 4808
rect 3476 4768 4684 4808
rect 4724 4768 4733 4808
rect 5731 4768 5740 4808
rect 5780 4768 8564 4808
rect 10147 4768 10156 4808
rect 10196 4768 11212 4808
rect 11252 4768 12460 4808
rect 12500 4768 12509 4808
rect 0 4748 80 4768
rect 4675 4767 4733 4768
rect 8524 4724 8564 4768
rect 2500 4684 7372 4724
rect 7412 4684 7421 4724
rect 8524 4684 13708 4724
rect 13748 4684 13757 4724
rect 2500 4640 2540 4684
rect 1699 4600 1708 4640
rect 1748 4600 2540 4640
rect 2947 4640 3005 4641
rect 3427 4640 3485 4641
rect 2947 4600 2956 4640
rect 2996 4600 3052 4640
rect 3092 4600 3101 4640
rect 3235 4600 3244 4640
rect 3284 4600 3436 4640
rect 3476 4600 3485 4640
rect 5923 4600 5932 4640
rect 5972 4600 7852 4640
rect 7892 4600 8620 4640
rect 8660 4600 8669 4640
rect 9667 4600 9676 4640
rect 9716 4600 12364 4640
rect 12404 4600 12413 4640
rect 2947 4599 3005 4600
rect 3427 4599 3485 4600
rect 13987 4556 14045 4557
rect 3679 4516 3688 4556
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 4056 4516 4065 4556
rect 7075 4516 7084 4556
rect 7124 4516 7756 4556
rect 7796 4516 7805 4556
rect 13027 4516 13036 4556
rect 13076 4516 13996 4556
rect 14036 4516 14045 4556
rect 18799 4516 18808 4556
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 19176 4516 19185 4556
rect 13987 4515 14045 4516
rect 0 4472 80 4492
rect 14467 4472 14525 4473
rect 0 4432 1420 4472
rect 1460 4432 1469 4472
rect 6883 4432 6892 4472
rect 6932 4432 7468 4472
rect 7508 4432 7517 4472
rect 13123 4432 13132 4472
rect 13172 4432 14476 4472
rect 14516 4432 14525 4472
rect 0 4412 80 4432
rect 14467 4431 14525 4432
rect 1987 4348 1996 4388
rect 2036 4348 10924 4388
rect 10964 4348 10973 4388
rect 3619 4264 3628 4304
rect 3668 4264 11596 4304
rect 11636 4264 11645 4304
rect 2467 4180 2476 4220
rect 2516 4180 11500 4220
rect 11540 4180 11549 4220
rect 14179 4180 14188 4220
rect 14228 4180 14956 4220
rect 14996 4180 16108 4220
rect 16148 4180 16157 4220
rect 0 4136 80 4156
rect 8899 4136 8957 4137
rect 0 4096 2284 4136
rect 2324 4096 2333 4136
rect 3427 4096 3436 4136
rect 3476 4096 8908 4136
rect 8948 4096 8957 4136
rect 9763 4096 9772 4136
rect 9812 4096 10060 4136
rect 10100 4096 10109 4136
rect 10435 4096 10444 4136
rect 10484 4096 10636 4136
rect 10676 4096 10685 4136
rect 11779 4096 11788 4136
rect 11828 4096 11980 4136
rect 12020 4096 12556 4136
rect 12596 4096 12605 4136
rect 13699 4096 13708 4136
rect 13748 4096 14764 4136
rect 14804 4096 14813 4136
rect 15235 4096 15244 4136
rect 15284 4096 15820 4136
rect 15860 4096 15869 4136
rect 0 4076 80 4096
rect 8899 4095 8957 4096
rect 2476 4012 6124 4052
rect 6164 4012 6173 4052
rect 8611 4012 8620 4052
rect 8660 4012 10196 4052
rect 2476 3968 2516 4012
rect 3139 3968 3197 3969
rect 10156 3968 10196 4012
rect 13315 3968 13373 3969
rect 2467 3928 2476 3968
rect 2516 3928 2525 3968
rect 3054 3928 3148 3968
rect 3188 3928 3197 3968
rect 4579 3928 4588 3968
rect 4628 3928 4876 3968
rect 4916 3928 4925 3968
rect 7651 3928 7660 3968
rect 7700 3928 8236 3968
rect 8276 3928 8285 3968
rect 10147 3928 10156 3968
rect 10196 3928 13324 3968
rect 13364 3928 13373 3968
rect 3139 3927 3197 3928
rect 13315 3927 13373 3928
rect 2179 3884 2237 3885
rect 7651 3884 7709 3885
rect 2179 3844 2188 3884
rect 2228 3844 2572 3884
rect 2612 3844 2621 3884
rect 7651 3844 7660 3884
rect 7700 3844 9676 3884
rect 9716 3844 9725 3884
rect 2179 3843 2237 3844
rect 7651 3843 7709 3844
rect 0 3800 80 3820
rect 5731 3800 5789 3801
rect 10819 3800 10877 3801
rect 0 3760 2668 3800
rect 2708 3760 2717 3800
rect 4919 3760 4928 3800
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 5296 3760 5305 3800
rect 5646 3760 5740 3800
rect 5780 3760 6124 3800
rect 6164 3760 6173 3800
rect 6307 3760 6316 3800
rect 6356 3760 10828 3800
rect 10868 3760 10877 3800
rect 20039 3760 20048 3800
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20416 3760 20425 3800
rect 0 3740 80 3760
rect 5731 3759 5789 3760
rect 10819 3759 10877 3760
rect 3619 3676 3628 3716
rect 3668 3676 11360 3716
rect 11320 3632 11360 3676
rect 4963 3592 4972 3632
rect 5012 3592 5356 3632
rect 5396 3592 5405 3632
rect 8227 3592 8236 3632
rect 8276 3592 10732 3632
rect 10772 3592 11212 3632
rect 11252 3592 11261 3632
rect 11320 3592 13804 3632
rect 13844 3592 13853 3632
rect 2284 3508 2476 3548
rect 2516 3508 2525 3548
rect 7459 3508 7468 3548
rect 7508 3508 7756 3548
rect 7796 3508 7805 3548
rect 8620 3508 10828 3548
rect 10868 3508 11116 3548
rect 11156 3508 11165 3548
rect 0 3464 80 3484
rect 2284 3464 2324 3508
rect 8620 3464 8660 3508
rect 11011 3464 11069 3465
rect 0 3424 1420 3464
rect 1460 3424 1469 3464
rect 2275 3424 2284 3464
rect 2324 3424 2333 3464
rect 5059 3424 5068 3464
rect 5108 3424 5644 3464
rect 5684 3424 5693 3464
rect 6211 3424 6220 3464
rect 6260 3424 8140 3464
rect 8180 3424 8189 3464
rect 8611 3424 8620 3464
rect 8660 3424 8669 3464
rect 10915 3424 10924 3464
rect 10964 3424 11020 3464
rect 11060 3424 11069 3464
rect 13411 3424 13420 3464
rect 13460 3424 15244 3464
rect 15284 3424 15293 3464
rect 0 3404 80 3424
rect 11011 3423 11069 3424
rect 2371 3380 2429 3381
rect 7651 3380 7709 3381
rect 2179 3340 2188 3380
rect 2228 3340 2380 3380
rect 2420 3340 2429 3380
rect 7566 3340 7660 3380
rect 7700 3340 7709 3380
rect 2371 3339 2429 3340
rect 7651 3339 7709 3340
rect 7756 3340 11732 3380
rect 12355 3340 12364 3380
rect 12404 3340 14188 3380
rect 14228 3340 14237 3380
rect 1603 3256 1612 3296
rect 1652 3256 7564 3296
rect 7604 3256 7613 3296
rect 1699 3172 1708 3212
rect 1748 3172 5164 3212
rect 5204 3172 5213 3212
rect 0 3128 80 3148
rect 7756 3128 7796 3340
rect 11692 3296 11732 3340
rect 10147 3256 10156 3296
rect 10196 3256 10540 3296
rect 10580 3256 10589 3296
rect 10819 3256 10828 3296
rect 10868 3256 11212 3296
rect 11252 3256 11261 3296
rect 11692 3256 14572 3296
rect 14612 3256 14621 3296
rect 7843 3172 7852 3212
rect 7892 3172 8044 3212
rect 8084 3172 8093 3212
rect 9859 3172 9868 3212
rect 9908 3172 10732 3212
rect 10772 3172 10781 3212
rect 11107 3172 11116 3212
rect 11156 3172 14860 3212
rect 14900 3172 14909 3212
rect 0 3088 1940 3128
rect 2947 3088 2956 3128
rect 2996 3088 7796 3128
rect 11299 3088 11308 3128
rect 11348 3088 13228 3128
rect 13268 3088 13277 3128
rect 0 3068 80 3088
rect 1900 3044 1940 3088
rect 11107 3044 11165 3045
rect 1891 3004 1900 3044
rect 1940 3004 1949 3044
rect 2563 3004 2572 3044
rect 2612 3004 3532 3044
rect 3572 3004 3581 3044
rect 3679 3004 3688 3044
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 4056 3004 4065 3044
rect 4195 3004 4204 3044
rect 4244 3004 10156 3044
rect 10196 3004 11116 3044
rect 11156 3004 11165 3044
rect 18799 3004 18808 3044
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 19176 3004 19185 3044
rect 11107 3003 11165 3004
rect 1795 2920 1804 2960
rect 1844 2920 5164 2960
rect 5204 2920 5213 2960
rect 11320 2920 13996 2960
rect 14036 2920 15436 2960
rect 15476 2920 15485 2960
rect 11320 2876 11360 2920
rect 931 2836 940 2876
rect 980 2836 3244 2876
rect 3284 2836 3293 2876
rect 3523 2836 3532 2876
rect 3572 2836 11360 2876
rect 0 2792 80 2812
rect 0 2752 3052 2792
rect 3092 2752 3101 2792
rect 4972 2752 8428 2792
rect 8468 2752 8477 2792
rect 9379 2752 9388 2792
rect 9428 2752 9964 2792
rect 10004 2752 15052 2792
rect 15092 2752 15532 2792
rect 15572 2752 16684 2792
rect 16724 2752 16733 2792
rect 0 2732 80 2752
rect 4972 2708 5012 2752
rect 5347 2708 5405 2709
rect 10531 2708 10589 2709
rect 11299 2708 11357 2709
rect 1612 2668 5012 2708
rect 5059 2668 5068 2708
rect 5108 2668 5356 2708
rect 5396 2668 5405 2708
rect 10435 2668 10444 2708
rect 10484 2668 10540 2708
rect 10580 2668 10589 2708
rect 10915 2668 10924 2708
rect 10964 2668 10973 2708
rect 11214 2668 11308 2708
rect 11348 2668 11357 2708
rect 12931 2668 12940 2708
rect 12980 2668 13228 2708
rect 13268 2668 13277 2708
rect 1612 2540 1652 2668
rect 5347 2667 5405 2668
rect 10531 2667 10589 2668
rect 10924 2624 10964 2668
rect 11299 2667 11357 2668
rect 2851 2584 2860 2624
rect 2900 2584 4204 2624
rect 4244 2584 4253 2624
rect 4675 2584 4684 2624
rect 4724 2584 4972 2624
rect 5012 2584 5021 2624
rect 5251 2584 5260 2624
rect 5300 2584 5309 2624
rect 5443 2584 5452 2624
rect 5492 2584 5932 2624
rect 5972 2584 5981 2624
rect 10051 2584 10060 2624
rect 10100 2584 10964 2624
rect 12067 2624 12125 2625
rect 12067 2584 12076 2624
rect 12116 2584 13268 2624
rect 14179 2584 14188 2624
rect 14228 2584 16876 2624
rect 16916 2584 16925 2624
rect 1603 2500 1612 2540
rect 1652 2500 1661 2540
rect 0 2456 80 2476
rect 5260 2456 5300 2584
rect 10444 2540 10484 2584
rect 12067 2583 12125 2584
rect 13228 2540 13268 2584
rect 10435 2500 10444 2540
rect 10484 2500 10493 2540
rect 13219 2500 13228 2540
rect 13268 2500 13277 2540
rect 5539 2456 5597 2457
rect 0 2416 2380 2456
rect 2420 2416 2429 2456
rect 5155 2416 5164 2456
rect 5204 2416 5213 2456
rect 5260 2416 5548 2456
rect 5588 2416 5597 2456
rect 0 2396 80 2416
rect 355 2372 413 2373
rect 5164 2372 5204 2416
rect 5539 2415 5597 2416
rect 10243 2456 10301 2457
rect 10243 2416 10252 2456
rect 10292 2416 14668 2456
rect 14708 2416 14717 2456
rect 10243 2415 10301 2416
rect 355 2332 364 2372
rect 404 2332 4396 2372
rect 4436 2332 4445 2372
rect 5164 2332 5548 2372
rect 5588 2332 5597 2372
rect 5644 2332 6700 2372
rect 6740 2332 6749 2372
rect 9379 2332 9388 2372
rect 9428 2332 9580 2372
rect 9620 2332 9629 2372
rect 12835 2332 12844 2372
rect 12884 2332 13708 2372
rect 13748 2332 13757 2372
rect 355 2331 413 2332
rect 1123 2288 1181 2289
rect 5644 2288 5684 2332
rect 1123 2248 1132 2288
rect 1172 2248 4492 2288
rect 4532 2248 4541 2288
rect 4919 2248 4928 2288
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 5296 2248 5305 2288
rect 5443 2248 5452 2288
rect 5492 2248 5684 2288
rect 5731 2288 5789 2289
rect 10531 2288 10589 2289
rect 5731 2248 5740 2288
rect 5780 2248 5874 2288
rect 6412 2248 10540 2288
rect 10580 2248 10589 2288
rect 20039 2248 20048 2288
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20416 2248 20425 2288
rect 1123 2247 1181 2248
rect 5731 2247 5789 2248
rect 6412 2204 6452 2248
rect 10531 2247 10589 2248
rect 6595 2204 6653 2205
rect 2083 2164 2092 2204
rect 2132 2164 6452 2204
rect 6510 2164 6604 2204
rect 6644 2164 6653 2204
rect 6595 2163 6653 2164
rect 8131 2204 8189 2205
rect 8131 2164 8140 2204
rect 8180 2164 11308 2204
rect 11348 2164 11357 2204
rect 8131 2163 8189 2164
rect 0 2120 80 2140
rect 5347 2120 5405 2121
rect 0 2080 1900 2120
rect 1940 2080 1949 2120
rect 5251 2080 5260 2120
rect 5300 2080 5356 2120
rect 5396 2080 5405 2120
rect 0 2060 80 2080
rect 5347 2079 5405 2080
rect 6691 2120 6749 2121
rect 16867 2120 16925 2121
rect 6691 2080 6700 2120
rect 6740 2080 6988 2120
rect 7028 2080 7037 2120
rect 10915 2080 10924 2120
rect 10964 2080 16876 2120
rect 16916 2080 16925 2120
rect 6691 2079 6749 2080
rect 16867 2079 16925 2080
rect 16579 2036 16637 2037
rect 9772 1996 10060 2036
rect 10100 1996 10109 2036
rect 10531 1996 10540 2036
rect 10580 1996 16588 2036
rect 16628 1996 16637 2036
rect 163 1952 221 1953
rect 5539 1952 5597 1953
rect 9772 1952 9812 1996
rect 16579 1995 16637 1996
rect 163 1912 172 1952
rect 212 1912 4204 1952
rect 4244 1912 4253 1952
rect 4963 1912 4972 1952
rect 5012 1912 5548 1952
rect 5588 1912 5597 1952
rect 163 1911 221 1912
rect 5539 1911 5597 1912
rect 5740 1912 9812 1952
rect 9859 1912 9868 1952
rect 9908 1912 11212 1952
rect 11252 1912 11261 1952
rect 2467 1868 2525 1869
rect 5740 1868 5780 1912
rect 2382 1828 2476 1868
rect 2516 1828 2525 1868
rect 4291 1828 4300 1868
rect 4340 1828 5780 1868
rect 5827 1868 5885 1869
rect 12259 1868 12317 1869
rect 12931 1868 12989 1869
rect 14083 1868 14141 1869
rect 5827 1828 5836 1868
rect 5876 1828 7852 1868
rect 7892 1828 7901 1868
rect 8227 1828 8236 1868
rect 8276 1828 8812 1868
rect 8852 1828 8861 1868
rect 12174 1828 12268 1868
rect 12308 1828 12317 1868
rect 12846 1828 12940 1868
rect 12980 1828 12989 1868
rect 13891 1828 13900 1868
rect 13940 1828 14092 1868
rect 14132 1828 14141 1868
rect 2467 1827 2525 1828
rect 5827 1827 5885 1828
rect 12259 1827 12317 1828
rect 12931 1827 12989 1828
rect 14083 1827 14141 1828
rect 14275 1868 14333 1869
rect 15235 1868 15293 1869
rect 14275 1828 14284 1868
rect 14324 1828 14418 1868
rect 15150 1828 15244 1868
rect 15284 1828 15293 1868
rect 14275 1827 14333 1828
rect 15235 1827 15293 1828
rect 15523 1868 15581 1869
rect 16003 1868 16061 1869
rect 15523 1828 15532 1868
rect 15572 1828 15628 1868
rect 15668 1828 15677 1868
rect 15918 1828 16012 1868
rect 16052 1828 16061 1868
rect 16387 1828 16396 1868
rect 16436 1828 20524 1868
rect 20564 1828 20573 1868
rect 15523 1827 15581 1828
rect 16003 1827 16061 1828
rect 0 1784 80 1804
rect 0 1744 1516 1784
rect 1556 1744 1565 1784
rect 1987 1744 1996 1784
rect 2036 1744 12844 1784
rect 12884 1744 12893 1784
rect 0 1724 80 1744
rect 3331 1660 3340 1700
rect 3380 1660 3389 1700
rect 4483 1660 4492 1700
rect 4532 1660 9004 1700
rect 9044 1660 9484 1700
rect 9524 1660 9533 1700
rect 9580 1660 10924 1700
rect 10964 1660 10973 1700
rect 11491 1660 11500 1700
rect 11540 1660 12364 1700
rect 12404 1660 12413 1700
rect 3340 1616 3380 1660
rect 3340 1576 9524 1616
rect 931 1532 989 1533
rect 9484 1532 9524 1576
rect 931 1492 940 1532
rect 980 1492 2540 1532
rect 3679 1492 3688 1532
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 4056 1492 4065 1532
rect 4387 1492 4396 1532
rect 4436 1492 7988 1532
rect 8419 1492 8428 1532
rect 8468 1492 9196 1532
rect 9236 1492 9245 1532
rect 9475 1492 9484 1532
rect 9524 1492 9533 1532
rect 931 1491 989 1492
rect 0 1448 80 1468
rect 2500 1448 2540 1492
rect 7948 1448 7988 1492
rect 9580 1448 9620 1660
rect 11491 1616 11549 1617
rect 14659 1616 14717 1617
rect 10531 1576 10540 1616
rect 10580 1576 11500 1616
rect 11540 1576 11549 1616
rect 13315 1576 13324 1616
rect 13364 1576 14668 1616
rect 14708 1576 14717 1616
rect 11491 1575 11549 1576
rect 14659 1575 14717 1576
rect 9859 1492 9868 1532
rect 9908 1492 12748 1532
rect 12788 1492 12797 1532
rect 18799 1492 18808 1532
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 19176 1492 19185 1532
rect 0 1408 2284 1448
rect 2324 1408 2333 1448
rect 2500 1408 4684 1448
rect 4724 1408 4733 1448
rect 5347 1408 5356 1448
rect 5396 1408 5548 1448
rect 5588 1408 5597 1448
rect 6787 1408 6796 1448
rect 6836 1408 7852 1448
rect 7892 1408 7901 1448
rect 7948 1408 9620 1448
rect 10723 1408 10732 1448
rect 10772 1408 11980 1448
rect 12020 1408 12029 1448
rect 14275 1408 14284 1448
rect 14324 1408 15436 1448
rect 15476 1408 15485 1448
rect 0 1388 80 1408
rect 2275 1364 2333 1365
rect 2275 1324 2284 1364
rect 2324 1324 6220 1364
rect 6260 1324 6269 1364
rect 7171 1324 7180 1364
rect 7220 1324 8044 1364
rect 8084 1324 8093 1364
rect 10627 1324 10636 1364
rect 10676 1324 11692 1364
rect 11732 1324 11741 1364
rect 2275 1323 2333 1324
rect 5443 1280 5501 1281
rect 6691 1280 6749 1281
rect 7363 1280 7421 1281
rect 7747 1280 7805 1281
rect 12739 1280 12797 1281
rect 13891 1280 13949 1281
rect 15619 1280 15677 1281
rect 17347 1280 17405 1281
rect 17731 1280 17789 1281
rect 18115 1280 18173 1281
rect 18499 1280 18557 1281
rect 19267 1280 19325 1281
rect 1027 1240 1036 1280
rect 1076 1240 3148 1280
rect 3188 1240 3197 1280
rect 3907 1240 3916 1280
rect 3956 1240 5452 1280
rect 5492 1240 5501 1280
rect 6606 1240 6700 1280
rect 6740 1240 6749 1280
rect 7278 1240 7372 1280
rect 7412 1240 7421 1280
rect 7662 1240 7756 1280
rect 7796 1240 7805 1280
rect 8131 1240 8140 1280
rect 8180 1240 8716 1280
rect 8756 1240 8765 1280
rect 11107 1240 11116 1280
rect 11156 1240 12172 1280
rect 12212 1240 12221 1280
rect 12654 1240 12748 1280
rect 12788 1240 12797 1280
rect 13806 1240 13900 1280
rect 13940 1240 13949 1280
rect 15534 1240 15628 1280
rect 15668 1240 15677 1280
rect 17262 1240 17356 1280
rect 17396 1240 17405 1280
rect 17539 1240 17548 1280
rect 17588 1240 17740 1280
rect 17780 1240 17789 1280
rect 18030 1240 18124 1280
rect 18164 1240 18173 1280
rect 18414 1240 18508 1280
rect 18548 1240 18557 1280
rect 19182 1240 19276 1280
rect 19316 1240 19325 1280
rect 5443 1239 5501 1240
rect 6691 1239 6749 1240
rect 7363 1239 7421 1240
rect 7747 1239 7805 1240
rect 12739 1239 12797 1240
rect 13891 1239 13949 1240
rect 15619 1239 15677 1240
rect 17347 1239 17405 1240
rect 17731 1239 17789 1240
rect 18115 1239 18173 1240
rect 18499 1239 18557 1240
rect 19267 1239 19325 1240
rect 19459 1280 19517 1281
rect 19459 1240 19468 1280
rect 19508 1240 19602 1280
rect 19459 1239 19517 1240
rect 8803 1196 8861 1197
rect 16771 1196 16829 1197
rect 19651 1196 19709 1197
rect 1123 1156 1132 1196
rect 1172 1156 4108 1196
rect 4148 1156 4157 1196
rect 6115 1156 6124 1196
rect 6164 1156 7180 1196
rect 7220 1156 7229 1196
rect 7939 1156 7948 1196
rect 7988 1156 8524 1196
rect 8564 1156 8573 1196
rect 8803 1156 8812 1196
rect 8852 1156 9004 1196
rect 9044 1156 9053 1196
rect 10147 1156 10156 1196
rect 10196 1156 10828 1196
rect 10868 1156 10877 1196
rect 15139 1156 15148 1196
rect 15188 1156 16780 1196
rect 16820 1156 16829 1196
rect 19075 1156 19084 1196
rect 19124 1156 19660 1196
rect 19700 1156 19709 1196
rect 8803 1155 8861 1156
rect 16771 1155 16829 1156
rect 19651 1155 19709 1156
rect 0 1112 80 1132
rect 6883 1112 6941 1113
rect 12547 1112 12605 1113
rect 20707 1112 20765 1113
rect 0 1072 1516 1112
rect 1556 1072 1565 1112
rect 6211 1072 6220 1112
rect 6260 1072 6892 1112
rect 6932 1072 6941 1112
rect 12462 1072 12556 1112
rect 12596 1072 12605 1112
rect 0 1052 80 1072
rect 6883 1071 6941 1072
rect 12547 1071 12605 1072
rect 14668 1072 14956 1112
rect 14996 1072 15005 1112
rect 18883 1072 18892 1112
rect 18932 1072 20716 1112
rect 20756 1072 20765 1112
rect 6211 1028 6269 1029
rect 14668 1028 14708 1072
rect 20707 1071 20765 1072
rect 20515 1028 20573 1029
rect 1795 988 1804 1028
rect 1844 988 6220 1028
rect 6260 988 6269 1028
rect 6403 988 6412 1028
rect 6452 988 7756 1028
rect 7796 988 7805 1028
rect 7852 988 14708 1028
rect 14851 988 14860 1028
rect 14900 988 15436 1028
rect 15476 988 15485 1028
rect 16003 988 16012 1028
rect 16052 988 16300 1028
rect 16340 988 16349 1028
rect 17923 988 17932 1028
rect 17972 988 20524 1028
rect 20564 988 20573 1028
rect 6211 987 6269 988
rect 1219 944 1277 945
rect 6307 944 6365 945
rect 7075 944 7133 945
rect 1219 904 1228 944
rect 1268 904 5932 944
rect 5972 904 5981 944
rect 6222 904 6316 944
rect 6356 904 6365 944
rect 6787 904 6796 944
rect 6836 904 7084 944
rect 7124 904 7133 944
rect 1219 903 1277 904
rect 6307 903 6365 904
rect 7075 903 7133 904
rect 7852 860 7892 988
rect 20515 987 20573 988
rect 18307 944 18365 945
rect 9187 904 9196 944
rect 9236 904 10060 944
rect 10100 904 10109 944
rect 11107 904 11116 944
rect 11156 904 11788 944
rect 11828 904 11837 944
rect 14467 904 14476 944
rect 14516 904 14956 944
rect 14996 904 15005 944
rect 18222 904 18316 944
rect 18356 904 18365 944
rect 18307 903 18365 904
rect 15043 860 15101 861
rect 20611 860 20669 861
rect 2083 820 2092 860
rect 2132 820 2540 860
rect 5827 820 5836 860
rect 5876 820 7892 860
rect 8803 820 8812 860
rect 8852 820 10252 860
rect 10292 820 10301 860
rect 13699 820 13708 860
rect 13748 820 15052 860
rect 15092 820 15101 860
rect 15235 820 15244 860
rect 15284 820 16204 860
rect 16244 820 16253 860
rect 17731 820 17740 860
rect 17780 820 20620 860
rect 20660 820 20669 860
rect 0 776 80 796
rect 0 736 2284 776
rect 2324 736 2333 776
rect 0 716 80 736
rect 2500 692 2540 820
rect 15043 819 15101 820
rect 20611 819 20669 820
rect 6403 776 6461 777
rect 6979 776 7037 777
rect 4919 736 4928 776
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 5296 736 5305 776
rect 6318 736 6412 776
rect 6452 736 6461 776
rect 6894 736 6988 776
rect 7028 736 7037 776
rect 9091 736 9100 776
rect 9140 736 11212 776
rect 11252 736 11261 776
rect 13411 736 13420 776
rect 13460 736 14092 776
rect 14132 736 14141 776
rect 15100 736 15724 776
rect 15764 736 15773 776
rect 20039 736 20048 776
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20416 736 20425 776
rect 6403 735 6461 736
rect 6979 735 7037 736
rect 14179 692 14237 693
rect 1315 652 1324 692
rect 1364 652 2188 692
rect 2228 652 2237 692
rect 2500 652 8620 692
rect 8660 652 8669 692
rect 13507 652 13516 692
rect 13556 652 14188 692
rect 14228 652 14237 692
rect 14179 651 14237 652
rect 15100 608 15140 736
rect 4195 568 4204 608
rect 4244 568 4876 608
rect 4916 568 4925 608
rect 5059 568 5068 608
rect 5108 568 5588 608
rect 6499 568 6508 608
rect 6548 568 7372 608
rect 7412 568 7421 608
rect 7555 568 7564 608
rect 7604 568 8140 608
rect 8180 568 8189 608
rect 9091 568 9100 608
rect 9140 568 15140 608
rect 17923 608 17981 609
rect 17923 568 17932 608
rect 17972 568 18700 608
rect 18740 568 18749 608
rect 2083 524 2141 525
rect 5548 524 5588 568
rect 17923 567 17981 568
rect 9859 524 9917 525
rect 2083 484 2092 524
rect 2132 484 5452 524
rect 5492 484 5501 524
rect 5548 484 9868 524
rect 9908 484 9917 524
rect 10723 484 10732 524
rect 10772 484 11596 524
rect 11636 484 11645 524
rect 15043 484 15052 524
rect 15092 484 15820 524
rect 15860 484 15869 524
rect 2083 483 2141 484
rect 9859 483 9917 484
rect 0 440 80 460
rect 9283 440 9341 441
rect 0 400 2668 440
rect 2708 400 2717 440
rect 5635 400 5644 440
rect 5684 400 6604 440
rect 6644 400 6653 440
rect 6883 400 6892 440
rect 6932 400 7564 440
rect 7604 400 7613 440
rect 7660 400 9292 440
rect 9332 400 9341 440
rect 9955 400 9964 440
rect 10004 400 10828 440
rect 10868 400 10877 440
rect 0 380 80 400
rect 3715 356 3773 357
rect 7660 356 7700 400
rect 9283 399 9341 400
rect 3630 316 3724 356
rect 3764 316 3773 356
rect 3715 315 3773 316
rect 3820 316 7700 356
rect 8899 316 8908 356
rect 8948 316 14956 356
rect 14996 316 15005 356
rect 15523 316 15532 356
rect 15572 316 15820 356
rect 15860 316 15869 356
rect 2947 272 3005 273
rect 3820 272 3860 316
rect 2862 232 2956 272
rect 2996 232 3005 272
rect 3523 232 3532 272
rect 3572 232 3860 272
rect 6019 232 6028 272
rect 6068 232 12076 272
rect 12116 232 12125 272
rect 2947 231 3005 232
rect 5251 188 5309 189
rect 13699 188 13757 189
rect 1891 148 1900 188
rect 1940 148 1949 188
rect 5166 148 5260 188
rect 5300 148 5309 188
rect 6595 148 6604 188
rect 6644 148 13708 188
rect 13748 148 13757 188
rect 0 104 80 124
rect 1900 104 1940 148
rect 5251 147 5309 148
rect 13699 147 13757 148
rect 11779 104 11837 105
rect 0 64 1940 104
rect 4483 64 4492 104
rect 4532 64 11788 104
rect 11828 64 11837 104
rect 0 44 80 64
rect 11779 63 11837 64
<< via3 >>
rect 15724 85576 15764 85616
rect 4780 85408 4820 85448
rect 1324 85072 1364 85112
rect 8236 84904 8276 84944
rect 15916 84904 15956 84944
rect 76 84736 116 84776
rect 3688 84652 3728 84692
rect 3770 84652 3810 84692
rect 3852 84652 3892 84692
rect 3934 84652 3974 84692
rect 4016 84652 4056 84692
rect 18808 84652 18848 84692
rect 18890 84652 18930 84692
rect 18972 84652 19012 84692
rect 19054 84652 19094 84692
rect 19136 84652 19176 84692
rect 5548 84484 5588 84524
rect 7372 84484 7412 84524
rect 12364 84484 12404 84524
rect 12844 84484 12884 84524
rect 5836 84400 5876 84440
rect 6124 84400 6164 84440
rect 6412 84400 6452 84440
rect 6700 84400 6740 84440
rect 7180 84400 7220 84440
rect 9676 84400 9716 84440
rect 10252 84400 10292 84440
rect 10444 84400 10484 84440
rect 11788 84400 11828 84440
rect 12940 84400 12980 84440
rect 13324 84400 13364 84440
rect 14092 84400 14132 84440
rect 16396 84400 16436 84440
rect 16876 84400 16916 84440
rect 3244 84316 3284 84356
rect 1228 84232 1268 84272
rect 4928 83896 4968 83936
rect 5010 83896 5050 83936
rect 5092 83896 5132 83936
rect 5174 83896 5214 83936
rect 5256 83896 5296 83936
rect 20048 83896 20088 83936
rect 20130 83896 20170 83936
rect 20212 83896 20252 83936
rect 20294 83896 20334 83936
rect 20376 83896 20416 83936
rect 2956 83476 2996 83516
rect 4396 83476 4436 83516
rect 6028 83476 6068 83516
rect 7756 83476 7796 83516
rect 9772 83476 9812 83516
rect 11020 83476 11060 83516
rect 11692 83476 11732 83516
rect 18316 83476 18356 83516
rect 18604 83476 18644 83516
rect 19084 83476 19124 83516
rect 19564 83476 19604 83516
rect 7084 83392 7124 83432
rect 2572 83308 2612 83348
rect 13132 83308 13172 83348
rect 13996 83308 14036 83348
rect 14476 83308 14516 83348
rect 14668 83308 14708 83348
rect 15052 83308 15092 83348
rect 7660 83224 7700 83264
rect 3688 83140 3728 83180
rect 3770 83140 3810 83180
rect 3852 83140 3892 83180
rect 3934 83140 3974 83180
rect 4016 83140 4056 83180
rect 10828 83140 10868 83180
rect 12748 83140 12788 83180
rect 18808 83140 18848 83180
rect 18890 83140 18930 83180
rect 18972 83140 19012 83180
rect 19054 83140 19094 83180
rect 19136 83140 19176 83180
rect 1900 83056 1940 83096
rect 2476 82720 2516 82760
rect 1900 82636 1940 82676
rect 14188 82552 14228 82592
rect 17356 82552 17396 82592
rect 17740 82552 17780 82592
rect 19468 82552 19508 82592
rect 4300 82384 4340 82424
rect 4928 82384 4968 82424
rect 5010 82384 5050 82424
rect 5092 82384 5132 82424
rect 5174 82384 5214 82424
rect 5256 82384 5296 82424
rect 20048 82384 20088 82424
rect 20130 82384 20170 82424
rect 20212 82384 20252 82424
rect 20294 82384 20334 82424
rect 20376 82384 20416 82424
rect 18412 81964 18452 82004
rect 18124 81880 18164 81920
rect 18508 81880 18548 81920
rect 19276 81880 19316 81920
rect 7564 81796 7604 81836
rect 13900 81796 13940 81836
rect 3688 81628 3728 81668
rect 3770 81628 3810 81668
rect 3852 81628 3892 81668
rect 3934 81628 3974 81668
rect 4016 81628 4056 81668
rect 18808 81628 18848 81668
rect 18890 81628 18930 81668
rect 18972 81628 19012 81668
rect 19054 81628 19094 81668
rect 19136 81628 19176 81668
rect 1612 81040 1652 81080
rect 4928 80872 4968 80912
rect 5010 80872 5050 80912
rect 5092 80872 5132 80912
rect 5174 80872 5214 80912
rect 5256 80872 5296 80912
rect 20048 80872 20088 80912
rect 20130 80872 20170 80912
rect 20212 80872 20252 80912
rect 20294 80872 20334 80912
rect 20376 80872 20416 80912
rect 2764 80704 2804 80744
rect 1612 80536 1652 80576
rect 2284 80536 2324 80576
rect 2476 80536 2516 80576
rect 5452 80452 5492 80492
rect 1516 80368 1556 80408
rect 6796 80368 6836 80408
rect 3688 80116 3728 80156
rect 3770 80116 3810 80156
rect 3852 80116 3892 80156
rect 3934 80116 3974 80156
rect 4016 80116 4056 80156
rect 18808 80116 18848 80156
rect 18890 80116 18930 80156
rect 18972 80116 19012 80156
rect 19054 80116 19094 80156
rect 19136 80116 19176 80156
rect 844 79948 884 79988
rect 5356 79780 5396 79820
rect 2284 79696 2324 79736
rect 4684 79696 4724 79736
rect 9004 79612 9044 79652
rect 12172 79528 12212 79568
rect 3148 79360 3188 79400
rect 4928 79360 4968 79400
rect 5010 79360 5050 79400
rect 5092 79360 5132 79400
rect 5174 79360 5214 79400
rect 5256 79360 5296 79400
rect 20048 79360 20088 79400
rect 20130 79360 20170 79400
rect 20212 79360 20252 79400
rect 20294 79360 20334 79400
rect 20376 79360 20416 79400
rect 1900 78940 1940 78980
rect 1516 78856 1556 78896
rect 3688 78604 3728 78644
rect 3770 78604 3810 78644
rect 3852 78604 3892 78644
rect 3934 78604 3974 78644
rect 4016 78604 4056 78644
rect 18808 78604 18848 78644
rect 18890 78604 18930 78644
rect 18972 78604 19012 78644
rect 19054 78604 19094 78644
rect 19136 78604 19176 78644
rect 3148 78184 3188 78224
rect 7468 78100 7508 78140
rect 4204 77932 4244 77972
rect 4928 77848 4968 77888
rect 5010 77848 5050 77888
rect 5092 77848 5132 77888
rect 5174 77848 5214 77888
rect 5256 77848 5296 77888
rect 20048 77848 20088 77888
rect 20130 77848 20170 77888
rect 20212 77848 20252 77888
rect 20294 77848 20334 77888
rect 20376 77848 20416 77888
rect 21196 77848 21236 77888
rect 3340 77680 3380 77720
rect 2956 77512 2996 77552
rect 4780 77512 4820 77552
rect 3436 77428 3476 77468
rect 21388 77176 21428 77216
rect 3688 77092 3728 77132
rect 3770 77092 3810 77132
rect 3852 77092 3892 77132
rect 3934 77092 3974 77132
rect 4016 77092 4056 77132
rect 18808 77092 18848 77132
rect 18890 77092 18930 77132
rect 18972 77092 19012 77132
rect 19054 77092 19094 77132
rect 19136 77092 19176 77132
rect 6508 76924 6548 76964
rect 4588 76840 4628 76880
rect 1996 76672 2036 76712
rect 8812 76588 8852 76628
rect 3532 76504 3572 76544
rect 4928 76336 4968 76376
rect 5010 76336 5050 76376
rect 5092 76336 5132 76376
rect 5174 76336 5214 76376
rect 5256 76336 5296 76376
rect 20048 76336 20088 76376
rect 20130 76336 20170 76376
rect 20212 76336 20252 76376
rect 20294 76336 20334 76376
rect 20376 76336 20416 76376
rect 364 76000 404 76040
rect 1804 76000 1844 76040
rect 4588 75916 4628 75956
rect 4780 75916 4820 75956
rect 8524 75916 8564 75956
rect 7468 75664 7508 75704
rect 3688 75580 3728 75620
rect 3770 75580 3810 75620
rect 3852 75580 3892 75620
rect 3934 75580 3974 75620
rect 4016 75580 4056 75620
rect 6508 75580 6548 75620
rect 9580 75580 9620 75620
rect 10636 75580 10676 75620
rect 18808 75580 18848 75620
rect 18890 75580 18930 75620
rect 18972 75580 19012 75620
rect 19054 75580 19094 75620
rect 19136 75580 19176 75620
rect 11308 75412 11348 75452
rect 3148 75244 3188 75284
rect 9196 75244 9236 75284
rect 10444 75244 10484 75284
rect 11020 75160 11060 75200
rect 6028 75076 6068 75116
rect 8908 74908 8948 74948
rect 9196 74908 9236 74948
rect 4928 74824 4968 74864
rect 5010 74824 5050 74864
rect 5092 74824 5132 74864
rect 5174 74824 5214 74864
rect 5256 74824 5296 74864
rect 20048 74824 20088 74864
rect 20130 74824 20170 74864
rect 20212 74824 20252 74864
rect 20294 74824 20334 74864
rect 20376 74824 20416 74864
rect 10156 74740 10196 74780
rect 9388 74656 9428 74696
rect 8812 74572 8852 74612
rect 9292 74572 9332 74612
rect 6028 74488 6068 74528
rect 8812 74404 8852 74444
rect 6988 74320 7028 74360
rect 8908 74320 8948 74360
rect 10636 74320 10676 74360
rect 4108 74236 4148 74276
rect 3688 74068 3728 74108
rect 3770 74068 3810 74108
rect 3852 74068 3892 74108
rect 3934 74068 3974 74108
rect 4016 74068 4056 74108
rect 18808 74068 18848 74108
rect 18890 74068 18930 74108
rect 18972 74068 19012 74108
rect 19054 74068 19094 74108
rect 19136 74068 19176 74108
rect 2476 73816 2516 73856
rect 9964 73816 10004 73856
rect 16300 73816 16340 73856
rect 6988 73648 7028 73688
rect 6508 73480 6548 73520
rect 4928 73312 4968 73352
rect 5010 73312 5050 73352
rect 5092 73312 5132 73352
rect 5174 73312 5214 73352
rect 5256 73312 5296 73352
rect 20048 73312 20088 73352
rect 20130 73312 20170 73352
rect 20212 73312 20252 73352
rect 20294 73312 20334 73352
rect 20376 73312 20416 73352
rect 1708 72976 1748 73016
rect 2284 72976 2324 73016
rect 3532 73060 3572 73100
rect 2476 72976 2516 73016
rect 3148 72976 3188 73016
rect 10732 72724 10772 72764
rect 3532 72556 3572 72596
rect 3688 72556 3728 72596
rect 3770 72556 3810 72596
rect 3852 72556 3892 72596
rect 3934 72556 3974 72596
rect 4016 72556 4056 72596
rect 460 72472 500 72512
rect 18808 72556 18848 72596
rect 18890 72556 18930 72596
rect 18972 72556 19012 72596
rect 19054 72556 19094 72596
rect 19136 72556 19176 72596
rect 7756 72472 7796 72512
rect 8908 72472 8948 72512
rect 8428 72388 8468 72428
rect 8812 72304 8852 72344
rect 6028 72220 6068 72260
rect 6220 72220 6260 72260
rect 3052 71968 3092 72008
rect 5644 71968 5684 72008
rect 6220 71968 6260 72008
rect 6604 71968 6644 72008
rect 12460 72136 12500 72176
rect 9100 72052 9140 72092
rect 15244 72052 15284 72092
rect 13804 71968 13844 72008
rect 2476 71884 2516 71924
rect 4928 71800 4968 71840
rect 5010 71800 5050 71840
rect 5092 71800 5132 71840
rect 5174 71800 5214 71840
rect 5256 71800 5296 71840
rect 6604 71800 6644 71840
rect 11596 71800 11636 71840
rect 12364 71800 12404 71840
rect 20048 71800 20088 71840
rect 20130 71800 20170 71840
rect 20212 71800 20252 71840
rect 20294 71800 20334 71840
rect 20376 71800 20416 71840
rect 3340 71716 3380 71756
rect 1900 71464 1940 71504
rect 12172 71464 12212 71504
rect 19372 71464 19412 71504
rect 3532 71380 3572 71420
rect 2092 71212 2132 71252
rect 15820 71212 15860 71252
rect 9868 71128 9908 71168
rect 3688 71044 3728 71084
rect 3770 71044 3810 71084
rect 3852 71044 3892 71084
rect 3934 71044 3974 71084
rect 4016 71044 4056 71084
rect 18808 71044 18848 71084
rect 18890 71044 18930 71084
rect 18972 71044 19012 71084
rect 19054 71044 19094 71084
rect 19136 71044 19176 71084
rect 16012 70960 16052 71000
rect 3148 70792 3188 70832
rect 10540 70792 10580 70832
rect 15628 70792 15668 70832
rect 1420 70708 1460 70748
rect 4108 70708 4148 70748
rect 6988 70708 7028 70748
rect 2188 70624 2228 70664
rect 4780 70624 4820 70664
rect 8140 70624 8180 70664
rect 9292 70624 9332 70664
rect 7756 70456 7796 70496
rect 9964 70372 10004 70412
rect 4928 70288 4968 70328
rect 5010 70288 5050 70328
rect 5092 70288 5132 70328
rect 5174 70288 5214 70328
rect 5256 70288 5296 70328
rect 15820 70372 15860 70412
rect 15628 70288 15668 70328
rect 20048 70288 20088 70328
rect 20130 70288 20170 70328
rect 20212 70288 20252 70328
rect 20294 70288 20334 70328
rect 20376 70288 20416 70328
rect 14956 70204 14996 70244
rect 19660 70120 19700 70160
rect 2860 70036 2900 70076
rect 1324 69952 1364 69992
rect 4300 69952 4340 69992
rect 11692 69952 11732 69992
rect 12556 69952 12596 69992
rect 2668 69700 2708 69740
rect 3148 69700 3188 69740
rect 5740 69868 5780 69908
rect 11884 69868 11924 69908
rect 11500 69784 11540 69824
rect 3436 69700 3476 69740
rect 16012 69616 16052 69656
rect 3688 69532 3728 69572
rect 3770 69532 3810 69572
rect 3852 69532 3892 69572
rect 3934 69532 3974 69572
rect 4016 69532 4056 69572
rect 4780 69532 4820 69572
rect 10156 69532 10196 69572
rect 18808 69532 18848 69572
rect 18890 69532 18930 69572
rect 18972 69532 19012 69572
rect 19054 69532 19094 69572
rect 19136 69532 19176 69572
rect 16012 69448 16052 69488
rect 16780 69448 16820 69488
rect 3244 69364 3284 69404
rect 8812 69280 8852 69320
rect 9196 69280 9236 69320
rect 9676 69280 9716 69320
rect 10348 69280 10388 69320
rect 13612 69280 13652 69320
rect 2764 69196 2804 69236
rect 19372 69196 19412 69236
rect 9772 69112 9812 69152
rect 11020 69112 11060 69152
rect 2764 68944 2804 68984
rect 7276 68944 7316 68984
rect 4928 68776 4968 68816
rect 5010 68776 5050 68816
rect 5092 68776 5132 68816
rect 5174 68776 5214 68816
rect 5256 68776 5296 68816
rect 20048 68776 20088 68816
rect 20130 68776 20170 68816
rect 20212 68776 20252 68816
rect 20294 68776 20334 68816
rect 20376 68776 20416 68816
rect 5548 68608 5588 68648
rect 3436 68524 3476 68564
rect 3628 68524 3668 68564
rect 4876 68524 4916 68564
rect 17164 68356 17204 68396
rect 4780 68272 4820 68312
rect 4108 68188 4148 68228
rect 7084 68272 7124 68312
rect 8620 68272 8660 68312
rect 1708 68104 1748 68144
rect 3688 68020 3728 68060
rect 3770 68020 3810 68060
rect 3852 68020 3892 68060
rect 3934 68020 3974 68060
rect 4016 68020 4056 68060
rect 7948 68020 7988 68060
rect 18808 68020 18848 68060
rect 18890 68020 18930 68060
rect 18972 68020 19012 68060
rect 19054 68020 19094 68060
rect 19136 68020 19176 68060
rect 15148 67852 15188 67892
rect 20140 67768 20180 67808
rect 1612 67684 1652 67724
rect 10156 67684 10196 67724
rect 13228 67600 13268 67640
rect 15340 67516 15380 67556
rect 3820 67432 3860 67472
rect 11404 67432 11444 67472
rect 3436 67264 3476 67304
rect 4928 67264 4968 67304
rect 5010 67264 5050 67304
rect 5092 67264 5132 67304
rect 5174 67264 5214 67304
rect 5256 67264 5296 67304
rect 20048 67264 20088 67304
rect 20130 67264 20170 67304
rect 20212 67264 20252 67304
rect 20294 67264 20334 67304
rect 20376 67264 20416 67304
rect 13516 67180 13556 67220
rect 76 67096 116 67136
rect 9196 67096 9236 67136
rect 12460 67096 12500 67136
rect 2764 66928 2804 66968
rect 364 66844 404 66884
rect 748 66760 788 66800
rect 2956 66760 2996 66800
rect 4780 66760 4820 66800
rect 17548 66760 17588 66800
rect 19948 66760 19988 66800
rect 7468 66676 7508 66716
rect 1132 66592 1172 66632
rect 6028 66592 6068 66632
rect 6316 66592 6356 66632
rect 12652 66592 12692 66632
rect 3688 66508 3728 66548
rect 3770 66508 3810 66548
rect 3852 66508 3892 66548
rect 3934 66508 3974 66548
rect 4016 66508 4056 66548
rect 4588 66508 4628 66548
rect 13132 66508 13172 66548
rect 18808 66508 18848 66548
rect 18890 66508 18930 66548
rect 18972 66508 19012 66548
rect 19054 66508 19094 66548
rect 19136 66508 19176 66548
rect 13036 66424 13076 66464
rect 16108 66424 16148 66464
rect 6892 66340 6932 66380
rect 13804 66340 13844 66380
rect 4588 66256 4628 66296
rect 8044 66088 8084 66128
rect 16012 66088 16052 66128
rect 5548 66004 5588 66044
rect 2860 65920 2900 65960
rect 10348 65920 10388 65960
rect 14380 65920 14420 65960
rect 13612 65836 13652 65876
rect 4928 65752 4968 65792
rect 5010 65752 5050 65792
rect 5092 65752 5132 65792
rect 5174 65752 5214 65792
rect 5256 65752 5296 65792
rect 7852 65752 7892 65792
rect 13420 65752 13460 65792
rect 20048 65752 20088 65792
rect 20130 65752 20170 65792
rect 20212 65752 20252 65792
rect 20294 65752 20334 65792
rect 20376 65752 20416 65792
rect 6028 65668 6068 65708
rect 3148 65584 3188 65624
rect 3436 65584 3476 65624
rect 17452 65584 17492 65624
rect 556 65500 596 65540
rect 17644 65500 17684 65540
rect 2092 65416 2132 65456
rect 15916 65416 15956 65456
rect 1612 65332 1652 65372
rect 1804 65332 1844 65372
rect 9484 65332 9524 65372
rect 6316 65248 6356 65288
rect 5548 65164 5588 65204
rect 3688 64996 3728 65036
rect 3770 64996 3810 65036
rect 3852 64996 3892 65036
rect 3934 64996 3974 65036
rect 4016 64996 4056 65036
rect 18808 64996 18848 65036
rect 18890 64996 18930 65036
rect 18972 64996 19012 65036
rect 19054 64996 19094 65036
rect 19136 64996 19176 65036
rect 940 64828 980 64868
rect 5932 64828 5972 64868
rect 13132 64828 13172 64868
rect 1324 64660 1364 64700
rect 8620 64660 8660 64700
rect 9484 64660 9524 64700
rect 11116 64408 11156 64448
rect 13612 64408 13652 64448
rect 5932 64324 5972 64364
rect 2668 64240 2708 64280
rect 4928 64240 4968 64280
rect 5010 64240 5050 64280
rect 5092 64240 5132 64280
rect 5174 64240 5214 64280
rect 5256 64240 5296 64280
rect 13420 64240 13460 64280
rect 15436 64240 15476 64280
rect 20048 64240 20088 64280
rect 20130 64240 20170 64280
rect 20212 64240 20252 64280
rect 20294 64240 20334 64280
rect 20376 64240 20416 64280
rect 11116 64156 11156 64196
rect 4108 64072 4148 64112
rect 5548 64072 5588 64112
rect 6028 64072 6068 64112
rect 6892 64072 6932 64112
rect 7564 64072 7604 64112
rect 8332 64072 8372 64112
rect 10636 64072 10676 64112
rect 12364 64156 12404 64196
rect 10156 63988 10196 64028
rect 13036 63988 13076 64028
rect 1420 63904 1460 63944
rect 9100 63904 9140 63944
rect 10924 63904 10964 63944
rect 8044 63652 8084 63692
rect 16972 63652 17012 63692
rect 3688 63484 3728 63524
rect 3770 63484 3810 63524
rect 3852 63484 3892 63524
rect 3934 63484 3974 63524
rect 4016 63484 4056 63524
rect 7468 63484 7508 63524
rect 1996 63400 2036 63440
rect 7564 63400 7604 63440
rect 11116 63484 11156 63524
rect 18808 63484 18848 63524
rect 18890 63484 18930 63524
rect 18972 63484 19012 63524
rect 19054 63484 19094 63524
rect 19136 63484 19176 63524
rect 12652 63400 12692 63440
rect 19852 63400 19892 63440
rect 3148 63316 3188 63356
rect 8332 63316 8372 63356
rect 10060 63232 10100 63272
rect 1708 62980 1748 63020
rect 2860 63064 2900 63104
rect 3148 63064 3188 63104
rect 21292 63064 21332 63104
rect 2956 62980 2996 63020
rect 4492 62980 4532 63020
rect 7852 62980 7892 63020
rect 9964 62980 10004 63020
rect 11308 62980 11348 63020
rect 19564 62980 19604 63020
rect 1612 62896 1652 62936
rect 5932 62896 5972 62936
rect 10924 62896 10964 62936
rect 2380 62812 2420 62852
rect 6124 62812 6164 62852
rect 7564 62812 7604 62852
rect 2668 62728 2708 62768
rect 4928 62728 4968 62768
rect 5010 62728 5050 62768
rect 5092 62728 5132 62768
rect 5174 62728 5214 62768
rect 5256 62728 5296 62768
rect 9196 62728 9236 62768
rect 20048 62728 20088 62768
rect 20130 62728 20170 62768
rect 20212 62728 20252 62768
rect 20294 62728 20334 62768
rect 20376 62728 20416 62768
rect 4780 62644 4820 62684
rect 9676 62644 9716 62684
rect 13516 62560 13556 62600
rect 8332 62476 8372 62516
rect 1516 62392 1556 62432
rect 10636 62392 10676 62432
rect 7948 62224 7988 62264
rect 10156 62224 10196 62264
rect 3148 62140 3188 62180
rect 11692 62140 11732 62180
rect 12172 62140 12212 62180
rect 9772 62056 9812 62096
rect 17548 62056 17588 62096
rect 3688 61972 3728 62012
rect 3770 61972 3810 62012
rect 3852 61972 3892 62012
rect 3934 61972 3974 62012
rect 4016 61972 4056 62012
rect 18808 61972 18848 62012
rect 18890 61972 18930 62012
rect 18972 61972 19012 62012
rect 19054 61972 19094 62012
rect 19136 61972 19176 62012
rect 2668 61888 2708 61928
rect 6412 61804 6452 61844
rect 7948 61804 7988 61844
rect 15532 61804 15572 61844
rect 3916 61720 3956 61760
rect 7756 61720 7796 61760
rect 15916 61636 15956 61676
rect 13036 61300 13076 61340
rect 16012 61300 16052 61340
rect 2188 61216 2228 61256
rect 4928 61216 4968 61256
rect 5010 61216 5050 61256
rect 5092 61216 5132 61256
rect 5174 61216 5214 61256
rect 5256 61216 5296 61256
rect 20048 61216 20088 61256
rect 20130 61216 20170 61256
rect 20212 61216 20252 61256
rect 20294 61216 20334 61256
rect 20376 61216 20416 61256
rect 3340 61132 3380 61172
rect 15532 61132 15572 61172
rect 4780 61048 4820 61088
rect 4588 60964 4628 61004
rect 5740 60880 5780 60920
rect 10828 61048 10868 61088
rect 11116 61048 11156 61088
rect 12268 61048 12308 61088
rect 13036 61048 13076 61088
rect 13420 60796 13460 60836
rect 15532 60628 15572 60668
rect 3688 60460 3728 60500
rect 3770 60460 3810 60500
rect 3852 60460 3892 60500
rect 3934 60460 3974 60500
rect 4016 60460 4056 60500
rect 6316 60460 6356 60500
rect 8620 60460 8660 60500
rect 18808 60460 18848 60500
rect 18890 60460 18930 60500
rect 18972 60460 19012 60500
rect 19054 60460 19094 60500
rect 19136 60460 19176 60500
rect 11692 60376 11732 60416
rect 21004 60376 21044 60416
rect 2764 60292 2804 60332
rect 4684 60292 4724 60332
rect 5548 60292 5588 60332
rect 13228 60292 13268 60332
rect 7468 60208 7508 60248
rect 8236 60124 8276 60164
rect 12268 60124 12308 60164
rect 12364 60040 12404 60080
rect 9580 59788 9620 59828
rect 4928 59704 4968 59744
rect 5010 59704 5050 59744
rect 5092 59704 5132 59744
rect 5174 59704 5214 59744
rect 5256 59704 5296 59744
rect 20048 59704 20088 59744
rect 20130 59704 20170 59744
rect 20212 59704 20252 59744
rect 20294 59704 20334 59744
rect 20376 59704 20416 59744
rect 16588 59452 16628 59492
rect 9484 59368 9524 59408
rect 12652 59368 12692 59408
rect 13420 59368 13460 59408
rect 15628 59368 15668 59408
rect 5644 59284 5684 59324
rect 2668 59200 2708 59240
rect 6412 59200 6452 59240
rect 17548 59116 17588 59156
rect 3688 58948 3728 58988
rect 3770 58948 3810 58988
rect 3852 58948 3892 58988
rect 3934 58948 3974 58988
rect 4016 58948 4056 58988
rect 6412 58948 6452 58988
rect 18808 58948 18848 58988
rect 18890 58948 18930 58988
rect 18972 58948 19012 58988
rect 19054 58948 19094 58988
rect 19136 58948 19176 58988
rect 13420 58780 13460 58820
rect 4780 58696 4820 58736
rect 15340 58696 15380 58736
rect 11308 58444 11348 58484
rect 12268 58444 12308 58484
rect 4928 58192 4968 58232
rect 5010 58192 5050 58232
rect 5092 58192 5132 58232
rect 5174 58192 5214 58232
rect 5256 58192 5296 58232
rect 20048 58192 20088 58232
rect 20130 58192 20170 58232
rect 20212 58192 20252 58232
rect 20294 58192 20334 58232
rect 20376 58192 20416 58232
rect 9580 57940 9620 57980
rect 3148 57856 3188 57896
rect 6316 57856 6356 57896
rect 8524 57856 8564 57896
rect 9196 57772 9236 57812
rect 17260 57688 17300 57728
rect 6412 57604 6452 57644
rect 13036 57604 13076 57644
rect 3688 57436 3728 57476
rect 3770 57436 3810 57476
rect 3852 57436 3892 57476
rect 3934 57436 3974 57476
rect 4016 57436 4056 57476
rect 18808 57436 18848 57476
rect 18890 57436 18930 57476
rect 18972 57436 19012 57476
rect 19054 57436 19094 57476
rect 19136 57436 19176 57476
rect 15340 57352 15380 57392
rect 12940 57268 12980 57308
rect 16396 57268 16436 57308
rect 6220 57016 6260 57056
rect 13708 57016 13748 57056
rect 13420 56764 13460 56804
rect 18700 56764 18740 56804
rect 4928 56680 4968 56720
rect 5010 56680 5050 56720
rect 5092 56680 5132 56720
rect 5174 56680 5214 56720
rect 5256 56680 5296 56720
rect 20048 56680 20088 56720
rect 20130 56680 20170 56720
rect 20212 56680 20252 56720
rect 20294 56680 20334 56720
rect 20376 56680 20416 56720
rect 9484 56512 9524 56552
rect 16876 56512 16916 56552
rect 16012 56428 16052 56468
rect 2764 56344 2804 56384
rect 17548 56344 17588 56384
rect 3244 56260 3284 56300
rect 10828 56260 10868 56300
rect 10060 56176 10100 56216
rect 3688 55924 3728 55964
rect 3770 55924 3810 55964
rect 3852 55924 3892 55964
rect 3934 55924 3974 55964
rect 4016 55924 4056 55964
rect 18808 55924 18848 55964
rect 18890 55924 18930 55964
rect 18972 55924 19012 55964
rect 19054 55924 19094 55964
rect 19136 55924 19176 55964
rect 11308 55756 11348 55796
rect 3340 55588 3380 55628
rect 10156 55504 10196 55544
rect 2764 55336 2804 55376
rect 4928 55168 4968 55208
rect 5010 55168 5050 55208
rect 5092 55168 5132 55208
rect 5174 55168 5214 55208
rect 5256 55168 5296 55208
rect 20048 55168 20088 55208
rect 20130 55168 20170 55208
rect 20212 55168 20252 55208
rect 20294 55168 20334 55208
rect 20376 55168 20416 55208
rect 16588 55000 16628 55040
rect 2956 54916 2996 54956
rect 10828 54916 10868 54956
rect 4108 54832 4148 54872
rect 9196 54832 9236 54872
rect 14284 54832 14324 54872
rect 3436 54748 3476 54788
rect 3688 54412 3728 54452
rect 3770 54412 3810 54452
rect 3852 54412 3892 54452
rect 3934 54412 3974 54452
rect 4016 54412 4056 54452
rect 18808 54412 18848 54452
rect 18890 54412 18930 54452
rect 18972 54412 19012 54452
rect 19054 54412 19094 54452
rect 19136 54412 19176 54452
rect 10156 53992 10196 54032
rect 2284 53908 2324 53948
rect 4928 53656 4968 53696
rect 5010 53656 5050 53696
rect 5092 53656 5132 53696
rect 5174 53656 5214 53696
rect 5256 53656 5296 53696
rect 15916 53656 15956 53696
rect 20048 53656 20088 53696
rect 20130 53656 20170 53696
rect 20212 53656 20252 53696
rect 20294 53656 20334 53696
rect 20376 53656 20416 53696
rect 6316 53572 6356 53612
rect 8812 53404 8852 53444
rect 1516 53320 1556 53360
rect 14284 53152 14324 53192
rect 6316 52984 6356 53024
rect 3244 52900 3284 52940
rect 3688 52900 3728 52940
rect 3770 52900 3810 52940
rect 3852 52900 3892 52940
rect 3934 52900 3974 52940
rect 4016 52900 4056 52940
rect 5644 52900 5684 52940
rect 18808 52900 18848 52940
rect 18890 52900 18930 52940
rect 18972 52900 19012 52940
rect 19054 52900 19094 52940
rect 19136 52900 19176 52940
rect 17548 52816 17588 52856
rect 18316 52816 18356 52856
rect 20620 52816 20660 52856
rect 2572 52732 2612 52772
rect 3436 52732 3476 52772
rect 3340 52480 3380 52520
rect 6412 52396 6452 52436
rect 4928 52144 4968 52184
rect 5010 52144 5050 52184
rect 5092 52144 5132 52184
rect 5174 52144 5214 52184
rect 5256 52144 5296 52184
rect 20048 52144 20088 52184
rect 20130 52144 20170 52184
rect 20212 52144 20252 52184
rect 20294 52144 20334 52184
rect 20376 52144 20416 52184
rect 2572 51892 2612 51932
rect 2764 51724 2804 51764
rect 8140 51724 8180 51764
rect 6508 51640 6548 51680
rect 6604 51472 6644 51512
rect 3688 51388 3728 51428
rect 3770 51388 3810 51428
rect 3852 51388 3892 51428
rect 3934 51388 3974 51428
rect 4016 51388 4056 51428
rect 18808 51388 18848 51428
rect 18890 51388 18930 51428
rect 18972 51388 19012 51428
rect 19054 51388 19094 51428
rect 19136 51388 19176 51428
rect 12652 51220 12692 51260
rect 13516 51220 13556 51260
rect 1516 50884 1556 50924
rect 4928 50632 4968 50672
rect 5010 50632 5050 50672
rect 5092 50632 5132 50672
rect 5174 50632 5214 50672
rect 5256 50632 5296 50672
rect 20048 50632 20088 50672
rect 20130 50632 20170 50672
rect 20212 50632 20252 50672
rect 20294 50632 20334 50672
rect 20376 50632 20416 50672
rect 2572 50548 2612 50588
rect 1516 50380 1556 50420
rect 18316 50464 18356 50504
rect 2572 50380 2612 50420
rect 13132 50380 13172 50420
rect 17932 50380 17972 50420
rect 6604 50044 6644 50084
rect 5644 49960 5684 50000
rect 3688 49876 3728 49916
rect 3770 49876 3810 49916
rect 3852 49876 3892 49916
rect 3934 49876 3974 49916
rect 4016 49876 4056 49916
rect 18808 49876 18848 49916
rect 18890 49876 18930 49916
rect 18972 49876 19012 49916
rect 19054 49876 19094 49916
rect 19136 49876 19176 49916
rect 17548 49708 17588 49748
rect 13708 49540 13748 49580
rect 4928 49120 4968 49160
rect 5010 49120 5050 49160
rect 5092 49120 5132 49160
rect 5174 49120 5214 49160
rect 5256 49120 5296 49160
rect 20048 49120 20088 49160
rect 20130 49120 20170 49160
rect 20212 49120 20252 49160
rect 20294 49120 20334 49160
rect 20376 49120 20416 49160
rect 6220 48784 6260 48824
rect 8908 48784 8948 48824
rect 9388 48784 9428 48824
rect 13132 48784 13172 48824
rect 13708 48616 13748 48656
rect 6220 48448 6260 48488
rect 3688 48364 3728 48404
rect 3770 48364 3810 48404
rect 3852 48364 3892 48404
rect 3934 48364 3974 48404
rect 4016 48364 4056 48404
rect 6124 48364 6164 48404
rect 18808 48364 18848 48404
rect 18890 48364 18930 48404
rect 18972 48364 19012 48404
rect 19054 48364 19094 48404
rect 19136 48364 19176 48404
rect 5932 47944 5972 47984
rect 6124 47944 6164 47984
rect 2764 47860 2804 47900
rect 4928 47608 4968 47648
rect 5010 47608 5050 47648
rect 5092 47608 5132 47648
rect 5174 47608 5214 47648
rect 5256 47608 5296 47648
rect 6124 47608 6164 47648
rect 20048 47608 20088 47648
rect 20130 47608 20170 47648
rect 20212 47608 20252 47648
rect 20294 47608 20334 47648
rect 20376 47608 20416 47648
rect 4108 47356 4148 47396
rect 13036 47356 13076 47396
rect 17068 47188 17108 47228
rect 3688 46852 3728 46892
rect 3770 46852 3810 46892
rect 3852 46852 3892 46892
rect 3934 46852 3974 46892
rect 4016 46852 4056 46892
rect 13516 46852 13556 46892
rect 18808 46852 18848 46892
rect 18890 46852 18930 46892
rect 18972 46852 19012 46892
rect 19054 46852 19094 46892
rect 19136 46852 19176 46892
rect 18316 46684 18356 46724
rect 5932 46600 5972 46640
rect 13036 46432 13076 46472
rect 18316 46432 18356 46472
rect 2284 46264 2324 46304
rect 4928 46096 4968 46136
rect 5010 46096 5050 46136
rect 5092 46096 5132 46136
rect 5174 46096 5214 46136
rect 5256 46096 5296 46136
rect 20048 46096 20088 46136
rect 20130 46096 20170 46136
rect 20212 46096 20252 46136
rect 20294 46096 20334 46136
rect 20376 46096 20416 46136
rect 10060 45676 10100 45716
rect 3340 45592 3380 45632
rect 16396 45508 16436 45548
rect 2284 45340 2324 45380
rect 3688 45340 3728 45380
rect 3770 45340 3810 45380
rect 3852 45340 3892 45380
rect 3934 45340 3974 45380
rect 4016 45340 4056 45380
rect 18808 45340 18848 45380
rect 18890 45340 18930 45380
rect 18972 45340 19012 45380
rect 19054 45340 19094 45380
rect 19136 45340 19176 45380
rect 2860 44920 2900 44960
rect 4928 44584 4968 44624
rect 5010 44584 5050 44624
rect 5092 44584 5132 44624
rect 5174 44584 5214 44624
rect 5256 44584 5296 44624
rect 20048 44584 20088 44624
rect 20130 44584 20170 44624
rect 20212 44584 20252 44624
rect 20294 44584 20334 44624
rect 20376 44584 20416 44624
rect 16396 44500 16436 44540
rect 16204 44332 16244 44372
rect 6220 44248 6260 44288
rect 17068 44248 17108 44288
rect 6220 44080 6260 44120
rect 9388 43996 9428 44036
rect 8908 43912 8948 43952
rect 3688 43828 3728 43868
rect 3770 43828 3810 43868
rect 3852 43828 3892 43868
rect 3934 43828 3974 43868
rect 4016 43828 4056 43868
rect 18808 43828 18848 43868
rect 18890 43828 18930 43868
rect 18972 43828 19012 43868
rect 19054 43828 19094 43868
rect 19136 43828 19176 43868
rect 21196 43660 21236 43700
rect 9388 43324 9428 43364
rect 12172 43324 12212 43364
rect 8908 43240 8948 43280
rect 9868 43240 9908 43280
rect 4928 43072 4968 43112
rect 5010 43072 5050 43112
rect 5092 43072 5132 43112
rect 5174 43072 5214 43112
rect 5256 43072 5296 43112
rect 20048 43072 20088 43112
rect 20130 43072 20170 43112
rect 20212 43072 20252 43112
rect 20294 43072 20334 43112
rect 20376 43072 20416 43112
rect 4396 42736 4436 42776
rect 6028 42736 6068 42776
rect 15724 42820 15764 42860
rect 16396 42820 16436 42860
rect 17644 42820 17684 42860
rect 21388 42568 21428 42608
rect 10252 42484 10292 42524
rect 18796 42484 18836 42524
rect 3688 42316 3728 42356
rect 3770 42316 3810 42356
rect 3852 42316 3892 42356
rect 3934 42316 3974 42356
rect 4016 42316 4056 42356
rect 18808 42316 18848 42356
rect 18890 42316 18930 42356
rect 18972 42316 19012 42356
rect 19054 42316 19094 42356
rect 19136 42316 19176 42356
rect 14956 42148 14996 42188
rect 18700 42148 18740 42188
rect 13804 42064 13844 42104
rect 2956 41812 2996 41852
rect 8620 41812 8660 41852
rect 19660 41728 19700 41768
rect 7564 41644 7604 41684
rect 11308 41644 11348 41684
rect 4396 41560 4436 41600
rect 4928 41560 4968 41600
rect 5010 41560 5050 41600
rect 5092 41560 5132 41600
rect 5174 41560 5214 41600
rect 5256 41560 5296 41600
rect 10732 41560 10772 41600
rect 11596 41560 11636 41600
rect 20048 41560 20088 41600
rect 20130 41560 20170 41600
rect 20212 41560 20252 41600
rect 20294 41560 20334 41600
rect 20376 41560 20416 41600
rect 11884 41476 11924 41516
rect 13228 41392 13268 41432
rect 19852 41392 19892 41432
rect 5452 41224 5492 41264
rect 6796 41224 6836 41264
rect 11500 41224 11540 41264
rect 5740 41140 5780 41180
rect 10924 41140 10964 41180
rect 19756 41056 19796 41096
rect 19468 40972 19508 41012
rect 4492 40888 4532 40928
rect 5932 40888 5972 40928
rect 8140 40888 8180 40928
rect 3688 40804 3728 40844
rect 3770 40804 3810 40844
rect 3852 40804 3892 40844
rect 3934 40804 3974 40844
rect 4016 40804 4056 40844
rect 18808 40804 18848 40844
rect 18890 40804 18930 40844
rect 18972 40804 19012 40844
rect 19054 40804 19094 40844
rect 19136 40804 19176 40844
rect 2284 40636 2324 40676
rect 17164 40636 17204 40676
rect 19468 40636 19508 40676
rect 9580 40468 9620 40508
rect 4780 40384 4820 40424
rect 8428 40384 8468 40424
rect 9868 40384 9908 40424
rect 10444 40384 10484 40424
rect 16876 40216 16916 40256
rect 4928 40048 4968 40088
rect 5010 40048 5050 40088
rect 5092 40048 5132 40088
rect 5174 40048 5214 40088
rect 5256 40048 5296 40088
rect 20048 40048 20088 40088
rect 20130 40048 20170 40088
rect 20212 40048 20252 40088
rect 20294 40048 20334 40088
rect 20376 40048 20416 40088
rect 16588 39964 16628 40004
rect 21004 39964 21044 40004
rect 652 39628 692 39668
rect 9292 39544 9332 39584
rect 13612 39544 13652 39584
rect 172 39376 212 39416
rect 364 39292 404 39332
rect 652 39292 692 39332
rect 3688 39292 3728 39332
rect 3770 39292 3810 39332
rect 3852 39292 3892 39332
rect 3934 39292 3974 39332
rect 4016 39292 4056 39332
rect 18808 39292 18848 39332
rect 18890 39292 18930 39332
rect 18972 39292 19012 39332
rect 19054 39292 19094 39332
rect 19136 39292 19176 39332
rect 3340 39208 3380 39248
rect 18412 39040 18452 39080
rect 20716 39040 20756 39080
rect 3244 38872 3284 38912
rect 11692 38872 11732 38912
rect 13420 38872 13460 38912
rect 4780 38788 4820 38828
rect 2476 38704 2516 38744
rect 10444 38704 10484 38744
rect 7084 38620 7124 38660
rect 14092 38620 14132 38660
rect 4928 38536 4968 38576
rect 5010 38536 5050 38576
rect 5092 38536 5132 38576
rect 5174 38536 5214 38576
rect 5256 38536 5296 38576
rect 20048 38536 20088 38576
rect 20130 38536 20170 38576
rect 20212 38536 20252 38576
rect 20294 38536 20334 38576
rect 20376 38536 20416 38576
rect 1420 38368 1460 38408
rect 7084 38452 7124 38492
rect 5836 38116 5876 38156
rect 8716 38032 8756 38072
rect 3688 37780 3728 37820
rect 3770 37780 3810 37820
rect 3852 37780 3892 37820
rect 3934 37780 3974 37820
rect 4016 37780 4056 37820
rect 11596 37780 11636 37820
rect 18808 37780 18848 37820
rect 18890 37780 18930 37820
rect 18972 37780 19012 37820
rect 19054 37780 19094 37820
rect 19136 37780 19176 37820
rect 13612 37696 13652 37736
rect 11116 37612 11156 37652
rect 16108 37612 16148 37652
rect 12076 37444 12116 37484
rect 19564 37444 19604 37484
rect 3052 37360 3092 37400
rect 1324 37276 1364 37316
rect 844 37192 884 37232
rect 8044 37192 8084 37232
rect 11116 37192 11156 37232
rect 11596 37192 11636 37232
rect 7468 37108 7508 37148
rect 4928 37024 4968 37064
rect 5010 37024 5050 37064
rect 5092 37024 5132 37064
rect 5174 37024 5214 37064
rect 5256 37024 5296 37064
rect 20048 37024 20088 37064
rect 20130 37024 20170 37064
rect 20212 37024 20252 37064
rect 20294 37024 20334 37064
rect 20376 37024 20416 37064
rect 5356 36772 5396 36812
rect 6892 36940 6932 36980
rect 8428 36856 8468 36896
rect 13228 36856 13268 36896
rect 10252 36772 10292 36812
rect 17452 36772 17492 36812
rect 6892 36688 6932 36728
rect 12940 36688 12980 36728
rect 11692 36604 11732 36644
rect 11980 36604 12020 36644
rect 18604 36520 18644 36560
rect 20524 36520 20564 36560
rect 13612 36436 13652 36476
rect 1612 36352 1652 36392
rect 7852 36352 7892 36392
rect 10444 36352 10484 36392
rect 3688 36268 3728 36308
rect 3770 36268 3810 36308
rect 3852 36268 3892 36308
rect 3934 36268 3974 36308
rect 4016 36268 4056 36308
rect 18808 36268 18848 36308
rect 18890 36268 18930 36308
rect 18972 36268 19012 36308
rect 19054 36268 19094 36308
rect 19136 36268 19176 36308
rect 2092 36100 2132 36140
rect 10828 36100 10868 36140
rect 3244 35848 3284 35888
rect 1324 35680 1364 35720
rect 13516 35680 13556 35720
rect 3148 35596 3188 35636
rect 11500 35596 11540 35636
rect 12268 35596 12308 35636
rect 4928 35512 4968 35552
rect 5010 35512 5050 35552
rect 5092 35512 5132 35552
rect 5174 35512 5214 35552
rect 5256 35512 5296 35552
rect 18028 35512 18068 35552
rect 20048 35512 20088 35552
rect 20130 35512 20170 35552
rect 20212 35512 20252 35552
rect 20294 35512 20334 35552
rect 20376 35512 20416 35552
rect 10828 35428 10868 35468
rect 1324 35344 1364 35384
rect 5836 35260 5876 35300
rect 7660 35260 7700 35300
rect 5548 35092 5588 35132
rect 6796 35092 6836 35132
rect 13420 35260 13460 35300
rect 11788 35176 11828 35216
rect 13804 35092 13844 35132
rect 3820 35008 3860 35048
rect 11116 35008 11156 35048
rect 21292 35008 21332 35048
rect 9580 34840 9620 34880
rect 3688 34756 3728 34796
rect 3770 34756 3810 34796
rect 3852 34756 3892 34796
rect 3934 34756 3974 34796
rect 4016 34756 4056 34796
rect 8428 34756 8468 34796
rect 18808 34756 18848 34796
rect 18890 34756 18930 34796
rect 18972 34756 19012 34796
rect 19054 34756 19094 34796
rect 19136 34756 19176 34796
rect 9580 34672 9620 34712
rect 10252 34588 10292 34628
rect 13132 34588 13172 34628
rect 13804 34588 13844 34628
rect 17260 34588 17300 34628
rect 2188 34336 2228 34376
rect 6028 34336 6068 34376
rect 8332 34336 8372 34376
rect 9100 34336 9140 34376
rect 3916 34252 3956 34292
rect 4396 34168 4436 34208
rect 12652 34168 12692 34208
rect 4928 34000 4968 34040
rect 5010 34000 5050 34040
rect 5092 34000 5132 34040
rect 5174 34000 5214 34040
rect 5256 34000 5296 34040
rect 13612 34000 13652 34040
rect 19372 34000 19412 34040
rect 20048 34000 20088 34040
rect 20130 34000 20170 34040
rect 20212 34000 20252 34040
rect 20294 34000 20334 34040
rect 20376 34000 20416 34040
rect 7756 33916 7796 33956
rect 4396 33580 4436 33620
rect 10540 33580 10580 33620
rect 3688 33244 3728 33284
rect 3770 33244 3810 33284
rect 3852 33244 3892 33284
rect 3934 33244 3974 33284
rect 4016 33244 4056 33284
rect 8236 33244 8276 33284
rect 12076 33244 12116 33284
rect 18808 33244 18848 33284
rect 18890 33244 18930 33284
rect 18972 33244 19012 33284
rect 19054 33244 19094 33284
rect 19136 33244 19176 33284
rect 1420 33160 1460 33200
rect 7564 33160 7604 33200
rect 19372 32824 19412 32864
rect 19948 32824 19988 32864
rect 3244 32740 3284 32780
rect 5356 32740 5396 32780
rect 7660 32656 7700 32696
rect 13228 32656 13268 32696
rect 4928 32488 4968 32528
rect 5010 32488 5050 32528
rect 5092 32488 5132 32528
rect 5174 32488 5214 32528
rect 5256 32488 5296 32528
rect 7756 32488 7796 32528
rect 20048 32488 20088 32528
rect 20130 32488 20170 32528
rect 20212 32488 20252 32528
rect 20294 32488 20334 32528
rect 20376 32488 20416 32528
rect 15724 32320 15764 32360
rect 6028 32236 6068 32276
rect 7468 32152 7508 32192
rect 16972 32152 17012 32192
rect 6796 32068 6836 32108
rect 7660 31984 7700 32024
rect 4108 31900 4148 31940
rect 2476 31816 2516 31856
rect 3688 31732 3728 31772
rect 3770 31732 3810 31772
rect 3852 31732 3892 31772
rect 3934 31732 3974 31772
rect 4016 31732 4056 31772
rect 18808 31732 18848 31772
rect 18890 31732 18930 31772
rect 18972 31732 19012 31772
rect 19054 31732 19094 31772
rect 19136 31732 19176 31772
rect 10348 31648 10388 31688
rect 9004 31564 9044 31604
rect 11596 31564 11636 31604
rect 2188 31480 2228 31520
rect 15340 31480 15380 31520
rect 14380 31396 14420 31436
rect 16684 31396 16724 31436
rect 11404 31312 11444 31352
rect 12268 31312 12308 31352
rect 9964 31228 10004 31268
rect 15436 31228 15476 31268
rect 19948 31144 19988 31184
rect 9484 31060 9524 31100
rect 4928 30976 4968 31016
rect 5010 30976 5050 31016
rect 5092 30976 5132 31016
rect 5174 30976 5214 31016
rect 5256 30976 5296 31016
rect 8812 30976 8852 31016
rect 11116 30976 11156 31016
rect 18700 30976 18740 31016
rect 20048 30976 20088 31016
rect 20130 30976 20170 31016
rect 20212 30976 20252 31016
rect 20294 30976 20334 31016
rect 20376 30976 20416 31016
rect 2188 30808 2228 30848
rect 6988 30808 7028 30848
rect 5836 30724 5876 30764
rect 11788 30724 11828 30764
rect 12364 30640 12404 30680
rect 15724 30388 15764 30428
rect 3148 30304 3188 30344
rect 8812 30304 8852 30344
rect 9484 30304 9524 30344
rect 3688 30220 3728 30260
rect 3770 30220 3810 30260
rect 3852 30220 3892 30260
rect 3934 30220 3974 30260
rect 4016 30220 4056 30260
rect 18808 30220 18848 30260
rect 18890 30220 18930 30260
rect 18972 30220 19012 30260
rect 19054 30220 19094 30260
rect 19136 30220 19176 30260
rect 19948 30220 19988 30260
rect 2188 30136 2228 30176
rect 1612 30052 1652 30092
rect 1996 30052 2036 30092
rect 9772 30052 9812 30092
rect 15340 30052 15380 30092
rect 4108 29800 4148 29840
rect 11308 29716 11348 29756
rect 8236 29632 8276 29672
rect 10252 29632 10292 29672
rect 13132 29632 13172 29672
rect 4928 29464 4968 29504
rect 5010 29464 5050 29504
rect 5092 29464 5132 29504
rect 5174 29464 5214 29504
rect 5256 29464 5296 29504
rect 20048 29464 20088 29504
rect 20130 29464 20170 29504
rect 20212 29464 20252 29504
rect 20294 29464 20334 29504
rect 20376 29464 20416 29504
rect 20812 29464 20852 29504
rect 15244 29296 15284 29336
rect 17068 29296 17108 29336
rect 10732 29212 10772 29252
rect 4204 29128 4244 29168
rect 5548 29128 5588 29168
rect 6892 29128 6932 29168
rect 1324 29044 1364 29084
rect 4780 29044 4820 29084
rect 1996 28960 2036 29000
rect 2956 28960 2996 29000
rect 17452 29044 17492 29084
rect 2764 28876 2804 28916
rect 10732 28876 10772 28916
rect 17068 28876 17108 28916
rect 7276 28792 7316 28832
rect 3688 28708 3728 28748
rect 3770 28708 3810 28748
rect 3852 28708 3892 28748
rect 3934 28708 3974 28748
rect 4016 28708 4056 28748
rect 18808 28708 18848 28748
rect 18890 28708 18930 28748
rect 18972 28708 19012 28748
rect 19054 28708 19094 28748
rect 19136 28708 19176 28748
rect 13324 28456 13364 28496
rect 19564 28456 19604 28496
rect 556 28372 596 28412
rect 19948 28288 19988 28328
rect 3148 28204 3188 28244
rect 10828 28204 10868 28244
rect 13516 28204 13556 28244
rect 4300 28120 4340 28160
rect 2284 27952 2324 27992
rect 4928 27952 4968 27992
rect 5010 27952 5050 27992
rect 5092 27952 5132 27992
rect 5174 27952 5214 27992
rect 5256 27952 5296 27992
rect 18700 27952 18740 27992
rect 20048 27952 20088 27992
rect 20130 27952 20170 27992
rect 20212 27952 20252 27992
rect 20294 27952 20334 27992
rect 20376 27952 20416 27992
rect 12460 27868 12500 27908
rect 6988 27784 7028 27824
rect 2284 27700 2324 27740
rect 11116 27700 11156 27740
rect 16012 27700 16052 27740
rect 7084 27532 7124 27572
rect 15820 27532 15860 27572
rect 4300 27448 4340 27488
rect 6988 27364 7028 27404
rect 3688 27196 3728 27236
rect 3770 27196 3810 27236
rect 3852 27196 3892 27236
rect 3934 27196 3974 27236
rect 4016 27196 4056 27236
rect 13804 27196 13844 27236
rect 18808 27196 18848 27236
rect 18890 27196 18930 27236
rect 18972 27196 19012 27236
rect 19054 27196 19094 27236
rect 19136 27196 19176 27236
rect 4204 27112 4244 27152
rect 3436 27028 3476 27068
rect 9484 27028 9524 27068
rect 2476 26944 2516 26984
rect 11596 26944 11636 26984
rect 12460 26944 12500 26984
rect 2188 26860 2228 26900
rect 2572 26776 2612 26816
rect 3532 26776 3572 26816
rect 6604 26776 6644 26816
rect 8812 26776 8852 26816
rect 9580 26776 9620 26816
rect 748 26692 788 26732
rect 4588 26608 4628 26648
rect 7084 26608 7124 26648
rect 12460 26776 12500 26816
rect 11596 26692 11636 26732
rect 12940 26608 12980 26648
rect 19948 26608 19988 26648
rect 19852 26524 19892 26564
rect 4396 26440 4436 26480
rect 4928 26440 4968 26480
rect 5010 26440 5050 26480
rect 5092 26440 5132 26480
rect 5174 26440 5214 26480
rect 5256 26440 5296 26480
rect 19564 26440 19604 26480
rect 20048 26440 20088 26480
rect 20130 26440 20170 26480
rect 20212 26440 20252 26480
rect 20294 26440 20334 26480
rect 20376 26440 20416 26480
rect 4684 26272 4724 26312
rect 7468 26272 7508 26312
rect 9676 26272 9716 26312
rect 11212 26272 11252 26312
rect 2476 26188 2516 26228
rect 3532 26104 3572 26144
rect 6124 26104 6164 26144
rect 7564 26104 7604 26144
rect 17644 26104 17684 26144
rect 14572 26020 14612 26060
rect 2860 25936 2900 25976
rect 3340 25936 3380 25976
rect 5932 25852 5972 25892
rect 8428 25852 8468 25892
rect 2668 25768 2708 25808
rect 3688 25684 3728 25724
rect 3770 25684 3810 25724
rect 3852 25684 3892 25724
rect 3934 25684 3974 25724
rect 4016 25684 4056 25724
rect 4780 25684 4820 25724
rect 18808 25684 18848 25724
rect 18890 25684 18930 25724
rect 18972 25684 19012 25724
rect 19054 25684 19094 25724
rect 19136 25684 19176 25724
rect 4972 25600 5012 25640
rect 11116 25432 11156 25472
rect 2668 25348 2708 25388
rect 3436 25348 3476 25388
rect 11308 25348 11348 25388
rect 4780 25180 4820 25220
rect 7084 25264 7124 25304
rect 9004 25264 9044 25304
rect 5068 25180 5108 25220
rect 6316 25180 6356 25220
rect 5260 25096 5300 25136
rect 12460 25096 12500 25136
rect 4396 25012 4436 25052
rect 844 24928 884 24968
rect 4928 24928 4968 24968
rect 5010 24928 5050 24968
rect 5092 24928 5132 24968
rect 5174 24928 5214 24968
rect 5256 24928 5296 24968
rect 20048 24928 20088 24968
rect 20130 24928 20170 24968
rect 20212 24928 20252 24968
rect 20294 24928 20334 24968
rect 20376 24928 20416 24968
rect 5740 24844 5780 24884
rect 4588 24760 4628 24800
rect 5644 24760 5684 24800
rect 8716 24760 8756 24800
rect 9196 24760 9236 24800
rect 9772 24760 9812 24800
rect 15148 24760 15188 24800
rect 2284 24676 2324 24716
rect 1324 24508 1364 24548
rect 3340 24508 3380 24548
rect 5548 24508 5588 24548
rect 7756 24508 7796 24548
rect 9676 24592 9716 24632
rect 10444 24592 10484 24632
rect 11212 24592 11252 24632
rect 15436 24592 15476 24632
rect 16972 24592 17012 24632
rect 8620 24508 8660 24548
rect 6124 24424 6164 24464
rect 6508 24340 6548 24380
rect 7468 24340 7508 24380
rect 9196 24340 9236 24380
rect 12364 24340 12404 24380
rect 6028 24256 6068 24296
rect 6796 24256 6836 24296
rect 3688 24172 3728 24212
rect 3770 24172 3810 24212
rect 3852 24172 3892 24212
rect 3934 24172 3974 24212
rect 4016 24172 4056 24212
rect 10444 24172 10484 24212
rect 11884 24172 11924 24212
rect 18808 24172 18848 24212
rect 18890 24172 18930 24212
rect 18972 24172 19012 24212
rect 19054 24172 19094 24212
rect 19136 24172 19176 24212
rect 12460 24088 12500 24128
rect 7756 23920 7796 23960
rect 12652 23920 12692 23960
rect 3436 23836 3476 23876
rect 7276 23836 7316 23876
rect 14092 23752 14132 23792
rect 12364 23584 12404 23624
rect 6508 23500 6548 23540
rect 8716 23500 8756 23540
rect 4928 23416 4968 23456
rect 5010 23416 5050 23456
rect 5092 23416 5132 23456
rect 5174 23416 5214 23456
rect 5256 23416 5296 23456
rect 20048 23416 20088 23456
rect 20130 23416 20170 23456
rect 20212 23416 20252 23456
rect 20294 23416 20334 23456
rect 20376 23416 20416 23456
rect 7276 23248 7316 23288
rect 7660 23248 7700 23288
rect 8716 23248 8756 23288
rect 4204 23164 4244 23204
rect 4204 22996 4244 23036
rect 15436 22996 15476 23036
rect 9964 22912 10004 22952
rect 15820 22828 15860 22868
rect 20140 22828 20180 22868
rect 2572 22744 2612 22784
rect 3688 22660 3728 22700
rect 3770 22660 3810 22700
rect 3852 22660 3892 22700
rect 3934 22660 3974 22700
rect 4016 22660 4056 22700
rect 18808 22660 18848 22700
rect 18890 22660 18930 22700
rect 18972 22660 19012 22700
rect 19054 22660 19094 22700
rect 19136 22660 19176 22700
rect 12460 22324 12500 22364
rect 3340 22240 3380 22280
rect 4492 22240 4532 22280
rect 13324 22240 13364 22280
rect 12172 21988 12212 22028
rect 4928 21904 4968 21944
rect 5010 21904 5050 21944
rect 5092 21904 5132 21944
rect 5174 21904 5214 21944
rect 5256 21904 5296 21944
rect 7756 21904 7796 21944
rect 20048 21904 20088 21944
rect 20130 21904 20170 21944
rect 20212 21904 20252 21944
rect 20294 21904 20334 21944
rect 20376 21904 20416 21944
rect 3436 21652 3476 21692
rect 1324 21568 1364 21608
rect 460 21484 500 21524
rect 8428 21652 8468 21692
rect 9196 21568 9236 21608
rect 19372 21568 19412 21608
rect 10156 21484 10196 21524
rect 6604 21316 6644 21356
rect 9772 21316 9812 21356
rect 2092 21232 2132 21272
rect 3688 21148 3728 21188
rect 3770 21148 3810 21188
rect 3852 21148 3892 21188
rect 3934 21148 3974 21188
rect 4016 21148 4056 21188
rect 18808 21148 18848 21188
rect 18890 21148 18930 21188
rect 18972 21148 19012 21188
rect 19054 21148 19094 21188
rect 19136 21148 19176 21188
rect 18412 21064 18452 21104
rect 12652 20980 12692 21020
rect 7852 20812 7892 20852
rect 3148 20728 3188 20768
rect 3436 20728 3476 20768
rect 4780 20728 4820 20768
rect 9484 20728 9524 20768
rect 12172 20728 12212 20768
rect 2764 20644 2804 20684
rect 4928 20392 4968 20432
rect 5010 20392 5050 20432
rect 5092 20392 5132 20432
rect 5174 20392 5214 20432
rect 5256 20392 5296 20432
rect 6508 20392 6548 20432
rect 18412 20392 18452 20432
rect 20048 20392 20088 20432
rect 20130 20392 20170 20432
rect 20212 20392 20252 20432
rect 20294 20392 20334 20432
rect 20376 20392 20416 20432
rect 3052 20224 3092 20264
rect 4780 20140 4820 20180
rect 3532 20056 3572 20096
rect 10156 20056 10196 20096
rect 18028 20056 18068 20096
rect 5644 19972 5684 20012
rect 8716 19972 8756 20012
rect 11884 19972 11924 20012
rect 12172 19972 12212 20012
rect 12556 19804 12596 19844
rect 6124 19720 6164 19760
rect 3688 19636 3728 19676
rect 3770 19636 3810 19676
rect 3852 19636 3892 19676
rect 3934 19636 3974 19676
rect 4016 19636 4056 19676
rect 8812 19636 8852 19676
rect 9196 19636 9236 19676
rect 18808 19636 18848 19676
rect 18890 19636 18930 19676
rect 18972 19636 19012 19676
rect 19054 19636 19094 19676
rect 19136 19636 19176 19676
rect 3148 19384 3188 19424
rect 10060 19384 10100 19424
rect 4204 19300 4244 19340
rect 6316 19300 6356 19340
rect 6508 19300 6548 19340
rect 4396 19216 4436 19256
rect 6988 19216 7028 19256
rect 10348 19048 10388 19088
rect 14764 19048 14804 19088
rect 5356 18964 5396 19004
rect 8812 18964 8852 19004
rect 3052 18880 3092 18920
rect 4928 18880 4968 18920
rect 5010 18880 5050 18920
rect 5092 18880 5132 18920
rect 5174 18880 5214 18920
rect 5256 18880 5296 18920
rect 5932 18880 5972 18920
rect 8044 18880 8084 18920
rect 20048 18880 20088 18920
rect 20130 18880 20170 18920
rect 20212 18880 20252 18920
rect 20294 18880 20334 18920
rect 20376 18880 20416 18920
rect 6796 18796 6836 18836
rect 11116 18796 11156 18836
rect 13804 18796 13844 18836
rect 15436 18796 15476 18836
rect 7852 18628 7892 18668
rect 4588 18544 4628 18584
rect 12172 18628 12212 18668
rect 17452 18628 17492 18668
rect 16972 18544 17012 18584
rect 10156 18208 10196 18248
rect 3688 18124 3728 18164
rect 3770 18124 3810 18164
rect 3852 18124 3892 18164
rect 3934 18124 3974 18164
rect 4016 18124 4056 18164
rect 16684 18124 16724 18164
rect 18808 18124 18848 18164
rect 18890 18124 18930 18164
rect 18972 18124 19012 18164
rect 19054 18124 19094 18164
rect 19136 18124 19176 18164
rect 7468 18040 7508 18080
rect 10060 18040 10100 18080
rect 3148 17788 3188 17828
rect 4492 17788 4532 17828
rect 10060 17788 10100 17828
rect 8716 17704 8756 17744
rect 3052 17620 3092 17660
rect 4396 17536 4436 17576
rect 4588 17536 4628 17576
rect 5740 17536 5780 17576
rect 2956 17452 2996 17492
rect 5356 17452 5396 17492
rect 3436 17368 3476 17408
rect 4928 17368 4968 17408
rect 5010 17368 5050 17408
rect 5092 17368 5132 17408
rect 5174 17368 5214 17408
rect 5256 17368 5296 17408
rect 16492 17368 16532 17408
rect 20048 17368 20088 17408
rect 20130 17368 20170 17408
rect 20212 17368 20252 17408
rect 20294 17368 20334 17408
rect 20376 17368 20416 17408
rect 8908 17284 8948 17324
rect 15436 17200 15476 17240
rect 3052 17032 3092 17072
rect 4108 17032 4148 17072
rect 5356 17032 5396 17072
rect 7660 17032 7700 17072
rect 7852 17032 7892 17072
rect 14764 17032 14804 17072
rect 6796 16948 6836 16988
rect 16684 16864 16724 16904
rect 6316 16780 6356 16820
rect 6604 16780 6644 16820
rect 5548 16696 5588 16736
rect 3688 16612 3728 16652
rect 3770 16612 3810 16652
rect 3852 16612 3892 16652
rect 3934 16612 3974 16652
rect 4016 16612 4056 16652
rect 8044 16612 8084 16652
rect 18808 16612 18848 16652
rect 18890 16612 18930 16652
rect 18972 16612 19012 16652
rect 19054 16612 19094 16652
rect 19136 16612 19176 16652
rect 2476 16360 2516 16400
rect 3340 16360 3380 16400
rect 12844 16192 12884 16232
rect 8908 16108 8948 16148
rect 10156 16024 10196 16064
rect 4928 15856 4968 15896
rect 5010 15856 5050 15896
rect 5092 15856 5132 15896
rect 5174 15856 5214 15896
rect 5256 15856 5296 15896
rect 20048 15856 20088 15896
rect 20130 15856 20170 15896
rect 20212 15856 20252 15896
rect 20294 15856 20334 15896
rect 20376 15856 20416 15896
rect 4300 15688 4340 15728
rect 15724 15520 15764 15560
rect 12844 15436 12884 15476
rect 3436 15268 3476 15308
rect 9196 15268 9236 15308
rect 3688 15100 3728 15140
rect 3770 15100 3810 15140
rect 3852 15100 3892 15140
rect 3934 15100 3974 15140
rect 4016 15100 4056 15140
rect 6508 15100 6548 15140
rect 18808 15100 18848 15140
rect 18890 15100 18930 15140
rect 18972 15100 19012 15140
rect 19054 15100 19094 15140
rect 19136 15100 19176 15140
rect 8044 15016 8084 15056
rect 3244 14932 3284 14972
rect 4204 14680 4244 14720
rect 13036 14596 13076 14636
rect 3340 14512 3380 14552
rect 9484 14428 9524 14468
rect 4928 14344 4968 14384
rect 5010 14344 5050 14384
rect 5092 14344 5132 14384
rect 5174 14344 5214 14384
rect 5256 14344 5296 14384
rect 20048 14344 20088 14384
rect 20130 14344 20170 14384
rect 20212 14344 20252 14384
rect 20294 14344 20334 14384
rect 20376 14344 20416 14384
rect 16492 14176 16532 14216
rect 4204 14092 4244 14132
rect 8908 14092 8948 14132
rect 9388 14008 9428 14048
rect 11212 13924 11252 13964
rect 7468 13840 7508 13880
rect 10348 13840 10388 13880
rect 13132 13840 13172 13880
rect 3688 13588 3728 13628
rect 3770 13588 3810 13628
rect 3852 13588 3892 13628
rect 3934 13588 3974 13628
rect 4016 13588 4056 13628
rect 18808 13588 18848 13628
rect 18890 13588 18930 13628
rect 18972 13588 19012 13628
rect 19054 13588 19094 13628
rect 19136 13588 19176 13628
rect 6220 13336 6260 13376
rect 5644 13252 5684 13292
rect 15820 13252 15860 13292
rect 4108 13168 4148 13208
rect 11020 13177 11060 13208
rect 11020 13168 11060 13177
rect 6796 13084 6836 13124
rect 6316 12916 6356 12956
rect 4928 12832 4968 12872
rect 5010 12832 5050 12872
rect 5092 12832 5132 12872
rect 5174 12832 5214 12872
rect 5256 12832 5296 12872
rect 20048 12832 20088 12872
rect 20130 12832 20170 12872
rect 20212 12832 20252 12872
rect 20294 12832 20334 12872
rect 20376 12832 20416 12872
rect 16204 12664 16244 12704
rect 11020 12580 11060 12620
rect 13132 12580 13172 12620
rect 15244 12580 15284 12620
rect 7180 12496 7220 12536
rect 7756 12496 7796 12536
rect 11020 12244 11060 12284
rect 11212 12244 11252 12284
rect 3688 12076 3728 12116
rect 3770 12076 3810 12116
rect 3852 12076 3892 12116
rect 3934 12076 3974 12116
rect 4016 12076 4056 12116
rect 18808 12076 18848 12116
rect 18890 12076 18930 12116
rect 18972 12076 19012 12116
rect 19054 12076 19094 12116
rect 19136 12076 19176 12116
rect 15820 11824 15860 11864
rect 16396 11740 16436 11780
rect 13132 11656 13172 11696
rect 4300 11488 4340 11528
rect 4928 11320 4968 11360
rect 5010 11320 5050 11360
rect 5092 11320 5132 11360
rect 5174 11320 5214 11360
rect 5256 11320 5296 11360
rect 20048 11320 20088 11360
rect 20130 11320 20170 11360
rect 20212 11320 20252 11360
rect 20294 11320 20334 11360
rect 20376 11320 20416 11360
rect 4108 11236 4148 11276
rect 6220 11236 6260 11276
rect 14380 11152 14420 11192
rect 4588 11068 4628 11108
rect 10156 10984 10196 11024
rect 2572 10564 2612 10604
rect 3688 10564 3728 10604
rect 3770 10564 3810 10604
rect 3852 10564 3892 10604
rect 3934 10564 3974 10604
rect 4016 10564 4056 10604
rect 18808 10564 18848 10604
rect 18890 10564 18930 10604
rect 18972 10564 19012 10604
rect 19054 10564 19094 10604
rect 19136 10564 19176 10604
rect 2860 9976 2900 10016
rect 14380 9892 14420 9932
rect 2956 9808 2996 9848
rect 4684 9808 4724 9848
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 7660 9724 7700 9764
rect 6796 9640 6836 9680
rect 8620 9640 8660 9680
rect 15724 9556 15764 9596
rect 7660 9220 7700 9260
rect 8620 9220 8660 9260
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 8908 9052 8948 9092
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 7852 8716 7892 8756
rect 13036 8632 13076 8672
rect 5356 8464 5396 8504
rect 2572 8380 2612 8420
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 11020 8296 11060 8336
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 7084 8128 7124 8168
rect 11020 8128 11060 8168
rect 5356 8044 5396 8084
rect 16108 7960 16148 8000
rect 10828 7876 10868 7916
rect 5548 7792 5588 7832
rect 6220 7624 6260 7664
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 13036 7540 13076 7580
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 11404 7456 11444 7496
rect 14764 7288 14804 7328
rect 4780 7204 4820 7244
rect 2380 7120 2420 7160
rect 11404 6952 11444 6992
rect 11212 6868 11252 6908
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 11596 6616 11636 6656
rect 4684 6448 4724 6488
rect 11020 6280 11060 6320
rect 11212 6280 11252 6320
rect 12172 6196 12212 6236
rect 2380 6112 2420 6152
rect 11596 6112 11636 6152
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 9100 5692 9140 5732
rect 2860 5608 2900 5648
rect 4780 5608 4820 5648
rect 8332 5608 8372 5648
rect 2380 5524 2420 5564
rect 16108 5440 16148 5480
rect 6988 5356 7028 5396
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 6988 5104 7028 5144
rect 2956 4936 2996 4976
rect 13036 4936 13076 4976
rect 4684 4768 4724 4808
rect 2956 4600 2996 4640
rect 3436 4600 3476 4640
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 13996 4516 14036 4556
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 14476 4432 14516 4472
rect 8908 4096 8948 4136
rect 3148 3928 3188 3968
rect 13324 3928 13364 3968
rect 2188 3844 2228 3884
rect 7660 3844 7700 3884
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 5740 3760 5780 3800
rect 10828 3760 10868 3800
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 11020 3424 11060 3464
rect 2380 3340 2420 3380
rect 7660 3340 7700 3380
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 11116 3004 11156 3044
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 5356 2668 5396 2708
rect 10540 2668 10580 2708
rect 11308 2668 11348 2708
rect 12076 2584 12116 2624
rect 5548 2416 5588 2456
rect 10252 2416 10292 2456
rect 364 2332 404 2372
rect 1132 2248 1172 2288
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 5740 2248 5780 2288
rect 10540 2248 10580 2288
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 6604 2164 6644 2204
rect 8140 2164 8180 2204
rect 5356 2080 5396 2120
rect 6700 2080 6740 2120
rect 16876 2080 16916 2120
rect 16588 1996 16628 2036
rect 172 1912 212 1952
rect 5548 1912 5588 1952
rect 2476 1828 2516 1868
rect 5836 1828 5876 1868
rect 12268 1828 12308 1868
rect 12940 1828 12980 1868
rect 14092 1828 14132 1868
rect 14284 1828 14324 1868
rect 15244 1828 15284 1868
rect 15532 1828 15572 1868
rect 16012 1828 16052 1868
rect 940 1492 980 1532
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 11500 1576 11540 1616
rect 14668 1576 14708 1616
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 2284 1324 2324 1364
rect 5452 1240 5492 1280
rect 6700 1240 6740 1280
rect 7372 1240 7412 1280
rect 7756 1240 7796 1280
rect 12748 1240 12788 1280
rect 13900 1240 13940 1280
rect 15628 1240 15668 1280
rect 17356 1240 17396 1280
rect 17740 1240 17780 1280
rect 18124 1240 18164 1280
rect 18508 1240 18548 1280
rect 19276 1240 19316 1280
rect 19468 1240 19508 1280
rect 8812 1156 8852 1196
rect 16780 1156 16820 1196
rect 19660 1156 19700 1196
rect 6892 1072 6932 1112
rect 12556 1072 12596 1112
rect 20716 1072 20756 1112
rect 6220 988 6260 1028
rect 20524 988 20564 1028
rect 1228 904 1268 944
rect 6316 904 6356 944
rect 7084 904 7124 944
rect 18316 904 18356 944
rect 15052 820 15092 860
rect 20620 820 20660 860
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 6412 736 6452 776
rect 6988 736 7028 776
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
rect 14188 652 14228 692
rect 17932 568 17972 608
rect 2092 484 2132 524
rect 9868 484 9908 524
rect 9292 400 9332 440
rect 3724 316 3764 356
rect 2956 232 2996 272
rect 5260 148 5300 188
rect 13708 148 13748 188
rect 11788 64 11828 104
<< metal4 >>
rect 15724 85616 15764 85625
rect 4780 85448 4820 85457
rect 1324 85112 1364 85121
rect 76 84776 116 84785
rect 76 67136 116 84736
rect 1228 84272 1268 84281
rect 844 79988 884 79997
rect 76 67087 116 67096
rect 364 76040 404 76049
rect 364 66884 404 76000
rect 364 66835 404 66844
rect 460 72512 500 72521
rect 172 39416 212 39425
rect 172 1952 212 39376
rect 364 39332 404 39341
rect 364 2372 404 39292
rect 460 21524 500 72472
rect 748 66800 788 66809
rect 556 65540 596 65549
rect 556 28412 596 65500
rect 651 63020 693 63029
rect 651 62980 652 63020
rect 692 62980 693 63020
rect 651 62971 693 62980
rect 652 39668 692 62971
rect 652 39332 692 39628
rect 652 39283 692 39292
rect 556 28363 596 28372
rect 748 26732 788 66760
rect 844 37232 884 79948
rect 1035 67472 1077 67481
rect 1035 67432 1036 67472
rect 1076 67432 1077 67472
rect 1035 67423 1077 67432
rect 940 64868 980 64877
rect 940 59240 980 64828
rect 1036 63356 1076 67423
rect 1132 66632 1172 66641
rect 1132 66389 1172 66592
rect 1131 66380 1173 66389
rect 1131 66340 1132 66380
rect 1172 66340 1173 66380
rect 1131 66331 1173 66340
rect 1036 63316 1172 63356
rect 940 59200 1076 59240
rect 844 37183 884 37192
rect 939 35048 981 35057
rect 939 35008 940 35048
rect 980 35008 981 35048
rect 939 34999 981 35008
rect 748 26683 788 26692
rect 843 25136 885 25145
rect 843 25096 844 25136
rect 884 25096 885 25136
rect 843 25087 885 25096
rect 844 24968 884 25087
rect 844 24919 884 24928
rect 460 21475 500 21484
rect 364 2323 404 2332
rect 172 1903 212 1912
rect 940 1532 980 34999
rect 940 1483 980 1492
rect 1036 953 1076 59200
rect 1132 2288 1172 63316
rect 1132 2239 1172 2248
rect 1035 944 1077 953
rect 1035 904 1036 944
rect 1076 904 1077 944
rect 1035 895 1077 904
rect 1228 944 1268 84232
rect 1324 69992 1364 85072
rect 3688 84692 4056 84701
rect 3728 84652 3770 84692
rect 3810 84652 3852 84692
rect 3892 84652 3934 84692
rect 3974 84652 4016 84692
rect 3688 84643 4056 84652
rect 3244 84356 3284 84365
rect 2956 83516 2996 83525
rect 2572 83348 2612 83357
rect 1900 83096 1940 83105
rect 1900 82676 1940 83056
rect 1612 81080 1652 81089
rect 1612 80576 1652 81040
rect 1516 80408 1556 80417
rect 1516 78896 1556 80368
rect 1324 64700 1364 69952
rect 1324 64651 1364 64660
rect 1420 70748 1460 70757
rect 1420 63944 1460 70708
rect 1420 63895 1460 63904
rect 1516 62432 1556 78856
rect 1612 67724 1652 80536
rect 1900 78980 1940 82636
rect 2476 82760 2516 82769
rect 1804 76040 1844 76049
rect 1612 67675 1652 67684
rect 1708 73016 1748 73025
rect 1708 68144 1748 72976
rect 1612 65372 1652 65381
rect 1612 62936 1652 65332
rect 1708 63020 1748 68104
rect 1804 65372 1844 76000
rect 1900 71504 1940 78940
rect 2284 80576 2324 80585
rect 2284 79736 2324 80536
rect 2476 80576 2516 82720
rect 2476 80527 2516 80536
rect 1900 71455 1940 71464
rect 1996 76712 2036 76721
rect 1804 65323 1844 65332
rect 1996 63440 2036 76672
rect 2284 73016 2324 79696
rect 2284 72967 2324 72976
rect 2476 73856 2516 73865
rect 2476 73016 2516 73816
rect 2476 71924 2516 72976
rect 2476 71875 2516 71884
rect 2092 71252 2132 71261
rect 2092 65456 2132 71212
rect 2092 65407 2132 65416
rect 2188 70664 2228 70673
rect 1996 63391 2036 63400
rect 1708 62971 1748 62980
rect 1612 62887 1652 62896
rect 1516 53360 1556 62392
rect 2188 61256 2228 70624
rect 2188 61207 2228 61216
rect 2380 62852 2420 62861
rect 1516 50924 1556 53320
rect 1516 50420 1556 50884
rect 1516 50371 1556 50380
rect 2284 53948 2324 53957
rect 2284 46304 2324 53908
rect 2284 45380 2324 46264
rect 2284 45331 2324 45340
rect 2284 40676 2324 40685
rect 1420 38408 1460 38417
rect 1324 37316 1364 37325
rect 1324 35720 1364 37276
rect 1324 35671 1364 35680
rect 1324 35384 1364 35393
rect 1324 29084 1364 35344
rect 1420 33200 1460 38368
rect 1420 33151 1460 33160
rect 1612 36392 1652 36401
rect 1612 30092 1652 36352
rect 2092 36140 2132 36149
rect 1612 30043 1652 30052
rect 1996 30092 2036 30101
rect 1324 29035 1364 29044
rect 1996 29000 2036 30052
rect 1996 28951 2036 28960
rect 1324 24548 1364 24557
rect 1324 21608 1364 24508
rect 1324 21559 1364 21568
rect 2092 21272 2132 36100
rect 2188 34376 2228 34385
rect 2188 31520 2228 34336
rect 2188 31471 2228 31480
rect 2188 30848 2228 30857
rect 2188 30176 2228 30808
rect 2188 30127 2228 30136
rect 2284 27992 2324 40636
rect 2284 27740 2324 27952
rect 2284 27691 2324 27700
rect 2092 21223 2132 21232
rect 2188 26900 2228 26909
rect 2091 10688 2133 10697
rect 2091 10648 2092 10688
rect 2132 10648 2133 10688
rect 2091 10639 2133 10648
rect 1228 895 1268 904
rect 2092 524 2132 10639
rect 2188 3884 2228 26860
rect 2284 24716 2324 24725
rect 2284 10697 2324 24676
rect 2283 10688 2325 10697
rect 2283 10648 2284 10688
rect 2324 10648 2325 10688
rect 2283 10639 2325 10648
rect 2380 7832 2420 62812
rect 2572 61769 2612 83308
rect 2764 80744 2804 80753
rect 2668 69740 2708 69749
rect 2668 64280 2708 69700
rect 2764 69236 2804 80704
rect 2956 77552 2996 83476
rect 2764 69187 2804 69196
rect 2860 70076 2900 70085
rect 2764 68984 2804 68993
rect 2764 66968 2804 68944
rect 2764 66919 2804 66928
rect 2860 66128 2900 70036
rect 2956 66800 2996 77512
rect 3148 79400 3188 79409
rect 3148 78224 3188 79360
rect 3148 75284 3188 78184
rect 3148 75235 3188 75244
rect 3148 73016 3188 73025
rect 2956 66751 2996 66760
rect 3052 72008 3092 72017
rect 2668 64231 2708 64240
rect 2764 66088 2900 66128
rect 2668 62768 2708 62777
rect 2668 61928 2708 62728
rect 2571 61760 2613 61769
rect 2571 61720 2572 61760
rect 2612 61720 2613 61760
rect 2571 61711 2613 61720
rect 2475 61004 2517 61013
rect 2475 60964 2476 61004
rect 2516 60964 2517 61004
rect 2475 60955 2517 60964
rect 2476 41273 2516 60955
rect 2668 59240 2708 61888
rect 2764 60332 2804 66088
rect 2860 65960 2900 65969
rect 2860 63104 2900 65920
rect 2860 63055 2900 63064
rect 2764 60283 2804 60292
rect 2956 63020 2996 63029
rect 2668 59191 2708 59200
rect 2764 56384 2804 56393
rect 2764 55376 2804 56344
rect 2764 55327 2804 55336
rect 2956 54956 2996 62980
rect 2956 54907 2996 54916
rect 2572 52772 2612 52781
rect 2572 51932 2612 52732
rect 2572 51883 2612 51892
rect 2764 51764 2804 51773
rect 2572 50588 2612 50597
rect 2572 50420 2612 50548
rect 2572 50371 2612 50380
rect 2764 47900 2804 51724
rect 2764 47851 2804 47860
rect 3052 46640 3092 71968
rect 3148 70832 3188 72976
rect 3148 70783 3188 70792
rect 3148 69740 3188 69749
rect 3148 65624 3188 69700
rect 3244 69404 3284 84316
rect 4396 83516 4436 83525
rect 3688 83180 4056 83189
rect 3728 83140 3770 83180
rect 3810 83140 3852 83180
rect 3892 83140 3934 83180
rect 3974 83140 4016 83180
rect 3688 83131 4056 83140
rect 4300 82424 4340 82433
rect 3688 81668 4056 81677
rect 3728 81628 3770 81668
rect 3810 81628 3852 81668
rect 3892 81628 3934 81668
rect 3974 81628 4016 81668
rect 3688 81619 4056 81628
rect 3688 80156 4056 80165
rect 3728 80116 3770 80156
rect 3810 80116 3852 80156
rect 3892 80116 3934 80156
rect 3974 80116 4016 80156
rect 3688 80107 4056 80116
rect 3688 78644 4056 78653
rect 3728 78604 3770 78644
rect 3810 78604 3852 78644
rect 3892 78604 3934 78644
rect 3974 78604 4016 78644
rect 3688 78595 4056 78604
rect 4204 77972 4244 77981
rect 3244 69355 3284 69364
rect 3340 77720 3380 77729
rect 3340 71756 3380 77680
rect 3148 65575 3188 65584
rect 3148 63356 3188 63365
rect 3148 63104 3188 63316
rect 3148 63055 3188 63064
rect 3148 62180 3188 62189
rect 3148 57896 3188 62140
rect 3148 57847 3188 57856
rect 3340 61172 3380 71716
rect 3436 77468 3476 77477
rect 3436 71000 3476 77428
rect 3688 77132 4056 77141
rect 3728 77092 3770 77132
rect 3810 77092 3852 77132
rect 3892 77092 3934 77132
rect 3974 77092 4016 77132
rect 3688 77083 4056 77092
rect 3532 76544 3572 76553
rect 3532 73100 3572 76504
rect 3688 75620 4056 75629
rect 3728 75580 3770 75620
rect 3810 75580 3852 75620
rect 3892 75580 3934 75620
rect 3974 75580 4016 75620
rect 3688 75571 4056 75580
rect 4108 74276 4148 74285
rect 3688 74108 4056 74117
rect 3728 74068 3770 74108
rect 3810 74068 3852 74108
rect 3892 74068 3934 74108
rect 3974 74068 4016 74108
rect 3688 74059 4056 74068
rect 3532 73051 3572 73060
rect 3532 72596 3572 72605
rect 3532 71420 3572 72556
rect 3688 72596 4056 72605
rect 3728 72556 3770 72596
rect 3810 72556 3852 72596
rect 3892 72556 3934 72596
rect 3974 72556 4016 72596
rect 3688 72547 4056 72556
rect 3532 71371 3572 71380
rect 3688 71084 4056 71093
rect 3728 71044 3770 71084
rect 3810 71044 3852 71084
rect 3892 71044 3934 71084
rect 3974 71044 4016 71084
rect 3688 71035 4056 71044
rect 3436 70960 3572 71000
rect 3436 69740 3476 69749
rect 3436 68564 3476 69700
rect 3436 68515 3476 68524
rect 3436 67304 3476 67313
rect 3436 65624 3476 67264
rect 3436 65575 3476 65584
rect 3244 56300 3284 56309
rect 3244 52940 3284 56260
rect 3244 52891 3284 52900
rect 3340 55628 3380 61132
rect 3340 52520 3380 55588
rect 3436 54788 3476 54797
rect 3436 52772 3476 54748
rect 3436 52723 3476 52732
rect 3052 46600 3188 46640
rect 2860 44960 2900 44969
rect 2475 41264 2517 41273
rect 2475 41224 2476 41264
rect 2516 41224 2517 41264
rect 2475 41215 2517 41224
rect 2476 38744 2516 38753
rect 2476 31856 2516 38704
rect 2476 31807 2516 31816
rect 2764 28916 2804 28925
rect 2476 26984 2516 26993
rect 2476 26228 2516 26944
rect 2476 26179 2516 26188
rect 2572 26816 2612 26825
rect 2572 22784 2612 26776
rect 2668 25808 2708 25817
rect 2668 25388 2708 25768
rect 2668 25339 2708 25348
rect 2572 22735 2612 22744
rect 2764 20684 2804 28876
rect 2860 28832 2900 44920
rect 2956 41852 2996 41861
rect 2956 29000 2996 41812
rect 2956 28951 2996 28960
rect 3052 37400 3092 37409
rect 2860 28792 2996 28832
rect 2860 25976 2900 25985
rect 2860 23801 2900 25936
rect 2859 23792 2901 23801
rect 2859 23752 2860 23792
rect 2900 23752 2901 23792
rect 2859 23743 2901 23752
rect 2956 22877 2996 28792
rect 2955 22868 2997 22877
rect 2955 22828 2956 22868
rect 2996 22828 2997 22868
rect 2955 22819 2997 22828
rect 2764 20635 2804 20644
rect 3052 20264 3092 37360
rect 3148 35636 3188 46600
rect 3340 45632 3380 52480
rect 3340 45583 3380 45592
rect 3340 39248 3380 39257
rect 3244 38912 3284 38921
rect 3244 35888 3284 38872
rect 3244 35839 3284 35848
rect 3148 35587 3188 35596
rect 3244 32780 3284 32789
rect 3148 30344 3188 30353
rect 3148 28421 3188 30304
rect 3147 28412 3189 28421
rect 3147 28372 3148 28412
rect 3188 28372 3189 28412
rect 3147 28363 3189 28372
rect 3148 28244 3188 28253
rect 3148 20768 3188 28204
rect 3148 20719 3188 20728
rect 3052 20180 3092 20224
rect 3052 20140 3188 20180
rect 3148 19424 3188 20140
rect 3148 19375 3188 19384
rect 3052 18920 3092 18929
rect 3052 17660 3092 18880
rect 2956 17492 2996 17501
rect 2956 16829 2996 17452
rect 3052 17072 3092 17620
rect 3052 17023 3092 17032
rect 3148 17828 3188 17837
rect 2955 16820 2997 16829
rect 2955 16780 2956 16820
rect 2996 16780 2997 16820
rect 2955 16771 2997 16780
rect 2188 3835 2228 3844
rect 2284 7792 2420 7832
rect 2476 16400 2516 16409
rect 2284 1364 2324 7792
rect 2380 7160 2420 7169
rect 2380 6152 2420 7120
rect 2380 6103 2420 6112
rect 2380 5564 2420 5573
rect 2380 3380 2420 5524
rect 2380 3331 2420 3340
rect 2476 1868 2516 16360
rect 2572 10604 2612 10613
rect 2572 8420 2612 10564
rect 2572 8371 2612 8380
rect 2860 10016 2900 10025
rect 2860 5648 2900 9976
rect 2860 5599 2900 5608
rect 2956 9848 2996 9857
rect 2956 4976 2996 9808
rect 2956 4640 2996 4936
rect 2956 4591 2996 4600
rect 3148 3968 3188 17788
rect 3244 14972 3284 32740
rect 3340 26144 3380 39208
rect 3435 28412 3477 28421
rect 3435 28372 3436 28412
rect 3476 28372 3477 28412
rect 3435 28363 3477 28372
rect 3436 27068 3476 28363
rect 3436 27019 3476 27028
rect 3532 26816 3572 70960
rect 4108 70748 4148 74236
rect 4108 70699 4148 70708
rect 3688 69572 4056 69581
rect 3728 69532 3770 69572
rect 3810 69532 3852 69572
rect 3892 69532 3934 69572
rect 3974 69532 4016 69572
rect 3688 69523 4056 69532
rect 3627 68564 3669 68573
rect 3627 68524 3628 68564
rect 3668 68524 3669 68564
rect 3627 68515 3669 68524
rect 3628 68430 3668 68515
rect 4108 68228 4148 68237
rect 3688 68060 4056 68069
rect 3728 68020 3770 68060
rect 3810 68020 3852 68060
rect 3892 68020 3934 68060
rect 3974 68020 4016 68060
rect 3688 68011 4056 68020
rect 3819 67472 3861 67481
rect 3819 67432 3820 67472
rect 3860 67432 3861 67472
rect 3819 67423 3861 67432
rect 3820 67338 3860 67423
rect 3688 66548 4056 66557
rect 3728 66508 3770 66548
rect 3810 66508 3852 66548
rect 3892 66508 3934 66548
rect 3974 66508 4016 66548
rect 3688 66499 4056 66508
rect 3688 65036 4056 65045
rect 3728 64996 3770 65036
rect 3810 64996 3852 65036
rect 3892 64996 3934 65036
rect 3974 64996 4016 65036
rect 3688 64987 4056 64996
rect 4108 64112 4148 68188
rect 4108 64063 4148 64072
rect 3688 63524 4056 63533
rect 3728 63484 3770 63524
rect 3810 63484 3852 63524
rect 3892 63484 3934 63524
rect 3974 63484 4016 63524
rect 3688 63475 4056 63484
rect 3688 62012 4056 62021
rect 3728 61972 3770 62012
rect 3810 61972 3852 62012
rect 3892 61972 3934 62012
rect 3974 61972 4016 62012
rect 3688 61963 4056 61972
rect 3915 61760 3957 61769
rect 3915 61720 3916 61760
rect 3956 61720 3957 61760
rect 3915 61711 3957 61720
rect 3916 61626 3956 61711
rect 3688 60500 4056 60509
rect 3728 60460 3770 60500
rect 3810 60460 3852 60500
rect 3892 60460 3934 60500
rect 3974 60460 4016 60500
rect 3688 60451 4056 60460
rect 3688 58988 4056 58997
rect 3728 58948 3770 58988
rect 3810 58948 3852 58988
rect 3892 58948 3934 58988
rect 3974 58948 4016 58988
rect 3688 58939 4056 58948
rect 3688 57476 4056 57485
rect 3728 57436 3770 57476
rect 3810 57436 3852 57476
rect 3892 57436 3934 57476
rect 3974 57436 4016 57476
rect 3688 57427 4056 57436
rect 3688 55964 4056 55973
rect 3728 55924 3770 55964
rect 3810 55924 3852 55964
rect 3892 55924 3934 55964
rect 3974 55924 4016 55964
rect 3688 55915 4056 55924
rect 4108 54872 4148 54881
rect 3688 54452 4056 54461
rect 3728 54412 3770 54452
rect 3810 54412 3852 54452
rect 3892 54412 3934 54452
rect 3974 54412 4016 54452
rect 3688 54403 4056 54412
rect 3688 52940 4056 52949
rect 3728 52900 3770 52940
rect 3810 52900 3852 52940
rect 3892 52900 3934 52940
rect 3974 52900 4016 52940
rect 3688 52891 4056 52900
rect 3688 51428 4056 51437
rect 3728 51388 3770 51428
rect 3810 51388 3852 51428
rect 3892 51388 3934 51428
rect 3974 51388 4016 51428
rect 3688 51379 4056 51388
rect 3688 49916 4056 49925
rect 3728 49876 3770 49916
rect 3810 49876 3852 49916
rect 3892 49876 3934 49916
rect 3974 49876 4016 49916
rect 3688 49867 4056 49876
rect 3688 48404 4056 48413
rect 3728 48364 3770 48404
rect 3810 48364 3852 48404
rect 3892 48364 3934 48404
rect 3974 48364 4016 48404
rect 3688 48355 4056 48364
rect 4108 47396 4148 54832
rect 4108 47347 4148 47356
rect 3688 46892 4056 46901
rect 3728 46852 3770 46892
rect 3810 46852 3852 46892
rect 3892 46852 3934 46892
rect 3974 46852 4016 46892
rect 3688 46843 4056 46852
rect 3688 45380 4056 45389
rect 3728 45340 3770 45380
rect 3810 45340 3852 45380
rect 3892 45340 3934 45380
rect 3974 45340 4016 45380
rect 3688 45331 4056 45340
rect 3688 43868 4056 43877
rect 3728 43828 3770 43868
rect 3810 43828 3852 43868
rect 3892 43828 3934 43868
rect 3974 43828 4016 43868
rect 3688 43819 4056 43828
rect 3688 42356 4056 42365
rect 3728 42316 3770 42356
rect 3810 42316 3852 42356
rect 3892 42316 3934 42356
rect 3974 42316 4016 42356
rect 3688 42307 4056 42316
rect 3688 40844 4056 40853
rect 3728 40804 3770 40844
rect 3810 40804 3852 40844
rect 3892 40804 3934 40844
rect 3974 40804 4016 40844
rect 3688 40795 4056 40804
rect 3688 39332 4056 39341
rect 3728 39292 3770 39332
rect 3810 39292 3852 39332
rect 3892 39292 3934 39332
rect 3974 39292 4016 39332
rect 3688 39283 4056 39292
rect 3688 37820 4056 37829
rect 3728 37780 3770 37820
rect 3810 37780 3852 37820
rect 3892 37780 3934 37820
rect 3974 37780 4016 37820
rect 3688 37771 4056 37780
rect 3688 36308 4056 36317
rect 3728 36268 3770 36308
rect 3810 36268 3852 36308
rect 3892 36268 3934 36308
rect 3974 36268 4016 36308
rect 3688 36259 4056 36268
rect 3819 35048 3861 35057
rect 3819 35008 3820 35048
rect 3860 35008 3861 35048
rect 3819 34999 3861 35008
rect 3820 34914 3860 34999
rect 3688 34796 4056 34805
rect 3728 34756 3770 34796
rect 3810 34756 3852 34796
rect 3892 34756 3934 34796
rect 3974 34756 4016 34796
rect 3688 34747 4056 34756
rect 3915 34292 3957 34301
rect 3915 34252 3916 34292
rect 3956 34252 3957 34292
rect 3915 34243 3957 34252
rect 3916 34158 3956 34243
rect 3688 33284 4056 33293
rect 3728 33244 3770 33284
rect 3810 33244 3852 33284
rect 3892 33244 3934 33284
rect 3974 33244 4016 33284
rect 3688 33235 4056 33244
rect 4108 31940 4148 31949
rect 3688 31772 4056 31781
rect 3728 31732 3770 31772
rect 3810 31732 3852 31772
rect 3892 31732 3934 31772
rect 3974 31732 4016 31772
rect 3688 31723 4056 31732
rect 3688 30260 4056 30269
rect 3728 30220 3770 30260
rect 3810 30220 3852 30260
rect 3892 30220 3934 30260
rect 3974 30220 4016 30260
rect 3688 30211 4056 30220
rect 4108 29840 4148 31900
rect 4108 29791 4148 29800
rect 4204 29168 4244 77932
rect 4300 69992 4340 82384
rect 4300 69943 4340 69952
rect 4396 42776 4436 83476
rect 4684 79736 4724 79745
rect 4588 76880 4628 76889
rect 4588 75956 4628 76840
rect 4588 66548 4628 75916
rect 4588 66296 4628 66508
rect 4588 66247 4628 66256
rect 4491 63020 4533 63029
rect 4491 62980 4492 63020
rect 4532 62980 4533 63020
rect 4491 62971 4533 62980
rect 4492 62886 4532 62971
rect 4587 61004 4629 61013
rect 4587 60964 4588 61004
rect 4628 60964 4629 61004
rect 4587 60955 4629 60964
rect 4588 60870 4628 60955
rect 4684 60332 4724 79696
rect 4780 77552 4820 85408
rect 8236 84944 8276 84953
rect 5548 84524 5588 84533
rect 4928 83936 5296 83945
rect 4968 83896 5010 83936
rect 5050 83896 5092 83936
rect 5132 83896 5174 83936
rect 5214 83896 5256 83936
rect 4928 83887 5296 83896
rect 4928 82424 5296 82433
rect 4968 82384 5010 82424
rect 5050 82384 5092 82424
rect 5132 82384 5174 82424
rect 5214 82384 5256 82424
rect 4928 82375 5296 82384
rect 4928 80912 5296 80921
rect 4968 80872 5010 80912
rect 5050 80872 5092 80912
rect 5132 80872 5174 80912
rect 5214 80872 5256 80912
rect 4928 80863 5296 80872
rect 5452 80492 5492 80501
rect 5356 79820 5396 79829
rect 4928 79400 5296 79409
rect 4968 79360 5010 79400
rect 5050 79360 5092 79400
rect 5132 79360 5174 79400
rect 5214 79360 5256 79400
rect 4928 79351 5296 79360
rect 4928 77888 5296 77897
rect 4968 77848 5010 77888
rect 5050 77848 5092 77888
rect 5132 77848 5174 77888
rect 5214 77848 5256 77888
rect 4928 77839 5296 77848
rect 4780 77503 4820 77512
rect 4928 76376 5296 76385
rect 4968 76336 5010 76376
rect 5050 76336 5092 76376
rect 5132 76336 5174 76376
rect 5214 76336 5256 76376
rect 4928 76327 5296 76336
rect 4780 75956 4820 75965
rect 4780 70664 4820 75916
rect 4928 74864 5296 74873
rect 4968 74824 5010 74864
rect 5050 74824 5092 74864
rect 5132 74824 5174 74864
rect 5214 74824 5256 74864
rect 4928 74815 5296 74824
rect 4928 73352 5296 73361
rect 4968 73312 5010 73352
rect 5050 73312 5092 73352
rect 5132 73312 5174 73352
rect 5214 73312 5256 73352
rect 4928 73303 5296 73312
rect 4928 71840 5296 71849
rect 4968 71800 5010 71840
rect 5050 71800 5092 71840
rect 5132 71800 5174 71840
rect 5214 71800 5256 71840
rect 4928 71791 5296 71800
rect 4780 70615 4820 70624
rect 4928 70328 5296 70337
rect 4968 70288 5010 70328
rect 5050 70288 5092 70328
rect 5132 70288 5174 70328
rect 5214 70288 5256 70328
rect 4928 70279 5296 70288
rect 4780 69572 4820 69581
rect 4780 68312 4820 69532
rect 4928 68816 5296 68825
rect 4968 68776 5010 68816
rect 5050 68776 5092 68816
rect 5132 68776 5174 68816
rect 5214 68776 5256 68816
rect 4928 68767 5296 68776
rect 4875 68564 4917 68573
rect 4875 68524 4876 68564
rect 4916 68524 4917 68564
rect 4875 68515 4917 68524
rect 4876 68430 4916 68515
rect 4780 68263 4820 68272
rect 4928 67304 5296 67313
rect 4968 67264 5010 67304
rect 5050 67264 5092 67304
rect 5132 67264 5174 67304
rect 5214 67264 5256 67304
rect 4928 67255 5296 67264
rect 4780 66800 4820 66809
rect 4780 62684 4820 66760
rect 4928 65792 5296 65801
rect 4968 65752 5010 65792
rect 5050 65752 5092 65792
rect 5132 65752 5174 65792
rect 5214 65752 5256 65792
rect 4928 65743 5296 65752
rect 4928 64280 5296 64289
rect 4968 64240 5010 64280
rect 5050 64240 5092 64280
rect 5132 64240 5174 64280
rect 5214 64240 5256 64280
rect 4928 64231 5296 64240
rect 4928 62768 5296 62777
rect 4968 62728 5010 62768
rect 5050 62728 5092 62768
rect 5132 62728 5174 62768
rect 5214 62728 5256 62768
rect 4928 62719 5296 62728
rect 4780 62635 4820 62644
rect 4928 61256 5296 61265
rect 4968 61216 5010 61256
rect 5050 61216 5092 61256
rect 5132 61216 5174 61256
rect 5214 61216 5256 61256
rect 4928 61207 5296 61216
rect 4684 60283 4724 60292
rect 4780 61088 4820 61097
rect 4780 58736 4820 61048
rect 4928 59744 5296 59753
rect 4968 59704 5010 59744
rect 5050 59704 5092 59744
rect 5132 59704 5174 59744
rect 5214 59704 5256 59744
rect 4928 59695 5296 59704
rect 4780 58687 4820 58696
rect 4928 58232 5296 58241
rect 4968 58192 5010 58232
rect 5050 58192 5092 58232
rect 5132 58192 5174 58232
rect 5214 58192 5256 58232
rect 4928 58183 5296 58192
rect 4928 56720 5296 56729
rect 4968 56680 5010 56720
rect 5050 56680 5092 56720
rect 5132 56680 5174 56720
rect 5214 56680 5256 56720
rect 4928 56671 5296 56680
rect 4928 55208 5296 55217
rect 4968 55168 5010 55208
rect 5050 55168 5092 55208
rect 5132 55168 5174 55208
rect 5214 55168 5256 55208
rect 4928 55159 5296 55168
rect 4928 53696 5296 53705
rect 4968 53656 5010 53696
rect 5050 53656 5092 53696
rect 5132 53656 5174 53696
rect 5214 53656 5256 53696
rect 4928 53647 5296 53656
rect 4928 52184 5296 52193
rect 4968 52144 5010 52184
rect 5050 52144 5092 52184
rect 5132 52144 5174 52184
rect 5214 52144 5256 52184
rect 4928 52135 5296 52144
rect 4928 50672 5296 50681
rect 4968 50632 5010 50672
rect 5050 50632 5092 50672
rect 5132 50632 5174 50672
rect 5214 50632 5256 50672
rect 4928 50623 5296 50632
rect 4928 49160 5296 49169
rect 4968 49120 5010 49160
rect 5050 49120 5092 49160
rect 5132 49120 5174 49160
rect 5214 49120 5256 49160
rect 4928 49111 5296 49120
rect 4928 47648 5296 47657
rect 4968 47608 5010 47648
rect 5050 47608 5092 47648
rect 5132 47608 5174 47648
rect 5214 47608 5256 47648
rect 4928 47599 5296 47608
rect 4928 46136 5296 46145
rect 4968 46096 5010 46136
rect 5050 46096 5092 46136
rect 5132 46096 5174 46136
rect 5214 46096 5256 46136
rect 4928 46087 5296 46096
rect 4928 44624 5296 44633
rect 4968 44584 5010 44624
rect 5050 44584 5092 44624
rect 5132 44584 5174 44624
rect 5214 44584 5256 44624
rect 4928 44575 5296 44584
rect 4928 43112 5296 43121
rect 4968 43072 5010 43112
rect 5050 43072 5092 43112
rect 5132 43072 5174 43112
rect 5214 43072 5256 43112
rect 4928 43063 5296 43072
rect 4396 41600 4436 42736
rect 4396 41551 4436 41560
rect 4928 41600 5296 41609
rect 4968 41560 5010 41600
rect 5050 41560 5092 41600
rect 5132 41560 5174 41600
rect 5214 41560 5256 41600
rect 4928 41551 5296 41560
rect 4492 40928 4532 40937
rect 4204 29119 4244 29128
rect 4396 34208 4436 34217
rect 4396 33620 4436 34168
rect 3688 28748 4056 28757
rect 3728 28708 3770 28748
rect 3810 28708 3852 28748
rect 3892 28708 3934 28748
rect 3974 28708 4016 28748
rect 3688 28699 4056 28708
rect 4300 28160 4340 28169
rect 4300 27488 4340 28120
rect 4300 27439 4340 27448
rect 3688 27236 4056 27245
rect 3728 27196 3770 27236
rect 3810 27196 3852 27236
rect 3892 27196 3934 27236
rect 3974 27196 4016 27236
rect 3688 27187 4056 27196
rect 3532 26767 3572 26776
rect 4204 27152 4244 27161
rect 3532 26144 3572 26153
rect 3340 26104 3532 26144
rect 3340 25976 3380 25985
rect 3340 24548 3380 25936
rect 3340 22280 3380 24508
rect 3340 22231 3380 22240
rect 3436 25388 3476 25397
rect 3436 23876 3476 25348
rect 3436 21692 3476 23836
rect 3436 21643 3476 21652
rect 3436 20768 3476 20777
rect 3436 17408 3476 20728
rect 3532 20096 3572 26104
rect 3688 25724 4056 25733
rect 3728 25684 3770 25724
rect 3810 25684 3852 25724
rect 3892 25684 3934 25724
rect 3974 25684 4016 25724
rect 3688 25675 4056 25684
rect 3688 24212 4056 24221
rect 3728 24172 3770 24212
rect 3810 24172 3852 24212
rect 3892 24172 3934 24212
rect 3974 24172 4016 24212
rect 3688 24163 4056 24172
rect 4204 23204 4244 27112
rect 4396 26480 4436 33580
rect 4396 26431 4436 26440
rect 4204 23155 4244 23164
rect 4396 25052 4436 25061
rect 4204 23036 4244 23045
rect 3688 22700 4056 22709
rect 3728 22660 3770 22700
rect 3810 22660 3852 22700
rect 3892 22660 3934 22700
rect 3974 22660 4016 22700
rect 3688 22651 4056 22660
rect 3688 21188 4056 21197
rect 3728 21148 3770 21188
rect 3810 21148 3852 21188
rect 3892 21148 3934 21188
rect 3974 21148 4016 21188
rect 3688 21139 4056 21148
rect 3532 20047 3572 20056
rect 3688 19676 4056 19685
rect 3728 19636 3770 19676
rect 3810 19636 3852 19676
rect 3892 19636 3934 19676
rect 3974 19636 4016 19676
rect 3688 19627 4056 19636
rect 4204 19340 4244 22996
rect 4204 19291 4244 19300
rect 4396 19256 4436 25012
rect 4396 19207 4436 19216
rect 4492 22280 4532 40888
rect 4780 40424 4820 40433
rect 4780 38828 4820 40384
rect 4928 40088 5296 40097
rect 4968 40048 5010 40088
rect 5050 40048 5092 40088
rect 5132 40048 5174 40088
rect 5214 40048 5256 40088
rect 4928 40039 5296 40048
rect 4780 38779 4820 38788
rect 4928 38576 5296 38585
rect 4968 38536 5010 38576
rect 5050 38536 5092 38576
rect 5132 38536 5174 38576
rect 5214 38536 5256 38576
rect 4928 38527 5296 38536
rect 4928 37064 5296 37073
rect 4968 37024 5010 37064
rect 5050 37024 5092 37064
rect 5132 37024 5174 37064
rect 5214 37024 5256 37064
rect 4928 37015 5296 37024
rect 5356 36812 5396 79780
rect 5356 36737 5396 36772
rect 5452 41264 5492 80452
rect 5548 79400 5588 84484
rect 7372 84524 7412 84533
rect 5836 84440 5876 84449
rect 5836 81920 5876 84400
rect 6124 84440 6164 84449
rect 6028 83516 6068 83525
rect 5836 81880 5972 81920
rect 5548 79360 5876 79400
rect 5644 72008 5684 72017
rect 5548 68648 5588 68657
rect 5548 66044 5588 68608
rect 5548 65995 5588 66004
rect 5548 65204 5588 65213
rect 5548 64112 5588 65164
rect 5548 64063 5588 64072
rect 5355 36728 5397 36737
rect 5355 36688 5356 36728
rect 5396 36688 5397 36728
rect 5355 36679 5397 36688
rect 5356 36677 5396 36679
rect 4928 35552 5296 35561
rect 4968 35512 5010 35552
rect 5050 35512 5092 35552
rect 5132 35512 5174 35552
rect 5214 35512 5256 35552
rect 4928 35503 5296 35512
rect 4928 34040 5296 34049
rect 4968 34000 5010 34040
rect 5050 34000 5092 34040
rect 5132 34000 5174 34040
rect 5214 34000 5256 34040
rect 4928 33991 5296 34000
rect 5356 32780 5396 32789
rect 4928 32528 5296 32537
rect 4968 32488 5010 32528
rect 5050 32488 5092 32528
rect 5132 32488 5174 32528
rect 5214 32488 5256 32528
rect 4928 32479 5296 32488
rect 4928 31016 5296 31025
rect 4968 30976 5010 31016
rect 5050 30976 5092 31016
rect 5132 30976 5174 31016
rect 5214 30976 5256 31016
rect 4928 30967 5296 30976
rect 4928 29504 5296 29513
rect 4968 29464 5010 29504
rect 5050 29464 5092 29504
rect 5132 29464 5174 29504
rect 5214 29464 5256 29504
rect 4928 29455 5296 29464
rect 4780 29084 4820 29093
rect 3688 18164 4056 18173
rect 3728 18124 3770 18164
rect 3810 18124 3852 18164
rect 3892 18124 3934 18164
rect 3974 18124 4016 18164
rect 3688 18115 4056 18124
rect 4492 17828 4532 22240
rect 4588 26648 4628 26657
rect 4588 24800 4628 26608
rect 4684 26312 4724 26321
rect 4684 26069 4724 26272
rect 4683 26060 4725 26069
rect 4683 26020 4684 26060
rect 4724 26020 4725 26060
rect 4683 26011 4725 26020
rect 4780 25724 4820 29044
rect 4928 27992 5296 28001
rect 4968 27952 5010 27992
rect 5050 27952 5092 27992
rect 5132 27952 5174 27992
rect 5214 27952 5256 27992
rect 4928 27943 5296 27952
rect 4928 26480 5296 26489
rect 4968 26440 5010 26480
rect 5050 26440 5092 26480
rect 5132 26440 5174 26480
rect 5214 26440 5256 26480
rect 4928 26431 5296 26440
rect 4780 25675 4820 25684
rect 4972 25640 5012 25649
rect 4876 25600 4972 25640
rect 4780 25220 4820 25229
rect 4876 25220 4916 25600
rect 4972 25591 5012 25600
rect 4820 25180 4916 25220
rect 5067 25220 5109 25229
rect 5067 25180 5068 25220
rect 5108 25180 5109 25220
rect 4780 25171 4820 25180
rect 5067 25171 5109 25180
rect 5068 25086 5108 25171
rect 5260 25145 5300 25230
rect 5259 25136 5301 25145
rect 5259 25096 5260 25136
rect 5300 25096 5301 25136
rect 5259 25087 5301 25096
rect 4928 24968 5296 24977
rect 4968 24928 5010 24968
rect 5050 24928 5092 24968
rect 5132 24928 5174 24968
rect 5214 24928 5256 24968
rect 4928 24919 5296 24928
rect 4588 18584 4628 24760
rect 4928 23456 5296 23465
rect 4968 23416 5010 23456
rect 5050 23416 5092 23456
rect 5132 23416 5174 23456
rect 5214 23416 5256 23456
rect 4928 23407 5296 23416
rect 4928 21944 5296 21953
rect 4968 21904 5010 21944
rect 5050 21904 5092 21944
rect 5132 21904 5174 21944
rect 5214 21904 5256 21944
rect 4928 21895 5296 21904
rect 4780 20768 4820 20777
rect 4780 20180 4820 20728
rect 4928 20432 5296 20441
rect 4968 20392 5010 20432
rect 5050 20392 5092 20432
rect 5132 20392 5174 20432
rect 5214 20392 5256 20432
rect 4928 20383 5296 20392
rect 4780 20131 4820 20140
rect 5356 19004 5396 32740
rect 5356 18955 5396 18964
rect 4928 18920 5296 18929
rect 4968 18880 5010 18920
rect 5050 18880 5092 18920
rect 5132 18880 5174 18920
rect 5214 18880 5256 18920
rect 4928 18871 5296 18880
rect 4588 18535 4628 18544
rect 4492 17779 4532 17788
rect 4395 17576 4437 17585
rect 4395 17536 4396 17576
rect 4436 17536 4437 17576
rect 4395 17527 4437 17536
rect 4588 17576 4628 17585
rect 4396 17442 4436 17527
rect 3436 17359 3476 17368
rect 4108 17072 4148 17081
rect 3688 16652 4056 16661
rect 3728 16612 3770 16652
rect 3810 16612 3852 16652
rect 3892 16612 3934 16652
rect 3974 16612 4016 16652
rect 3688 16603 4056 16612
rect 3244 14923 3284 14932
rect 3340 16400 3380 16409
rect 3340 14552 3380 16360
rect 3340 14503 3380 14512
rect 3436 15308 3476 15317
rect 3436 4640 3476 15268
rect 3688 15140 4056 15149
rect 3728 15100 3770 15140
rect 3810 15100 3852 15140
rect 3892 15100 3934 15140
rect 3974 15100 4016 15140
rect 3688 15091 4056 15100
rect 3688 13628 4056 13637
rect 3728 13588 3770 13628
rect 3810 13588 3852 13628
rect 3892 13588 3934 13628
rect 3974 13588 4016 13628
rect 3688 13579 4056 13588
rect 4108 13208 4148 17032
rect 4300 15728 4340 15737
rect 4204 14720 4244 14729
rect 4204 14132 4244 14680
rect 4204 14083 4244 14092
rect 3688 12116 4056 12125
rect 3728 12076 3770 12116
rect 3810 12076 3852 12116
rect 3892 12076 3934 12116
rect 3974 12076 4016 12116
rect 3688 12067 4056 12076
rect 4108 11276 4148 13168
rect 4300 11528 4340 15688
rect 4300 11479 4340 11488
rect 4108 11227 4148 11236
rect 4588 11108 4628 17536
rect 5356 17492 5396 17501
rect 4928 17408 5296 17417
rect 4968 17368 5010 17408
rect 5050 17368 5092 17408
rect 5132 17368 5174 17408
rect 5214 17368 5256 17408
rect 4928 17359 5296 17368
rect 5356 17072 5396 17452
rect 5356 17023 5396 17032
rect 4928 15896 5296 15905
rect 4968 15856 5010 15896
rect 5050 15856 5092 15896
rect 5132 15856 5174 15896
rect 5214 15856 5256 15896
rect 4928 15847 5296 15856
rect 4928 14384 5296 14393
rect 4968 14344 5010 14384
rect 5050 14344 5092 14384
rect 5132 14344 5174 14384
rect 5214 14344 5256 14384
rect 4928 14335 5296 14344
rect 4928 12872 5296 12881
rect 4968 12832 5010 12872
rect 5050 12832 5092 12872
rect 5132 12832 5174 12872
rect 5214 12832 5256 12872
rect 4928 12823 5296 12832
rect 4928 11360 5296 11369
rect 4968 11320 5010 11360
rect 5050 11320 5092 11360
rect 5132 11320 5174 11360
rect 5214 11320 5256 11360
rect 4928 11311 5296 11320
rect 4588 11059 4628 11068
rect 3688 10604 4056 10613
rect 3728 10564 3770 10604
rect 3810 10564 3852 10604
rect 3892 10564 3934 10604
rect 3974 10564 4016 10604
rect 3688 10555 4056 10564
rect 4684 9848 4724 9857
rect 3688 9092 4056 9101
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 3688 9043 4056 9052
rect 3688 7580 4056 7589
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 3688 7531 4056 7540
rect 4684 6488 4724 9808
rect 4928 9848 5296 9857
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 4928 9799 5296 9808
rect 5356 8504 5396 8513
rect 4928 8336 5296 8345
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 4928 8287 5296 8296
rect 5356 8084 5396 8464
rect 5356 8035 5396 8044
rect 3688 6068 4056 6077
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 3688 6019 4056 6028
rect 4684 4808 4724 6448
rect 4780 7244 4820 7253
rect 4780 5648 4820 7204
rect 4928 6824 5296 6833
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 4928 6775 5296 6784
rect 4780 5599 4820 5608
rect 4928 5312 5296 5321
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 4928 5263 5296 5272
rect 4684 4759 4724 4768
rect 3436 4591 3476 4600
rect 3688 4556 4056 4565
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 3688 4507 4056 4516
rect 3148 3919 3188 3928
rect 4928 3800 5296 3809
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 4928 3751 5296 3760
rect 3688 3044 4056 3053
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 3688 2995 4056 3004
rect 5356 2708 5396 2717
rect 4928 2288 5296 2297
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 4928 2239 5296 2248
rect 5356 2120 5396 2668
rect 5356 2071 5396 2080
rect 2476 1819 2516 1828
rect 3688 1532 4056 1541
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 3688 1483 4056 1492
rect 2284 1315 2324 1324
rect 5452 1280 5492 41224
rect 5548 60332 5588 60341
rect 5548 35132 5588 60292
rect 5644 59324 5684 71968
rect 5740 69908 5780 69917
rect 5740 60920 5780 69868
rect 5836 64457 5876 79360
rect 5932 64868 5972 81880
rect 6028 75116 6068 83476
rect 6028 75067 6068 75076
rect 6028 74528 6068 74537
rect 6028 72260 6068 74488
rect 6028 72211 6068 72220
rect 5932 64819 5972 64828
rect 6028 66632 6068 66641
rect 6028 65708 6068 66592
rect 5835 64448 5877 64457
rect 5835 64408 5836 64448
rect 5876 64408 5877 64448
rect 5835 64399 5877 64408
rect 5932 64364 5972 64373
rect 5932 62936 5972 64324
rect 6028 64112 6068 65668
rect 6028 64063 6068 64072
rect 5932 62887 5972 62896
rect 6124 62852 6164 84400
rect 6412 84440 6452 84449
rect 6220 72260 6260 72269
rect 6220 72008 6260 72220
rect 6220 71959 6260 71968
rect 6316 66632 6356 66641
rect 6316 65288 6356 66592
rect 6316 65239 6356 65248
rect 6124 62803 6164 62812
rect 6412 61844 6452 84400
rect 6700 84440 6740 84449
rect 6508 76964 6548 76973
rect 6508 75620 6548 76924
rect 6508 75571 6548 75580
rect 6412 61795 6452 61804
rect 6508 73520 6548 73529
rect 5740 60871 5780 60880
rect 5644 59275 5684 59284
rect 6316 60500 6356 60509
rect 6316 57896 6356 60460
rect 6220 57056 6260 57065
rect 5644 52940 5684 52949
rect 5644 50000 5684 52900
rect 5644 49951 5684 49960
rect 6220 48824 6260 57016
rect 6316 53612 6356 57856
rect 6412 59240 6452 59249
rect 6412 58988 6452 59200
rect 6412 57644 6452 58948
rect 6412 57595 6452 57604
rect 6316 53024 6356 53572
rect 6316 52975 6356 52984
rect 6220 48775 6260 48784
rect 6412 52436 6452 52445
rect 6220 48488 6260 48497
rect 6124 48404 6164 48413
rect 5932 47984 5972 47993
rect 5932 46640 5972 47944
rect 6124 47984 6164 48364
rect 6124 47648 6164 47944
rect 6124 47599 6164 47608
rect 5932 46591 5972 46600
rect 6220 44288 6260 48448
rect 6220 44120 6260 44248
rect 6220 44071 6260 44080
rect 6027 42776 6069 42785
rect 6027 42736 6028 42776
rect 6068 42736 6069 42776
rect 6027 42727 6069 42736
rect 6028 42642 6068 42727
rect 5931 41264 5973 41273
rect 5931 41224 5932 41264
rect 5972 41224 5973 41264
rect 5931 41215 5973 41224
rect 5548 35083 5588 35092
rect 5740 41180 5780 41189
rect 5548 29168 5588 29177
rect 5548 24548 5588 29128
rect 5740 24884 5780 41140
rect 5932 40928 5972 41215
rect 5932 40879 5972 40888
rect 5836 38156 5876 38165
rect 5836 35300 5876 38116
rect 5836 35251 5876 35260
rect 6028 34376 6068 34385
rect 6028 32276 6068 34336
rect 5740 24835 5780 24844
rect 5836 30764 5876 30773
rect 5548 16736 5588 24508
rect 5644 24800 5684 24809
rect 5644 20012 5684 24760
rect 5644 19963 5684 19972
rect 5739 17576 5781 17585
rect 5739 17536 5740 17576
rect 5780 17536 5781 17576
rect 5739 17527 5781 17536
rect 5740 17442 5780 17527
rect 5643 16820 5685 16829
rect 5643 16780 5644 16820
rect 5684 16780 5685 16820
rect 5643 16771 5685 16780
rect 5548 7832 5588 16696
rect 5644 13292 5684 16771
rect 5644 13243 5684 13252
rect 5548 7783 5588 7792
rect 5740 3800 5780 3809
rect 5548 2456 5588 2465
rect 5548 1952 5588 2416
rect 5740 2288 5780 3760
rect 5740 2239 5780 2248
rect 5548 1903 5588 1912
rect 5836 1868 5876 30724
rect 5932 25892 5972 25901
rect 5932 18920 5972 25852
rect 6028 24296 6068 32236
rect 6028 24247 6068 24256
rect 6124 26144 6164 26153
rect 6124 24464 6164 26104
rect 6124 19760 6164 24424
rect 6124 19711 6164 19720
rect 6316 25220 6356 25229
rect 6316 19340 6356 25180
rect 6316 19291 6356 19300
rect 5932 18871 5972 18880
rect 6316 16820 6356 16829
rect 6220 13376 6260 13385
rect 6220 11276 6260 13336
rect 6316 12956 6356 16780
rect 6316 12907 6356 12916
rect 6220 11227 6260 11236
rect 5836 1819 5876 1828
rect 6220 7664 6260 7673
rect 5452 1231 5492 1240
rect 6220 1028 6260 7624
rect 6220 979 6260 988
rect 6315 944 6357 953
rect 6315 904 6316 944
rect 6356 904 6357 944
rect 6315 895 6357 904
rect 6316 810 6356 895
rect 4928 776 5296 785
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 4928 727 5296 736
rect 6412 776 6452 52396
rect 6508 51680 6548 73480
rect 6604 72008 6644 72017
rect 6604 71840 6644 71968
rect 6604 71791 6644 71800
rect 6508 51631 6548 51640
rect 6604 51512 6644 51521
rect 6604 50084 6644 51472
rect 6604 50035 6644 50044
rect 6604 26816 6644 26825
rect 6508 24380 6548 24389
rect 6508 23540 6548 24340
rect 6508 20432 6548 23500
rect 6604 21356 6644 26776
rect 6604 21307 6644 21316
rect 6508 20383 6548 20392
rect 6508 19340 6548 19349
rect 6508 15140 6548 19300
rect 6603 16820 6645 16829
rect 6603 16780 6604 16820
rect 6644 16780 6645 16820
rect 6603 16771 6645 16780
rect 6604 16686 6644 16771
rect 6508 15091 6548 15100
rect 6603 2204 6645 2213
rect 6603 2164 6604 2204
rect 6644 2164 6645 2204
rect 6603 2155 6645 2164
rect 6604 2070 6644 2155
rect 6700 2120 6740 84400
rect 7180 84440 7220 84449
rect 7084 83432 7124 83441
rect 6796 80408 6836 80417
rect 6796 41264 6836 80368
rect 6988 74360 7028 74369
rect 6988 73688 7028 74320
rect 6988 73639 7028 73648
rect 6988 70748 7028 70757
rect 6892 66380 6932 66389
rect 6892 64112 6932 66340
rect 6892 64063 6932 64072
rect 6796 41215 6836 41224
rect 6892 36980 6932 36989
rect 6892 36728 6932 36940
rect 6892 36679 6932 36688
rect 6796 35132 6836 35141
rect 6796 32108 6836 35092
rect 6796 32059 6836 32068
rect 6988 30848 7028 70708
rect 7084 68312 7124 83392
rect 7084 68263 7124 68272
rect 6988 30799 7028 30808
rect 7084 38660 7124 38669
rect 7084 38492 7124 38620
rect 6892 29168 6932 29177
rect 6796 24296 6836 24305
rect 6796 18836 6836 24256
rect 6796 18787 6836 18796
rect 6796 16988 6836 16997
rect 6796 13124 6836 16948
rect 6796 9680 6836 13084
rect 6796 9631 6836 9640
rect 6700 2071 6740 2080
rect 6699 1280 6741 1289
rect 6699 1240 6700 1280
rect 6740 1240 6741 1280
rect 6699 1231 6741 1240
rect 6700 1146 6740 1231
rect 6892 1112 6932 29128
rect 6988 27824 7028 27833
rect 6988 27404 7028 27784
rect 6988 27355 7028 27364
rect 7084 27572 7124 38452
rect 7084 26648 7124 27532
rect 7084 26599 7124 26608
rect 7084 25304 7124 25313
rect 6988 25264 7084 25304
rect 6988 19256 7028 25264
rect 7084 25255 7124 25264
rect 6988 19207 7028 19216
rect 7180 12536 7220 84400
rect 7276 68984 7316 68993
rect 7276 28832 7316 68944
rect 7276 28783 7316 28792
rect 7276 23876 7316 23885
rect 7276 23288 7316 23836
rect 7276 23239 7316 23248
rect 7180 12487 7220 12496
rect 7084 8168 7124 8177
rect 6988 5396 7028 5405
rect 6988 5144 7028 5356
rect 6988 5095 7028 5104
rect 6987 4808 7029 4817
rect 6987 4768 6988 4808
rect 7028 4768 7029 4808
rect 6987 4759 7029 4768
rect 6892 1063 6932 1072
rect 6412 727 6452 736
rect 6988 776 7028 4759
rect 7084 944 7124 8128
rect 7372 1280 7412 84484
rect 7755 83516 7797 83525
rect 7755 83476 7756 83516
rect 7796 83476 7797 83516
rect 7755 83467 7797 83476
rect 7756 83382 7796 83467
rect 7660 83264 7700 83273
rect 7564 81836 7604 81845
rect 7468 78140 7508 78149
rect 7468 75704 7508 78100
rect 7468 75655 7508 75664
rect 7468 66716 7508 66725
rect 7468 63524 7508 66676
rect 7564 64112 7604 81796
rect 7564 64063 7604 64072
rect 7468 60248 7508 63484
rect 7564 63440 7604 63449
rect 7564 62852 7604 63400
rect 7564 62803 7604 62812
rect 7468 60199 7508 60208
rect 7564 41684 7604 41693
rect 7468 37148 7508 37157
rect 7468 32192 7508 37108
rect 7468 32143 7508 32152
rect 7564 33200 7604 41644
rect 7660 35300 7700 83224
rect 7756 72512 7796 72521
rect 7756 70496 7796 72472
rect 7756 61760 7796 70456
rect 8140 70664 8180 70673
rect 7948 68060 7988 68069
rect 7852 65792 7892 65801
rect 7852 63020 7892 65752
rect 7852 62971 7892 62980
rect 7948 62264 7988 68020
rect 8044 66128 8084 66137
rect 8044 63692 8084 66088
rect 8044 63643 8084 63652
rect 7948 62215 7988 62224
rect 7756 61711 7796 61720
rect 7948 61844 7988 61853
rect 7660 35251 7700 35260
rect 7852 36392 7892 36401
rect 7468 26312 7508 26321
rect 7468 24380 7508 26272
rect 7564 26144 7604 33160
rect 7756 33956 7796 33965
rect 7660 32696 7700 32705
rect 7660 32024 7700 32656
rect 7756 32528 7796 33916
rect 7756 32479 7796 32488
rect 7660 31975 7700 31984
rect 7564 26095 7604 26104
rect 7468 24331 7508 24340
rect 7756 24548 7796 24557
rect 7756 23960 7796 24508
rect 7660 23288 7700 23297
rect 7468 18080 7508 18089
rect 7468 13880 7508 18040
rect 7660 17072 7700 23248
rect 7756 21944 7796 23920
rect 7756 21895 7796 21904
rect 7852 20852 7892 36352
rect 7852 18668 7892 20812
rect 7852 18619 7892 18628
rect 7660 17023 7700 17032
rect 7852 17072 7892 17081
rect 7468 13831 7508 13840
rect 7756 12536 7796 12545
rect 7660 9764 7700 9773
rect 7660 9260 7700 9724
rect 7660 9211 7700 9220
rect 7660 3884 7700 3893
rect 7660 3380 7700 3844
rect 7660 3331 7700 3340
rect 7372 1231 7412 1240
rect 7756 1280 7796 12496
rect 7852 8756 7892 17032
rect 7852 8707 7892 8716
rect 7948 2213 7988 61804
rect 8140 51764 8180 70624
rect 8236 60164 8276 84904
rect 12364 84524 12404 84533
rect 9676 84440 9716 84449
rect 9004 79652 9044 79661
rect 8812 76628 8852 76637
rect 8524 75956 8564 75965
rect 8428 72428 8468 72437
rect 8332 64112 8372 64121
rect 8332 63356 8372 64072
rect 8332 63307 8372 63316
rect 8236 60115 8276 60124
rect 8332 62516 8372 62525
rect 8140 51715 8180 51724
rect 8332 42533 8372 62476
rect 8331 42524 8373 42533
rect 8331 42484 8332 42524
rect 8372 42484 8373 42524
rect 8331 42475 8373 42484
rect 8428 41021 8468 72388
rect 8524 57896 8564 75916
rect 8812 74612 8852 76588
rect 8812 74563 8852 74572
rect 8908 74948 8948 74957
rect 8812 74444 8852 74453
rect 8812 72344 8852 74404
rect 8908 74360 8948 74908
rect 8908 74311 8948 74320
rect 8812 72295 8852 72304
rect 8908 72512 8948 72521
rect 8812 69320 8852 69329
rect 8620 68312 8660 68321
rect 8620 64700 8660 68272
rect 8715 67808 8757 67817
rect 8715 67768 8716 67808
rect 8756 67768 8757 67808
rect 8715 67759 8757 67768
rect 8620 60500 8660 64660
rect 8620 60451 8660 60460
rect 8427 41012 8469 41021
rect 8427 40972 8428 41012
rect 8468 40972 8469 41012
rect 8427 40963 8469 40972
rect 8140 40928 8180 40937
rect 8044 37232 8084 37241
rect 8044 18920 8084 37192
rect 8044 18871 8084 18880
rect 8044 16652 8084 16661
rect 8044 15056 8084 16612
rect 8044 15007 8084 15016
rect 7947 2204 7989 2213
rect 7947 2164 7948 2204
rect 7988 2164 7989 2204
rect 7947 2155 7989 2164
rect 8140 2204 8180 40888
rect 8428 40424 8468 40433
rect 8428 36896 8468 40384
rect 8428 36847 8468 36856
rect 8428 34796 8468 34805
rect 8332 34376 8372 34385
rect 8236 33284 8276 33293
rect 8236 29672 8276 33244
rect 8236 29623 8276 29632
rect 8332 5648 8372 34336
rect 8428 25892 8468 34756
rect 8428 21692 8468 25852
rect 8428 21643 8468 21652
rect 8332 5599 8372 5608
rect 8524 4817 8564 57856
rect 8620 41852 8660 41861
rect 8620 24548 8660 41812
rect 8716 38072 8756 67759
rect 8812 53444 8852 69280
rect 8812 53395 8852 53404
rect 8908 48824 8948 72472
rect 8908 48775 8948 48784
rect 8716 38023 8756 38032
rect 8908 43952 8948 43961
rect 8908 43280 8948 43912
rect 8812 31016 8852 31025
rect 8812 30344 8852 30976
rect 8812 30295 8852 30304
rect 8812 26816 8852 26825
rect 8620 24499 8660 24508
rect 8716 24800 8756 24809
rect 8716 23540 8756 24760
rect 8716 23288 8756 23500
rect 8716 23239 8756 23248
rect 8716 20012 8756 20021
rect 8716 17744 8756 19972
rect 8812 19676 8852 26776
rect 8812 19627 8852 19636
rect 8716 17695 8756 17704
rect 8812 19004 8852 19013
rect 8620 9680 8660 9689
rect 8620 9260 8660 9640
rect 8620 9211 8660 9220
rect 8523 4808 8565 4817
rect 8523 4768 8524 4808
rect 8564 4768 8565 4808
rect 8523 4759 8565 4768
rect 8140 2155 8180 2164
rect 7756 1231 7796 1240
rect 8812 1196 8852 18964
rect 8908 17324 8948 43240
rect 9004 34301 9044 79612
rect 9580 75620 9620 75629
rect 9196 75284 9236 75293
rect 9196 74948 9236 75244
rect 9100 72092 9140 72101
rect 9100 63944 9140 72052
rect 9196 69320 9236 74908
rect 9388 74696 9428 74705
rect 9292 74612 9332 74621
rect 9292 70664 9332 74572
rect 9292 70615 9332 70624
rect 9196 69271 9236 69280
rect 9100 63895 9140 63904
rect 9196 67136 9236 67145
rect 9196 62768 9236 67096
rect 9196 62719 9236 62728
rect 9196 57812 9236 57821
rect 9196 54872 9236 57772
rect 9196 54823 9236 54832
rect 9388 48824 9428 74656
rect 9484 65372 9524 65381
rect 9484 64700 9524 65332
rect 9484 59408 9524 64660
rect 9580 59828 9620 75580
rect 9676 69320 9716 84400
rect 10252 84440 10292 84449
rect 9676 69271 9716 69280
rect 9772 83516 9812 83525
rect 9772 69152 9812 83476
rect 10156 74780 10196 74789
rect 9964 73856 10004 73865
rect 9772 69103 9812 69112
rect 9868 71168 9908 71177
rect 9580 59779 9620 59788
rect 9676 62684 9716 62693
rect 9484 56552 9524 59368
rect 9484 56503 9524 56512
rect 9580 57980 9620 57989
rect 9388 48775 9428 48784
rect 9388 44036 9428 44045
rect 9388 43364 9428 43996
rect 9292 39584 9332 39593
rect 9100 34376 9140 34385
rect 9003 34292 9045 34301
rect 9003 34252 9004 34292
rect 9044 34252 9045 34292
rect 9003 34243 9045 34252
rect 8908 17275 8948 17284
rect 9004 31604 9044 31613
rect 9004 25304 9044 31564
rect 8908 16148 8948 16157
rect 8908 14132 8948 16108
rect 8908 14083 8948 14092
rect 8908 9092 8948 9101
rect 9004 9092 9044 25264
rect 8948 9052 9044 9092
rect 8908 4136 8948 9052
rect 9100 5732 9140 34336
rect 9196 24800 9236 24809
rect 9196 24380 9236 24760
rect 9196 21608 9236 24340
rect 9196 21559 9236 21568
rect 9196 19676 9236 19685
rect 9196 15308 9236 19636
rect 9196 15259 9236 15268
rect 9100 5683 9140 5692
rect 8908 4087 8948 4096
rect 8812 1147 8852 1156
rect 7084 895 7124 904
rect 6988 727 7028 736
rect 2092 475 2132 484
rect 9292 440 9332 39544
rect 9388 14048 9428 43324
rect 9580 40508 9620 57940
rect 9676 41777 9716 62644
rect 9772 62096 9812 62105
rect 9675 41768 9717 41777
rect 9675 41728 9676 41768
rect 9716 41728 9717 41768
rect 9675 41719 9717 41728
rect 9580 40459 9620 40468
rect 9580 34880 9620 34889
rect 9580 34712 9620 34840
rect 9484 31100 9524 31109
rect 9484 30344 9524 31060
rect 9484 30295 9524 30304
rect 9484 27068 9524 27077
rect 9484 20768 9524 27028
rect 9580 26816 9620 34672
rect 9772 30092 9812 62056
rect 9868 43280 9908 71128
rect 9964 70412 10004 73816
rect 9964 70363 10004 70372
rect 10156 69572 10196 74740
rect 10156 67724 10196 69532
rect 10156 67675 10196 67684
rect 10156 64028 10196 64037
rect 10060 63272 10100 63281
rect 9963 63020 10005 63029
rect 9963 62980 9964 63020
rect 10004 62980 10005 63020
rect 9963 62971 10005 62980
rect 9964 62886 10004 62971
rect 10060 56216 10100 63232
rect 10156 62264 10196 63988
rect 10156 62215 10196 62224
rect 10060 56167 10100 56176
rect 10156 55544 10196 55553
rect 10156 54032 10196 55504
rect 10156 53983 10196 53992
rect 9868 43231 9908 43240
rect 10060 45716 10100 45725
rect 9772 30043 9812 30052
rect 9868 40424 9908 40433
rect 9580 26767 9620 26776
rect 9676 26312 9716 26321
rect 9676 24632 9716 26272
rect 9676 24583 9716 24592
rect 9772 24800 9812 24809
rect 9772 21356 9812 24760
rect 9772 21307 9812 21316
rect 9484 14468 9524 20728
rect 9484 14419 9524 14428
rect 9388 13999 9428 14008
rect 9868 524 9908 40384
rect 9964 31268 10004 31277
rect 9964 22952 10004 31228
rect 9964 22903 10004 22912
rect 10060 19424 10100 45676
rect 10252 42524 10292 84400
rect 10444 84440 10484 84449
rect 10444 75284 10484 84400
rect 11788 84440 11828 84449
rect 11020 83516 11060 83525
rect 10828 83180 10868 83189
rect 10347 69320 10389 69329
rect 10347 69280 10348 69320
rect 10388 69280 10389 69320
rect 10347 69271 10389 69280
rect 10348 69186 10388 69271
rect 10252 42475 10292 42484
rect 10348 65960 10388 65969
rect 10252 36812 10292 36821
rect 10252 34628 10292 36772
rect 10156 34588 10252 34628
rect 10156 21524 10196 34588
rect 10252 34579 10292 34588
rect 10348 31688 10388 65920
rect 10444 40424 10484 75244
rect 10636 75620 10676 75629
rect 10636 74360 10676 75580
rect 10444 40375 10484 40384
rect 10540 70832 10580 70841
rect 10444 38744 10484 38753
rect 10444 36392 10484 38704
rect 10444 36343 10484 36352
rect 10540 33620 10580 70792
rect 10636 64280 10676 74320
rect 10731 72764 10773 72773
rect 10731 72724 10732 72764
rect 10772 72724 10773 72764
rect 10731 72715 10773 72724
rect 10732 72630 10772 72715
rect 10636 64240 10772 64280
rect 10636 64112 10676 64121
rect 10636 62432 10676 64072
rect 10636 62383 10676 62392
rect 10732 41600 10772 64240
rect 10828 61088 10868 83140
rect 11020 75200 11060 83476
rect 11692 83516 11732 83525
rect 11020 73100 11060 75160
rect 11308 75452 11348 75461
rect 11020 73060 11252 73100
rect 11020 69152 11060 69161
rect 10924 63944 10964 63953
rect 10924 62936 10964 63904
rect 10924 62887 10964 62896
rect 10828 61039 10868 61048
rect 10828 56300 10868 56309
rect 10828 54956 10868 56260
rect 10828 54907 10868 54916
rect 10732 41551 10772 41560
rect 10924 41180 10964 41189
rect 10828 36140 10868 36149
rect 10828 35468 10868 36100
rect 10828 35419 10868 35428
rect 10540 33571 10580 33580
rect 10348 31639 10388 31648
rect 10156 21475 10196 21484
rect 10252 29672 10292 29681
rect 10060 19375 10100 19384
rect 10156 20096 10196 20105
rect 10156 18248 10196 20056
rect 10156 18199 10196 18208
rect 10060 18080 10100 18089
rect 10060 17828 10100 18040
rect 10060 17779 10100 17788
rect 10156 16064 10196 16073
rect 10156 11024 10196 16024
rect 10156 10975 10196 10984
rect 10252 2456 10292 29632
rect 10732 29252 10772 29261
rect 10732 28916 10772 29212
rect 10732 28867 10772 28876
rect 10828 28244 10868 28253
rect 10828 25145 10868 28204
rect 10827 25136 10869 25145
rect 10827 25096 10828 25136
rect 10868 25096 10869 25136
rect 10827 25087 10869 25096
rect 10444 24632 10484 24641
rect 10444 24212 10484 24592
rect 10444 24163 10484 24172
rect 10348 19088 10388 19097
rect 10348 13880 10388 19048
rect 10348 13831 10388 13840
rect 10828 7916 10868 7925
rect 10828 3800 10868 7876
rect 10828 3751 10868 3760
rect 10252 2407 10292 2416
rect 10540 2708 10580 2717
rect 10540 2288 10580 2668
rect 10924 2540 10964 41140
rect 11020 15812 11060 69112
rect 11116 64448 11156 64457
rect 11116 64196 11156 64408
rect 11116 64147 11156 64156
rect 11116 63524 11156 63533
rect 11116 61088 11156 63484
rect 11116 61039 11156 61048
rect 11116 37652 11156 37661
rect 11116 37232 11156 37612
rect 11116 35048 11156 37192
rect 11116 34999 11156 35008
rect 11116 31016 11156 31025
rect 11116 27740 11156 30976
rect 11116 27691 11156 27700
rect 11212 26312 11252 73060
rect 11308 63020 11348 75412
rect 11596 71840 11636 71849
rect 11500 69824 11540 69833
rect 11308 58484 11348 62980
rect 11308 55796 11348 58444
rect 11308 55747 11348 55756
rect 11404 67472 11444 67481
rect 11308 41684 11348 41693
rect 11308 41441 11348 41644
rect 11307 41432 11349 41441
rect 11307 41392 11308 41432
rect 11348 41392 11349 41432
rect 11307 41383 11349 41392
rect 11404 31352 11444 67432
rect 11500 41264 11540 69784
rect 11596 46640 11636 71800
rect 11692 69992 11732 83476
rect 11692 69943 11732 69952
rect 11692 62180 11732 62189
rect 11692 60416 11732 62140
rect 11692 60367 11732 60376
rect 11596 46600 11732 46640
rect 11596 41600 11636 41609
rect 11596 41441 11636 41560
rect 11595 41432 11637 41441
rect 11595 41392 11596 41432
rect 11636 41392 11637 41432
rect 11595 41383 11637 41392
rect 11500 41215 11540 41224
rect 11692 38912 11732 46600
rect 11788 42785 11828 84400
rect 12172 79568 12212 79577
rect 12172 71504 12212 79528
rect 12364 71840 12404 84484
rect 12844 84524 12884 84533
rect 12748 83180 12788 83189
rect 12459 72176 12501 72185
rect 12459 72136 12460 72176
rect 12500 72136 12501 72176
rect 12459 72127 12501 72136
rect 12460 72042 12500 72127
rect 12364 71791 12404 71800
rect 11884 69908 11924 69917
rect 11787 42776 11829 42785
rect 11787 42736 11788 42776
rect 11828 42736 11829 42776
rect 11787 42727 11829 42736
rect 11884 41516 11924 69868
rect 12172 62180 12212 71464
rect 12556 69992 12596 70001
rect 12460 67136 12500 67145
rect 12172 62131 12212 62140
rect 12364 64196 12404 64205
rect 12268 61088 12308 61097
rect 12268 60164 12308 61048
rect 12268 60115 12308 60124
rect 12364 60080 12404 64156
rect 12364 60031 12404 60040
rect 12268 58484 12308 58493
rect 11884 41467 11924 41476
rect 12172 43364 12212 43373
rect 11692 38863 11732 38872
rect 11596 37820 11636 37829
rect 11636 37780 11732 37820
rect 11596 37771 11636 37780
rect 11596 37232 11636 37241
rect 11404 31303 11444 31312
rect 11500 35636 11540 35645
rect 11212 26263 11252 26272
rect 11308 29756 11348 29765
rect 11116 25472 11156 25481
rect 11116 18836 11156 25432
rect 11308 25388 11348 29716
rect 11308 25339 11348 25348
rect 11307 25136 11349 25145
rect 11307 25096 11308 25136
rect 11348 25096 11349 25136
rect 11307 25087 11349 25096
rect 11116 18787 11156 18796
rect 11212 24632 11252 24641
rect 11020 15772 11156 15812
rect 11020 13208 11060 13217
rect 11020 12620 11060 13168
rect 11020 12571 11060 12580
rect 11020 12284 11060 12293
rect 11020 8336 11060 12244
rect 11020 8287 11060 8296
rect 11020 8168 11060 8177
rect 11020 6320 11060 8128
rect 11020 6271 11060 6280
rect 11019 3464 11061 3473
rect 11019 3424 11020 3464
rect 11060 3424 11061 3464
rect 11019 3415 11061 3424
rect 11020 3330 11060 3415
rect 11116 3044 11156 15772
rect 11212 13964 11252 24592
rect 11212 12284 11252 13924
rect 11212 12235 11252 12244
rect 11212 6908 11252 6917
rect 11212 6320 11252 6868
rect 11212 6271 11252 6280
rect 11116 2995 11156 3004
rect 11308 2708 11348 25087
rect 11404 7496 11444 7505
rect 11404 6992 11444 7456
rect 11404 6943 11444 6952
rect 11308 2659 11348 2668
rect 10540 2239 10580 2248
rect 10828 2500 10964 2540
rect 9868 475 9908 484
rect 9292 391 9332 400
rect 3723 356 3765 365
rect 3723 316 3724 356
rect 3764 316 3765 356
rect 3723 307 3765 316
rect 2955 272 2997 281
rect 2955 232 2956 272
rect 2996 232 2997 272
rect 2955 223 2997 232
rect 2956 138 2996 223
rect 3724 222 3764 307
rect 10828 197 10868 2500
rect 11500 1616 11540 35596
rect 11596 31604 11636 37192
rect 11692 36644 11732 37780
rect 12076 37484 12116 37493
rect 11787 36728 11829 36737
rect 11787 36688 11788 36728
rect 11828 36688 11829 36728
rect 11787 36679 11829 36688
rect 11692 36595 11732 36604
rect 11788 35216 11828 36679
rect 11788 35167 11828 35176
rect 11980 36644 12020 36653
rect 11980 34217 12020 36604
rect 11979 34208 12021 34217
rect 11979 34168 11980 34208
rect 12020 34168 12021 34208
rect 11979 34159 12021 34168
rect 11596 31555 11636 31564
rect 11788 30764 11828 30773
rect 11596 26984 11636 26993
rect 11596 26732 11636 26944
rect 11596 26683 11636 26692
rect 11596 6656 11636 6665
rect 11596 6152 11636 6616
rect 11596 6103 11636 6112
rect 11500 1567 11540 1576
rect 5259 188 5301 197
rect 5259 148 5260 188
rect 5300 148 5301 188
rect 5259 139 5301 148
rect 10827 188 10869 197
rect 10827 148 10828 188
rect 10868 148 10869 188
rect 10827 139 10869 148
rect 5260 54 5300 139
rect 11788 104 11828 30724
rect 11884 24212 11924 24221
rect 11884 20012 11924 24172
rect 11884 19963 11924 19972
rect 11980 365 12020 34159
rect 12076 33284 12116 37444
rect 12076 33235 12116 33244
rect 12075 26480 12117 26489
rect 12075 26440 12076 26480
rect 12116 26440 12117 26480
rect 12075 26431 12117 26440
rect 12076 2624 12116 26431
rect 12172 22028 12212 43324
rect 12268 35636 12308 58444
rect 12460 37820 12500 67096
rect 12364 37780 12500 37820
rect 12364 37493 12404 37780
rect 12363 37484 12405 37493
rect 12363 37444 12364 37484
rect 12404 37444 12405 37484
rect 12363 37435 12405 37444
rect 12268 35587 12308 35596
rect 12172 21979 12212 21988
rect 12268 31352 12308 31361
rect 12172 20768 12212 20777
rect 12172 20012 12212 20728
rect 12172 19963 12212 19972
rect 12172 18668 12212 18677
rect 12172 6236 12212 18628
rect 12172 6187 12212 6196
rect 12076 2575 12116 2584
rect 12268 1868 12308 31312
rect 12363 30680 12405 30689
rect 12363 30640 12364 30680
rect 12404 30640 12405 30680
rect 12363 30631 12405 30640
rect 12364 30546 12404 30631
rect 12460 27908 12500 27917
rect 12460 26984 12500 27868
rect 12460 26935 12500 26944
rect 12460 26816 12500 26825
rect 12363 26312 12405 26321
rect 12363 26272 12364 26312
rect 12404 26272 12405 26312
rect 12363 26263 12405 26272
rect 12364 24380 12404 26263
rect 12460 25136 12500 26776
rect 12460 25087 12500 25096
rect 12364 24331 12404 24340
rect 12460 24128 12500 24137
rect 12364 23624 12404 23633
rect 12364 7001 12404 23584
rect 12460 22364 12500 24088
rect 12460 22315 12500 22324
rect 12556 19844 12596 69952
rect 12652 66632 12692 66641
rect 12652 63440 12692 66592
rect 12652 63391 12692 63400
rect 12652 59408 12692 59417
rect 12652 51260 12692 59368
rect 12652 51211 12692 51220
rect 12651 34208 12693 34217
rect 12651 34168 12652 34208
rect 12692 34168 12693 34208
rect 12651 34159 12693 34168
rect 12652 34074 12692 34159
rect 12652 23960 12692 23969
rect 12652 21020 12692 23920
rect 12652 20971 12692 20980
rect 12556 19795 12596 19804
rect 12363 6992 12405 7001
rect 12363 6952 12364 6992
rect 12404 6952 12405 6992
rect 12363 6943 12405 6952
rect 12268 1819 12308 1828
rect 12748 1280 12788 83140
rect 12844 16232 12884 84484
rect 12940 84440 12980 84449
rect 12940 57308 12980 84400
rect 13324 84440 13364 84449
rect 13131 83348 13173 83357
rect 13131 83308 13132 83348
rect 13172 83308 13173 83348
rect 13131 83299 13173 83308
rect 13132 83214 13172 83299
rect 13228 67640 13268 67649
rect 13132 66548 13172 66557
rect 13036 66464 13076 66473
rect 13036 64028 13076 66424
rect 13132 64868 13172 66508
rect 13132 64819 13172 64828
rect 13228 64280 13268 67600
rect 13036 63979 13076 63988
rect 13132 64240 13268 64280
rect 13035 61340 13077 61349
rect 13035 61300 13036 61340
rect 13076 61300 13077 61340
rect 13035 61291 13077 61300
rect 13036 61206 13076 61291
rect 13036 61088 13076 61097
rect 13036 57644 13076 61048
rect 13036 57595 13076 57604
rect 12940 57259 12980 57268
rect 13132 50420 13172 64240
rect 13132 48824 13172 50380
rect 13132 48775 13172 48784
rect 13228 60332 13268 60341
rect 13036 47396 13076 47405
rect 13036 46472 13076 47356
rect 12939 36728 12981 36737
rect 12939 36688 12940 36728
rect 12980 36688 12981 36728
rect 12939 36679 12981 36688
rect 12940 36594 12980 36679
rect 12844 15476 12884 16192
rect 12844 15427 12884 15436
rect 12940 26648 12980 26657
rect 12940 1868 12980 26608
rect 13036 14636 13076 46432
rect 13228 41432 13268 60292
rect 13228 41383 13268 41392
rect 13228 36896 13268 36905
rect 13132 34628 13172 34637
rect 13132 29672 13172 34588
rect 13228 32696 13268 36856
rect 13228 32647 13268 32656
rect 13132 29623 13172 29632
rect 13324 28496 13364 84400
rect 14092 84440 14132 84449
rect 13996 83348 14036 83357
rect 13900 81836 13940 81845
rect 13804 72008 13844 72017
rect 13708 71968 13804 72008
rect 13612 69320 13652 69329
rect 13516 67220 13556 67229
rect 13420 65792 13460 65801
rect 13420 64280 13460 65752
rect 13420 64231 13460 64240
rect 13516 62600 13556 67180
rect 13612 65876 13652 69280
rect 13612 65827 13652 65836
rect 13516 62551 13556 62560
rect 13612 64448 13652 64457
rect 13420 60836 13460 60845
rect 13420 59408 13460 60796
rect 13420 59359 13460 59368
rect 13420 58820 13460 58829
rect 13420 56804 13460 58780
rect 13420 56755 13460 56764
rect 13516 51260 13556 51269
rect 13516 46892 13556 51220
rect 13516 46843 13556 46852
rect 13612 39584 13652 64408
rect 13708 64280 13748 71968
rect 13804 71959 13844 71968
rect 13803 66380 13845 66389
rect 13803 66340 13804 66380
rect 13844 66340 13845 66380
rect 13803 66331 13845 66340
rect 13804 66246 13844 66331
rect 13708 64240 13844 64280
rect 13708 57056 13748 57065
rect 13708 49580 13748 57016
rect 13708 49531 13748 49540
rect 13612 39535 13652 39544
rect 13708 48656 13748 48665
rect 13420 38912 13460 38921
rect 13420 35300 13460 38872
rect 13612 37736 13652 37745
rect 13612 36476 13652 37696
rect 13420 35251 13460 35260
rect 13516 35720 13556 35729
rect 13324 28447 13364 28456
rect 13516 28244 13556 35680
rect 13612 34040 13652 36436
rect 13612 33991 13652 34000
rect 13516 28195 13556 28204
rect 13036 14587 13076 14596
rect 13324 22280 13364 22289
rect 13132 13880 13172 13889
rect 13132 12620 13172 13840
rect 13132 11696 13172 12580
rect 13132 11647 13172 11656
rect 13036 8672 13076 8681
rect 13036 7580 13076 8632
rect 13036 4976 13076 7540
rect 13036 4927 13076 4936
rect 13324 3968 13364 22240
rect 13324 3919 13364 3928
rect 12940 1819 12980 1828
rect 12748 1231 12788 1240
rect 12555 1112 12597 1121
rect 12555 1072 12556 1112
rect 12596 1072 12597 1112
rect 12555 1063 12597 1072
rect 12556 978 12596 1063
rect 11979 356 12021 365
rect 11979 316 11980 356
rect 12020 316 12021 356
rect 11979 307 12021 316
rect 13708 188 13748 48616
rect 13804 42104 13844 64240
rect 13804 42055 13844 42064
rect 13804 35132 13844 35141
rect 13804 34628 13844 35092
rect 13804 34579 13844 34588
rect 13804 27236 13844 27245
rect 13804 18836 13844 27196
rect 13804 18787 13844 18796
rect 13900 1280 13940 81796
rect 13996 4556 14036 83308
rect 14092 38660 14132 84400
rect 14476 83348 14516 83357
rect 14092 38611 14132 38620
rect 14188 82592 14228 82601
rect 14091 23792 14133 23801
rect 14091 23752 14092 23792
rect 14132 23752 14133 23792
rect 14091 23743 14133 23752
rect 14092 23658 14132 23743
rect 14091 17660 14133 17669
rect 14091 17620 14092 17660
rect 14132 17620 14133 17660
rect 14091 17611 14133 17620
rect 13996 4507 14036 4516
rect 14092 1868 14132 17611
rect 14092 1819 14132 1828
rect 13900 1231 13940 1240
rect 14188 692 14228 82552
rect 14380 65960 14420 65969
rect 14284 54872 14324 54881
rect 14284 53192 14324 54832
rect 14284 53143 14324 53152
rect 14380 31436 14420 65920
rect 14380 31387 14420 31396
rect 14380 11192 14420 11201
rect 14380 9932 14420 11152
rect 14380 9883 14420 9892
rect 14283 6992 14325 7001
rect 14283 6952 14284 6992
rect 14324 6952 14325 6992
rect 14283 6943 14325 6952
rect 14284 1868 14324 6943
rect 14476 4472 14516 83308
rect 14668 83348 14708 83357
rect 14571 26060 14613 26069
rect 14571 26020 14572 26060
rect 14612 26020 14613 26060
rect 14571 26011 14613 26020
rect 14572 25926 14612 26011
rect 14476 4423 14516 4432
rect 14284 1819 14324 1828
rect 14668 1616 14708 83308
rect 15052 83348 15092 83357
rect 14956 70244 14996 70253
rect 14956 42188 14996 70204
rect 14956 42139 14996 42148
rect 14764 19088 14804 19097
rect 14764 17072 14804 19048
rect 14764 7328 14804 17032
rect 14764 7279 14804 7288
rect 14668 1567 14708 1576
rect 15052 860 15092 83308
rect 15244 72092 15284 72101
rect 15148 67892 15188 67901
rect 15148 24800 15188 67852
rect 15244 29336 15284 72052
rect 15628 70832 15668 70841
rect 15628 70328 15668 70792
rect 15628 70279 15668 70288
rect 15340 67556 15380 67565
rect 15340 58913 15380 67516
rect 15436 64280 15476 64289
rect 15339 58904 15381 58913
rect 15339 58864 15340 58904
rect 15380 58864 15381 58904
rect 15339 58855 15381 58864
rect 15340 58736 15380 58745
rect 15340 57392 15380 58696
rect 15340 57343 15380 57352
rect 15340 31520 15380 31529
rect 15340 30092 15380 31480
rect 15436 31268 15476 64240
rect 15532 61844 15572 61853
rect 15532 61172 15572 61804
rect 15532 61123 15572 61132
rect 15436 31219 15476 31228
rect 15532 60668 15572 60677
rect 15340 30043 15380 30052
rect 15244 29287 15284 29296
rect 15148 24751 15188 24760
rect 15436 24632 15476 24641
rect 15436 23036 15476 24592
rect 15436 22987 15476 22996
rect 15436 18836 15476 18845
rect 15436 17240 15476 18796
rect 15436 17191 15476 17200
rect 15244 12620 15284 12629
rect 15244 1868 15284 12580
rect 15244 1819 15284 1828
rect 15532 1868 15572 60628
rect 15532 1819 15572 1828
rect 15628 59408 15668 59417
rect 15628 1280 15668 59368
rect 15724 42860 15764 85576
rect 15916 84944 15956 84953
rect 15820 71252 15860 71261
rect 15820 70412 15860 71212
rect 15820 70363 15860 70372
rect 15916 65456 15956 84904
rect 18808 84692 19176 84701
rect 18848 84652 18890 84692
rect 18930 84652 18972 84692
rect 19012 84652 19054 84692
rect 19094 84652 19136 84692
rect 18808 84643 19176 84652
rect 16396 84440 16436 84449
rect 16300 73856 16340 73865
rect 16012 71000 16052 71009
rect 16012 69656 16052 70960
rect 16012 69607 16052 69616
rect 16012 69488 16052 69497
rect 16012 66128 16052 69448
rect 16012 66079 16052 66088
rect 16108 66464 16148 66473
rect 15916 65407 15956 65416
rect 15916 61676 15956 61685
rect 15916 53696 15956 61636
rect 16011 61340 16053 61349
rect 16011 61300 16012 61340
rect 16052 61300 16053 61340
rect 16011 61291 16053 61300
rect 16012 61206 16052 61291
rect 16011 58904 16053 58913
rect 16011 58864 16012 58904
rect 16052 58864 16053 58904
rect 16011 58855 16053 58864
rect 16012 56468 16052 58855
rect 16012 56419 16052 56428
rect 15916 53647 15956 53656
rect 15724 42811 15764 42820
rect 16108 37652 16148 66424
rect 16108 37603 16148 37612
rect 16204 44372 16244 44381
rect 15724 32360 15764 32369
rect 15724 30428 15764 32320
rect 15724 15560 15764 30388
rect 16012 27740 16052 27749
rect 15724 9596 15764 15520
rect 15820 27572 15860 27581
rect 15820 22868 15860 27532
rect 15820 13292 15860 22828
rect 15820 11864 15860 13252
rect 15820 11815 15860 11824
rect 15724 9547 15764 9556
rect 16012 1868 16052 27700
rect 16204 12704 16244 44332
rect 16300 40685 16340 73816
rect 16396 57308 16436 84400
rect 16876 84440 16916 84449
rect 16780 69488 16820 69497
rect 16396 57259 16436 57268
rect 16588 59492 16628 59501
rect 16588 55040 16628 59452
rect 16588 54991 16628 55000
rect 16396 45548 16436 45557
rect 16396 44540 16436 45508
rect 16396 44491 16436 44500
rect 16396 42860 16436 42869
rect 16299 40676 16341 40685
rect 16299 40636 16300 40676
rect 16340 40636 16341 40676
rect 16299 40627 16341 40636
rect 16204 12655 16244 12664
rect 16396 11780 16436 42820
rect 16588 40004 16628 40013
rect 16492 17408 16532 17417
rect 16492 14216 16532 17368
rect 16492 14167 16532 14176
rect 16396 11731 16436 11740
rect 16108 8000 16148 8009
rect 16108 5480 16148 7960
rect 16108 5431 16148 5440
rect 16588 2036 16628 39964
rect 16684 31436 16724 31445
rect 16684 29681 16724 31396
rect 16683 29672 16725 29681
rect 16683 29632 16684 29672
rect 16724 29632 16725 29672
rect 16683 29623 16725 29632
rect 16684 18164 16724 18173
rect 16684 16904 16724 18124
rect 16684 16855 16724 16864
rect 16588 1987 16628 1996
rect 16012 1819 16052 1828
rect 15628 1231 15668 1240
rect 16780 1196 16820 69448
rect 16876 56552 16916 84400
rect 20048 83936 20416 83945
rect 20088 83896 20130 83936
rect 20170 83896 20212 83936
rect 20252 83896 20294 83936
rect 20334 83896 20376 83936
rect 20048 83887 20416 83896
rect 18316 83516 18356 83525
rect 17356 82592 17396 82601
rect 17164 68396 17204 68405
rect 16876 56503 16916 56512
rect 16972 63692 17012 63701
rect 16876 40256 16916 40265
rect 16876 2120 16916 40216
rect 16972 32192 17012 63652
rect 17068 47228 17108 47237
rect 17068 44288 17108 47188
rect 17068 44239 17108 44248
rect 17164 40676 17204 68356
rect 17164 40627 17204 40636
rect 17260 57728 17300 57737
rect 17260 34628 17300 57688
rect 17260 34579 17300 34588
rect 16972 32143 17012 32152
rect 17068 29336 17108 29345
rect 17068 28916 17108 29296
rect 17068 28867 17108 28876
rect 16972 24632 17012 24641
rect 16972 18584 17012 24592
rect 16972 18535 17012 18544
rect 16876 2071 16916 2080
rect 17356 1280 17396 82552
rect 17740 82592 17780 82601
rect 17548 66800 17588 66809
rect 17452 65624 17492 65633
rect 17452 36812 17492 65584
rect 17548 62096 17588 66760
rect 17548 62047 17588 62056
rect 17644 65540 17684 65549
rect 17548 59156 17588 59165
rect 17548 56384 17588 59116
rect 17548 56335 17588 56344
rect 17548 52856 17588 52865
rect 17548 49748 17588 52816
rect 17548 49699 17588 49708
rect 17644 42860 17684 65500
rect 17644 42811 17684 42820
rect 17452 36763 17492 36772
rect 17452 29084 17492 29093
rect 17452 18668 17492 29044
rect 17644 26144 17684 26153
rect 17644 25229 17684 26104
rect 17643 25220 17685 25229
rect 17643 25180 17644 25220
rect 17684 25180 17685 25220
rect 17643 25171 17685 25180
rect 17452 18619 17492 18628
rect 17356 1231 17396 1240
rect 17740 1280 17780 82552
rect 18124 81920 18164 81929
rect 17740 1231 17780 1240
rect 17932 50420 17972 50429
rect 16780 1147 16820 1156
rect 15052 811 15092 820
rect 14188 643 14228 652
rect 17932 608 17972 50380
rect 18028 35552 18068 35561
rect 18028 20096 18068 35512
rect 18028 20047 18068 20056
rect 18124 1280 18164 81880
rect 18316 52856 18356 83476
rect 18604 83516 18644 83525
rect 18316 52807 18356 52816
rect 18412 82004 18452 82013
rect 18316 50504 18356 50513
rect 18316 46724 18356 50464
rect 18316 46472 18356 46684
rect 18316 46423 18356 46432
rect 18412 39080 18452 81964
rect 18412 39031 18452 39040
rect 18508 81920 18548 81929
rect 18412 21104 18452 21113
rect 18412 20432 18452 21064
rect 18412 20383 18452 20392
rect 18315 6320 18357 6329
rect 18315 6280 18316 6320
rect 18356 6280 18357 6320
rect 18315 6271 18357 6280
rect 18124 1231 18164 1240
rect 18316 944 18356 6271
rect 18508 1280 18548 81880
rect 18604 36560 18644 83476
rect 19083 83516 19125 83525
rect 19083 83476 19084 83516
rect 19124 83476 19125 83516
rect 19083 83467 19125 83476
rect 19564 83516 19604 83525
rect 19084 83382 19124 83467
rect 18808 83180 19176 83189
rect 18848 83140 18890 83180
rect 18930 83140 18972 83180
rect 19012 83140 19054 83180
rect 19094 83140 19136 83180
rect 18808 83131 19176 83140
rect 19468 82592 19508 82601
rect 19276 81920 19316 81929
rect 18808 81668 19176 81677
rect 18848 81628 18890 81668
rect 18930 81628 18972 81668
rect 19012 81628 19054 81668
rect 19094 81628 19136 81668
rect 18808 81619 19176 81628
rect 18808 80156 19176 80165
rect 18848 80116 18890 80156
rect 18930 80116 18972 80156
rect 19012 80116 19054 80156
rect 19094 80116 19136 80156
rect 18808 80107 19176 80116
rect 18808 78644 19176 78653
rect 18848 78604 18890 78644
rect 18930 78604 18972 78644
rect 19012 78604 19054 78644
rect 19094 78604 19136 78644
rect 18808 78595 19176 78604
rect 18808 77132 19176 77141
rect 18848 77092 18890 77132
rect 18930 77092 18972 77132
rect 19012 77092 19054 77132
rect 19094 77092 19136 77132
rect 18808 77083 19176 77092
rect 18808 75620 19176 75629
rect 18848 75580 18890 75620
rect 18930 75580 18972 75620
rect 19012 75580 19054 75620
rect 19094 75580 19136 75620
rect 18808 75571 19176 75580
rect 18808 74108 19176 74117
rect 18848 74068 18890 74108
rect 18930 74068 18972 74108
rect 19012 74068 19054 74108
rect 19094 74068 19136 74108
rect 18808 74059 19176 74068
rect 18808 72596 19176 72605
rect 18848 72556 18890 72596
rect 18930 72556 18972 72596
rect 19012 72556 19054 72596
rect 19094 72556 19136 72596
rect 18808 72547 19176 72556
rect 18808 71084 19176 71093
rect 18848 71044 18890 71084
rect 18930 71044 18972 71084
rect 19012 71044 19054 71084
rect 19094 71044 19136 71084
rect 18808 71035 19176 71044
rect 18808 69572 19176 69581
rect 18848 69532 18890 69572
rect 18930 69532 18972 69572
rect 19012 69532 19054 69572
rect 19094 69532 19136 69572
rect 18808 69523 19176 69532
rect 18808 68060 19176 68069
rect 18848 68020 18890 68060
rect 18930 68020 18972 68060
rect 19012 68020 19054 68060
rect 19094 68020 19136 68060
rect 18808 68011 19176 68020
rect 18808 66548 19176 66557
rect 18848 66508 18890 66548
rect 18930 66508 18972 66548
rect 19012 66508 19054 66548
rect 19094 66508 19136 66548
rect 18808 66499 19176 66508
rect 18808 65036 19176 65045
rect 18848 64996 18890 65036
rect 18930 64996 18972 65036
rect 19012 64996 19054 65036
rect 19094 64996 19136 65036
rect 18808 64987 19176 64996
rect 18808 63524 19176 63533
rect 18848 63484 18890 63524
rect 18930 63484 18972 63524
rect 19012 63484 19054 63524
rect 19094 63484 19136 63524
rect 18808 63475 19176 63484
rect 18808 62012 19176 62021
rect 18848 61972 18890 62012
rect 18930 61972 18972 62012
rect 19012 61972 19054 62012
rect 19094 61972 19136 62012
rect 18808 61963 19176 61972
rect 18808 60500 19176 60509
rect 18848 60460 18890 60500
rect 18930 60460 18972 60500
rect 19012 60460 19054 60500
rect 19094 60460 19136 60500
rect 18808 60451 19176 60460
rect 18808 58988 19176 58997
rect 18848 58948 18890 58988
rect 18930 58948 18972 58988
rect 19012 58948 19054 58988
rect 19094 58948 19136 58988
rect 18808 58939 19176 58948
rect 18808 57476 19176 57485
rect 18848 57436 18890 57476
rect 18930 57436 18972 57476
rect 19012 57436 19054 57476
rect 19094 57436 19136 57476
rect 18808 57427 19176 57436
rect 18700 56804 18740 56813
rect 18700 42188 18740 56764
rect 18808 55964 19176 55973
rect 18848 55924 18890 55964
rect 18930 55924 18972 55964
rect 19012 55924 19054 55964
rect 19094 55924 19136 55964
rect 18808 55915 19176 55924
rect 18808 54452 19176 54461
rect 18848 54412 18890 54452
rect 18930 54412 18972 54452
rect 19012 54412 19054 54452
rect 19094 54412 19136 54452
rect 18808 54403 19176 54412
rect 18808 52940 19176 52949
rect 18848 52900 18890 52940
rect 18930 52900 18972 52940
rect 19012 52900 19054 52940
rect 19094 52900 19136 52940
rect 18808 52891 19176 52900
rect 18808 51428 19176 51437
rect 18848 51388 18890 51428
rect 18930 51388 18972 51428
rect 19012 51388 19054 51428
rect 19094 51388 19136 51428
rect 18808 51379 19176 51388
rect 18808 49916 19176 49925
rect 18848 49876 18890 49916
rect 18930 49876 18972 49916
rect 19012 49876 19054 49916
rect 19094 49876 19136 49916
rect 18808 49867 19176 49876
rect 18808 48404 19176 48413
rect 18848 48364 18890 48404
rect 18930 48364 18972 48404
rect 19012 48364 19054 48404
rect 19094 48364 19136 48404
rect 18808 48355 19176 48364
rect 18808 46892 19176 46901
rect 18848 46852 18890 46892
rect 18930 46852 18972 46892
rect 19012 46852 19054 46892
rect 19094 46852 19136 46892
rect 18808 46843 19176 46852
rect 18808 45380 19176 45389
rect 18848 45340 18890 45380
rect 18930 45340 18972 45380
rect 19012 45340 19054 45380
rect 19094 45340 19136 45380
rect 18808 45331 19176 45340
rect 18808 43868 19176 43877
rect 18848 43828 18890 43868
rect 18930 43828 18972 43868
rect 19012 43828 19054 43868
rect 19094 43828 19136 43868
rect 18808 43819 19176 43828
rect 18796 42533 18836 42618
rect 18795 42524 18837 42533
rect 18795 42484 18796 42524
rect 18836 42484 18837 42524
rect 18795 42475 18837 42484
rect 18808 42356 19176 42365
rect 18848 42316 18890 42356
rect 18930 42316 18972 42356
rect 19012 42316 19054 42356
rect 19094 42316 19136 42356
rect 18808 42307 19176 42316
rect 18700 42139 18740 42148
rect 18808 40844 19176 40853
rect 18848 40804 18890 40844
rect 18930 40804 18972 40844
rect 19012 40804 19054 40844
rect 19094 40804 19136 40844
rect 18808 40795 19176 40804
rect 18808 39332 19176 39341
rect 18848 39292 18890 39332
rect 18930 39292 18972 39332
rect 19012 39292 19054 39332
rect 19094 39292 19136 39332
rect 18808 39283 19176 39292
rect 18808 37820 19176 37829
rect 18848 37780 18890 37820
rect 18930 37780 18972 37820
rect 19012 37780 19054 37820
rect 19094 37780 19136 37820
rect 18808 37771 19176 37780
rect 18604 36511 18644 36520
rect 18808 36308 19176 36317
rect 18848 36268 18890 36308
rect 18930 36268 18972 36308
rect 19012 36268 19054 36308
rect 19094 36268 19136 36308
rect 18808 36259 19176 36268
rect 18808 34796 19176 34805
rect 18848 34756 18890 34796
rect 18930 34756 18972 34796
rect 19012 34756 19054 34796
rect 19094 34756 19136 34796
rect 18808 34747 19176 34756
rect 18808 33284 19176 33293
rect 18848 33244 18890 33284
rect 18930 33244 18972 33284
rect 19012 33244 19054 33284
rect 19094 33244 19136 33284
rect 18808 33235 19176 33244
rect 18808 31772 19176 31781
rect 18848 31732 18890 31772
rect 18930 31732 18972 31772
rect 19012 31732 19054 31772
rect 19094 31732 19136 31772
rect 18808 31723 19176 31732
rect 18700 31016 18740 31025
rect 18700 27992 18740 30976
rect 18808 30260 19176 30269
rect 18848 30220 18890 30260
rect 18930 30220 18972 30260
rect 19012 30220 19054 30260
rect 19094 30220 19136 30260
rect 18808 30211 19176 30220
rect 18808 28748 19176 28757
rect 18848 28708 18890 28748
rect 18930 28708 18972 28748
rect 19012 28708 19054 28748
rect 19094 28708 19136 28748
rect 18808 28699 19176 28708
rect 18700 27943 18740 27952
rect 18808 27236 19176 27245
rect 18848 27196 18890 27236
rect 18930 27196 18972 27236
rect 19012 27196 19054 27236
rect 19094 27196 19136 27236
rect 18808 27187 19176 27196
rect 18808 25724 19176 25733
rect 18848 25684 18890 25724
rect 18930 25684 18972 25724
rect 19012 25684 19054 25724
rect 19094 25684 19136 25724
rect 18808 25675 19176 25684
rect 18808 24212 19176 24221
rect 18848 24172 18890 24212
rect 18930 24172 18972 24212
rect 19012 24172 19054 24212
rect 19094 24172 19136 24212
rect 18808 24163 19176 24172
rect 18808 22700 19176 22709
rect 18848 22660 18890 22700
rect 18930 22660 18972 22700
rect 19012 22660 19054 22700
rect 19094 22660 19136 22700
rect 18808 22651 19176 22660
rect 18808 21188 19176 21197
rect 18848 21148 18890 21188
rect 18930 21148 18972 21188
rect 19012 21148 19054 21188
rect 19094 21148 19136 21188
rect 18808 21139 19176 21148
rect 18808 19676 19176 19685
rect 18848 19636 18890 19676
rect 18930 19636 18972 19676
rect 19012 19636 19054 19676
rect 19094 19636 19136 19676
rect 18808 19627 19176 19636
rect 18808 18164 19176 18173
rect 18848 18124 18890 18164
rect 18930 18124 18972 18164
rect 19012 18124 19054 18164
rect 19094 18124 19136 18164
rect 18808 18115 19176 18124
rect 18808 16652 19176 16661
rect 18848 16612 18890 16652
rect 18930 16612 18972 16652
rect 19012 16612 19054 16652
rect 19094 16612 19136 16652
rect 18808 16603 19176 16612
rect 18808 15140 19176 15149
rect 18848 15100 18890 15140
rect 18930 15100 18972 15140
rect 19012 15100 19054 15140
rect 19094 15100 19136 15140
rect 18808 15091 19176 15100
rect 18808 13628 19176 13637
rect 18848 13588 18890 13628
rect 18930 13588 18972 13628
rect 19012 13588 19054 13628
rect 19094 13588 19136 13628
rect 18808 13579 19176 13588
rect 18808 12116 19176 12125
rect 18848 12076 18890 12116
rect 18930 12076 18972 12116
rect 19012 12076 19054 12116
rect 19094 12076 19136 12116
rect 18808 12067 19176 12076
rect 18808 10604 19176 10613
rect 18848 10564 18890 10604
rect 18930 10564 18972 10604
rect 19012 10564 19054 10604
rect 19094 10564 19136 10604
rect 18808 10555 19176 10564
rect 18808 9092 19176 9101
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 18808 9043 19176 9052
rect 18808 7580 19176 7589
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 18808 7531 19176 7540
rect 18808 6068 19176 6077
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 18808 6019 19176 6028
rect 18808 4556 19176 4565
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 18808 4507 19176 4516
rect 18808 3044 19176 3053
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 18808 2995 19176 3004
rect 18808 1532 19176 1541
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 18808 1483 19176 1492
rect 18508 1231 18548 1240
rect 19276 1280 19316 81880
rect 19372 71504 19412 71513
rect 19372 69236 19412 71464
rect 19372 69187 19412 69196
rect 19468 46640 19508 82552
rect 19564 63020 19604 83476
rect 20048 82424 20416 82433
rect 20088 82384 20130 82424
rect 20170 82384 20212 82424
rect 20252 82384 20294 82424
rect 20334 82384 20376 82424
rect 20048 82375 20416 82384
rect 20048 80912 20416 80921
rect 20088 80872 20130 80912
rect 20170 80872 20212 80912
rect 20252 80872 20294 80912
rect 20334 80872 20376 80912
rect 20048 80863 20416 80872
rect 20048 79400 20416 79409
rect 20088 79360 20130 79400
rect 20170 79360 20212 79400
rect 20252 79360 20294 79400
rect 20334 79360 20376 79400
rect 20048 79351 20416 79360
rect 20048 77888 20416 77897
rect 20088 77848 20130 77888
rect 20170 77848 20212 77888
rect 20252 77848 20294 77888
rect 20334 77848 20376 77888
rect 20048 77839 20416 77848
rect 21196 77888 21236 77897
rect 20048 76376 20416 76385
rect 20088 76336 20130 76376
rect 20170 76336 20212 76376
rect 20252 76336 20294 76376
rect 20334 76336 20376 76376
rect 20048 76327 20416 76336
rect 20048 74864 20416 74873
rect 20088 74824 20130 74864
rect 20170 74824 20212 74864
rect 20252 74824 20294 74864
rect 20334 74824 20376 74864
rect 20048 74815 20416 74824
rect 20048 73352 20416 73361
rect 20088 73312 20130 73352
rect 20170 73312 20212 73352
rect 20252 73312 20294 73352
rect 20334 73312 20376 73352
rect 20048 73303 20416 73312
rect 20048 71840 20416 71849
rect 20088 71800 20130 71840
rect 20170 71800 20212 71840
rect 20252 71800 20294 71840
rect 20334 71800 20376 71840
rect 20048 71791 20416 71800
rect 20048 70328 20416 70337
rect 20088 70288 20130 70328
rect 20170 70288 20212 70328
rect 20252 70288 20294 70328
rect 20334 70288 20376 70328
rect 20048 70279 20416 70288
rect 19564 62971 19604 62980
rect 19660 70160 19700 70169
rect 19660 46640 19700 70120
rect 20048 68816 20416 68825
rect 20088 68776 20130 68816
rect 20170 68776 20212 68816
rect 20252 68776 20294 68816
rect 20334 68776 20376 68816
rect 20048 68767 20416 68776
rect 20139 67808 20181 67817
rect 20139 67768 20140 67808
rect 20180 67768 20181 67808
rect 20139 67759 20181 67768
rect 20140 67674 20180 67759
rect 20048 67304 20416 67313
rect 20088 67264 20130 67304
rect 20170 67264 20212 67304
rect 20252 67264 20294 67304
rect 20334 67264 20376 67304
rect 20048 67255 20416 67264
rect 19948 66800 19988 66809
rect 19372 46600 19508 46640
rect 19564 46600 19700 46640
rect 19852 63440 19892 63449
rect 19372 37820 19412 46600
rect 19467 41012 19509 41021
rect 19467 40972 19468 41012
rect 19508 40972 19509 41012
rect 19467 40963 19509 40972
rect 19468 40878 19508 40963
rect 19467 40676 19509 40685
rect 19467 40636 19468 40676
rect 19508 40636 19509 40676
rect 19467 40627 19509 40636
rect 19468 40542 19508 40627
rect 19564 37820 19604 46600
rect 19659 41768 19701 41777
rect 19659 41728 19660 41768
rect 19700 41728 19701 41768
rect 19659 41719 19701 41728
rect 19660 41634 19700 41719
rect 19852 41432 19892 63400
rect 19852 41383 19892 41392
rect 19756 41096 19796 41105
rect 19372 37780 19508 37820
rect 19564 37780 19700 37820
rect 19372 34040 19412 34049
rect 19372 32864 19412 34000
rect 19372 21608 19412 32824
rect 19372 21559 19412 21568
rect 19276 1231 19316 1240
rect 19468 1280 19508 37780
rect 19563 37484 19605 37493
rect 19563 37444 19564 37484
rect 19604 37444 19605 37484
rect 19563 37435 19605 37444
rect 19564 37350 19604 37435
rect 19564 28496 19604 28505
rect 19564 26480 19604 28456
rect 19564 26431 19604 26440
rect 19468 1231 19508 1240
rect 19660 1196 19700 37780
rect 19756 29000 19796 41056
rect 19948 32864 19988 66760
rect 20048 65792 20416 65801
rect 20088 65752 20130 65792
rect 20170 65752 20212 65792
rect 20252 65752 20294 65792
rect 20334 65752 20376 65792
rect 20048 65743 20416 65752
rect 20048 64280 20416 64289
rect 20088 64240 20130 64280
rect 20170 64240 20212 64280
rect 20252 64240 20294 64280
rect 20334 64240 20376 64280
rect 20048 64231 20416 64240
rect 20048 62768 20416 62777
rect 20088 62728 20130 62768
rect 20170 62728 20212 62768
rect 20252 62728 20294 62768
rect 20334 62728 20376 62768
rect 20048 62719 20416 62728
rect 20048 61256 20416 61265
rect 20088 61216 20130 61256
rect 20170 61216 20212 61256
rect 20252 61216 20294 61256
rect 20334 61216 20376 61256
rect 20048 61207 20416 61216
rect 21004 60416 21044 60425
rect 20048 59744 20416 59753
rect 20088 59704 20130 59744
rect 20170 59704 20212 59744
rect 20252 59704 20294 59744
rect 20334 59704 20376 59744
rect 20048 59695 20416 59704
rect 20048 58232 20416 58241
rect 20088 58192 20130 58232
rect 20170 58192 20212 58232
rect 20252 58192 20294 58232
rect 20334 58192 20376 58232
rect 20048 58183 20416 58192
rect 20048 56720 20416 56729
rect 20088 56680 20130 56720
rect 20170 56680 20212 56720
rect 20252 56680 20294 56720
rect 20334 56680 20376 56720
rect 20048 56671 20416 56680
rect 20048 55208 20416 55217
rect 20088 55168 20130 55208
rect 20170 55168 20212 55208
rect 20252 55168 20294 55208
rect 20334 55168 20376 55208
rect 20048 55159 20416 55168
rect 20048 53696 20416 53705
rect 20088 53656 20130 53696
rect 20170 53656 20212 53696
rect 20252 53656 20294 53696
rect 20334 53656 20376 53696
rect 20048 53647 20416 53656
rect 20620 52856 20660 52865
rect 20048 52184 20416 52193
rect 20088 52144 20130 52184
rect 20170 52144 20212 52184
rect 20252 52144 20294 52184
rect 20334 52144 20376 52184
rect 20048 52135 20416 52144
rect 20048 50672 20416 50681
rect 20088 50632 20130 50672
rect 20170 50632 20212 50672
rect 20252 50632 20294 50672
rect 20334 50632 20376 50672
rect 20048 50623 20416 50632
rect 20048 49160 20416 49169
rect 20088 49120 20130 49160
rect 20170 49120 20212 49160
rect 20252 49120 20294 49160
rect 20334 49120 20376 49160
rect 20048 49111 20416 49120
rect 20048 47648 20416 47657
rect 20088 47608 20130 47648
rect 20170 47608 20212 47648
rect 20252 47608 20294 47648
rect 20334 47608 20376 47648
rect 20048 47599 20416 47608
rect 20048 46136 20416 46145
rect 20088 46096 20130 46136
rect 20170 46096 20212 46136
rect 20252 46096 20294 46136
rect 20334 46096 20376 46136
rect 20048 46087 20416 46096
rect 20048 44624 20416 44633
rect 20088 44584 20130 44624
rect 20170 44584 20212 44624
rect 20252 44584 20294 44624
rect 20334 44584 20376 44624
rect 20048 44575 20416 44584
rect 20048 43112 20416 43121
rect 20088 43072 20130 43112
rect 20170 43072 20212 43112
rect 20252 43072 20294 43112
rect 20334 43072 20376 43112
rect 20048 43063 20416 43072
rect 20048 41600 20416 41609
rect 20088 41560 20130 41600
rect 20170 41560 20212 41600
rect 20252 41560 20294 41600
rect 20334 41560 20376 41600
rect 20048 41551 20416 41560
rect 20048 40088 20416 40097
rect 20088 40048 20130 40088
rect 20170 40048 20212 40088
rect 20252 40048 20294 40088
rect 20334 40048 20376 40088
rect 20048 40039 20416 40048
rect 20048 38576 20416 38585
rect 20088 38536 20130 38576
rect 20170 38536 20212 38576
rect 20252 38536 20294 38576
rect 20334 38536 20376 38576
rect 20048 38527 20416 38536
rect 20048 37064 20416 37073
rect 20088 37024 20130 37064
rect 20170 37024 20212 37064
rect 20252 37024 20294 37064
rect 20334 37024 20376 37064
rect 20048 37015 20416 37024
rect 20524 36560 20564 36569
rect 20048 35552 20416 35561
rect 20088 35512 20130 35552
rect 20170 35512 20212 35552
rect 20252 35512 20294 35552
rect 20334 35512 20376 35552
rect 20048 35503 20416 35512
rect 20048 34040 20416 34049
rect 20088 34000 20130 34040
rect 20170 34000 20212 34040
rect 20252 34000 20294 34040
rect 20334 34000 20376 34040
rect 20048 33991 20416 34000
rect 19948 32815 19988 32824
rect 20048 32528 20416 32537
rect 20088 32488 20130 32528
rect 20170 32488 20212 32528
rect 20252 32488 20294 32528
rect 20334 32488 20376 32528
rect 20048 32479 20416 32488
rect 19948 31184 19988 31193
rect 19948 30260 19988 31144
rect 20048 31016 20416 31025
rect 20088 30976 20130 31016
rect 20170 30976 20212 31016
rect 20252 30976 20294 31016
rect 20334 30976 20376 31016
rect 20048 30967 20416 30976
rect 19948 30211 19988 30220
rect 20048 29504 20416 29513
rect 20088 29464 20130 29504
rect 20170 29464 20212 29504
rect 20252 29464 20294 29504
rect 20334 29464 20376 29504
rect 20048 29455 20416 29464
rect 19756 28960 19892 29000
rect 19852 26564 19892 28960
rect 19948 28328 19988 28337
rect 19948 26648 19988 28288
rect 20048 27992 20416 28001
rect 20088 27952 20130 27992
rect 20170 27952 20212 27992
rect 20252 27952 20294 27992
rect 20334 27952 20376 27992
rect 20048 27943 20416 27952
rect 19948 26599 19988 26608
rect 19852 26515 19892 26524
rect 20048 26480 20416 26489
rect 20088 26440 20130 26480
rect 20170 26440 20212 26480
rect 20252 26440 20294 26480
rect 20334 26440 20376 26480
rect 20048 26431 20416 26440
rect 20048 24968 20416 24977
rect 20088 24928 20130 24968
rect 20170 24928 20212 24968
rect 20252 24928 20294 24968
rect 20334 24928 20376 24968
rect 20048 24919 20416 24928
rect 20048 23456 20416 23465
rect 20088 23416 20130 23456
rect 20170 23416 20212 23456
rect 20252 23416 20294 23456
rect 20334 23416 20376 23456
rect 20048 23407 20416 23416
rect 20139 22868 20181 22877
rect 20139 22828 20140 22868
rect 20180 22828 20181 22868
rect 20139 22819 20181 22828
rect 20140 22734 20180 22819
rect 20048 21944 20416 21953
rect 20088 21904 20130 21944
rect 20170 21904 20212 21944
rect 20252 21904 20294 21944
rect 20334 21904 20376 21944
rect 20048 21895 20416 21904
rect 20048 20432 20416 20441
rect 20088 20392 20130 20432
rect 20170 20392 20212 20432
rect 20252 20392 20294 20432
rect 20334 20392 20376 20432
rect 20048 20383 20416 20392
rect 20048 18920 20416 18929
rect 20088 18880 20130 18920
rect 20170 18880 20212 18920
rect 20252 18880 20294 18920
rect 20334 18880 20376 18920
rect 20048 18871 20416 18880
rect 20048 17408 20416 17417
rect 20088 17368 20130 17408
rect 20170 17368 20212 17408
rect 20252 17368 20294 17408
rect 20334 17368 20376 17408
rect 20048 17359 20416 17368
rect 20048 15896 20416 15905
rect 20088 15856 20130 15896
rect 20170 15856 20212 15896
rect 20252 15856 20294 15896
rect 20334 15856 20376 15896
rect 20048 15847 20416 15856
rect 20048 14384 20416 14393
rect 20088 14344 20130 14384
rect 20170 14344 20212 14384
rect 20252 14344 20294 14384
rect 20334 14344 20376 14384
rect 20048 14335 20416 14344
rect 20048 12872 20416 12881
rect 20088 12832 20130 12872
rect 20170 12832 20212 12872
rect 20252 12832 20294 12872
rect 20334 12832 20376 12872
rect 20048 12823 20416 12832
rect 20048 11360 20416 11369
rect 20088 11320 20130 11360
rect 20170 11320 20212 11360
rect 20252 11320 20294 11360
rect 20334 11320 20376 11360
rect 20048 11311 20416 11320
rect 20048 9848 20416 9857
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20048 9799 20416 9808
rect 20048 8336 20416 8345
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20048 8287 20416 8296
rect 20048 6824 20416 6833
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20048 6775 20416 6784
rect 20048 5312 20416 5321
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20048 5263 20416 5272
rect 20048 3800 20416 3809
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20048 3751 20416 3760
rect 20048 2288 20416 2297
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20048 2239 20416 2248
rect 19660 1147 19700 1156
rect 20524 1028 20564 36520
rect 20524 979 20564 988
rect 18316 895 18356 904
rect 20620 860 20660 52816
rect 21004 40004 21044 60376
rect 21196 43700 21236 77848
rect 21388 77216 21428 77225
rect 21196 43651 21236 43660
rect 21292 63104 21332 63113
rect 21004 39955 21044 39964
rect 20716 39080 20756 39089
rect 20716 1112 20756 39040
rect 21292 35048 21332 63064
rect 21388 42608 21428 77176
rect 21388 42559 21428 42568
rect 21292 34999 21332 35008
rect 20811 29672 20853 29681
rect 20811 29632 20812 29672
rect 20852 29632 20853 29672
rect 20811 29623 20853 29632
rect 20812 29504 20852 29623
rect 20812 29455 20852 29464
rect 20716 1063 20756 1072
rect 20620 811 20660 820
rect 20048 776 20416 785
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20048 727 20416 736
rect 17932 559 17972 568
rect 13708 139 13748 148
rect 11788 55 11828 64
<< via4 >>
rect 652 62980 692 63020
rect 1036 67432 1076 67472
rect 1132 66340 1172 66380
rect 940 35008 980 35048
rect 844 25096 884 25136
rect 1036 904 1076 944
rect 3688 84652 3728 84692
rect 3770 84652 3810 84692
rect 3852 84652 3892 84692
rect 3934 84652 3974 84692
rect 4016 84652 4056 84692
rect 2092 10648 2132 10688
rect 2284 10648 2324 10688
rect 2572 61720 2612 61760
rect 2476 60964 2516 61004
rect 3688 83140 3728 83180
rect 3770 83140 3810 83180
rect 3852 83140 3892 83180
rect 3934 83140 3974 83180
rect 4016 83140 4056 83180
rect 3688 81628 3728 81668
rect 3770 81628 3810 81668
rect 3852 81628 3892 81668
rect 3934 81628 3974 81668
rect 4016 81628 4056 81668
rect 3688 80116 3728 80156
rect 3770 80116 3810 80156
rect 3852 80116 3892 80156
rect 3934 80116 3974 80156
rect 4016 80116 4056 80156
rect 3688 78604 3728 78644
rect 3770 78604 3810 78644
rect 3852 78604 3892 78644
rect 3934 78604 3974 78644
rect 4016 78604 4056 78644
rect 3688 77092 3728 77132
rect 3770 77092 3810 77132
rect 3852 77092 3892 77132
rect 3934 77092 3974 77132
rect 4016 77092 4056 77132
rect 3688 75580 3728 75620
rect 3770 75580 3810 75620
rect 3852 75580 3892 75620
rect 3934 75580 3974 75620
rect 4016 75580 4056 75620
rect 3688 74068 3728 74108
rect 3770 74068 3810 74108
rect 3852 74068 3892 74108
rect 3934 74068 3974 74108
rect 4016 74068 4056 74108
rect 3688 72556 3728 72596
rect 3770 72556 3810 72596
rect 3852 72556 3892 72596
rect 3934 72556 3974 72596
rect 4016 72556 4056 72596
rect 3688 71044 3728 71084
rect 3770 71044 3810 71084
rect 3852 71044 3892 71084
rect 3934 71044 3974 71084
rect 4016 71044 4056 71084
rect 2476 41224 2516 41264
rect 2860 23752 2900 23792
rect 2956 22828 2996 22868
rect 3148 28372 3188 28412
rect 2956 16780 2996 16820
rect 3436 28372 3476 28412
rect 3688 69532 3728 69572
rect 3770 69532 3810 69572
rect 3852 69532 3892 69572
rect 3934 69532 3974 69572
rect 4016 69532 4056 69572
rect 3628 68524 3668 68564
rect 3688 68020 3728 68060
rect 3770 68020 3810 68060
rect 3852 68020 3892 68060
rect 3934 68020 3974 68060
rect 4016 68020 4056 68060
rect 3820 67432 3860 67472
rect 3688 66508 3728 66548
rect 3770 66508 3810 66548
rect 3852 66508 3892 66548
rect 3934 66508 3974 66548
rect 4016 66508 4056 66548
rect 3688 64996 3728 65036
rect 3770 64996 3810 65036
rect 3852 64996 3892 65036
rect 3934 64996 3974 65036
rect 4016 64996 4056 65036
rect 3688 63484 3728 63524
rect 3770 63484 3810 63524
rect 3852 63484 3892 63524
rect 3934 63484 3974 63524
rect 4016 63484 4056 63524
rect 3688 61972 3728 62012
rect 3770 61972 3810 62012
rect 3852 61972 3892 62012
rect 3934 61972 3974 62012
rect 4016 61972 4056 62012
rect 3916 61720 3956 61760
rect 3688 60460 3728 60500
rect 3770 60460 3810 60500
rect 3852 60460 3892 60500
rect 3934 60460 3974 60500
rect 4016 60460 4056 60500
rect 3688 58948 3728 58988
rect 3770 58948 3810 58988
rect 3852 58948 3892 58988
rect 3934 58948 3974 58988
rect 4016 58948 4056 58988
rect 3688 57436 3728 57476
rect 3770 57436 3810 57476
rect 3852 57436 3892 57476
rect 3934 57436 3974 57476
rect 4016 57436 4056 57476
rect 3688 55924 3728 55964
rect 3770 55924 3810 55964
rect 3852 55924 3892 55964
rect 3934 55924 3974 55964
rect 4016 55924 4056 55964
rect 3688 54412 3728 54452
rect 3770 54412 3810 54452
rect 3852 54412 3892 54452
rect 3934 54412 3974 54452
rect 4016 54412 4056 54452
rect 3688 52900 3728 52940
rect 3770 52900 3810 52940
rect 3852 52900 3892 52940
rect 3934 52900 3974 52940
rect 4016 52900 4056 52940
rect 3688 51388 3728 51428
rect 3770 51388 3810 51428
rect 3852 51388 3892 51428
rect 3934 51388 3974 51428
rect 4016 51388 4056 51428
rect 3688 49876 3728 49916
rect 3770 49876 3810 49916
rect 3852 49876 3892 49916
rect 3934 49876 3974 49916
rect 4016 49876 4056 49916
rect 3688 48364 3728 48404
rect 3770 48364 3810 48404
rect 3852 48364 3892 48404
rect 3934 48364 3974 48404
rect 4016 48364 4056 48404
rect 3688 46852 3728 46892
rect 3770 46852 3810 46892
rect 3852 46852 3892 46892
rect 3934 46852 3974 46892
rect 4016 46852 4056 46892
rect 3688 45340 3728 45380
rect 3770 45340 3810 45380
rect 3852 45340 3892 45380
rect 3934 45340 3974 45380
rect 4016 45340 4056 45380
rect 3688 43828 3728 43868
rect 3770 43828 3810 43868
rect 3852 43828 3892 43868
rect 3934 43828 3974 43868
rect 4016 43828 4056 43868
rect 3688 42316 3728 42356
rect 3770 42316 3810 42356
rect 3852 42316 3892 42356
rect 3934 42316 3974 42356
rect 4016 42316 4056 42356
rect 3688 40804 3728 40844
rect 3770 40804 3810 40844
rect 3852 40804 3892 40844
rect 3934 40804 3974 40844
rect 4016 40804 4056 40844
rect 3688 39292 3728 39332
rect 3770 39292 3810 39332
rect 3852 39292 3892 39332
rect 3934 39292 3974 39332
rect 4016 39292 4056 39332
rect 3688 37780 3728 37820
rect 3770 37780 3810 37820
rect 3852 37780 3892 37820
rect 3934 37780 3974 37820
rect 4016 37780 4056 37820
rect 3688 36268 3728 36308
rect 3770 36268 3810 36308
rect 3852 36268 3892 36308
rect 3934 36268 3974 36308
rect 4016 36268 4056 36308
rect 3820 35008 3860 35048
rect 3688 34756 3728 34796
rect 3770 34756 3810 34796
rect 3852 34756 3892 34796
rect 3934 34756 3974 34796
rect 4016 34756 4056 34796
rect 3916 34252 3956 34292
rect 3688 33244 3728 33284
rect 3770 33244 3810 33284
rect 3852 33244 3892 33284
rect 3934 33244 3974 33284
rect 4016 33244 4056 33284
rect 3688 31732 3728 31772
rect 3770 31732 3810 31772
rect 3852 31732 3892 31772
rect 3934 31732 3974 31772
rect 4016 31732 4056 31772
rect 3688 30220 3728 30260
rect 3770 30220 3810 30260
rect 3852 30220 3892 30260
rect 3934 30220 3974 30260
rect 4016 30220 4056 30260
rect 4492 62980 4532 63020
rect 4588 60964 4628 61004
rect 4928 83896 4968 83936
rect 5010 83896 5050 83936
rect 5092 83896 5132 83936
rect 5174 83896 5214 83936
rect 5256 83896 5296 83936
rect 4928 82384 4968 82424
rect 5010 82384 5050 82424
rect 5092 82384 5132 82424
rect 5174 82384 5214 82424
rect 5256 82384 5296 82424
rect 4928 80872 4968 80912
rect 5010 80872 5050 80912
rect 5092 80872 5132 80912
rect 5174 80872 5214 80912
rect 5256 80872 5296 80912
rect 4928 79360 4968 79400
rect 5010 79360 5050 79400
rect 5092 79360 5132 79400
rect 5174 79360 5214 79400
rect 5256 79360 5296 79400
rect 4928 77848 4968 77888
rect 5010 77848 5050 77888
rect 5092 77848 5132 77888
rect 5174 77848 5214 77888
rect 5256 77848 5296 77888
rect 4928 76336 4968 76376
rect 5010 76336 5050 76376
rect 5092 76336 5132 76376
rect 5174 76336 5214 76376
rect 5256 76336 5296 76376
rect 4928 74824 4968 74864
rect 5010 74824 5050 74864
rect 5092 74824 5132 74864
rect 5174 74824 5214 74864
rect 5256 74824 5296 74864
rect 4928 73312 4968 73352
rect 5010 73312 5050 73352
rect 5092 73312 5132 73352
rect 5174 73312 5214 73352
rect 5256 73312 5296 73352
rect 4928 71800 4968 71840
rect 5010 71800 5050 71840
rect 5092 71800 5132 71840
rect 5174 71800 5214 71840
rect 5256 71800 5296 71840
rect 4928 70288 4968 70328
rect 5010 70288 5050 70328
rect 5092 70288 5132 70328
rect 5174 70288 5214 70328
rect 5256 70288 5296 70328
rect 4928 68776 4968 68816
rect 5010 68776 5050 68816
rect 5092 68776 5132 68816
rect 5174 68776 5214 68816
rect 5256 68776 5296 68816
rect 4876 68524 4916 68564
rect 4928 67264 4968 67304
rect 5010 67264 5050 67304
rect 5092 67264 5132 67304
rect 5174 67264 5214 67304
rect 5256 67264 5296 67304
rect 4928 65752 4968 65792
rect 5010 65752 5050 65792
rect 5092 65752 5132 65792
rect 5174 65752 5214 65792
rect 5256 65752 5296 65792
rect 4928 64240 4968 64280
rect 5010 64240 5050 64280
rect 5092 64240 5132 64280
rect 5174 64240 5214 64280
rect 5256 64240 5296 64280
rect 4928 62728 4968 62768
rect 5010 62728 5050 62768
rect 5092 62728 5132 62768
rect 5174 62728 5214 62768
rect 5256 62728 5296 62768
rect 4928 61216 4968 61256
rect 5010 61216 5050 61256
rect 5092 61216 5132 61256
rect 5174 61216 5214 61256
rect 5256 61216 5296 61256
rect 4928 59704 4968 59744
rect 5010 59704 5050 59744
rect 5092 59704 5132 59744
rect 5174 59704 5214 59744
rect 5256 59704 5296 59744
rect 4928 58192 4968 58232
rect 5010 58192 5050 58232
rect 5092 58192 5132 58232
rect 5174 58192 5214 58232
rect 5256 58192 5296 58232
rect 4928 56680 4968 56720
rect 5010 56680 5050 56720
rect 5092 56680 5132 56720
rect 5174 56680 5214 56720
rect 5256 56680 5296 56720
rect 4928 55168 4968 55208
rect 5010 55168 5050 55208
rect 5092 55168 5132 55208
rect 5174 55168 5214 55208
rect 5256 55168 5296 55208
rect 4928 53656 4968 53696
rect 5010 53656 5050 53696
rect 5092 53656 5132 53696
rect 5174 53656 5214 53696
rect 5256 53656 5296 53696
rect 4928 52144 4968 52184
rect 5010 52144 5050 52184
rect 5092 52144 5132 52184
rect 5174 52144 5214 52184
rect 5256 52144 5296 52184
rect 4928 50632 4968 50672
rect 5010 50632 5050 50672
rect 5092 50632 5132 50672
rect 5174 50632 5214 50672
rect 5256 50632 5296 50672
rect 4928 49120 4968 49160
rect 5010 49120 5050 49160
rect 5092 49120 5132 49160
rect 5174 49120 5214 49160
rect 5256 49120 5296 49160
rect 4928 47608 4968 47648
rect 5010 47608 5050 47648
rect 5092 47608 5132 47648
rect 5174 47608 5214 47648
rect 5256 47608 5296 47648
rect 4928 46096 4968 46136
rect 5010 46096 5050 46136
rect 5092 46096 5132 46136
rect 5174 46096 5214 46136
rect 5256 46096 5296 46136
rect 4928 44584 4968 44624
rect 5010 44584 5050 44624
rect 5092 44584 5132 44624
rect 5174 44584 5214 44624
rect 5256 44584 5296 44624
rect 4928 43072 4968 43112
rect 5010 43072 5050 43112
rect 5092 43072 5132 43112
rect 5174 43072 5214 43112
rect 5256 43072 5296 43112
rect 4928 41560 4968 41600
rect 5010 41560 5050 41600
rect 5092 41560 5132 41600
rect 5174 41560 5214 41600
rect 5256 41560 5296 41600
rect 3688 28708 3728 28748
rect 3770 28708 3810 28748
rect 3852 28708 3892 28748
rect 3934 28708 3974 28748
rect 4016 28708 4056 28748
rect 3688 27196 3728 27236
rect 3770 27196 3810 27236
rect 3852 27196 3892 27236
rect 3934 27196 3974 27236
rect 4016 27196 4056 27236
rect 3688 25684 3728 25724
rect 3770 25684 3810 25724
rect 3852 25684 3892 25724
rect 3934 25684 3974 25724
rect 4016 25684 4056 25724
rect 3688 24172 3728 24212
rect 3770 24172 3810 24212
rect 3852 24172 3892 24212
rect 3934 24172 3974 24212
rect 4016 24172 4056 24212
rect 3688 22660 3728 22700
rect 3770 22660 3810 22700
rect 3852 22660 3892 22700
rect 3934 22660 3974 22700
rect 4016 22660 4056 22700
rect 3688 21148 3728 21188
rect 3770 21148 3810 21188
rect 3852 21148 3892 21188
rect 3934 21148 3974 21188
rect 4016 21148 4056 21188
rect 3688 19636 3728 19676
rect 3770 19636 3810 19676
rect 3852 19636 3892 19676
rect 3934 19636 3974 19676
rect 4016 19636 4056 19676
rect 4928 40048 4968 40088
rect 5010 40048 5050 40088
rect 5092 40048 5132 40088
rect 5174 40048 5214 40088
rect 5256 40048 5296 40088
rect 4928 38536 4968 38576
rect 5010 38536 5050 38576
rect 5092 38536 5132 38576
rect 5174 38536 5214 38576
rect 5256 38536 5296 38576
rect 4928 37024 4968 37064
rect 5010 37024 5050 37064
rect 5092 37024 5132 37064
rect 5174 37024 5214 37064
rect 5256 37024 5296 37064
rect 5356 36688 5396 36728
rect 4928 35512 4968 35552
rect 5010 35512 5050 35552
rect 5092 35512 5132 35552
rect 5174 35512 5214 35552
rect 5256 35512 5296 35552
rect 4928 34000 4968 34040
rect 5010 34000 5050 34040
rect 5092 34000 5132 34040
rect 5174 34000 5214 34040
rect 5256 34000 5296 34040
rect 4928 32488 4968 32528
rect 5010 32488 5050 32528
rect 5092 32488 5132 32528
rect 5174 32488 5214 32528
rect 5256 32488 5296 32528
rect 4928 30976 4968 31016
rect 5010 30976 5050 31016
rect 5092 30976 5132 31016
rect 5174 30976 5214 31016
rect 5256 30976 5296 31016
rect 4928 29464 4968 29504
rect 5010 29464 5050 29504
rect 5092 29464 5132 29504
rect 5174 29464 5214 29504
rect 5256 29464 5296 29504
rect 3688 18124 3728 18164
rect 3770 18124 3810 18164
rect 3852 18124 3892 18164
rect 3934 18124 3974 18164
rect 4016 18124 4056 18164
rect 4684 26020 4724 26060
rect 4928 27952 4968 27992
rect 5010 27952 5050 27992
rect 5092 27952 5132 27992
rect 5174 27952 5214 27992
rect 5256 27952 5296 27992
rect 4928 26440 4968 26480
rect 5010 26440 5050 26480
rect 5092 26440 5132 26480
rect 5174 26440 5214 26480
rect 5256 26440 5296 26480
rect 5068 25180 5108 25220
rect 5260 25096 5300 25136
rect 4928 24928 4968 24968
rect 5010 24928 5050 24968
rect 5092 24928 5132 24968
rect 5174 24928 5214 24968
rect 5256 24928 5296 24968
rect 4928 23416 4968 23456
rect 5010 23416 5050 23456
rect 5092 23416 5132 23456
rect 5174 23416 5214 23456
rect 5256 23416 5296 23456
rect 4928 21904 4968 21944
rect 5010 21904 5050 21944
rect 5092 21904 5132 21944
rect 5174 21904 5214 21944
rect 5256 21904 5296 21944
rect 4928 20392 4968 20432
rect 5010 20392 5050 20432
rect 5092 20392 5132 20432
rect 5174 20392 5214 20432
rect 5256 20392 5296 20432
rect 4928 18880 4968 18920
rect 5010 18880 5050 18920
rect 5092 18880 5132 18920
rect 5174 18880 5214 18920
rect 5256 18880 5296 18920
rect 4396 17536 4436 17576
rect 3688 16612 3728 16652
rect 3770 16612 3810 16652
rect 3852 16612 3892 16652
rect 3934 16612 3974 16652
rect 4016 16612 4056 16652
rect 3688 15100 3728 15140
rect 3770 15100 3810 15140
rect 3852 15100 3892 15140
rect 3934 15100 3974 15140
rect 4016 15100 4056 15140
rect 3688 13588 3728 13628
rect 3770 13588 3810 13628
rect 3852 13588 3892 13628
rect 3934 13588 3974 13628
rect 4016 13588 4056 13628
rect 3688 12076 3728 12116
rect 3770 12076 3810 12116
rect 3852 12076 3892 12116
rect 3934 12076 3974 12116
rect 4016 12076 4056 12116
rect 4928 17368 4968 17408
rect 5010 17368 5050 17408
rect 5092 17368 5132 17408
rect 5174 17368 5214 17408
rect 5256 17368 5296 17408
rect 4928 15856 4968 15896
rect 5010 15856 5050 15896
rect 5092 15856 5132 15896
rect 5174 15856 5214 15896
rect 5256 15856 5296 15896
rect 4928 14344 4968 14384
rect 5010 14344 5050 14384
rect 5092 14344 5132 14384
rect 5174 14344 5214 14384
rect 5256 14344 5296 14384
rect 4928 12832 4968 12872
rect 5010 12832 5050 12872
rect 5092 12832 5132 12872
rect 5174 12832 5214 12872
rect 5256 12832 5296 12872
rect 4928 11320 4968 11360
rect 5010 11320 5050 11360
rect 5092 11320 5132 11360
rect 5174 11320 5214 11360
rect 5256 11320 5296 11360
rect 3688 10564 3728 10604
rect 3770 10564 3810 10604
rect 3852 10564 3892 10604
rect 3934 10564 3974 10604
rect 4016 10564 4056 10604
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 5836 64408 5876 64448
rect 6028 42736 6068 42776
rect 5932 41224 5972 41264
rect 5740 17536 5780 17576
rect 5644 16780 5684 16820
rect 6316 904 6356 944
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 6604 16780 6644 16820
rect 6604 2164 6644 2204
rect 6700 1240 6740 1280
rect 6988 4768 7028 4808
rect 7756 83476 7796 83516
rect 8332 42484 8372 42524
rect 8716 67768 8756 67808
rect 8428 40972 8468 41012
rect 7948 2164 7988 2204
rect 8524 4768 8564 4808
rect 9004 34252 9044 34292
rect 9676 41728 9716 41768
rect 9964 62980 10004 63020
rect 10348 69280 10388 69320
rect 10732 72724 10772 72764
rect 10828 25096 10868 25136
rect 11308 41392 11348 41432
rect 11596 41392 11636 41432
rect 12460 72136 12500 72176
rect 11788 42736 11828 42776
rect 11308 25096 11348 25136
rect 11020 3424 11060 3464
rect 3724 316 3764 356
rect 2956 232 2996 272
rect 11788 36688 11828 36728
rect 11980 34168 12020 34208
rect 5260 148 5300 188
rect 10828 148 10868 188
rect 12076 26440 12116 26480
rect 12364 37444 12404 37484
rect 12364 30640 12404 30680
rect 12364 26272 12404 26312
rect 12652 34168 12692 34208
rect 12364 6952 12404 6992
rect 13132 83308 13172 83348
rect 13036 61300 13076 61340
rect 12940 36688 12980 36728
rect 13804 66340 13844 66380
rect 12556 1072 12596 1112
rect 11980 316 12020 356
rect 14092 23752 14132 23792
rect 14092 17620 14132 17660
rect 14284 6952 14324 6992
rect 14572 26020 14612 26060
rect 15340 58864 15380 58904
rect 18808 84652 18848 84692
rect 18890 84652 18930 84692
rect 18972 84652 19012 84692
rect 19054 84652 19094 84692
rect 19136 84652 19176 84692
rect 16012 61300 16052 61340
rect 16012 58864 16052 58904
rect 16300 40636 16340 40676
rect 16684 29632 16724 29672
rect 20048 83896 20088 83936
rect 20130 83896 20170 83936
rect 20212 83896 20252 83936
rect 20294 83896 20334 83936
rect 20376 83896 20416 83936
rect 17644 25180 17684 25220
rect 18316 6280 18356 6320
rect 19084 83476 19124 83516
rect 18808 83140 18848 83180
rect 18890 83140 18930 83180
rect 18972 83140 19012 83180
rect 19054 83140 19094 83180
rect 19136 83140 19176 83180
rect 18808 81628 18848 81668
rect 18890 81628 18930 81668
rect 18972 81628 19012 81668
rect 19054 81628 19094 81668
rect 19136 81628 19176 81668
rect 18808 80116 18848 80156
rect 18890 80116 18930 80156
rect 18972 80116 19012 80156
rect 19054 80116 19094 80156
rect 19136 80116 19176 80156
rect 18808 78604 18848 78644
rect 18890 78604 18930 78644
rect 18972 78604 19012 78644
rect 19054 78604 19094 78644
rect 19136 78604 19176 78644
rect 18808 77092 18848 77132
rect 18890 77092 18930 77132
rect 18972 77092 19012 77132
rect 19054 77092 19094 77132
rect 19136 77092 19176 77132
rect 18808 75580 18848 75620
rect 18890 75580 18930 75620
rect 18972 75580 19012 75620
rect 19054 75580 19094 75620
rect 19136 75580 19176 75620
rect 18808 74068 18848 74108
rect 18890 74068 18930 74108
rect 18972 74068 19012 74108
rect 19054 74068 19094 74108
rect 19136 74068 19176 74108
rect 18808 72556 18848 72596
rect 18890 72556 18930 72596
rect 18972 72556 19012 72596
rect 19054 72556 19094 72596
rect 19136 72556 19176 72596
rect 18808 71044 18848 71084
rect 18890 71044 18930 71084
rect 18972 71044 19012 71084
rect 19054 71044 19094 71084
rect 19136 71044 19176 71084
rect 18808 69532 18848 69572
rect 18890 69532 18930 69572
rect 18972 69532 19012 69572
rect 19054 69532 19094 69572
rect 19136 69532 19176 69572
rect 18808 68020 18848 68060
rect 18890 68020 18930 68060
rect 18972 68020 19012 68060
rect 19054 68020 19094 68060
rect 19136 68020 19176 68060
rect 18808 66508 18848 66548
rect 18890 66508 18930 66548
rect 18972 66508 19012 66548
rect 19054 66508 19094 66548
rect 19136 66508 19176 66548
rect 18808 64996 18848 65036
rect 18890 64996 18930 65036
rect 18972 64996 19012 65036
rect 19054 64996 19094 65036
rect 19136 64996 19176 65036
rect 18808 63484 18848 63524
rect 18890 63484 18930 63524
rect 18972 63484 19012 63524
rect 19054 63484 19094 63524
rect 19136 63484 19176 63524
rect 18808 61972 18848 62012
rect 18890 61972 18930 62012
rect 18972 61972 19012 62012
rect 19054 61972 19094 62012
rect 19136 61972 19176 62012
rect 18808 60460 18848 60500
rect 18890 60460 18930 60500
rect 18972 60460 19012 60500
rect 19054 60460 19094 60500
rect 19136 60460 19176 60500
rect 18808 58948 18848 58988
rect 18890 58948 18930 58988
rect 18972 58948 19012 58988
rect 19054 58948 19094 58988
rect 19136 58948 19176 58988
rect 18808 57436 18848 57476
rect 18890 57436 18930 57476
rect 18972 57436 19012 57476
rect 19054 57436 19094 57476
rect 19136 57436 19176 57476
rect 18808 55924 18848 55964
rect 18890 55924 18930 55964
rect 18972 55924 19012 55964
rect 19054 55924 19094 55964
rect 19136 55924 19176 55964
rect 18808 54412 18848 54452
rect 18890 54412 18930 54452
rect 18972 54412 19012 54452
rect 19054 54412 19094 54452
rect 19136 54412 19176 54452
rect 18808 52900 18848 52940
rect 18890 52900 18930 52940
rect 18972 52900 19012 52940
rect 19054 52900 19094 52940
rect 19136 52900 19176 52940
rect 18808 51388 18848 51428
rect 18890 51388 18930 51428
rect 18972 51388 19012 51428
rect 19054 51388 19094 51428
rect 19136 51388 19176 51428
rect 18808 49876 18848 49916
rect 18890 49876 18930 49916
rect 18972 49876 19012 49916
rect 19054 49876 19094 49916
rect 19136 49876 19176 49916
rect 18808 48364 18848 48404
rect 18890 48364 18930 48404
rect 18972 48364 19012 48404
rect 19054 48364 19094 48404
rect 19136 48364 19176 48404
rect 18808 46852 18848 46892
rect 18890 46852 18930 46892
rect 18972 46852 19012 46892
rect 19054 46852 19094 46892
rect 19136 46852 19176 46892
rect 18808 45340 18848 45380
rect 18890 45340 18930 45380
rect 18972 45340 19012 45380
rect 19054 45340 19094 45380
rect 19136 45340 19176 45380
rect 18808 43828 18848 43868
rect 18890 43828 18930 43868
rect 18972 43828 19012 43868
rect 19054 43828 19094 43868
rect 19136 43828 19176 43868
rect 18796 42484 18836 42524
rect 18808 42316 18848 42356
rect 18890 42316 18930 42356
rect 18972 42316 19012 42356
rect 19054 42316 19094 42356
rect 19136 42316 19176 42356
rect 18808 40804 18848 40844
rect 18890 40804 18930 40844
rect 18972 40804 19012 40844
rect 19054 40804 19094 40844
rect 19136 40804 19176 40844
rect 18808 39292 18848 39332
rect 18890 39292 18930 39332
rect 18972 39292 19012 39332
rect 19054 39292 19094 39332
rect 19136 39292 19176 39332
rect 18808 37780 18848 37820
rect 18890 37780 18930 37820
rect 18972 37780 19012 37820
rect 19054 37780 19094 37820
rect 19136 37780 19176 37820
rect 18808 36268 18848 36308
rect 18890 36268 18930 36308
rect 18972 36268 19012 36308
rect 19054 36268 19094 36308
rect 19136 36268 19176 36308
rect 18808 34756 18848 34796
rect 18890 34756 18930 34796
rect 18972 34756 19012 34796
rect 19054 34756 19094 34796
rect 19136 34756 19176 34796
rect 18808 33244 18848 33284
rect 18890 33244 18930 33284
rect 18972 33244 19012 33284
rect 19054 33244 19094 33284
rect 19136 33244 19176 33284
rect 18808 31732 18848 31772
rect 18890 31732 18930 31772
rect 18972 31732 19012 31772
rect 19054 31732 19094 31772
rect 19136 31732 19176 31772
rect 18808 30220 18848 30260
rect 18890 30220 18930 30260
rect 18972 30220 19012 30260
rect 19054 30220 19094 30260
rect 19136 30220 19176 30260
rect 18808 28708 18848 28748
rect 18890 28708 18930 28748
rect 18972 28708 19012 28748
rect 19054 28708 19094 28748
rect 19136 28708 19176 28748
rect 18808 27196 18848 27236
rect 18890 27196 18930 27236
rect 18972 27196 19012 27236
rect 19054 27196 19094 27236
rect 19136 27196 19176 27236
rect 18808 25684 18848 25724
rect 18890 25684 18930 25724
rect 18972 25684 19012 25724
rect 19054 25684 19094 25724
rect 19136 25684 19176 25724
rect 18808 24172 18848 24212
rect 18890 24172 18930 24212
rect 18972 24172 19012 24212
rect 19054 24172 19094 24212
rect 19136 24172 19176 24212
rect 18808 22660 18848 22700
rect 18890 22660 18930 22700
rect 18972 22660 19012 22700
rect 19054 22660 19094 22700
rect 19136 22660 19176 22700
rect 18808 21148 18848 21188
rect 18890 21148 18930 21188
rect 18972 21148 19012 21188
rect 19054 21148 19094 21188
rect 19136 21148 19176 21188
rect 18808 19636 18848 19676
rect 18890 19636 18930 19676
rect 18972 19636 19012 19676
rect 19054 19636 19094 19676
rect 19136 19636 19176 19676
rect 18808 18124 18848 18164
rect 18890 18124 18930 18164
rect 18972 18124 19012 18164
rect 19054 18124 19094 18164
rect 19136 18124 19176 18164
rect 18808 16612 18848 16652
rect 18890 16612 18930 16652
rect 18972 16612 19012 16652
rect 19054 16612 19094 16652
rect 19136 16612 19176 16652
rect 18808 15100 18848 15140
rect 18890 15100 18930 15140
rect 18972 15100 19012 15140
rect 19054 15100 19094 15140
rect 19136 15100 19176 15140
rect 18808 13588 18848 13628
rect 18890 13588 18930 13628
rect 18972 13588 19012 13628
rect 19054 13588 19094 13628
rect 19136 13588 19176 13628
rect 18808 12076 18848 12116
rect 18890 12076 18930 12116
rect 18972 12076 19012 12116
rect 19054 12076 19094 12116
rect 19136 12076 19176 12116
rect 18808 10564 18848 10604
rect 18890 10564 18930 10604
rect 18972 10564 19012 10604
rect 19054 10564 19094 10604
rect 19136 10564 19176 10604
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 20048 82384 20088 82424
rect 20130 82384 20170 82424
rect 20212 82384 20252 82424
rect 20294 82384 20334 82424
rect 20376 82384 20416 82424
rect 20048 80872 20088 80912
rect 20130 80872 20170 80912
rect 20212 80872 20252 80912
rect 20294 80872 20334 80912
rect 20376 80872 20416 80912
rect 20048 79360 20088 79400
rect 20130 79360 20170 79400
rect 20212 79360 20252 79400
rect 20294 79360 20334 79400
rect 20376 79360 20416 79400
rect 20048 77848 20088 77888
rect 20130 77848 20170 77888
rect 20212 77848 20252 77888
rect 20294 77848 20334 77888
rect 20376 77848 20416 77888
rect 20048 76336 20088 76376
rect 20130 76336 20170 76376
rect 20212 76336 20252 76376
rect 20294 76336 20334 76376
rect 20376 76336 20416 76376
rect 20048 74824 20088 74864
rect 20130 74824 20170 74864
rect 20212 74824 20252 74864
rect 20294 74824 20334 74864
rect 20376 74824 20416 74864
rect 20048 73312 20088 73352
rect 20130 73312 20170 73352
rect 20212 73312 20252 73352
rect 20294 73312 20334 73352
rect 20376 73312 20416 73352
rect 20048 71800 20088 71840
rect 20130 71800 20170 71840
rect 20212 71800 20252 71840
rect 20294 71800 20334 71840
rect 20376 71800 20416 71840
rect 20048 70288 20088 70328
rect 20130 70288 20170 70328
rect 20212 70288 20252 70328
rect 20294 70288 20334 70328
rect 20376 70288 20416 70328
rect 20048 68776 20088 68816
rect 20130 68776 20170 68816
rect 20212 68776 20252 68816
rect 20294 68776 20334 68816
rect 20376 68776 20416 68816
rect 20140 67768 20180 67808
rect 20048 67264 20088 67304
rect 20130 67264 20170 67304
rect 20212 67264 20252 67304
rect 20294 67264 20334 67304
rect 20376 67264 20416 67304
rect 19468 40972 19508 41012
rect 19468 40636 19508 40676
rect 19660 41728 19700 41768
rect 19564 37444 19604 37484
rect 20048 65752 20088 65792
rect 20130 65752 20170 65792
rect 20212 65752 20252 65792
rect 20294 65752 20334 65792
rect 20376 65752 20416 65792
rect 20048 64240 20088 64280
rect 20130 64240 20170 64280
rect 20212 64240 20252 64280
rect 20294 64240 20334 64280
rect 20376 64240 20416 64280
rect 20048 62728 20088 62768
rect 20130 62728 20170 62768
rect 20212 62728 20252 62768
rect 20294 62728 20334 62768
rect 20376 62728 20416 62768
rect 20048 61216 20088 61256
rect 20130 61216 20170 61256
rect 20212 61216 20252 61256
rect 20294 61216 20334 61256
rect 20376 61216 20416 61256
rect 20048 59704 20088 59744
rect 20130 59704 20170 59744
rect 20212 59704 20252 59744
rect 20294 59704 20334 59744
rect 20376 59704 20416 59744
rect 20048 58192 20088 58232
rect 20130 58192 20170 58232
rect 20212 58192 20252 58232
rect 20294 58192 20334 58232
rect 20376 58192 20416 58232
rect 20048 56680 20088 56720
rect 20130 56680 20170 56720
rect 20212 56680 20252 56720
rect 20294 56680 20334 56720
rect 20376 56680 20416 56720
rect 20048 55168 20088 55208
rect 20130 55168 20170 55208
rect 20212 55168 20252 55208
rect 20294 55168 20334 55208
rect 20376 55168 20416 55208
rect 20048 53656 20088 53696
rect 20130 53656 20170 53696
rect 20212 53656 20252 53696
rect 20294 53656 20334 53696
rect 20376 53656 20416 53696
rect 20048 52144 20088 52184
rect 20130 52144 20170 52184
rect 20212 52144 20252 52184
rect 20294 52144 20334 52184
rect 20376 52144 20416 52184
rect 20048 50632 20088 50672
rect 20130 50632 20170 50672
rect 20212 50632 20252 50672
rect 20294 50632 20334 50672
rect 20376 50632 20416 50672
rect 20048 49120 20088 49160
rect 20130 49120 20170 49160
rect 20212 49120 20252 49160
rect 20294 49120 20334 49160
rect 20376 49120 20416 49160
rect 20048 47608 20088 47648
rect 20130 47608 20170 47648
rect 20212 47608 20252 47648
rect 20294 47608 20334 47648
rect 20376 47608 20416 47648
rect 20048 46096 20088 46136
rect 20130 46096 20170 46136
rect 20212 46096 20252 46136
rect 20294 46096 20334 46136
rect 20376 46096 20416 46136
rect 20048 44584 20088 44624
rect 20130 44584 20170 44624
rect 20212 44584 20252 44624
rect 20294 44584 20334 44624
rect 20376 44584 20416 44624
rect 20048 43072 20088 43112
rect 20130 43072 20170 43112
rect 20212 43072 20252 43112
rect 20294 43072 20334 43112
rect 20376 43072 20416 43112
rect 20048 41560 20088 41600
rect 20130 41560 20170 41600
rect 20212 41560 20252 41600
rect 20294 41560 20334 41600
rect 20376 41560 20416 41600
rect 20048 40048 20088 40088
rect 20130 40048 20170 40088
rect 20212 40048 20252 40088
rect 20294 40048 20334 40088
rect 20376 40048 20416 40088
rect 20048 38536 20088 38576
rect 20130 38536 20170 38576
rect 20212 38536 20252 38576
rect 20294 38536 20334 38576
rect 20376 38536 20416 38576
rect 20048 37024 20088 37064
rect 20130 37024 20170 37064
rect 20212 37024 20252 37064
rect 20294 37024 20334 37064
rect 20376 37024 20416 37064
rect 20048 35512 20088 35552
rect 20130 35512 20170 35552
rect 20212 35512 20252 35552
rect 20294 35512 20334 35552
rect 20376 35512 20416 35552
rect 20048 34000 20088 34040
rect 20130 34000 20170 34040
rect 20212 34000 20252 34040
rect 20294 34000 20334 34040
rect 20376 34000 20416 34040
rect 20048 32488 20088 32528
rect 20130 32488 20170 32528
rect 20212 32488 20252 32528
rect 20294 32488 20334 32528
rect 20376 32488 20416 32528
rect 20048 30976 20088 31016
rect 20130 30976 20170 31016
rect 20212 30976 20252 31016
rect 20294 30976 20334 31016
rect 20376 30976 20416 31016
rect 20048 29464 20088 29504
rect 20130 29464 20170 29504
rect 20212 29464 20252 29504
rect 20294 29464 20334 29504
rect 20376 29464 20416 29504
rect 20048 27952 20088 27992
rect 20130 27952 20170 27992
rect 20212 27952 20252 27992
rect 20294 27952 20334 27992
rect 20376 27952 20416 27992
rect 20048 26440 20088 26480
rect 20130 26440 20170 26480
rect 20212 26440 20252 26480
rect 20294 26440 20334 26480
rect 20376 26440 20416 26480
rect 20048 24928 20088 24968
rect 20130 24928 20170 24968
rect 20212 24928 20252 24968
rect 20294 24928 20334 24968
rect 20376 24928 20416 24968
rect 20048 23416 20088 23456
rect 20130 23416 20170 23456
rect 20212 23416 20252 23456
rect 20294 23416 20334 23456
rect 20376 23416 20416 23456
rect 20140 22828 20180 22868
rect 20048 21904 20088 21944
rect 20130 21904 20170 21944
rect 20212 21904 20252 21944
rect 20294 21904 20334 21944
rect 20376 21904 20416 21944
rect 20048 20392 20088 20432
rect 20130 20392 20170 20432
rect 20212 20392 20252 20432
rect 20294 20392 20334 20432
rect 20376 20392 20416 20432
rect 20048 18880 20088 18920
rect 20130 18880 20170 18920
rect 20212 18880 20252 18920
rect 20294 18880 20334 18920
rect 20376 18880 20416 18920
rect 20048 17368 20088 17408
rect 20130 17368 20170 17408
rect 20212 17368 20252 17408
rect 20294 17368 20334 17408
rect 20376 17368 20416 17408
rect 20048 15856 20088 15896
rect 20130 15856 20170 15896
rect 20212 15856 20252 15896
rect 20294 15856 20334 15896
rect 20376 15856 20416 15896
rect 20048 14344 20088 14384
rect 20130 14344 20170 14384
rect 20212 14344 20252 14384
rect 20294 14344 20334 14384
rect 20376 14344 20416 14384
rect 20048 12832 20088 12872
rect 20130 12832 20170 12872
rect 20212 12832 20252 12872
rect 20294 12832 20334 12872
rect 20376 12832 20416 12872
rect 20048 11320 20088 11360
rect 20130 11320 20170 11360
rect 20212 11320 20252 11360
rect 20294 11320 20334 11360
rect 20376 11320 20416 11360
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 20812 29632 20852 29672
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
<< metal5 >>
rect 3679 84715 4065 84734
rect 3679 84692 3745 84715
rect 3831 84692 3913 84715
rect 3999 84692 4065 84715
rect 3679 84652 3688 84692
rect 3728 84652 3745 84692
rect 3831 84652 3852 84692
rect 3892 84652 3913 84692
rect 3999 84652 4016 84692
rect 4056 84652 4065 84692
rect 3679 84629 3745 84652
rect 3831 84629 3913 84652
rect 3999 84629 4065 84652
rect 3679 84610 4065 84629
rect 18799 84715 19185 84734
rect 18799 84692 18865 84715
rect 18951 84692 19033 84715
rect 19119 84692 19185 84715
rect 18799 84652 18808 84692
rect 18848 84652 18865 84692
rect 18951 84652 18972 84692
rect 19012 84652 19033 84692
rect 19119 84652 19136 84692
rect 19176 84652 19185 84692
rect 18799 84629 18865 84652
rect 18951 84629 19033 84652
rect 19119 84629 19185 84652
rect 18799 84610 19185 84629
rect 4919 83959 5305 83978
rect 4919 83936 4985 83959
rect 5071 83936 5153 83959
rect 5239 83936 5305 83959
rect 4919 83896 4928 83936
rect 4968 83896 4985 83936
rect 5071 83896 5092 83936
rect 5132 83896 5153 83936
rect 5239 83896 5256 83936
rect 5296 83896 5305 83936
rect 4919 83873 4985 83896
rect 5071 83873 5153 83896
rect 5239 83873 5305 83896
rect 4919 83854 5305 83873
rect 20039 83959 20425 83978
rect 20039 83936 20105 83959
rect 20191 83936 20273 83959
rect 20359 83936 20425 83959
rect 20039 83896 20048 83936
rect 20088 83896 20105 83936
rect 20191 83896 20212 83936
rect 20252 83896 20273 83936
rect 20359 83896 20376 83936
rect 20416 83896 20425 83936
rect 20039 83873 20105 83896
rect 20191 83873 20273 83896
rect 20359 83873 20425 83896
rect 20039 83854 20425 83873
rect 8018 83539 8142 83558
rect 8018 83516 8037 83539
rect 7747 83476 7756 83516
rect 7796 83476 8037 83516
rect 8018 83453 8037 83476
rect 8123 83453 8142 83539
rect 8018 83434 8142 83453
rect 17138 83539 17262 83558
rect 17138 83453 17157 83539
rect 17243 83516 17262 83539
rect 17243 83476 19084 83516
rect 19124 83476 19133 83516
rect 17243 83453 17262 83476
rect 17138 83434 17262 83453
rect 13490 83371 13614 83390
rect 13490 83348 13509 83371
rect 13123 83308 13132 83348
rect 13172 83308 13509 83348
rect 13490 83285 13509 83308
rect 13595 83285 13614 83371
rect 13490 83266 13614 83285
rect 3679 83203 4065 83222
rect 3679 83180 3745 83203
rect 3831 83180 3913 83203
rect 3999 83180 4065 83203
rect 3679 83140 3688 83180
rect 3728 83140 3745 83180
rect 3831 83140 3852 83180
rect 3892 83140 3913 83180
rect 3999 83140 4016 83180
rect 4056 83140 4065 83180
rect 3679 83117 3745 83140
rect 3831 83117 3913 83140
rect 3999 83117 4065 83140
rect 3679 83098 4065 83117
rect 18799 83203 19185 83222
rect 18799 83180 18865 83203
rect 18951 83180 19033 83203
rect 19119 83180 19185 83203
rect 18799 83140 18808 83180
rect 18848 83140 18865 83180
rect 18951 83140 18972 83180
rect 19012 83140 19033 83180
rect 19119 83140 19136 83180
rect 19176 83140 19185 83180
rect 18799 83117 18865 83140
rect 18951 83117 19033 83140
rect 19119 83117 19185 83140
rect 18799 83098 19185 83117
rect 4919 82447 5305 82466
rect 4919 82424 4985 82447
rect 5071 82424 5153 82447
rect 5239 82424 5305 82447
rect 4919 82384 4928 82424
rect 4968 82384 4985 82424
rect 5071 82384 5092 82424
rect 5132 82384 5153 82424
rect 5239 82384 5256 82424
rect 5296 82384 5305 82424
rect 4919 82361 4985 82384
rect 5071 82361 5153 82384
rect 5239 82361 5305 82384
rect 4919 82342 5305 82361
rect 20039 82447 20425 82466
rect 20039 82424 20105 82447
rect 20191 82424 20273 82447
rect 20359 82424 20425 82447
rect 20039 82384 20048 82424
rect 20088 82384 20105 82424
rect 20191 82384 20212 82424
rect 20252 82384 20273 82424
rect 20359 82384 20376 82424
rect 20416 82384 20425 82424
rect 20039 82361 20105 82384
rect 20191 82361 20273 82384
rect 20359 82361 20425 82384
rect 20039 82342 20425 82361
rect 3679 81691 4065 81710
rect 3679 81668 3745 81691
rect 3831 81668 3913 81691
rect 3999 81668 4065 81691
rect 3679 81628 3688 81668
rect 3728 81628 3745 81668
rect 3831 81628 3852 81668
rect 3892 81628 3913 81668
rect 3999 81628 4016 81668
rect 4056 81628 4065 81668
rect 3679 81605 3745 81628
rect 3831 81605 3913 81628
rect 3999 81605 4065 81628
rect 3679 81586 4065 81605
rect 18799 81691 19185 81710
rect 18799 81668 18865 81691
rect 18951 81668 19033 81691
rect 19119 81668 19185 81691
rect 18799 81628 18808 81668
rect 18848 81628 18865 81668
rect 18951 81628 18972 81668
rect 19012 81628 19033 81668
rect 19119 81628 19136 81668
rect 19176 81628 19185 81668
rect 18799 81605 18865 81628
rect 18951 81605 19033 81628
rect 19119 81605 19185 81628
rect 18799 81586 19185 81605
rect 4919 80935 5305 80954
rect 4919 80912 4985 80935
rect 5071 80912 5153 80935
rect 5239 80912 5305 80935
rect 4919 80872 4928 80912
rect 4968 80872 4985 80912
rect 5071 80872 5092 80912
rect 5132 80872 5153 80912
rect 5239 80872 5256 80912
rect 5296 80872 5305 80912
rect 4919 80849 4985 80872
rect 5071 80849 5153 80872
rect 5239 80849 5305 80872
rect 4919 80830 5305 80849
rect 20039 80935 20425 80954
rect 20039 80912 20105 80935
rect 20191 80912 20273 80935
rect 20359 80912 20425 80935
rect 20039 80872 20048 80912
rect 20088 80872 20105 80912
rect 20191 80872 20212 80912
rect 20252 80872 20273 80912
rect 20359 80872 20376 80912
rect 20416 80872 20425 80912
rect 20039 80849 20105 80872
rect 20191 80849 20273 80872
rect 20359 80849 20425 80872
rect 20039 80830 20425 80849
rect 3679 80179 4065 80198
rect 3679 80156 3745 80179
rect 3831 80156 3913 80179
rect 3999 80156 4065 80179
rect 3679 80116 3688 80156
rect 3728 80116 3745 80156
rect 3831 80116 3852 80156
rect 3892 80116 3913 80156
rect 3999 80116 4016 80156
rect 4056 80116 4065 80156
rect 3679 80093 3745 80116
rect 3831 80093 3913 80116
rect 3999 80093 4065 80116
rect 3679 80074 4065 80093
rect 18799 80179 19185 80198
rect 18799 80156 18865 80179
rect 18951 80156 19033 80179
rect 19119 80156 19185 80179
rect 18799 80116 18808 80156
rect 18848 80116 18865 80156
rect 18951 80116 18972 80156
rect 19012 80116 19033 80156
rect 19119 80116 19136 80156
rect 19176 80116 19185 80156
rect 18799 80093 18865 80116
rect 18951 80093 19033 80116
rect 19119 80093 19185 80116
rect 18799 80074 19185 80093
rect 4919 79423 5305 79442
rect 4919 79400 4985 79423
rect 5071 79400 5153 79423
rect 5239 79400 5305 79423
rect 4919 79360 4928 79400
rect 4968 79360 4985 79400
rect 5071 79360 5092 79400
rect 5132 79360 5153 79400
rect 5239 79360 5256 79400
rect 5296 79360 5305 79400
rect 4919 79337 4985 79360
rect 5071 79337 5153 79360
rect 5239 79337 5305 79360
rect 4919 79318 5305 79337
rect 20039 79423 20425 79442
rect 20039 79400 20105 79423
rect 20191 79400 20273 79423
rect 20359 79400 20425 79423
rect 20039 79360 20048 79400
rect 20088 79360 20105 79400
rect 20191 79360 20212 79400
rect 20252 79360 20273 79400
rect 20359 79360 20376 79400
rect 20416 79360 20425 79400
rect 20039 79337 20105 79360
rect 20191 79337 20273 79360
rect 20359 79337 20425 79360
rect 20039 79318 20425 79337
rect 3679 78667 4065 78686
rect 3679 78644 3745 78667
rect 3831 78644 3913 78667
rect 3999 78644 4065 78667
rect 3679 78604 3688 78644
rect 3728 78604 3745 78644
rect 3831 78604 3852 78644
rect 3892 78604 3913 78644
rect 3999 78604 4016 78644
rect 4056 78604 4065 78644
rect 3679 78581 3745 78604
rect 3831 78581 3913 78604
rect 3999 78581 4065 78604
rect 3679 78562 4065 78581
rect 18799 78667 19185 78686
rect 18799 78644 18865 78667
rect 18951 78644 19033 78667
rect 19119 78644 19185 78667
rect 18799 78604 18808 78644
rect 18848 78604 18865 78644
rect 18951 78604 18972 78644
rect 19012 78604 19033 78644
rect 19119 78604 19136 78644
rect 19176 78604 19185 78644
rect 18799 78581 18865 78604
rect 18951 78581 19033 78604
rect 19119 78581 19185 78604
rect 18799 78562 19185 78581
rect 4919 77911 5305 77930
rect 4919 77888 4985 77911
rect 5071 77888 5153 77911
rect 5239 77888 5305 77911
rect 4919 77848 4928 77888
rect 4968 77848 4985 77888
rect 5071 77848 5092 77888
rect 5132 77848 5153 77888
rect 5239 77848 5256 77888
rect 5296 77848 5305 77888
rect 4919 77825 4985 77848
rect 5071 77825 5153 77848
rect 5239 77825 5305 77848
rect 4919 77806 5305 77825
rect 20039 77911 20425 77930
rect 20039 77888 20105 77911
rect 20191 77888 20273 77911
rect 20359 77888 20425 77911
rect 20039 77848 20048 77888
rect 20088 77848 20105 77888
rect 20191 77848 20212 77888
rect 20252 77848 20273 77888
rect 20359 77848 20376 77888
rect 20416 77848 20425 77888
rect 20039 77825 20105 77848
rect 20191 77825 20273 77848
rect 20359 77825 20425 77848
rect 20039 77806 20425 77825
rect 3679 77155 4065 77174
rect 3679 77132 3745 77155
rect 3831 77132 3913 77155
rect 3999 77132 4065 77155
rect 3679 77092 3688 77132
rect 3728 77092 3745 77132
rect 3831 77092 3852 77132
rect 3892 77092 3913 77132
rect 3999 77092 4016 77132
rect 4056 77092 4065 77132
rect 3679 77069 3745 77092
rect 3831 77069 3913 77092
rect 3999 77069 4065 77092
rect 3679 77050 4065 77069
rect 18799 77155 19185 77174
rect 18799 77132 18865 77155
rect 18951 77132 19033 77155
rect 19119 77132 19185 77155
rect 18799 77092 18808 77132
rect 18848 77092 18865 77132
rect 18951 77092 18972 77132
rect 19012 77092 19033 77132
rect 19119 77092 19136 77132
rect 19176 77092 19185 77132
rect 18799 77069 18865 77092
rect 18951 77069 19033 77092
rect 19119 77069 19185 77092
rect 18799 77050 19185 77069
rect 4919 76399 5305 76418
rect 4919 76376 4985 76399
rect 5071 76376 5153 76399
rect 5239 76376 5305 76399
rect 4919 76336 4928 76376
rect 4968 76336 4985 76376
rect 5071 76336 5092 76376
rect 5132 76336 5153 76376
rect 5239 76336 5256 76376
rect 5296 76336 5305 76376
rect 4919 76313 4985 76336
rect 5071 76313 5153 76336
rect 5239 76313 5305 76336
rect 4919 76294 5305 76313
rect 20039 76399 20425 76418
rect 20039 76376 20105 76399
rect 20191 76376 20273 76399
rect 20359 76376 20425 76399
rect 20039 76336 20048 76376
rect 20088 76336 20105 76376
rect 20191 76336 20212 76376
rect 20252 76336 20273 76376
rect 20359 76336 20376 76376
rect 20416 76336 20425 76376
rect 20039 76313 20105 76336
rect 20191 76313 20273 76336
rect 20359 76313 20425 76336
rect 20039 76294 20425 76313
rect 3679 75643 4065 75662
rect 3679 75620 3745 75643
rect 3831 75620 3913 75643
rect 3999 75620 4065 75643
rect 3679 75580 3688 75620
rect 3728 75580 3745 75620
rect 3831 75580 3852 75620
rect 3892 75580 3913 75620
rect 3999 75580 4016 75620
rect 4056 75580 4065 75620
rect 3679 75557 3745 75580
rect 3831 75557 3913 75580
rect 3999 75557 4065 75580
rect 3679 75538 4065 75557
rect 18799 75643 19185 75662
rect 18799 75620 18865 75643
rect 18951 75620 19033 75643
rect 19119 75620 19185 75643
rect 18799 75580 18808 75620
rect 18848 75580 18865 75620
rect 18951 75580 18972 75620
rect 19012 75580 19033 75620
rect 19119 75580 19136 75620
rect 19176 75580 19185 75620
rect 18799 75557 18865 75580
rect 18951 75557 19033 75580
rect 19119 75557 19185 75580
rect 18799 75538 19185 75557
rect 4919 74887 5305 74906
rect 4919 74864 4985 74887
rect 5071 74864 5153 74887
rect 5239 74864 5305 74887
rect 4919 74824 4928 74864
rect 4968 74824 4985 74864
rect 5071 74824 5092 74864
rect 5132 74824 5153 74864
rect 5239 74824 5256 74864
rect 5296 74824 5305 74864
rect 4919 74801 4985 74824
rect 5071 74801 5153 74824
rect 5239 74801 5305 74824
rect 4919 74782 5305 74801
rect 20039 74887 20425 74906
rect 20039 74864 20105 74887
rect 20191 74864 20273 74887
rect 20359 74864 20425 74887
rect 20039 74824 20048 74864
rect 20088 74824 20105 74864
rect 20191 74824 20212 74864
rect 20252 74824 20273 74864
rect 20359 74824 20376 74864
rect 20416 74824 20425 74864
rect 20039 74801 20105 74824
rect 20191 74801 20273 74824
rect 20359 74801 20425 74824
rect 20039 74782 20425 74801
rect 3679 74131 4065 74150
rect 3679 74108 3745 74131
rect 3831 74108 3913 74131
rect 3999 74108 4065 74131
rect 3679 74068 3688 74108
rect 3728 74068 3745 74108
rect 3831 74068 3852 74108
rect 3892 74068 3913 74108
rect 3999 74068 4016 74108
rect 4056 74068 4065 74108
rect 3679 74045 3745 74068
rect 3831 74045 3913 74068
rect 3999 74045 4065 74068
rect 3679 74026 4065 74045
rect 18799 74131 19185 74150
rect 18799 74108 18865 74131
rect 18951 74108 19033 74131
rect 19119 74108 19185 74131
rect 18799 74068 18808 74108
rect 18848 74068 18865 74108
rect 18951 74068 18972 74108
rect 19012 74068 19033 74108
rect 19119 74068 19136 74108
rect 19176 74068 19185 74108
rect 18799 74045 18865 74068
rect 18951 74045 19033 74068
rect 19119 74045 19185 74068
rect 18799 74026 19185 74045
rect 4919 73375 5305 73394
rect 4919 73352 4985 73375
rect 5071 73352 5153 73375
rect 5239 73352 5305 73375
rect 4919 73312 4928 73352
rect 4968 73312 4985 73352
rect 5071 73312 5092 73352
rect 5132 73312 5153 73352
rect 5239 73312 5256 73352
rect 5296 73312 5305 73352
rect 4919 73289 4985 73312
rect 5071 73289 5153 73312
rect 5239 73289 5305 73312
rect 4919 73270 5305 73289
rect 20039 73375 20425 73394
rect 20039 73352 20105 73375
rect 20191 73352 20273 73375
rect 20359 73352 20425 73375
rect 20039 73312 20048 73352
rect 20088 73312 20105 73352
rect 20191 73312 20212 73352
rect 20252 73312 20273 73352
rect 20359 73312 20376 73352
rect 20416 73312 20425 73352
rect 20039 73289 20105 73312
rect 20191 73289 20273 73312
rect 20359 73289 20425 73312
rect 20039 73270 20425 73289
rect 15314 72787 15438 72806
rect 15314 72764 15333 72787
rect 10723 72724 10732 72764
rect 10772 72724 15333 72764
rect 15314 72701 15333 72724
rect 15419 72701 15438 72787
rect 15314 72682 15438 72701
rect 3679 72619 4065 72638
rect 3679 72596 3745 72619
rect 3831 72596 3913 72619
rect 3999 72596 4065 72619
rect 3679 72556 3688 72596
rect 3728 72556 3745 72596
rect 3831 72556 3852 72596
rect 3892 72556 3913 72596
rect 3999 72556 4016 72596
rect 4056 72556 4065 72596
rect 3679 72533 3745 72556
rect 3831 72533 3913 72556
rect 3999 72533 4065 72556
rect 3679 72514 4065 72533
rect 18799 72619 19185 72638
rect 18799 72596 18865 72619
rect 18951 72596 19033 72619
rect 19119 72596 19185 72619
rect 18799 72556 18808 72596
rect 18848 72556 18865 72596
rect 18951 72556 18972 72596
rect 19012 72556 19033 72596
rect 19119 72556 19136 72596
rect 19176 72556 19185 72596
rect 18799 72533 18865 72556
rect 18951 72533 19033 72556
rect 19119 72533 19185 72556
rect 18799 72514 19185 72533
rect 12122 72199 12246 72218
rect 12122 72113 12141 72199
rect 12227 72176 12246 72199
rect 12227 72136 12460 72176
rect 12500 72136 12509 72176
rect 12227 72113 12246 72136
rect 12122 72094 12246 72113
rect 4919 71863 5305 71882
rect 4919 71840 4985 71863
rect 5071 71840 5153 71863
rect 5239 71840 5305 71863
rect 4919 71800 4928 71840
rect 4968 71800 4985 71840
rect 5071 71800 5092 71840
rect 5132 71800 5153 71840
rect 5239 71800 5256 71840
rect 5296 71800 5305 71840
rect 4919 71777 4985 71800
rect 5071 71777 5153 71800
rect 5239 71777 5305 71800
rect 4919 71758 5305 71777
rect 20039 71863 20425 71882
rect 20039 71840 20105 71863
rect 20191 71840 20273 71863
rect 20359 71840 20425 71863
rect 20039 71800 20048 71840
rect 20088 71800 20105 71840
rect 20191 71800 20212 71840
rect 20252 71800 20273 71840
rect 20359 71800 20376 71840
rect 20416 71800 20425 71840
rect 20039 71777 20105 71800
rect 20191 71777 20273 71800
rect 20359 71777 20425 71800
rect 20039 71758 20425 71777
rect 3679 71107 4065 71126
rect 3679 71084 3745 71107
rect 3831 71084 3913 71107
rect 3999 71084 4065 71107
rect 3679 71044 3688 71084
rect 3728 71044 3745 71084
rect 3831 71044 3852 71084
rect 3892 71044 3913 71084
rect 3999 71044 4016 71084
rect 4056 71044 4065 71084
rect 3679 71021 3745 71044
rect 3831 71021 3913 71044
rect 3999 71021 4065 71044
rect 3679 71002 4065 71021
rect 18799 71107 19185 71126
rect 18799 71084 18865 71107
rect 18951 71084 19033 71107
rect 19119 71084 19185 71107
rect 18799 71044 18808 71084
rect 18848 71044 18865 71084
rect 18951 71044 18972 71084
rect 19012 71044 19033 71084
rect 19119 71044 19136 71084
rect 19176 71044 19185 71084
rect 18799 71021 18865 71044
rect 18951 71021 19033 71044
rect 19119 71021 19185 71044
rect 18799 71002 19185 71021
rect 4919 70351 5305 70370
rect 4919 70328 4985 70351
rect 5071 70328 5153 70351
rect 5239 70328 5305 70351
rect 4919 70288 4928 70328
rect 4968 70288 4985 70328
rect 5071 70288 5092 70328
rect 5132 70288 5153 70328
rect 5239 70288 5256 70328
rect 5296 70288 5305 70328
rect 4919 70265 4985 70288
rect 5071 70265 5153 70288
rect 5239 70265 5305 70288
rect 4919 70246 5305 70265
rect 20039 70351 20425 70370
rect 20039 70328 20105 70351
rect 20191 70328 20273 70351
rect 20359 70328 20425 70351
rect 20039 70288 20048 70328
rect 20088 70288 20105 70328
rect 20191 70288 20212 70328
rect 20252 70288 20273 70328
rect 20359 70288 20376 70328
rect 20416 70288 20425 70328
rect 20039 70265 20105 70288
rect 20191 70265 20273 70288
rect 20359 70265 20425 70288
rect 20039 70246 20425 70265
rect 3679 69595 4065 69614
rect 3679 69572 3745 69595
rect 3831 69572 3913 69595
rect 3999 69572 4065 69595
rect 3679 69532 3688 69572
rect 3728 69532 3745 69572
rect 3831 69532 3852 69572
rect 3892 69532 3913 69572
rect 3999 69532 4016 69572
rect 4056 69532 4065 69572
rect 3679 69509 3745 69532
rect 3831 69509 3913 69532
rect 3999 69509 4065 69532
rect 3679 69490 4065 69509
rect 18799 69595 19185 69614
rect 18799 69572 18865 69595
rect 18951 69572 19033 69595
rect 19119 69572 19185 69595
rect 18799 69532 18808 69572
rect 18848 69532 18865 69572
rect 18951 69532 18972 69572
rect 19012 69532 19033 69572
rect 19119 69532 19136 69572
rect 19176 69532 19185 69572
rect 18799 69509 18865 69532
rect 18951 69509 19033 69532
rect 19119 69509 19185 69532
rect 18799 69490 19185 69509
rect 11210 69343 11334 69362
rect 11210 69320 11229 69343
rect 10339 69280 10348 69320
rect 10388 69280 11229 69320
rect 11210 69257 11229 69280
rect 11315 69257 11334 69343
rect 11210 69238 11334 69257
rect 4919 68839 5305 68858
rect 4919 68816 4985 68839
rect 5071 68816 5153 68839
rect 5239 68816 5305 68839
rect 4919 68776 4928 68816
rect 4968 68776 4985 68816
rect 5071 68776 5092 68816
rect 5132 68776 5153 68816
rect 5239 68776 5256 68816
rect 5296 68776 5305 68816
rect 4919 68753 4985 68776
rect 5071 68753 5153 68776
rect 5239 68753 5305 68776
rect 4919 68734 5305 68753
rect 20039 68839 20425 68858
rect 20039 68816 20105 68839
rect 20191 68816 20273 68839
rect 20359 68816 20425 68839
rect 20039 68776 20048 68816
rect 20088 68776 20105 68816
rect 20191 68776 20212 68816
rect 20252 68776 20273 68816
rect 20359 68776 20376 68816
rect 20416 68776 20425 68816
rect 20039 68753 20105 68776
rect 20191 68753 20273 68776
rect 20359 68753 20425 68776
rect 20039 68734 20425 68753
rect 3619 68524 3628 68564
rect 3668 68524 4876 68564
rect 4916 68524 4925 68564
rect 3679 68083 4065 68102
rect 3679 68060 3745 68083
rect 3831 68060 3913 68083
rect 3999 68060 4065 68083
rect 3679 68020 3688 68060
rect 3728 68020 3745 68060
rect 3831 68020 3852 68060
rect 3892 68020 3913 68060
rect 3999 68020 4016 68060
rect 4056 68020 4065 68060
rect 3679 67997 3745 68020
rect 3831 67997 3913 68020
rect 3999 67997 4065 68020
rect 3679 67978 4065 67997
rect 18799 68083 19185 68102
rect 18799 68060 18865 68083
rect 18951 68060 19033 68083
rect 19119 68060 19185 68083
rect 18799 68020 18808 68060
rect 18848 68020 18865 68060
rect 18951 68020 18972 68060
rect 19012 68020 19033 68060
rect 19119 68020 19136 68060
rect 19176 68020 19185 68060
rect 18799 67997 18865 68020
rect 18951 67997 19033 68020
rect 19119 67997 19185 68020
rect 18799 67978 19185 67997
rect 8707 67768 8716 67808
rect 8756 67768 20140 67808
rect 20180 67768 20189 67808
rect 1027 67432 1036 67472
rect 1076 67432 3820 67472
rect 3860 67432 3869 67472
rect 4919 67327 5305 67346
rect 4919 67304 4985 67327
rect 5071 67304 5153 67327
rect 5239 67304 5305 67327
rect 4919 67264 4928 67304
rect 4968 67264 4985 67304
rect 5071 67264 5092 67304
rect 5132 67264 5153 67304
rect 5239 67264 5256 67304
rect 5296 67264 5305 67304
rect 4919 67241 4985 67264
rect 5071 67241 5153 67264
rect 5239 67241 5305 67264
rect 4919 67222 5305 67241
rect 20039 67327 20425 67346
rect 20039 67304 20105 67327
rect 20191 67304 20273 67327
rect 20359 67304 20425 67327
rect 20039 67264 20048 67304
rect 20088 67264 20105 67304
rect 20191 67264 20212 67304
rect 20252 67264 20273 67304
rect 20359 67264 20376 67304
rect 20416 67264 20425 67304
rect 20039 67241 20105 67264
rect 20191 67241 20273 67264
rect 20359 67241 20425 67264
rect 20039 67222 20425 67241
rect 3679 66571 4065 66590
rect 3679 66548 3745 66571
rect 3831 66548 3913 66571
rect 3999 66548 4065 66571
rect 3679 66508 3688 66548
rect 3728 66508 3745 66548
rect 3831 66508 3852 66548
rect 3892 66508 3913 66548
rect 3999 66508 4016 66548
rect 4056 66508 4065 66548
rect 3679 66485 3745 66508
rect 3831 66485 3913 66508
rect 3999 66485 4065 66508
rect 3679 66466 4065 66485
rect 18799 66571 19185 66590
rect 18799 66548 18865 66571
rect 18951 66548 19033 66571
rect 19119 66548 19185 66571
rect 18799 66508 18808 66548
rect 18848 66508 18865 66548
rect 18951 66508 18972 66548
rect 19012 66508 19033 66548
rect 19119 66508 19136 66548
rect 19176 66508 19185 66548
rect 18799 66485 18865 66508
rect 18951 66485 19033 66508
rect 19119 66485 19185 66508
rect 18799 66466 19185 66485
rect 1123 66340 1132 66380
rect 1172 66340 13804 66380
rect 13844 66340 13853 66380
rect 4919 65815 5305 65834
rect 4919 65792 4985 65815
rect 5071 65792 5153 65815
rect 5239 65792 5305 65815
rect 4919 65752 4928 65792
rect 4968 65752 4985 65792
rect 5071 65752 5092 65792
rect 5132 65752 5153 65792
rect 5239 65752 5256 65792
rect 5296 65752 5305 65792
rect 4919 65729 4985 65752
rect 5071 65729 5153 65752
rect 5239 65729 5305 65752
rect 4919 65710 5305 65729
rect 20039 65815 20425 65834
rect 20039 65792 20105 65815
rect 20191 65792 20273 65815
rect 20359 65792 20425 65815
rect 20039 65752 20048 65792
rect 20088 65752 20105 65792
rect 20191 65752 20212 65792
rect 20252 65752 20273 65792
rect 20359 65752 20376 65792
rect 20416 65752 20425 65792
rect 20039 65729 20105 65752
rect 20191 65729 20273 65752
rect 20359 65729 20425 65752
rect 20039 65710 20425 65729
rect 3679 65059 4065 65078
rect 3679 65036 3745 65059
rect 3831 65036 3913 65059
rect 3999 65036 4065 65059
rect 3679 64996 3688 65036
rect 3728 64996 3745 65036
rect 3831 64996 3852 65036
rect 3892 64996 3913 65036
rect 3999 64996 4016 65036
rect 4056 64996 4065 65036
rect 3679 64973 3745 64996
rect 3831 64973 3913 64996
rect 3999 64973 4065 64996
rect 3679 64954 4065 64973
rect 18799 65059 19185 65078
rect 18799 65036 18865 65059
rect 18951 65036 19033 65059
rect 19119 65036 19185 65059
rect 18799 64996 18808 65036
rect 18848 64996 18865 65036
rect 18951 64996 18972 65036
rect 19012 64996 19033 65036
rect 19119 64996 19136 65036
rect 19176 64996 19185 65036
rect 18799 64973 18865 64996
rect 18951 64973 19033 64996
rect 19119 64973 19185 64996
rect 18799 64954 19185 64973
rect 1178 64471 1302 64490
rect 1178 64385 1197 64471
rect 1283 64448 1302 64471
rect 1283 64408 5836 64448
rect 5876 64408 5885 64448
rect 1283 64385 1302 64408
rect 1178 64366 1302 64385
rect 4919 64303 5305 64322
rect 4919 64280 4985 64303
rect 5071 64280 5153 64303
rect 5239 64280 5305 64303
rect 4919 64240 4928 64280
rect 4968 64240 4985 64280
rect 5071 64240 5092 64280
rect 5132 64240 5153 64280
rect 5239 64240 5256 64280
rect 5296 64240 5305 64280
rect 4919 64217 4985 64240
rect 5071 64217 5153 64240
rect 5239 64217 5305 64240
rect 4919 64198 5305 64217
rect 20039 64303 20425 64322
rect 20039 64280 20105 64303
rect 20191 64280 20273 64303
rect 20359 64280 20425 64303
rect 20039 64240 20048 64280
rect 20088 64240 20105 64280
rect 20191 64240 20212 64280
rect 20252 64240 20273 64280
rect 20359 64240 20376 64280
rect 20416 64240 20425 64280
rect 20039 64217 20105 64240
rect 20191 64217 20273 64240
rect 20359 64217 20425 64240
rect 20039 64198 20425 64217
rect 3679 63547 4065 63566
rect 3679 63524 3745 63547
rect 3831 63524 3913 63547
rect 3999 63524 4065 63547
rect 3679 63484 3688 63524
rect 3728 63484 3745 63524
rect 3831 63484 3852 63524
rect 3892 63484 3913 63524
rect 3999 63484 4016 63524
rect 4056 63484 4065 63524
rect 3679 63461 3745 63484
rect 3831 63461 3913 63484
rect 3999 63461 4065 63484
rect 3679 63442 4065 63461
rect 18799 63547 19185 63566
rect 18799 63524 18865 63547
rect 18951 63524 19033 63547
rect 19119 63524 19185 63547
rect 18799 63484 18808 63524
rect 18848 63484 18865 63524
rect 18951 63484 18972 63524
rect 19012 63484 19033 63524
rect 19119 63484 19136 63524
rect 19176 63484 19185 63524
rect 18799 63461 18865 63484
rect 18951 63461 19033 63484
rect 19119 63461 19185 63484
rect 18799 63442 19185 63461
rect 9842 63043 9966 63062
rect 643 62980 652 63020
rect 692 62980 4492 63020
rect 4532 62980 4541 63020
rect 9842 62957 9861 63043
rect 9947 63020 9966 63043
rect 9947 62980 9964 63020
rect 10004 62980 10013 63020
rect 9947 62957 9966 62980
rect 9842 62938 9966 62957
rect 4919 62791 5305 62810
rect 4919 62768 4985 62791
rect 5071 62768 5153 62791
rect 5239 62768 5305 62791
rect 4919 62728 4928 62768
rect 4968 62728 4985 62768
rect 5071 62728 5092 62768
rect 5132 62728 5153 62768
rect 5239 62728 5256 62768
rect 5296 62728 5305 62768
rect 4919 62705 4985 62728
rect 5071 62705 5153 62728
rect 5239 62705 5305 62728
rect 4919 62686 5305 62705
rect 20039 62791 20425 62810
rect 20039 62768 20105 62791
rect 20191 62768 20273 62791
rect 20359 62768 20425 62791
rect 20039 62728 20048 62768
rect 20088 62728 20105 62768
rect 20191 62728 20212 62768
rect 20252 62728 20273 62768
rect 20359 62728 20376 62768
rect 20416 62728 20425 62768
rect 20039 62705 20105 62728
rect 20191 62705 20273 62728
rect 20359 62705 20425 62728
rect 20039 62686 20425 62705
rect 3679 62035 4065 62054
rect 3679 62012 3745 62035
rect 3831 62012 3913 62035
rect 3999 62012 4065 62035
rect 3679 61972 3688 62012
rect 3728 61972 3745 62012
rect 3831 61972 3852 62012
rect 3892 61972 3913 62012
rect 3999 61972 4016 62012
rect 4056 61972 4065 62012
rect 3679 61949 3745 61972
rect 3831 61949 3913 61972
rect 3999 61949 4065 61972
rect 3679 61930 4065 61949
rect 18799 62035 19185 62054
rect 18799 62012 18865 62035
rect 18951 62012 19033 62035
rect 19119 62012 19185 62035
rect 18799 61972 18808 62012
rect 18848 61972 18865 62012
rect 18951 61972 18972 62012
rect 19012 61972 19033 62012
rect 19119 61972 19136 62012
rect 19176 61972 19185 62012
rect 18799 61949 18865 61972
rect 18951 61949 19033 61972
rect 19119 61949 19185 61972
rect 18799 61930 19185 61949
rect 2563 61720 2572 61760
rect 2612 61720 3916 61760
rect 3956 61720 3965 61760
rect 13027 61300 13036 61340
rect 13076 61300 16012 61340
rect 16052 61300 16061 61340
rect 4919 61279 5305 61298
rect 4919 61256 4985 61279
rect 5071 61256 5153 61279
rect 5239 61256 5305 61279
rect 4919 61216 4928 61256
rect 4968 61216 4985 61256
rect 5071 61216 5092 61256
rect 5132 61216 5153 61256
rect 5239 61216 5256 61256
rect 5296 61216 5305 61256
rect 4919 61193 4985 61216
rect 5071 61193 5153 61216
rect 5239 61193 5305 61216
rect 4919 61174 5305 61193
rect 20039 61279 20425 61298
rect 20039 61256 20105 61279
rect 20191 61256 20273 61279
rect 20359 61256 20425 61279
rect 20039 61216 20048 61256
rect 20088 61216 20105 61256
rect 20191 61216 20212 61256
rect 20252 61216 20273 61256
rect 20359 61216 20376 61256
rect 20416 61216 20425 61256
rect 20039 61193 20105 61216
rect 20191 61193 20273 61216
rect 20359 61193 20425 61216
rect 20039 61174 20425 61193
rect 2467 60964 2476 61004
rect 2516 60964 4588 61004
rect 4628 60964 4637 61004
rect 3679 60523 4065 60542
rect 3679 60500 3745 60523
rect 3831 60500 3913 60523
rect 3999 60500 4065 60523
rect 3679 60460 3688 60500
rect 3728 60460 3745 60500
rect 3831 60460 3852 60500
rect 3892 60460 3913 60500
rect 3999 60460 4016 60500
rect 4056 60460 4065 60500
rect 3679 60437 3745 60460
rect 3831 60437 3913 60460
rect 3999 60437 4065 60460
rect 3679 60418 4065 60437
rect 18799 60523 19185 60542
rect 18799 60500 18865 60523
rect 18951 60500 19033 60523
rect 19119 60500 19185 60523
rect 18799 60460 18808 60500
rect 18848 60460 18865 60500
rect 18951 60460 18972 60500
rect 19012 60460 19033 60500
rect 19119 60460 19136 60500
rect 19176 60460 19185 60500
rect 18799 60437 18865 60460
rect 18951 60437 19033 60460
rect 19119 60437 19185 60460
rect 18799 60418 19185 60437
rect 4919 59767 5305 59786
rect 4919 59744 4985 59767
rect 5071 59744 5153 59767
rect 5239 59744 5305 59767
rect 4919 59704 4928 59744
rect 4968 59704 4985 59744
rect 5071 59704 5092 59744
rect 5132 59704 5153 59744
rect 5239 59704 5256 59744
rect 5296 59704 5305 59744
rect 4919 59681 4985 59704
rect 5071 59681 5153 59704
rect 5239 59681 5305 59704
rect 4919 59662 5305 59681
rect 20039 59767 20425 59786
rect 20039 59744 20105 59767
rect 20191 59744 20273 59767
rect 20359 59744 20425 59767
rect 20039 59704 20048 59744
rect 20088 59704 20105 59744
rect 20191 59704 20212 59744
rect 20252 59704 20273 59744
rect 20359 59704 20376 59744
rect 20416 59704 20425 59744
rect 20039 59681 20105 59704
rect 20191 59681 20273 59704
rect 20359 59681 20425 59704
rect 20039 59662 20425 59681
rect 3679 59011 4065 59030
rect 3679 58988 3745 59011
rect 3831 58988 3913 59011
rect 3999 58988 4065 59011
rect 3679 58948 3688 58988
rect 3728 58948 3745 58988
rect 3831 58948 3852 58988
rect 3892 58948 3913 58988
rect 3999 58948 4016 58988
rect 4056 58948 4065 58988
rect 3679 58925 3745 58948
rect 3831 58925 3913 58948
rect 3999 58925 4065 58948
rect 3679 58906 4065 58925
rect 18799 59011 19185 59030
rect 18799 58988 18865 59011
rect 18951 58988 19033 59011
rect 19119 58988 19185 59011
rect 18799 58948 18808 58988
rect 18848 58948 18865 58988
rect 18951 58948 18972 58988
rect 19012 58948 19033 58988
rect 19119 58948 19136 58988
rect 19176 58948 19185 58988
rect 18799 58925 18865 58948
rect 18951 58925 19033 58948
rect 19119 58925 19185 58948
rect 18799 58906 19185 58925
rect 15331 58864 15340 58904
rect 15380 58864 16012 58904
rect 16052 58864 16061 58904
rect 4919 58255 5305 58274
rect 4919 58232 4985 58255
rect 5071 58232 5153 58255
rect 5239 58232 5305 58255
rect 4919 58192 4928 58232
rect 4968 58192 4985 58232
rect 5071 58192 5092 58232
rect 5132 58192 5153 58232
rect 5239 58192 5256 58232
rect 5296 58192 5305 58232
rect 4919 58169 4985 58192
rect 5071 58169 5153 58192
rect 5239 58169 5305 58192
rect 4919 58150 5305 58169
rect 20039 58255 20425 58274
rect 20039 58232 20105 58255
rect 20191 58232 20273 58255
rect 20359 58232 20425 58255
rect 20039 58192 20048 58232
rect 20088 58192 20105 58232
rect 20191 58192 20212 58232
rect 20252 58192 20273 58232
rect 20359 58192 20376 58232
rect 20416 58192 20425 58232
rect 20039 58169 20105 58192
rect 20191 58169 20273 58192
rect 20359 58169 20425 58192
rect 20039 58150 20425 58169
rect 3679 57499 4065 57518
rect 3679 57476 3745 57499
rect 3831 57476 3913 57499
rect 3999 57476 4065 57499
rect 3679 57436 3688 57476
rect 3728 57436 3745 57476
rect 3831 57436 3852 57476
rect 3892 57436 3913 57476
rect 3999 57436 4016 57476
rect 4056 57436 4065 57476
rect 3679 57413 3745 57436
rect 3831 57413 3913 57436
rect 3999 57413 4065 57436
rect 3679 57394 4065 57413
rect 18799 57499 19185 57518
rect 18799 57476 18865 57499
rect 18951 57476 19033 57499
rect 19119 57476 19185 57499
rect 18799 57436 18808 57476
rect 18848 57436 18865 57476
rect 18951 57436 18972 57476
rect 19012 57436 19033 57476
rect 19119 57436 19136 57476
rect 19176 57436 19185 57476
rect 18799 57413 18865 57436
rect 18951 57413 19033 57436
rect 19119 57413 19185 57436
rect 18799 57394 19185 57413
rect 4919 56743 5305 56762
rect 4919 56720 4985 56743
rect 5071 56720 5153 56743
rect 5239 56720 5305 56743
rect 4919 56680 4928 56720
rect 4968 56680 4985 56720
rect 5071 56680 5092 56720
rect 5132 56680 5153 56720
rect 5239 56680 5256 56720
rect 5296 56680 5305 56720
rect 4919 56657 4985 56680
rect 5071 56657 5153 56680
rect 5239 56657 5305 56680
rect 4919 56638 5305 56657
rect 20039 56743 20425 56762
rect 20039 56720 20105 56743
rect 20191 56720 20273 56743
rect 20359 56720 20425 56743
rect 20039 56680 20048 56720
rect 20088 56680 20105 56720
rect 20191 56680 20212 56720
rect 20252 56680 20273 56720
rect 20359 56680 20376 56720
rect 20416 56680 20425 56720
rect 20039 56657 20105 56680
rect 20191 56657 20273 56680
rect 20359 56657 20425 56680
rect 20039 56638 20425 56657
rect 3679 55987 4065 56006
rect 3679 55964 3745 55987
rect 3831 55964 3913 55987
rect 3999 55964 4065 55987
rect 3679 55924 3688 55964
rect 3728 55924 3745 55964
rect 3831 55924 3852 55964
rect 3892 55924 3913 55964
rect 3999 55924 4016 55964
rect 4056 55924 4065 55964
rect 3679 55901 3745 55924
rect 3831 55901 3913 55924
rect 3999 55901 4065 55924
rect 3679 55882 4065 55901
rect 18799 55987 19185 56006
rect 18799 55964 18865 55987
rect 18951 55964 19033 55987
rect 19119 55964 19185 55987
rect 18799 55924 18808 55964
rect 18848 55924 18865 55964
rect 18951 55924 18972 55964
rect 19012 55924 19033 55964
rect 19119 55924 19136 55964
rect 19176 55924 19185 55964
rect 18799 55901 18865 55924
rect 18951 55901 19033 55924
rect 19119 55901 19185 55924
rect 18799 55882 19185 55901
rect 4919 55231 5305 55250
rect 4919 55208 4985 55231
rect 5071 55208 5153 55231
rect 5239 55208 5305 55231
rect 4919 55168 4928 55208
rect 4968 55168 4985 55208
rect 5071 55168 5092 55208
rect 5132 55168 5153 55208
rect 5239 55168 5256 55208
rect 5296 55168 5305 55208
rect 4919 55145 4985 55168
rect 5071 55145 5153 55168
rect 5239 55145 5305 55168
rect 4919 55126 5305 55145
rect 20039 55231 20425 55250
rect 20039 55208 20105 55231
rect 20191 55208 20273 55231
rect 20359 55208 20425 55231
rect 20039 55168 20048 55208
rect 20088 55168 20105 55208
rect 20191 55168 20212 55208
rect 20252 55168 20273 55208
rect 20359 55168 20376 55208
rect 20416 55168 20425 55208
rect 20039 55145 20105 55168
rect 20191 55145 20273 55168
rect 20359 55145 20425 55168
rect 20039 55126 20425 55145
rect 3679 54475 4065 54494
rect 3679 54452 3745 54475
rect 3831 54452 3913 54475
rect 3999 54452 4065 54475
rect 3679 54412 3688 54452
rect 3728 54412 3745 54452
rect 3831 54412 3852 54452
rect 3892 54412 3913 54452
rect 3999 54412 4016 54452
rect 4056 54412 4065 54452
rect 3679 54389 3745 54412
rect 3831 54389 3913 54412
rect 3999 54389 4065 54412
rect 3679 54370 4065 54389
rect 18799 54475 19185 54494
rect 18799 54452 18865 54475
rect 18951 54452 19033 54475
rect 19119 54452 19185 54475
rect 18799 54412 18808 54452
rect 18848 54412 18865 54452
rect 18951 54412 18972 54452
rect 19012 54412 19033 54452
rect 19119 54412 19136 54452
rect 19176 54412 19185 54452
rect 18799 54389 18865 54412
rect 18951 54389 19033 54412
rect 19119 54389 19185 54412
rect 18799 54370 19185 54389
rect 4919 53719 5305 53738
rect 4919 53696 4985 53719
rect 5071 53696 5153 53719
rect 5239 53696 5305 53719
rect 4919 53656 4928 53696
rect 4968 53656 4985 53696
rect 5071 53656 5092 53696
rect 5132 53656 5153 53696
rect 5239 53656 5256 53696
rect 5296 53656 5305 53696
rect 4919 53633 4985 53656
rect 5071 53633 5153 53656
rect 5239 53633 5305 53656
rect 4919 53614 5305 53633
rect 20039 53719 20425 53738
rect 20039 53696 20105 53719
rect 20191 53696 20273 53719
rect 20359 53696 20425 53719
rect 20039 53656 20048 53696
rect 20088 53656 20105 53696
rect 20191 53656 20212 53696
rect 20252 53656 20273 53696
rect 20359 53656 20376 53696
rect 20416 53656 20425 53696
rect 20039 53633 20105 53656
rect 20191 53633 20273 53656
rect 20359 53633 20425 53656
rect 20039 53614 20425 53633
rect 3679 52963 4065 52982
rect 3679 52940 3745 52963
rect 3831 52940 3913 52963
rect 3999 52940 4065 52963
rect 3679 52900 3688 52940
rect 3728 52900 3745 52940
rect 3831 52900 3852 52940
rect 3892 52900 3913 52940
rect 3999 52900 4016 52940
rect 4056 52900 4065 52940
rect 3679 52877 3745 52900
rect 3831 52877 3913 52900
rect 3999 52877 4065 52900
rect 3679 52858 4065 52877
rect 18799 52963 19185 52982
rect 18799 52940 18865 52963
rect 18951 52940 19033 52963
rect 19119 52940 19185 52963
rect 18799 52900 18808 52940
rect 18848 52900 18865 52940
rect 18951 52900 18972 52940
rect 19012 52900 19033 52940
rect 19119 52900 19136 52940
rect 19176 52900 19185 52940
rect 18799 52877 18865 52900
rect 18951 52877 19033 52900
rect 19119 52877 19185 52900
rect 18799 52858 19185 52877
rect 4919 52207 5305 52226
rect 4919 52184 4985 52207
rect 5071 52184 5153 52207
rect 5239 52184 5305 52207
rect 4919 52144 4928 52184
rect 4968 52144 4985 52184
rect 5071 52144 5092 52184
rect 5132 52144 5153 52184
rect 5239 52144 5256 52184
rect 5296 52144 5305 52184
rect 4919 52121 4985 52144
rect 5071 52121 5153 52144
rect 5239 52121 5305 52144
rect 4919 52102 5305 52121
rect 20039 52207 20425 52226
rect 20039 52184 20105 52207
rect 20191 52184 20273 52207
rect 20359 52184 20425 52207
rect 20039 52144 20048 52184
rect 20088 52144 20105 52184
rect 20191 52144 20212 52184
rect 20252 52144 20273 52184
rect 20359 52144 20376 52184
rect 20416 52144 20425 52184
rect 20039 52121 20105 52144
rect 20191 52121 20273 52144
rect 20359 52121 20425 52144
rect 20039 52102 20425 52121
rect 3679 51451 4065 51470
rect 3679 51428 3745 51451
rect 3831 51428 3913 51451
rect 3999 51428 4065 51451
rect 3679 51388 3688 51428
rect 3728 51388 3745 51428
rect 3831 51388 3852 51428
rect 3892 51388 3913 51428
rect 3999 51388 4016 51428
rect 4056 51388 4065 51428
rect 3679 51365 3745 51388
rect 3831 51365 3913 51388
rect 3999 51365 4065 51388
rect 3679 51346 4065 51365
rect 18799 51451 19185 51470
rect 18799 51428 18865 51451
rect 18951 51428 19033 51451
rect 19119 51428 19185 51451
rect 18799 51388 18808 51428
rect 18848 51388 18865 51428
rect 18951 51388 18972 51428
rect 19012 51388 19033 51428
rect 19119 51388 19136 51428
rect 19176 51388 19185 51428
rect 18799 51365 18865 51388
rect 18951 51365 19033 51388
rect 19119 51365 19185 51388
rect 18799 51346 19185 51365
rect 4919 50695 5305 50714
rect 4919 50672 4985 50695
rect 5071 50672 5153 50695
rect 5239 50672 5305 50695
rect 4919 50632 4928 50672
rect 4968 50632 4985 50672
rect 5071 50632 5092 50672
rect 5132 50632 5153 50672
rect 5239 50632 5256 50672
rect 5296 50632 5305 50672
rect 4919 50609 4985 50632
rect 5071 50609 5153 50632
rect 5239 50609 5305 50632
rect 4919 50590 5305 50609
rect 20039 50695 20425 50714
rect 20039 50672 20105 50695
rect 20191 50672 20273 50695
rect 20359 50672 20425 50695
rect 20039 50632 20048 50672
rect 20088 50632 20105 50672
rect 20191 50632 20212 50672
rect 20252 50632 20273 50672
rect 20359 50632 20376 50672
rect 20416 50632 20425 50672
rect 20039 50609 20105 50632
rect 20191 50609 20273 50632
rect 20359 50609 20425 50632
rect 20039 50590 20425 50609
rect 3679 49939 4065 49958
rect 3679 49916 3745 49939
rect 3831 49916 3913 49939
rect 3999 49916 4065 49939
rect 3679 49876 3688 49916
rect 3728 49876 3745 49916
rect 3831 49876 3852 49916
rect 3892 49876 3913 49916
rect 3999 49876 4016 49916
rect 4056 49876 4065 49916
rect 3679 49853 3745 49876
rect 3831 49853 3913 49876
rect 3999 49853 4065 49876
rect 3679 49834 4065 49853
rect 18799 49939 19185 49958
rect 18799 49916 18865 49939
rect 18951 49916 19033 49939
rect 19119 49916 19185 49939
rect 18799 49876 18808 49916
rect 18848 49876 18865 49916
rect 18951 49876 18972 49916
rect 19012 49876 19033 49916
rect 19119 49876 19136 49916
rect 19176 49876 19185 49916
rect 18799 49853 18865 49876
rect 18951 49853 19033 49876
rect 19119 49853 19185 49876
rect 18799 49834 19185 49853
rect 4919 49183 5305 49202
rect 4919 49160 4985 49183
rect 5071 49160 5153 49183
rect 5239 49160 5305 49183
rect 4919 49120 4928 49160
rect 4968 49120 4985 49160
rect 5071 49120 5092 49160
rect 5132 49120 5153 49160
rect 5239 49120 5256 49160
rect 5296 49120 5305 49160
rect 4919 49097 4985 49120
rect 5071 49097 5153 49120
rect 5239 49097 5305 49120
rect 4919 49078 5305 49097
rect 20039 49183 20425 49202
rect 20039 49160 20105 49183
rect 20191 49160 20273 49183
rect 20359 49160 20425 49183
rect 20039 49120 20048 49160
rect 20088 49120 20105 49160
rect 20191 49120 20212 49160
rect 20252 49120 20273 49160
rect 20359 49120 20376 49160
rect 20416 49120 20425 49160
rect 20039 49097 20105 49120
rect 20191 49097 20273 49120
rect 20359 49097 20425 49120
rect 20039 49078 20425 49097
rect 3679 48427 4065 48446
rect 3679 48404 3745 48427
rect 3831 48404 3913 48427
rect 3999 48404 4065 48427
rect 3679 48364 3688 48404
rect 3728 48364 3745 48404
rect 3831 48364 3852 48404
rect 3892 48364 3913 48404
rect 3999 48364 4016 48404
rect 4056 48364 4065 48404
rect 3679 48341 3745 48364
rect 3831 48341 3913 48364
rect 3999 48341 4065 48364
rect 3679 48322 4065 48341
rect 18799 48427 19185 48446
rect 18799 48404 18865 48427
rect 18951 48404 19033 48427
rect 19119 48404 19185 48427
rect 18799 48364 18808 48404
rect 18848 48364 18865 48404
rect 18951 48364 18972 48404
rect 19012 48364 19033 48404
rect 19119 48364 19136 48404
rect 19176 48364 19185 48404
rect 18799 48341 18865 48364
rect 18951 48341 19033 48364
rect 19119 48341 19185 48364
rect 18799 48322 19185 48341
rect 4919 47671 5305 47690
rect 4919 47648 4985 47671
rect 5071 47648 5153 47671
rect 5239 47648 5305 47671
rect 4919 47608 4928 47648
rect 4968 47608 4985 47648
rect 5071 47608 5092 47648
rect 5132 47608 5153 47648
rect 5239 47608 5256 47648
rect 5296 47608 5305 47648
rect 4919 47585 4985 47608
rect 5071 47585 5153 47608
rect 5239 47585 5305 47608
rect 4919 47566 5305 47585
rect 20039 47671 20425 47690
rect 20039 47648 20105 47671
rect 20191 47648 20273 47671
rect 20359 47648 20425 47671
rect 20039 47608 20048 47648
rect 20088 47608 20105 47648
rect 20191 47608 20212 47648
rect 20252 47608 20273 47648
rect 20359 47608 20376 47648
rect 20416 47608 20425 47648
rect 20039 47585 20105 47608
rect 20191 47585 20273 47608
rect 20359 47585 20425 47608
rect 20039 47566 20425 47585
rect 3679 46915 4065 46934
rect 3679 46892 3745 46915
rect 3831 46892 3913 46915
rect 3999 46892 4065 46915
rect 3679 46852 3688 46892
rect 3728 46852 3745 46892
rect 3831 46852 3852 46892
rect 3892 46852 3913 46892
rect 3999 46852 4016 46892
rect 4056 46852 4065 46892
rect 3679 46829 3745 46852
rect 3831 46829 3913 46852
rect 3999 46829 4065 46852
rect 3679 46810 4065 46829
rect 18799 46915 19185 46934
rect 18799 46892 18865 46915
rect 18951 46892 19033 46915
rect 19119 46892 19185 46915
rect 18799 46852 18808 46892
rect 18848 46852 18865 46892
rect 18951 46852 18972 46892
rect 19012 46852 19033 46892
rect 19119 46852 19136 46892
rect 19176 46852 19185 46892
rect 18799 46829 18865 46852
rect 18951 46829 19033 46852
rect 19119 46829 19185 46852
rect 18799 46810 19185 46829
rect 4919 46159 5305 46178
rect 4919 46136 4985 46159
rect 5071 46136 5153 46159
rect 5239 46136 5305 46159
rect 4919 46096 4928 46136
rect 4968 46096 4985 46136
rect 5071 46096 5092 46136
rect 5132 46096 5153 46136
rect 5239 46096 5256 46136
rect 5296 46096 5305 46136
rect 4919 46073 4985 46096
rect 5071 46073 5153 46096
rect 5239 46073 5305 46096
rect 4919 46054 5305 46073
rect 20039 46159 20425 46178
rect 20039 46136 20105 46159
rect 20191 46136 20273 46159
rect 20359 46136 20425 46159
rect 20039 46096 20048 46136
rect 20088 46096 20105 46136
rect 20191 46096 20212 46136
rect 20252 46096 20273 46136
rect 20359 46096 20376 46136
rect 20416 46096 20425 46136
rect 20039 46073 20105 46096
rect 20191 46073 20273 46096
rect 20359 46073 20425 46096
rect 20039 46054 20425 46073
rect 3679 45403 4065 45422
rect 3679 45380 3745 45403
rect 3831 45380 3913 45403
rect 3999 45380 4065 45403
rect 3679 45340 3688 45380
rect 3728 45340 3745 45380
rect 3831 45340 3852 45380
rect 3892 45340 3913 45380
rect 3999 45340 4016 45380
rect 4056 45340 4065 45380
rect 3679 45317 3745 45340
rect 3831 45317 3913 45340
rect 3999 45317 4065 45340
rect 3679 45298 4065 45317
rect 18799 45403 19185 45422
rect 18799 45380 18865 45403
rect 18951 45380 19033 45403
rect 19119 45380 19185 45403
rect 18799 45340 18808 45380
rect 18848 45340 18865 45380
rect 18951 45340 18972 45380
rect 19012 45340 19033 45380
rect 19119 45340 19136 45380
rect 19176 45340 19185 45380
rect 18799 45317 18865 45340
rect 18951 45317 19033 45340
rect 19119 45317 19185 45340
rect 18799 45298 19185 45317
rect 4919 44647 5305 44666
rect 4919 44624 4985 44647
rect 5071 44624 5153 44647
rect 5239 44624 5305 44647
rect 4919 44584 4928 44624
rect 4968 44584 4985 44624
rect 5071 44584 5092 44624
rect 5132 44584 5153 44624
rect 5239 44584 5256 44624
rect 5296 44584 5305 44624
rect 4919 44561 4985 44584
rect 5071 44561 5153 44584
rect 5239 44561 5305 44584
rect 4919 44542 5305 44561
rect 20039 44647 20425 44666
rect 20039 44624 20105 44647
rect 20191 44624 20273 44647
rect 20359 44624 20425 44647
rect 20039 44584 20048 44624
rect 20088 44584 20105 44624
rect 20191 44584 20212 44624
rect 20252 44584 20273 44624
rect 20359 44584 20376 44624
rect 20416 44584 20425 44624
rect 20039 44561 20105 44584
rect 20191 44561 20273 44584
rect 20359 44561 20425 44584
rect 20039 44542 20425 44561
rect 3679 43891 4065 43910
rect 3679 43868 3745 43891
rect 3831 43868 3913 43891
rect 3999 43868 4065 43891
rect 3679 43828 3688 43868
rect 3728 43828 3745 43868
rect 3831 43828 3852 43868
rect 3892 43828 3913 43868
rect 3999 43828 4016 43868
rect 4056 43828 4065 43868
rect 3679 43805 3745 43828
rect 3831 43805 3913 43828
rect 3999 43805 4065 43828
rect 3679 43786 4065 43805
rect 18799 43891 19185 43910
rect 18799 43868 18865 43891
rect 18951 43868 19033 43891
rect 19119 43868 19185 43891
rect 18799 43828 18808 43868
rect 18848 43828 18865 43868
rect 18951 43828 18972 43868
rect 19012 43828 19033 43868
rect 19119 43828 19136 43868
rect 19176 43828 19185 43868
rect 18799 43805 18865 43828
rect 18951 43805 19033 43828
rect 19119 43805 19185 43828
rect 18799 43786 19185 43805
rect 4919 43135 5305 43154
rect 4919 43112 4985 43135
rect 5071 43112 5153 43135
rect 5239 43112 5305 43135
rect 4919 43072 4928 43112
rect 4968 43072 4985 43112
rect 5071 43072 5092 43112
rect 5132 43072 5153 43112
rect 5239 43072 5256 43112
rect 5296 43072 5305 43112
rect 4919 43049 4985 43072
rect 5071 43049 5153 43072
rect 5239 43049 5305 43072
rect 4919 43030 5305 43049
rect 20039 43135 20425 43154
rect 20039 43112 20105 43135
rect 20191 43112 20273 43135
rect 20359 43112 20425 43135
rect 20039 43072 20048 43112
rect 20088 43072 20105 43112
rect 20191 43072 20212 43112
rect 20252 43072 20273 43112
rect 20359 43072 20376 43112
rect 20416 43072 20425 43112
rect 20039 43049 20105 43072
rect 20191 43049 20273 43072
rect 20359 43049 20425 43072
rect 20039 43030 20425 43049
rect 6019 42736 6028 42776
rect 6068 42736 11788 42776
rect 11828 42736 11837 42776
rect 8323 42484 8332 42524
rect 8372 42484 18796 42524
rect 18836 42484 18845 42524
rect 3679 42379 4065 42398
rect 3679 42356 3745 42379
rect 3831 42356 3913 42379
rect 3999 42356 4065 42379
rect 3679 42316 3688 42356
rect 3728 42316 3745 42356
rect 3831 42316 3852 42356
rect 3892 42316 3913 42356
rect 3999 42316 4016 42356
rect 4056 42316 4065 42356
rect 3679 42293 3745 42316
rect 3831 42293 3913 42316
rect 3999 42293 4065 42316
rect 3679 42274 4065 42293
rect 18799 42379 19185 42398
rect 18799 42356 18865 42379
rect 18951 42356 19033 42379
rect 19119 42356 19185 42379
rect 18799 42316 18808 42356
rect 18848 42316 18865 42356
rect 18951 42316 18972 42356
rect 19012 42316 19033 42356
rect 19119 42316 19136 42356
rect 19176 42316 19185 42356
rect 18799 42293 18865 42316
rect 18951 42293 19033 42316
rect 19119 42293 19185 42316
rect 18799 42274 19185 42293
rect 9667 41728 9676 41768
rect 9716 41728 19660 41768
rect 19700 41728 19709 41768
rect 4919 41623 5305 41642
rect 4919 41600 4985 41623
rect 5071 41600 5153 41623
rect 5239 41600 5305 41623
rect 4919 41560 4928 41600
rect 4968 41560 4985 41600
rect 5071 41560 5092 41600
rect 5132 41560 5153 41600
rect 5239 41560 5256 41600
rect 5296 41560 5305 41600
rect 4919 41537 4985 41560
rect 5071 41537 5153 41560
rect 5239 41537 5305 41560
rect 4919 41518 5305 41537
rect 20039 41623 20425 41642
rect 20039 41600 20105 41623
rect 20191 41600 20273 41623
rect 20359 41600 20425 41623
rect 20039 41560 20048 41600
rect 20088 41560 20105 41600
rect 20191 41560 20212 41600
rect 20252 41560 20273 41600
rect 20359 41560 20376 41600
rect 20416 41560 20425 41600
rect 20039 41537 20105 41560
rect 20191 41537 20273 41560
rect 20359 41537 20425 41560
rect 20039 41518 20425 41537
rect 11299 41392 11308 41432
rect 11348 41392 11596 41432
rect 11636 41392 11645 41432
rect 2467 41224 2476 41264
rect 2516 41224 5932 41264
rect 5972 41224 5981 41264
rect 8419 40972 8428 41012
rect 8468 40972 19468 41012
rect 19508 40972 19517 41012
rect 3679 40867 4065 40886
rect 3679 40844 3745 40867
rect 3831 40844 3913 40867
rect 3999 40844 4065 40867
rect 3679 40804 3688 40844
rect 3728 40804 3745 40844
rect 3831 40804 3852 40844
rect 3892 40804 3913 40844
rect 3999 40804 4016 40844
rect 4056 40804 4065 40844
rect 3679 40781 3745 40804
rect 3831 40781 3913 40804
rect 3999 40781 4065 40804
rect 3679 40762 4065 40781
rect 18799 40867 19185 40886
rect 18799 40844 18865 40867
rect 18951 40844 19033 40867
rect 19119 40844 19185 40867
rect 18799 40804 18808 40844
rect 18848 40804 18865 40844
rect 18951 40804 18972 40844
rect 19012 40804 19033 40844
rect 19119 40804 19136 40844
rect 19176 40804 19185 40844
rect 18799 40781 18865 40804
rect 18951 40781 19033 40804
rect 19119 40781 19185 40804
rect 18799 40762 19185 40781
rect 16291 40636 16300 40676
rect 16340 40636 19468 40676
rect 19508 40636 19517 40676
rect 4919 40111 5305 40130
rect 4919 40088 4985 40111
rect 5071 40088 5153 40111
rect 5239 40088 5305 40111
rect 4919 40048 4928 40088
rect 4968 40048 4985 40088
rect 5071 40048 5092 40088
rect 5132 40048 5153 40088
rect 5239 40048 5256 40088
rect 5296 40048 5305 40088
rect 4919 40025 4985 40048
rect 5071 40025 5153 40048
rect 5239 40025 5305 40048
rect 4919 40006 5305 40025
rect 20039 40111 20425 40130
rect 20039 40088 20105 40111
rect 20191 40088 20273 40111
rect 20359 40088 20425 40111
rect 20039 40048 20048 40088
rect 20088 40048 20105 40088
rect 20191 40048 20212 40088
rect 20252 40048 20273 40088
rect 20359 40048 20376 40088
rect 20416 40048 20425 40088
rect 20039 40025 20105 40048
rect 20191 40025 20273 40048
rect 20359 40025 20425 40048
rect 20039 40006 20425 40025
rect 3679 39355 4065 39374
rect 3679 39332 3745 39355
rect 3831 39332 3913 39355
rect 3999 39332 4065 39355
rect 3679 39292 3688 39332
rect 3728 39292 3745 39332
rect 3831 39292 3852 39332
rect 3892 39292 3913 39332
rect 3999 39292 4016 39332
rect 4056 39292 4065 39332
rect 3679 39269 3745 39292
rect 3831 39269 3913 39292
rect 3999 39269 4065 39292
rect 3679 39250 4065 39269
rect 18799 39355 19185 39374
rect 18799 39332 18865 39355
rect 18951 39332 19033 39355
rect 19119 39332 19185 39355
rect 18799 39292 18808 39332
rect 18848 39292 18865 39332
rect 18951 39292 18972 39332
rect 19012 39292 19033 39332
rect 19119 39292 19136 39332
rect 19176 39292 19185 39332
rect 18799 39269 18865 39292
rect 18951 39269 19033 39292
rect 19119 39269 19185 39292
rect 18799 39250 19185 39269
rect 4919 38599 5305 38618
rect 4919 38576 4985 38599
rect 5071 38576 5153 38599
rect 5239 38576 5305 38599
rect 4919 38536 4928 38576
rect 4968 38536 4985 38576
rect 5071 38536 5092 38576
rect 5132 38536 5153 38576
rect 5239 38536 5256 38576
rect 5296 38536 5305 38576
rect 4919 38513 4985 38536
rect 5071 38513 5153 38536
rect 5239 38513 5305 38536
rect 4919 38494 5305 38513
rect 20039 38599 20425 38618
rect 20039 38576 20105 38599
rect 20191 38576 20273 38599
rect 20359 38576 20425 38599
rect 20039 38536 20048 38576
rect 20088 38536 20105 38576
rect 20191 38536 20212 38576
rect 20252 38536 20273 38576
rect 20359 38536 20376 38576
rect 20416 38536 20425 38576
rect 20039 38513 20105 38536
rect 20191 38513 20273 38536
rect 20359 38513 20425 38536
rect 20039 38494 20425 38513
rect 3679 37843 4065 37862
rect 3679 37820 3745 37843
rect 3831 37820 3913 37843
rect 3999 37820 4065 37843
rect 3679 37780 3688 37820
rect 3728 37780 3745 37820
rect 3831 37780 3852 37820
rect 3892 37780 3913 37820
rect 3999 37780 4016 37820
rect 4056 37780 4065 37820
rect 3679 37757 3745 37780
rect 3831 37757 3913 37780
rect 3999 37757 4065 37780
rect 3679 37738 4065 37757
rect 18799 37843 19185 37862
rect 18799 37820 18865 37843
rect 18951 37820 19033 37843
rect 19119 37820 19185 37843
rect 18799 37780 18808 37820
rect 18848 37780 18865 37820
rect 18951 37780 18972 37820
rect 19012 37780 19033 37820
rect 19119 37780 19136 37820
rect 19176 37780 19185 37820
rect 18799 37757 18865 37780
rect 18951 37757 19033 37780
rect 19119 37757 19185 37780
rect 18799 37738 19185 37757
rect 12355 37444 12364 37484
rect 12404 37444 19564 37484
rect 19604 37444 19613 37484
rect 4919 37087 5305 37106
rect 4919 37064 4985 37087
rect 5071 37064 5153 37087
rect 5239 37064 5305 37087
rect 4919 37024 4928 37064
rect 4968 37024 4985 37064
rect 5071 37024 5092 37064
rect 5132 37024 5153 37064
rect 5239 37024 5256 37064
rect 5296 37024 5305 37064
rect 4919 37001 4985 37024
rect 5071 37001 5153 37024
rect 5239 37001 5305 37024
rect 4919 36982 5305 37001
rect 20039 37087 20425 37106
rect 20039 37064 20105 37087
rect 20191 37064 20273 37087
rect 20359 37064 20425 37087
rect 20039 37024 20048 37064
rect 20088 37024 20105 37064
rect 20191 37024 20212 37064
rect 20252 37024 20273 37064
rect 20359 37024 20376 37064
rect 20416 37024 20425 37064
rect 20039 37001 20105 37024
rect 20191 37001 20273 37024
rect 20359 37001 20425 37024
rect 20039 36982 20425 37001
rect 5347 36688 5356 36728
rect 5396 36688 11788 36728
rect 11828 36688 12940 36728
rect 12980 36688 12989 36728
rect 3679 36331 4065 36350
rect 3679 36308 3745 36331
rect 3831 36308 3913 36331
rect 3999 36308 4065 36331
rect 3679 36268 3688 36308
rect 3728 36268 3745 36308
rect 3831 36268 3852 36308
rect 3892 36268 3913 36308
rect 3999 36268 4016 36308
rect 4056 36268 4065 36308
rect 3679 36245 3745 36268
rect 3831 36245 3913 36268
rect 3999 36245 4065 36268
rect 3679 36226 4065 36245
rect 18799 36331 19185 36350
rect 18799 36308 18865 36331
rect 18951 36308 19033 36331
rect 19119 36308 19185 36331
rect 18799 36268 18808 36308
rect 18848 36268 18865 36308
rect 18951 36268 18972 36308
rect 19012 36268 19033 36308
rect 19119 36268 19136 36308
rect 19176 36268 19185 36308
rect 18799 36245 18865 36268
rect 18951 36245 19033 36268
rect 19119 36245 19185 36268
rect 18799 36226 19185 36245
rect 4919 35575 5305 35594
rect 4919 35552 4985 35575
rect 5071 35552 5153 35575
rect 5239 35552 5305 35575
rect 4919 35512 4928 35552
rect 4968 35512 4985 35552
rect 5071 35512 5092 35552
rect 5132 35512 5153 35552
rect 5239 35512 5256 35552
rect 5296 35512 5305 35552
rect 4919 35489 4985 35512
rect 5071 35489 5153 35512
rect 5239 35489 5305 35512
rect 4919 35470 5305 35489
rect 20039 35575 20425 35594
rect 20039 35552 20105 35575
rect 20191 35552 20273 35575
rect 20359 35552 20425 35575
rect 20039 35512 20048 35552
rect 20088 35512 20105 35552
rect 20191 35512 20212 35552
rect 20252 35512 20273 35552
rect 20359 35512 20376 35552
rect 20416 35512 20425 35552
rect 20039 35489 20105 35512
rect 20191 35489 20273 35512
rect 20359 35489 20425 35512
rect 20039 35470 20425 35489
rect 931 35008 940 35048
rect 980 35008 3820 35048
rect 3860 35008 3869 35048
rect 3679 34819 4065 34838
rect 3679 34796 3745 34819
rect 3831 34796 3913 34819
rect 3999 34796 4065 34819
rect 3679 34756 3688 34796
rect 3728 34756 3745 34796
rect 3831 34756 3852 34796
rect 3892 34756 3913 34796
rect 3999 34756 4016 34796
rect 4056 34756 4065 34796
rect 3679 34733 3745 34756
rect 3831 34733 3913 34756
rect 3999 34733 4065 34756
rect 3679 34714 4065 34733
rect 18799 34819 19185 34838
rect 18799 34796 18865 34819
rect 18951 34796 19033 34819
rect 19119 34796 19185 34819
rect 18799 34756 18808 34796
rect 18848 34756 18865 34796
rect 18951 34756 18972 34796
rect 19012 34756 19033 34796
rect 19119 34756 19136 34796
rect 19176 34756 19185 34796
rect 18799 34733 18865 34756
rect 18951 34733 19033 34756
rect 19119 34733 19185 34756
rect 18799 34714 19185 34733
rect 3907 34252 3916 34292
rect 3956 34252 9004 34292
rect 9044 34252 9053 34292
rect 11971 34168 11980 34208
rect 12020 34168 12652 34208
rect 12692 34168 12701 34208
rect 4919 34063 5305 34082
rect 4919 34040 4985 34063
rect 5071 34040 5153 34063
rect 5239 34040 5305 34063
rect 4919 34000 4928 34040
rect 4968 34000 4985 34040
rect 5071 34000 5092 34040
rect 5132 34000 5153 34040
rect 5239 34000 5256 34040
rect 5296 34000 5305 34040
rect 4919 33977 4985 34000
rect 5071 33977 5153 34000
rect 5239 33977 5305 34000
rect 4919 33958 5305 33977
rect 20039 34063 20425 34082
rect 20039 34040 20105 34063
rect 20191 34040 20273 34063
rect 20359 34040 20425 34063
rect 20039 34000 20048 34040
rect 20088 34000 20105 34040
rect 20191 34000 20212 34040
rect 20252 34000 20273 34040
rect 20359 34000 20376 34040
rect 20416 34000 20425 34040
rect 20039 33977 20105 34000
rect 20191 33977 20273 34000
rect 20359 33977 20425 34000
rect 20039 33958 20425 33977
rect 3679 33307 4065 33326
rect 3679 33284 3745 33307
rect 3831 33284 3913 33307
rect 3999 33284 4065 33307
rect 3679 33244 3688 33284
rect 3728 33244 3745 33284
rect 3831 33244 3852 33284
rect 3892 33244 3913 33284
rect 3999 33244 4016 33284
rect 4056 33244 4065 33284
rect 3679 33221 3745 33244
rect 3831 33221 3913 33244
rect 3999 33221 4065 33244
rect 3679 33202 4065 33221
rect 18799 33307 19185 33326
rect 18799 33284 18865 33307
rect 18951 33284 19033 33307
rect 19119 33284 19185 33307
rect 18799 33244 18808 33284
rect 18848 33244 18865 33284
rect 18951 33244 18972 33284
rect 19012 33244 19033 33284
rect 19119 33244 19136 33284
rect 19176 33244 19185 33284
rect 18799 33221 18865 33244
rect 18951 33221 19033 33244
rect 19119 33221 19185 33244
rect 18799 33202 19185 33221
rect 4919 32551 5305 32570
rect 4919 32528 4985 32551
rect 5071 32528 5153 32551
rect 5239 32528 5305 32551
rect 4919 32488 4928 32528
rect 4968 32488 4985 32528
rect 5071 32488 5092 32528
rect 5132 32488 5153 32528
rect 5239 32488 5256 32528
rect 5296 32488 5305 32528
rect 4919 32465 4985 32488
rect 5071 32465 5153 32488
rect 5239 32465 5305 32488
rect 4919 32446 5305 32465
rect 20039 32551 20425 32570
rect 20039 32528 20105 32551
rect 20191 32528 20273 32551
rect 20359 32528 20425 32551
rect 20039 32488 20048 32528
rect 20088 32488 20105 32528
rect 20191 32488 20212 32528
rect 20252 32488 20273 32528
rect 20359 32488 20376 32528
rect 20416 32488 20425 32528
rect 20039 32465 20105 32488
rect 20191 32465 20273 32488
rect 20359 32465 20425 32488
rect 20039 32446 20425 32465
rect 3679 31795 4065 31814
rect 3679 31772 3745 31795
rect 3831 31772 3913 31795
rect 3999 31772 4065 31795
rect 3679 31732 3688 31772
rect 3728 31732 3745 31772
rect 3831 31732 3852 31772
rect 3892 31732 3913 31772
rect 3999 31732 4016 31772
rect 4056 31732 4065 31772
rect 3679 31709 3745 31732
rect 3831 31709 3913 31732
rect 3999 31709 4065 31732
rect 3679 31690 4065 31709
rect 18799 31795 19185 31814
rect 18799 31772 18865 31795
rect 18951 31772 19033 31795
rect 19119 31772 19185 31795
rect 18799 31732 18808 31772
rect 18848 31732 18865 31772
rect 18951 31732 18972 31772
rect 19012 31732 19033 31772
rect 19119 31732 19136 31772
rect 19176 31732 19185 31772
rect 18799 31709 18865 31732
rect 18951 31709 19033 31732
rect 19119 31709 19185 31732
rect 18799 31690 19185 31709
rect 4919 31039 5305 31058
rect 4919 31016 4985 31039
rect 5071 31016 5153 31039
rect 5239 31016 5305 31039
rect 4919 30976 4928 31016
rect 4968 30976 4985 31016
rect 5071 30976 5092 31016
rect 5132 30976 5153 31016
rect 5239 30976 5256 31016
rect 5296 30976 5305 31016
rect 4919 30953 4985 30976
rect 5071 30953 5153 30976
rect 5239 30953 5305 30976
rect 4919 30934 5305 30953
rect 20039 31039 20425 31058
rect 20039 31016 20105 31039
rect 20191 31016 20273 31039
rect 20359 31016 20425 31039
rect 20039 30976 20048 31016
rect 20088 30976 20105 31016
rect 20191 30976 20212 31016
rect 20252 30976 20273 31016
rect 20359 30976 20376 31016
rect 20416 30976 20425 31016
rect 20039 30953 20105 30976
rect 20191 30953 20273 30976
rect 20359 30953 20425 30976
rect 20039 30934 20425 30953
rect 12122 30703 12246 30722
rect 12122 30617 12141 30703
rect 12227 30680 12246 30703
rect 12227 30640 12364 30680
rect 12404 30640 12413 30680
rect 12227 30617 12246 30640
rect 12122 30598 12246 30617
rect 3679 30283 4065 30302
rect 3679 30260 3745 30283
rect 3831 30260 3913 30283
rect 3999 30260 4065 30283
rect 3679 30220 3688 30260
rect 3728 30220 3745 30260
rect 3831 30220 3852 30260
rect 3892 30220 3913 30260
rect 3999 30220 4016 30260
rect 4056 30220 4065 30260
rect 3679 30197 3745 30220
rect 3831 30197 3913 30220
rect 3999 30197 4065 30220
rect 3679 30178 4065 30197
rect 18799 30283 19185 30302
rect 18799 30260 18865 30283
rect 18951 30260 19033 30283
rect 19119 30260 19185 30283
rect 18799 30220 18808 30260
rect 18848 30220 18865 30260
rect 18951 30220 18972 30260
rect 19012 30220 19033 30260
rect 19119 30220 19136 30260
rect 19176 30220 19185 30260
rect 18799 30197 18865 30220
rect 18951 30197 19033 30220
rect 19119 30197 19185 30220
rect 18799 30178 19185 30197
rect 16675 29632 16684 29672
rect 16724 29632 20812 29672
rect 20852 29632 20861 29672
rect 4919 29527 5305 29546
rect 4919 29504 4985 29527
rect 5071 29504 5153 29527
rect 5239 29504 5305 29527
rect 4919 29464 4928 29504
rect 4968 29464 4985 29504
rect 5071 29464 5092 29504
rect 5132 29464 5153 29504
rect 5239 29464 5256 29504
rect 5296 29464 5305 29504
rect 4919 29441 4985 29464
rect 5071 29441 5153 29464
rect 5239 29441 5305 29464
rect 4919 29422 5305 29441
rect 20039 29527 20425 29546
rect 20039 29504 20105 29527
rect 20191 29504 20273 29527
rect 20359 29504 20425 29527
rect 20039 29464 20048 29504
rect 20088 29464 20105 29504
rect 20191 29464 20212 29504
rect 20252 29464 20273 29504
rect 20359 29464 20376 29504
rect 20416 29464 20425 29504
rect 20039 29441 20105 29464
rect 20191 29441 20273 29464
rect 20359 29441 20425 29464
rect 20039 29422 20425 29441
rect 3679 28771 4065 28790
rect 3679 28748 3745 28771
rect 3831 28748 3913 28771
rect 3999 28748 4065 28771
rect 3679 28708 3688 28748
rect 3728 28708 3745 28748
rect 3831 28708 3852 28748
rect 3892 28708 3913 28748
rect 3999 28708 4016 28748
rect 4056 28708 4065 28748
rect 3679 28685 3745 28708
rect 3831 28685 3913 28708
rect 3999 28685 4065 28708
rect 3679 28666 4065 28685
rect 18799 28771 19185 28790
rect 18799 28748 18865 28771
rect 18951 28748 19033 28771
rect 19119 28748 19185 28771
rect 18799 28708 18808 28748
rect 18848 28708 18865 28748
rect 18951 28708 18972 28748
rect 19012 28708 19033 28748
rect 19119 28708 19136 28748
rect 19176 28708 19185 28748
rect 18799 28685 18865 28708
rect 18951 28685 19033 28708
rect 19119 28685 19185 28708
rect 18799 28666 19185 28685
rect 3139 28372 3148 28412
rect 3188 28372 3436 28412
rect 3476 28372 3485 28412
rect 4919 28015 5305 28034
rect 4919 27992 4985 28015
rect 5071 27992 5153 28015
rect 5239 27992 5305 28015
rect 4919 27952 4928 27992
rect 4968 27952 4985 27992
rect 5071 27952 5092 27992
rect 5132 27952 5153 27992
rect 5239 27952 5256 27992
rect 5296 27952 5305 27992
rect 4919 27929 4985 27952
rect 5071 27929 5153 27952
rect 5239 27929 5305 27952
rect 4919 27910 5305 27929
rect 20039 28015 20425 28034
rect 20039 27992 20105 28015
rect 20191 27992 20273 28015
rect 20359 27992 20425 28015
rect 20039 27952 20048 27992
rect 20088 27952 20105 27992
rect 20191 27952 20212 27992
rect 20252 27952 20273 27992
rect 20359 27952 20376 27992
rect 20416 27952 20425 27992
rect 20039 27929 20105 27952
rect 20191 27929 20273 27952
rect 20359 27929 20425 27952
rect 20039 27910 20425 27929
rect 3679 27259 4065 27278
rect 3679 27236 3745 27259
rect 3831 27236 3913 27259
rect 3999 27236 4065 27259
rect 3679 27196 3688 27236
rect 3728 27196 3745 27236
rect 3831 27196 3852 27236
rect 3892 27196 3913 27236
rect 3999 27196 4016 27236
rect 4056 27196 4065 27236
rect 3679 27173 3745 27196
rect 3831 27173 3913 27196
rect 3999 27173 4065 27196
rect 3679 27154 4065 27173
rect 18799 27259 19185 27278
rect 18799 27236 18865 27259
rect 18951 27236 19033 27259
rect 19119 27236 19185 27259
rect 18799 27196 18808 27236
rect 18848 27196 18865 27236
rect 18951 27196 18972 27236
rect 19012 27196 19033 27236
rect 19119 27196 19136 27236
rect 19176 27196 19185 27236
rect 18799 27173 18865 27196
rect 18951 27173 19033 27196
rect 19119 27173 19185 27196
rect 18799 27154 19185 27173
rect 4919 26503 5305 26522
rect 4919 26480 4985 26503
rect 5071 26480 5153 26503
rect 5239 26480 5305 26503
rect 4919 26440 4928 26480
rect 4968 26440 4985 26480
rect 5071 26440 5092 26480
rect 5132 26440 5153 26480
rect 5239 26440 5256 26480
rect 5296 26440 5305 26480
rect 4919 26417 4985 26440
rect 5071 26417 5153 26440
rect 5239 26417 5305 26440
rect 4919 26398 5305 26417
rect 9842 26503 9966 26522
rect 9842 26417 9861 26503
rect 9947 26480 9966 26503
rect 20039 26503 20425 26522
rect 20039 26480 20105 26503
rect 20191 26480 20273 26503
rect 20359 26480 20425 26503
rect 9947 26440 12076 26480
rect 12116 26440 12125 26480
rect 20039 26440 20048 26480
rect 20088 26440 20105 26480
rect 20191 26440 20212 26480
rect 20252 26440 20273 26480
rect 20359 26440 20376 26480
rect 20416 26440 20425 26480
rect 9947 26417 9966 26440
rect 9842 26398 9966 26417
rect 20039 26417 20105 26440
rect 20191 26417 20273 26440
rect 20359 26417 20425 26440
rect 20039 26398 20425 26417
rect 8018 26335 8142 26354
rect 8018 26249 8037 26335
rect 8123 26312 8142 26335
rect 8123 26272 12364 26312
rect 12404 26272 12413 26312
rect 8123 26249 8142 26272
rect 8018 26230 8142 26249
rect 4675 26020 4684 26060
rect 4724 26020 14572 26060
rect 14612 26020 14621 26060
rect 3679 25747 4065 25766
rect 3679 25724 3745 25747
rect 3831 25724 3913 25747
rect 3999 25724 4065 25747
rect 3679 25684 3688 25724
rect 3728 25684 3745 25724
rect 3831 25684 3852 25724
rect 3892 25684 3913 25724
rect 3999 25684 4016 25724
rect 4056 25684 4065 25724
rect 3679 25661 3745 25684
rect 3831 25661 3913 25684
rect 3999 25661 4065 25684
rect 3679 25642 4065 25661
rect 18799 25747 19185 25766
rect 18799 25724 18865 25747
rect 18951 25724 19033 25747
rect 19119 25724 19185 25747
rect 18799 25684 18808 25724
rect 18848 25684 18865 25724
rect 18951 25684 18972 25724
rect 19012 25684 19033 25724
rect 19119 25684 19136 25724
rect 19176 25684 19185 25724
rect 18799 25661 18865 25684
rect 18951 25661 19033 25684
rect 19119 25661 19185 25684
rect 18799 25642 19185 25661
rect 5059 25180 5068 25220
rect 5108 25180 17644 25220
rect 17684 25180 17693 25220
rect 835 25096 844 25136
rect 884 25096 5260 25136
rect 5300 25096 5309 25136
rect 10819 25096 10828 25136
rect 10868 25096 11308 25136
rect 11348 25096 11357 25136
rect 4919 24991 5305 25010
rect 4919 24968 4985 24991
rect 5071 24968 5153 24991
rect 5239 24968 5305 24991
rect 4919 24928 4928 24968
rect 4968 24928 4985 24968
rect 5071 24928 5092 24968
rect 5132 24928 5153 24968
rect 5239 24928 5256 24968
rect 5296 24928 5305 24968
rect 4919 24905 4985 24928
rect 5071 24905 5153 24928
rect 5239 24905 5305 24928
rect 4919 24886 5305 24905
rect 20039 24991 20425 25010
rect 20039 24968 20105 24991
rect 20191 24968 20273 24991
rect 20359 24968 20425 24991
rect 20039 24928 20048 24968
rect 20088 24928 20105 24968
rect 20191 24928 20212 24968
rect 20252 24928 20273 24968
rect 20359 24928 20376 24968
rect 20416 24928 20425 24968
rect 20039 24905 20105 24928
rect 20191 24905 20273 24928
rect 20359 24905 20425 24928
rect 20039 24886 20425 24905
rect 3679 24235 4065 24254
rect 3679 24212 3745 24235
rect 3831 24212 3913 24235
rect 3999 24212 4065 24235
rect 3679 24172 3688 24212
rect 3728 24172 3745 24212
rect 3831 24172 3852 24212
rect 3892 24172 3913 24212
rect 3999 24172 4016 24212
rect 4056 24172 4065 24212
rect 3679 24149 3745 24172
rect 3831 24149 3913 24172
rect 3999 24149 4065 24172
rect 3679 24130 4065 24149
rect 18799 24235 19185 24254
rect 18799 24212 18865 24235
rect 18951 24212 19033 24235
rect 19119 24212 19185 24235
rect 18799 24172 18808 24212
rect 18848 24172 18865 24212
rect 18951 24172 18972 24212
rect 19012 24172 19033 24212
rect 19119 24172 19136 24212
rect 19176 24172 19185 24212
rect 18799 24149 18865 24172
rect 18951 24149 19033 24172
rect 19119 24149 19185 24172
rect 18799 24130 19185 24149
rect 2851 23752 2860 23792
rect 2900 23752 14092 23792
rect 14132 23752 14141 23792
rect 4919 23479 5305 23498
rect 4919 23456 4985 23479
rect 5071 23456 5153 23479
rect 5239 23456 5305 23479
rect 4919 23416 4928 23456
rect 4968 23416 4985 23456
rect 5071 23416 5092 23456
rect 5132 23416 5153 23456
rect 5239 23416 5256 23456
rect 5296 23416 5305 23456
rect 4919 23393 4985 23416
rect 5071 23393 5153 23416
rect 5239 23393 5305 23416
rect 4919 23374 5305 23393
rect 20039 23479 20425 23498
rect 20039 23456 20105 23479
rect 20191 23456 20273 23479
rect 20359 23456 20425 23479
rect 20039 23416 20048 23456
rect 20088 23416 20105 23456
rect 20191 23416 20212 23456
rect 20252 23416 20273 23456
rect 20359 23416 20376 23456
rect 20416 23416 20425 23456
rect 20039 23393 20105 23416
rect 20191 23393 20273 23416
rect 20359 23393 20425 23416
rect 20039 23374 20425 23393
rect 2947 22828 2956 22868
rect 2996 22828 20140 22868
rect 20180 22828 20189 22868
rect 3679 22723 4065 22742
rect 3679 22700 3745 22723
rect 3831 22700 3913 22723
rect 3999 22700 4065 22723
rect 3679 22660 3688 22700
rect 3728 22660 3745 22700
rect 3831 22660 3852 22700
rect 3892 22660 3913 22700
rect 3999 22660 4016 22700
rect 4056 22660 4065 22700
rect 3679 22637 3745 22660
rect 3831 22637 3913 22660
rect 3999 22637 4065 22660
rect 3679 22618 4065 22637
rect 18799 22723 19185 22742
rect 18799 22700 18865 22723
rect 18951 22700 19033 22723
rect 19119 22700 19185 22723
rect 18799 22660 18808 22700
rect 18848 22660 18865 22700
rect 18951 22660 18972 22700
rect 19012 22660 19033 22700
rect 19119 22660 19136 22700
rect 19176 22660 19185 22700
rect 18799 22637 18865 22660
rect 18951 22637 19033 22660
rect 19119 22637 19185 22660
rect 18799 22618 19185 22637
rect 4919 21967 5305 21986
rect 4919 21944 4985 21967
rect 5071 21944 5153 21967
rect 5239 21944 5305 21967
rect 4919 21904 4928 21944
rect 4968 21904 4985 21944
rect 5071 21904 5092 21944
rect 5132 21904 5153 21944
rect 5239 21904 5256 21944
rect 5296 21904 5305 21944
rect 4919 21881 4985 21904
rect 5071 21881 5153 21904
rect 5239 21881 5305 21904
rect 4919 21862 5305 21881
rect 20039 21967 20425 21986
rect 20039 21944 20105 21967
rect 20191 21944 20273 21967
rect 20359 21944 20425 21967
rect 20039 21904 20048 21944
rect 20088 21904 20105 21944
rect 20191 21904 20212 21944
rect 20252 21904 20273 21944
rect 20359 21904 20376 21944
rect 20416 21904 20425 21944
rect 20039 21881 20105 21904
rect 20191 21881 20273 21904
rect 20359 21881 20425 21904
rect 20039 21862 20425 21881
rect 3679 21211 4065 21230
rect 3679 21188 3745 21211
rect 3831 21188 3913 21211
rect 3999 21188 4065 21211
rect 3679 21148 3688 21188
rect 3728 21148 3745 21188
rect 3831 21148 3852 21188
rect 3892 21148 3913 21188
rect 3999 21148 4016 21188
rect 4056 21148 4065 21188
rect 3679 21125 3745 21148
rect 3831 21125 3913 21148
rect 3999 21125 4065 21148
rect 3679 21106 4065 21125
rect 18799 21211 19185 21230
rect 18799 21188 18865 21211
rect 18951 21188 19033 21211
rect 19119 21188 19185 21211
rect 18799 21148 18808 21188
rect 18848 21148 18865 21188
rect 18951 21148 18972 21188
rect 19012 21148 19033 21188
rect 19119 21148 19136 21188
rect 19176 21148 19185 21188
rect 18799 21125 18865 21148
rect 18951 21125 19033 21148
rect 19119 21125 19185 21148
rect 18799 21106 19185 21125
rect 4919 20455 5305 20474
rect 4919 20432 4985 20455
rect 5071 20432 5153 20455
rect 5239 20432 5305 20455
rect 4919 20392 4928 20432
rect 4968 20392 4985 20432
rect 5071 20392 5092 20432
rect 5132 20392 5153 20432
rect 5239 20392 5256 20432
rect 5296 20392 5305 20432
rect 4919 20369 4985 20392
rect 5071 20369 5153 20392
rect 5239 20369 5305 20392
rect 4919 20350 5305 20369
rect 20039 20455 20425 20474
rect 20039 20432 20105 20455
rect 20191 20432 20273 20455
rect 20359 20432 20425 20455
rect 20039 20392 20048 20432
rect 20088 20392 20105 20432
rect 20191 20392 20212 20432
rect 20252 20392 20273 20432
rect 20359 20392 20376 20432
rect 20416 20392 20425 20432
rect 20039 20369 20105 20392
rect 20191 20369 20273 20392
rect 20359 20369 20425 20392
rect 20039 20350 20425 20369
rect 3679 19699 4065 19718
rect 3679 19676 3745 19699
rect 3831 19676 3913 19699
rect 3999 19676 4065 19699
rect 3679 19636 3688 19676
rect 3728 19636 3745 19676
rect 3831 19636 3852 19676
rect 3892 19636 3913 19676
rect 3999 19636 4016 19676
rect 4056 19636 4065 19676
rect 3679 19613 3745 19636
rect 3831 19613 3913 19636
rect 3999 19613 4065 19636
rect 3679 19594 4065 19613
rect 18799 19699 19185 19718
rect 18799 19676 18865 19699
rect 18951 19676 19033 19699
rect 19119 19676 19185 19699
rect 18799 19636 18808 19676
rect 18848 19636 18865 19676
rect 18951 19636 18972 19676
rect 19012 19636 19033 19676
rect 19119 19636 19136 19676
rect 19176 19636 19185 19676
rect 18799 19613 18865 19636
rect 18951 19613 19033 19636
rect 19119 19613 19185 19636
rect 18799 19594 19185 19613
rect 4919 18943 5305 18962
rect 4919 18920 4985 18943
rect 5071 18920 5153 18943
rect 5239 18920 5305 18943
rect 4919 18880 4928 18920
rect 4968 18880 4985 18920
rect 5071 18880 5092 18920
rect 5132 18880 5153 18920
rect 5239 18880 5256 18920
rect 5296 18880 5305 18920
rect 4919 18857 4985 18880
rect 5071 18857 5153 18880
rect 5239 18857 5305 18880
rect 4919 18838 5305 18857
rect 20039 18943 20425 18962
rect 20039 18920 20105 18943
rect 20191 18920 20273 18943
rect 20359 18920 20425 18943
rect 20039 18880 20048 18920
rect 20088 18880 20105 18920
rect 20191 18880 20212 18920
rect 20252 18880 20273 18920
rect 20359 18880 20376 18920
rect 20416 18880 20425 18920
rect 20039 18857 20105 18880
rect 20191 18857 20273 18880
rect 20359 18857 20425 18880
rect 20039 18838 20425 18857
rect 3679 18187 4065 18206
rect 3679 18164 3745 18187
rect 3831 18164 3913 18187
rect 3999 18164 4065 18187
rect 3679 18124 3688 18164
rect 3728 18124 3745 18164
rect 3831 18124 3852 18164
rect 3892 18124 3913 18164
rect 3999 18124 4016 18164
rect 4056 18124 4065 18164
rect 3679 18101 3745 18124
rect 3831 18101 3913 18124
rect 3999 18101 4065 18124
rect 3679 18082 4065 18101
rect 18799 18187 19185 18206
rect 18799 18164 18865 18187
rect 18951 18164 19033 18187
rect 19119 18164 19185 18187
rect 18799 18124 18808 18164
rect 18848 18124 18865 18164
rect 18951 18124 18972 18164
rect 19012 18124 19033 18164
rect 19119 18124 19136 18164
rect 19176 18124 19185 18164
rect 18799 18101 18865 18124
rect 18951 18101 19033 18124
rect 19119 18101 19185 18124
rect 18799 18082 19185 18101
rect 15314 17683 15438 17702
rect 15314 17660 15333 17683
rect 14083 17620 14092 17660
rect 14132 17620 15333 17660
rect 15314 17597 15333 17620
rect 15419 17597 15438 17683
rect 15314 17578 15438 17597
rect 4387 17536 4396 17576
rect 4436 17536 5740 17576
rect 5780 17536 5789 17576
rect 4919 17431 5305 17450
rect 4919 17408 4985 17431
rect 5071 17408 5153 17431
rect 5239 17408 5305 17431
rect 4919 17368 4928 17408
rect 4968 17368 4985 17408
rect 5071 17368 5092 17408
rect 5132 17368 5153 17408
rect 5239 17368 5256 17408
rect 5296 17368 5305 17408
rect 4919 17345 4985 17368
rect 5071 17345 5153 17368
rect 5239 17345 5305 17368
rect 4919 17326 5305 17345
rect 20039 17431 20425 17450
rect 20039 17408 20105 17431
rect 20191 17408 20273 17431
rect 20359 17408 20425 17431
rect 20039 17368 20048 17408
rect 20088 17368 20105 17408
rect 20191 17368 20212 17408
rect 20252 17368 20273 17408
rect 20359 17368 20376 17408
rect 20416 17368 20425 17408
rect 20039 17345 20105 17368
rect 20191 17345 20273 17368
rect 20359 17345 20425 17368
rect 20039 17326 20425 17345
rect 2947 16780 2956 16820
rect 2996 16780 5644 16820
rect 5684 16780 6604 16820
rect 6644 16780 6653 16820
rect 3679 16675 4065 16694
rect 3679 16652 3745 16675
rect 3831 16652 3913 16675
rect 3999 16652 4065 16675
rect 3679 16612 3688 16652
rect 3728 16612 3745 16652
rect 3831 16612 3852 16652
rect 3892 16612 3913 16652
rect 3999 16612 4016 16652
rect 4056 16612 4065 16652
rect 3679 16589 3745 16612
rect 3831 16589 3913 16612
rect 3999 16589 4065 16612
rect 3679 16570 4065 16589
rect 18799 16675 19185 16694
rect 18799 16652 18865 16675
rect 18951 16652 19033 16675
rect 19119 16652 19185 16675
rect 18799 16612 18808 16652
rect 18848 16612 18865 16652
rect 18951 16612 18972 16652
rect 19012 16612 19033 16652
rect 19119 16612 19136 16652
rect 19176 16612 19185 16652
rect 18799 16589 18865 16612
rect 18951 16589 19033 16612
rect 19119 16589 19185 16612
rect 18799 16570 19185 16589
rect 4919 15919 5305 15938
rect 4919 15896 4985 15919
rect 5071 15896 5153 15919
rect 5239 15896 5305 15919
rect 4919 15856 4928 15896
rect 4968 15856 4985 15896
rect 5071 15856 5092 15896
rect 5132 15856 5153 15896
rect 5239 15856 5256 15896
rect 5296 15856 5305 15896
rect 4919 15833 4985 15856
rect 5071 15833 5153 15856
rect 5239 15833 5305 15856
rect 4919 15814 5305 15833
rect 20039 15919 20425 15938
rect 20039 15896 20105 15919
rect 20191 15896 20273 15919
rect 20359 15896 20425 15919
rect 20039 15856 20048 15896
rect 20088 15856 20105 15896
rect 20191 15856 20212 15896
rect 20252 15856 20273 15896
rect 20359 15856 20376 15896
rect 20416 15856 20425 15896
rect 20039 15833 20105 15856
rect 20191 15833 20273 15856
rect 20359 15833 20425 15856
rect 20039 15814 20425 15833
rect 3679 15163 4065 15182
rect 3679 15140 3745 15163
rect 3831 15140 3913 15163
rect 3999 15140 4065 15163
rect 3679 15100 3688 15140
rect 3728 15100 3745 15140
rect 3831 15100 3852 15140
rect 3892 15100 3913 15140
rect 3999 15100 4016 15140
rect 4056 15100 4065 15140
rect 3679 15077 3745 15100
rect 3831 15077 3913 15100
rect 3999 15077 4065 15100
rect 3679 15058 4065 15077
rect 18799 15163 19185 15182
rect 18799 15140 18865 15163
rect 18951 15140 19033 15163
rect 19119 15140 19185 15163
rect 18799 15100 18808 15140
rect 18848 15100 18865 15140
rect 18951 15100 18972 15140
rect 19012 15100 19033 15140
rect 19119 15100 19136 15140
rect 19176 15100 19185 15140
rect 18799 15077 18865 15100
rect 18951 15077 19033 15100
rect 19119 15077 19185 15100
rect 18799 15058 19185 15077
rect 4919 14407 5305 14426
rect 4919 14384 4985 14407
rect 5071 14384 5153 14407
rect 5239 14384 5305 14407
rect 4919 14344 4928 14384
rect 4968 14344 4985 14384
rect 5071 14344 5092 14384
rect 5132 14344 5153 14384
rect 5239 14344 5256 14384
rect 5296 14344 5305 14384
rect 4919 14321 4985 14344
rect 5071 14321 5153 14344
rect 5239 14321 5305 14344
rect 4919 14302 5305 14321
rect 20039 14407 20425 14426
rect 20039 14384 20105 14407
rect 20191 14384 20273 14407
rect 20359 14384 20425 14407
rect 20039 14344 20048 14384
rect 20088 14344 20105 14384
rect 20191 14344 20212 14384
rect 20252 14344 20273 14384
rect 20359 14344 20376 14384
rect 20416 14344 20425 14384
rect 20039 14321 20105 14344
rect 20191 14321 20273 14344
rect 20359 14321 20425 14344
rect 20039 14302 20425 14321
rect 3679 13651 4065 13670
rect 3679 13628 3745 13651
rect 3831 13628 3913 13651
rect 3999 13628 4065 13651
rect 3679 13588 3688 13628
rect 3728 13588 3745 13628
rect 3831 13588 3852 13628
rect 3892 13588 3913 13628
rect 3999 13588 4016 13628
rect 4056 13588 4065 13628
rect 3679 13565 3745 13588
rect 3831 13565 3913 13588
rect 3999 13565 4065 13588
rect 3679 13546 4065 13565
rect 18799 13651 19185 13670
rect 18799 13628 18865 13651
rect 18951 13628 19033 13651
rect 19119 13628 19185 13651
rect 18799 13588 18808 13628
rect 18848 13588 18865 13628
rect 18951 13588 18972 13628
rect 19012 13588 19033 13628
rect 19119 13588 19136 13628
rect 19176 13588 19185 13628
rect 18799 13565 18865 13588
rect 18951 13565 19033 13588
rect 19119 13565 19185 13588
rect 18799 13546 19185 13565
rect 4919 12895 5305 12914
rect 4919 12872 4985 12895
rect 5071 12872 5153 12895
rect 5239 12872 5305 12895
rect 4919 12832 4928 12872
rect 4968 12832 4985 12872
rect 5071 12832 5092 12872
rect 5132 12832 5153 12872
rect 5239 12832 5256 12872
rect 5296 12832 5305 12872
rect 4919 12809 4985 12832
rect 5071 12809 5153 12832
rect 5239 12809 5305 12832
rect 4919 12790 5305 12809
rect 20039 12895 20425 12914
rect 20039 12872 20105 12895
rect 20191 12872 20273 12895
rect 20359 12872 20425 12895
rect 20039 12832 20048 12872
rect 20088 12832 20105 12872
rect 20191 12832 20212 12872
rect 20252 12832 20273 12872
rect 20359 12832 20376 12872
rect 20416 12832 20425 12872
rect 20039 12809 20105 12832
rect 20191 12809 20273 12832
rect 20359 12809 20425 12832
rect 20039 12790 20425 12809
rect 3679 12139 4065 12158
rect 3679 12116 3745 12139
rect 3831 12116 3913 12139
rect 3999 12116 4065 12139
rect 3679 12076 3688 12116
rect 3728 12076 3745 12116
rect 3831 12076 3852 12116
rect 3892 12076 3913 12116
rect 3999 12076 4016 12116
rect 4056 12076 4065 12116
rect 3679 12053 3745 12076
rect 3831 12053 3913 12076
rect 3999 12053 4065 12076
rect 3679 12034 4065 12053
rect 18799 12139 19185 12158
rect 18799 12116 18865 12139
rect 18951 12116 19033 12139
rect 19119 12116 19185 12139
rect 18799 12076 18808 12116
rect 18848 12076 18865 12116
rect 18951 12076 18972 12116
rect 19012 12076 19033 12116
rect 19119 12076 19136 12116
rect 19176 12076 19185 12116
rect 18799 12053 18865 12076
rect 18951 12053 19033 12076
rect 19119 12053 19185 12076
rect 18799 12034 19185 12053
rect 4919 11383 5305 11402
rect 4919 11360 4985 11383
rect 5071 11360 5153 11383
rect 5239 11360 5305 11383
rect 4919 11320 4928 11360
rect 4968 11320 4985 11360
rect 5071 11320 5092 11360
rect 5132 11320 5153 11360
rect 5239 11320 5256 11360
rect 5296 11320 5305 11360
rect 4919 11297 4985 11320
rect 5071 11297 5153 11320
rect 5239 11297 5305 11320
rect 4919 11278 5305 11297
rect 20039 11383 20425 11402
rect 20039 11360 20105 11383
rect 20191 11360 20273 11383
rect 20359 11360 20425 11383
rect 20039 11320 20048 11360
rect 20088 11320 20105 11360
rect 20191 11320 20212 11360
rect 20252 11320 20273 11360
rect 20359 11320 20376 11360
rect 20416 11320 20425 11360
rect 20039 11297 20105 11320
rect 20191 11297 20273 11320
rect 20359 11297 20425 11320
rect 20039 11278 20425 11297
rect 2083 10648 2092 10688
rect 2132 10648 2284 10688
rect 2324 10648 2333 10688
rect 3679 10627 4065 10646
rect 3679 10604 3745 10627
rect 3831 10604 3913 10627
rect 3999 10604 4065 10627
rect 3679 10564 3688 10604
rect 3728 10564 3745 10604
rect 3831 10564 3852 10604
rect 3892 10564 3913 10604
rect 3999 10564 4016 10604
rect 4056 10564 4065 10604
rect 3679 10541 3745 10564
rect 3831 10541 3913 10564
rect 3999 10541 4065 10564
rect 3679 10522 4065 10541
rect 18799 10627 19185 10646
rect 18799 10604 18865 10627
rect 18951 10604 19033 10627
rect 19119 10604 19185 10627
rect 18799 10564 18808 10604
rect 18848 10564 18865 10604
rect 18951 10564 18972 10604
rect 19012 10564 19033 10604
rect 19119 10564 19136 10604
rect 19176 10564 19185 10604
rect 18799 10541 18865 10564
rect 18951 10541 19033 10564
rect 19119 10541 19185 10564
rect 18799 10522 19185 10541
rect 4919 9871 5305 9890
rect 4919 9848 4985 9871
rect 5071 9848 5153 9871
rect 5239 9848 5305 9871
rect 4919 9808 4928 9848
rect 4968 9808 4985 9848
rect 5071 9808 5092 9848
rect 5132 9808 5153 9848
rect 5239 9808 5256 9848
rect 5296 9808 5305 9848
rect 4919 9785 4985 9808
rect 5071 9785 5153 9808
rect 5239 9785 5305 9808
rect 4919 9766 5305 9785
rect 20039 9871 20425 9890
rect 20039 9848 20105 9871
rect 20191 9848 20273 9871
rect 20359 9848 20425 9871
rect 20039 9808 20048 9848
rect 20088 9808 20105 9848
rect 20191 9808 20212 9848
rect 20252 9808 20273 9848
rect 20359 9808 20376 9848
rect 20416 9808 20425 9848
rect 20039 9785 20105 9808
rect 20191 9785 20273 9808
rect 20359 9785 20425 9808
rect 20039 9766 20425 9785
rect 3679 9115 4065 9134
rect 3679 9092 3745 9115
rect 3831 9092 3913 9115
rect 3999 9092 4065 9115
rect 3679 9052 3688 9092
rect 3728 9052 3745 9092
rect 3831 9052 3852 9092
rect 3892 9052 3913 9092
rect 3999 9052 4016 9092
rect 4056 9052 4065 9092
rect 3679 9029 3745 9052
rect 3831 9029 3913 9052
rect 3999 9029 4065 9052
rect 3679 9010 4065 9029
rect 18799 9115 19185 9134
rect 18799 9092 18865 9115
rect 18951 9092 19033 9115
rect 19119 9092 19185 9115
rect 18799 9052 18808 9092
rect 18848 9052 18865 9092
rect 18951 9052 18972 9092
rect 19012 9052 19033 9092
rect 19119 9052 19136 9092
rect 19176 9052 19185 9092
rect 18799 9029 18865 9052
rect 18951 9029 19033 9052
rect 19119 9029 19185 9052
rect 18799 9010 19185 9029
rect 4919 8359 5305 8378
rect 4919 8336 4985 8359
rect 5071 8336 5153 8359
rect 5239 8336 5305 8359
rect 4919 8296 4928 8336
rect 4968 8296 4985 8336
rect 5071 8296 5092 8336
rect 5132 8296 5153 8336
rect 5239 8296 5256 8336
rect 5296 8296 5305 8336
rect 4919 8273 4985 8296
rect 5071 8273 5153 8296
rect 5239 8273 5305 8296
rect 4919 8254 5305 8273
rect 20039 8359 20425 8378
rect 20039 8336 20105 8359
rect 20191 8336 20273 8359
rect 20359 8336 20425 8359
rect 20039 8296 20048 8336
rect 20088 8296 20105 8336
rect 20191 8296 20212 8336
rect 20252 8296 20273 8336
rect 20359 8296 20376 8336
rect 20416 8296 20425 8336
rect 20039 8273 20105 8296
rect 20191 8273 20273 8296
rect 20359 8273 20425 8296
rect 20039 8254 20425 8273
rect 3679 7603 4065 7622
rect 3679 7580 3745 7603
rect 3831 7580 3913 7603
rect 3999 7580 4065 7603
rect 3679 7540 3688 7580
rect 3728 7540 3745 7580
rect 3831 7540 3852 7580
rect 3892 7540 3913 7580
rect 3999 7540 4016 7580
rect 4056 7540 4065 7580
rect 3679 7517 3745 7540
rect 3831 7517 3913 7540
rect 3999 7517 4065 7540
rect 3679 7498 4065 7517
rect 18799 7603 19185 7622
rect 18799 7580 18865 7603
rect 18951 7580 19033 7603
rect 19119 7580 19185 7603
rect 18799 7540 18808 7580
rect 18848 7540 18865 7580
rect 18951 7540 18972 7580
rect 19012 7540 19033 7580
rect 19119 7540 19136 7580
rect 19176 7540 19185 7580
rect 18799 7517 18865 7540
rect 18951 7517 19033 7540
rect 19119 7517 19185 7540
rect 18799 7498 19185 7517
rect 12355 6952 12364 6992
rect 12404 6952 14284 6992
rect 14324 6952 14333 6992
rect 4919 6847 5305 6866
rect 4919 6824 4985 6847
rect 5071 6824 5153 6847
rect 5239 6824 5305 6847
rect 4919 6784 4928 6824
rect 4968 6784 4985 6824
rect 5071 6784 5092 6824
rect 5132 6784 5153 6824
rect 5239 6784 5256 6824
rect 5296 6784 5305 6824
rect 4919 6761 4985 6784
rect 5071 6761 5153 6784
rect 5239 6761 5305 6784
rect 4919 6742 5305 6761
rect 20039 6847 20425 6866
rect 20039 6824 20105 6847
rect 20191 6824 20273 6847
rect 20359 6824 20425 6847
rect 20039 6784 20048 6824
rect 20088 6784 20105 6824
rect 20191 6784 20212 6824
rect 20252 6784 20273 6824
rect 20359 6784 20376 6824
rect 20416 6784 20425 6824
rect 20039 6761 20105 6784
rect 20191 6761 20273 6784
rect 20359 6761 20425 6784
rect 20039 6742 20425 6761
rect 17138 6343 17262 6362
rect 17138 6257 17157 6343
rect 17243 6320 17262 6343
rect 17243 6280 18316 6320
rect 18356 6280 18365 6320
rect 17243 6257 17262 6280
rect 17138 6238 17262 6257
rect 3679 6091 4065 6110
rect 3679 6068 3745 6091
rect 3831 6068 3913 6091
rect 3999 6068 4065 6091
rect 3679 6028 3688 6068
rect 3728 6028 3745 6068
rect 3831 6028 3852 6068
rect 3892 6028 3913 6068
rect 3999 6028 4016 6068
rect 4056 6028 4065 6068
rect 3679 6005 3745 6028
rect 3831 6005 3913 6028
rect 3999 6005 4065 6028
rect 3679 5986 4065 6005
rect 18799 6091 19185 6110
rect 18799 6068 18865 6091
rect 18951 6068 19033 6091
rect 19119 6068 19185 6091
rect 18799 6028 18808 6068
rect 18848 6028 18865 6068
rect 18951 6028 18972 6068
rect 19012 6028 19033 6068
rect 19119 6028 19136 6068
rect 19176 6028 19185 6068
rect 18799 6005 18865 6028
rect 18951 6005 19033 6028
rect 19119 6005 19185 6028
rect 18799 5986 19185 6005
rect 4919 5335 5305 5354
rect 4919 5312 4985 5335
rect 5071 5312 5153 5335
rect 5239 5312 5305 5335
rect 4919 5272 4928 5312
rect 4968 5272 4985 5312
rect 5071 5272 5092 5312
rect 5132 5272 5153 5312
rect 5239 5272 5256 5312
rect 5296 5272 5305 5312
rect 4919 5249 4985 5272
rect 5071 5249 5153 5272
rect 5239 5249 5305 5272
rect 4919 5230 5305 5249
rect 20039 5335 20425 5354
rect 20039 5312 20105 5335
rect 20191 5312 20273 5335
rect 20359 5312 20425 5335
rect 20039 5272 20048 5312
rect 20088 5272 20105 5312
rect 20191 5272 20212 5312
rect 20252 5272 20273 5312
rect 20359 5272 20376 5312
rect 20416 5272 20425 5312
rect 20039 5249 20105 5272
rect 20191 5249 20273 5272
rect 20359 5249 20425 5272
rect 20039 5230 20425 5249
rect 6979 4768 6988 4808
rect 7028 4768 8524 4808
rect 8564 4768 8573 4808
rect 3679 4579 4065 4598
rect 3679 4556 3745 4579
rect 3831 4556 3913 4579
rect 3999 4556 4065 4579
rect 3679 4516 3688 4556
rect 3728 4516 3745 4556
rect 3831 4516 3852 4556
rect 3892 4516 3913 4556
rect 3999 4516 4016 4556
rect 4056 4516 4065 4556
rect 3679 4493 3745 4516
rect 3831 4493 3913 4516
rect 3999 4493 4065 4516
rect 3679 4474 4065 4493
rect 18799 4579 19185 4598
rect 18799 4556 18865 4579
rect 18951 4556 19033 4579
rect 19119 4556 19185 4579
rect 18799 4516 18808 4556
rect 18848 4516 18865 4556
rect 18951 4516 18972 4556
rect 19012 4516 19033 4556
rect 19119 4516 19136 4556
rect 19176 4516 19185 4556
rect 18799 4493 18865 4516
rect 18951 4493 19033 4516
rect 19119 4493 19185 4516
rect 18799 4474 19185 4493
rect 4919 3823 5305 3842
rect 4919 3800 4985 3823
rect 5071 3800 5153 3823
rect 5239 3800 5305 3823
rect 4919 3760 4928 3800
rect 4968 3760 4985 3800
rect 5071 3760 5092 3800
rect 5132 3760 5153 3800
rect 5239 3760 5256 3800
rect 5296 3760 5305 3800
rect 4919 3737 4985 3760
rect 5071 3737 5153 3760
rect 5239 3737 5305 3760
rect 4919 3718 5305 3737
rect 20039 3823 20425 3842
rect 20039 3800 20105 3823
rect 20191 3800 20273 3823
rect 20359 3800 20425 3823
rect 20039 3760 20048 3800
rect 20088 3760 20105 3800
rect 20191 3760 20212 3800
rect 20252 3760 20273 3800
rect 20359 3760 20376 3800
rect 20416 3760 20425 3800
rect 20039 3737 20105 3760
rect 20191 3737 20273 3760
rect 20359 3737 20425 3760
rect 20039 3718 20425 3737
rect 11210 3487 11334 3506
rect 11210 3464 11229 3487
rect 11011 3424 11020 3464
rect 11060 3424 11229 3464
rect 11210 3401 11229 3424
rect 11315 3401 11334 3487
rect 11210 3382 11334 3401
rect 3679 3067 4065 3086
rect 3679 3044 3745 3067
rect 3831 3044 3913 3067
rect 3999 3044 4065 3067
rect 3679 3004 3688 3044
rect 3728 3004 3745 3044
rect 3831 3004 3852 3044
rect 3892 3004 3913 3044
rect 3999 3004 4016 3044
rect 4056 3004 4065 3044
rect 3679 2981 3745 3004
rect 3831 2981 3913 3004
rect 3999 2981 4065 3004
rect 3679 2962 4065 2981
rect 18799 3067 19185 3086
rect 18799 3044 18865 3067
rect 18951 3044 19033 3067
rect 19119 3044 19185 3067
rect 18799 3004 18808 3044
rect 18848 3004 18865 3044
rect 18951 3004 18972 3044
rect 19012 3004 19033 3044
rect 19119 3004 19136 3044
rect 19176 3004 19185 3044
rect 18799 2981 18865 3004
rect 18951 2981 19033 3004
rect 19119 2981 19185 3004
rect 18799 2962 19185 2981
rect 4919 2311 5305 2330
rect 4919 2288 4985 2311
rect 5071 2288 5153 2311
rect 5239 2288 5305 2311
rect 4919 2248 4928 2288
rect 4968 2248 4985 2288
rect 5071 2248 5092 2288
rect 5132 2248 5153 2288
rect 5239 2248 5256 2288
rect 5296 2248 5305 2288
rect 4919 2225 4985 2248
rect 5071 2225 5153 2248
rect 5239 2225 5305 2248
rect 4919 2206 5305 2225
rect 20039 2311 20425 2330
rect 20039 2288 20105 2311
rect 20191 2288 20273 2311
rect 20359 2288 20425 2311
rect 20039 2248 20048 2288
rect 20088 2248 20105 2288
rect 20191 2248 20212 2288
rect 20252 2248 20273 2288
rect 20359 2248 20376 2288
rect 20416 2248 20425 2288
rect 20039 2225 20105 2248
rect 20191 2225 20273 2248
rect 20359 2225 20425 2248
rect 20039 2206 20425 2225
rect 6595 2164 6604 2204
rect 6644 2164 7948 2204
rect 7988 2164 7997 2204
rect 3679 1555 4065 1574
rect 3679 1532 3745 1555
rect 3831 1532 3913 1555
rect 3999 1532 4065 1555
rect 3679 1492 3688 1532
rect 3728 1492 3745 1532
rect 3831 1492 3852 1532
rect 3892 1492 3913 1532
rect 3999 1492 4016 1532
rect 4056 1492 4065 1532
rect 3679 1469 3745 1492
rect 3831 1469 3913 1492
rect 3999 1469 4065 1492
rect 3679 1450 4065 1469
rect 18799 1555 19185 1574
rect 18799 1532 18865 1555
rect 18951 1532 19033 1555
rect 19119 1532 19185 1555
rect 18799 1492 18808 1532
rect 18848 1492 18865 1532
rect 18951 1492 18972 1532
rect 19012 1492 19033 1532
rect 19119 1492 19136 1532
rect 19176 1492 19185 1532
rect 18799 1469 18865 1492
rect 18951 1469 19033 1492
rect 19119 1469 19185 1492
rect 18799 1450 19185 1469
rect 1178 1303 1302 1322
rect 1178 1217 1197 1303
rect 1283 1280 1302 1303
rect 1283 1240 6700 1280
rect 6740 1240 6749 1280
rect 1283 1217 1302 1240
rect 1178 1198 1302 1217
rect 13490 1135 13614 1154
rect 13490 1112 13509 1135
rect 12547 1072 12556 1112
rect 12596 1072 13509 1112
rect 13490 1049 13509 1072
rect 13595 1049 13614 1135
rect 13490 1030 13614 1049
rect 1027 904 1036 944
rect 1076 904 6316 944
rect 6356 904 6365 944
rect 4919 799 5305 818
rect 4919 776 4985 799
rect 5071 776 5153 799
rect 5239 776 5305 799
rect 4919 736 4928 776
rect 4968 736 4985 776
rect 5071 736 5092 776
rect 5132 736 5153 776
rect 5239 736 5256 776
rect 5296 736 5305 776
rect 4919 713 4985 736
rect 5071 713 5153 736
rect 5239 713 5305 736
rect 4919 694 5305 713
rect 20039 799 20425 818
rect 20039 776 20105 799
rect 20191 776 20273 799
rect 20359 776 20425 799
rect 20039 736 20048 776
rect 20088 736 20105 776
rect 20191 736 20212 776
rect 20252 736 20273 776
rect 20359 736 20376 776
rect 20416 736 20425 776
rect 20039 713 20105 736
rect 20191 713 20273 736
rect 20359 713 20425 736
rect 20039 694 20425 713
rect 3715 316 3724 356
rect 3764 316 11980 356
rect 12020 316 12029 356
rect 12122 295 12246 314
rect 12122 272 12141 295
rect 2947 232 2956 272
rect 2996 232 12141 272
rect 12122 209 12141 232
rect 12227 209 12246 295
rect 12122 190 12246 209
rect 5251 148 5260 188
rect 5300 148 10828 188
rect 10868 148 10877 188
<< via5 >>
rect 3745 84692 3831 84715
rect 3913 84692 3999 84715
rect 3745 84652 3770 84692
rect 3770 84652 3810 84692
rect 3810 84652 3831 84692
rect 3913 84652 3934 84692
rect 3934 84652 3974 84692
rect 3974 84652 3999 84692
rect 3745 84629 3831 84652
rect 3913 84629 3999 84652
rect 18865 84692 18951 84715
rect 19033 84692 19119 84715
rect 18865 84652 18890 84692
rect 18890 84652 18930 84692
rect 18930 84652 18951 84692
rect 19033 84652 19054 84692
rect 19054 84652 19094 84692
rect 19094 84652 19119 84692
rect 18865 84629 18951 84652
rect 19033 84629 19119 84652
rect 4985 83936 5071 83959
rect 5153 83936 5239 83959
rect 4985 83896 5010 83936
rect 5010 83896 5050 83936
rect 5050 83896 5071 83936
rect 5153 83896 5174 83936
rect 5174 83896 5214 83936
rect 5214 83896 5239 83936
rect 4985 83873 5071 83896
rect 5153 83873 5239 83896
rect 20105 83936 20191 83959
rect 20273 83936 20359 83959
rect 20105 83896 20130 83936
rect 20130 83896 20170 83936
rect 20170 83896 20191 83936
rect 20273 83896 20294 83936
rect 20294 83896 20334 83936
rect 20334 83896 20359 83936
rect 20105 83873 20191 83896
rect 20273 83873 20359 83896
rect 8037 83453 8123 83539
rect 17157 83453 17243 83539
rect 13509 83285 13595 83371
rect 3745 83180 3831 83203
rect 3913 83180 3999 83203
rect 3745 83140 3770 83180
rect 3770 83140 3810 83180
rect 3810 83140 3831 83180
rect 3913 83140 3934 83180
rect 3934 83140 3974 83180
rect 3974 83140 3999 83180
rect 3745 83117 3831 83140
rect 3913 83117 3999 83140
rect 18865 83180 18951 83203
rect 19033 83180 19119 83203
rect 18865 83140 18890 83180
rect 18890 83140 18930 83180
rect 18930 83140 18951 83180
rect 19033 83140 19054 83180
rect 19054 83140 19094 83180
rect 19094 83140 19119 83180
rect 18865 83117 18951 83140
rect 19033 83117 19119 83140
rect 4985 82424 5071 82447
rect 5153 82424 5239 82447
rect 4985 82384 5010 82424
rect 5010 82384 5050 82424
rect 5050 82384 5071 82424
rect 5153 82384 5174 82424
rect 5174 82384 5214 82424
rect 5214 82384 5239 82424
rect 4985 82361 5071 82384
rect 5153 82361 5239 82384
rect 20105 82424 20191 82447
rect 20273 82424 20359 82447
rect 20105 82384 20130 82424
rect 20130 82384 20170 82424
rect 20170 82384 20191 82424
rect 20273 82384 20294 82424
rect 20294 82384 20334 82424
rect 20334 82384 20359 82424
rect 20105 82361 20191 82384
rect 20273 82361 20359 82384
rect 3745 81668 3831 81691
rect 3913 81668 3999 81691
rect 3745 81628 3770 81668
rect 3770 81628 3810 81668
rect 3810 81628 3831 81668
rect 3913 81628 3934 81668
rect 3934 81628 3974 81668
rect 3974 81628 3999 81668
rect 3745 81605 3831 81628
rect 3913 81605 3999 81628
rect 18865 81668 18951 81691
rect 19033 81668 19119 81691
rect 18865 81628 18890 81668
rect 18890 81628 18930 81668
rect 18930 81628 18951 81668
rect 19033 81628 19054 81668
rect 19054 81628 19094 81668
rect 19094 81628 19119 81668
rect 18865 81605 18951 81628
rect 19033 81605 19119 81628
rect 4985 80912 5071 80935
rect 5153 80912 5239 80935
rect 4985 80872 5010 80912
rect 5010 80872 5050 80912
rect 5050 80872 5071 80912
rect 5153 80872 5174 80912
rect 5174 80872 5214 80912
rect 5214 80872 5239 80912
rect 4985 80849 5071 80872
rect 5153 80849 5239 80872
rect 20105 80912 20191 80935
rect 20273 80912 20359 80935
rect 20105 80872 20130 80912
rect 20130 80872 20170 80912
rect 20170 80872 20191 80912
rect 20273 80872 20294 80912
rect 20294 80872 20334 80912
rect 20334 80872 20359 80912
rect 20105 80849 20191 80872
rect 20273 80849 20359 80872
rect 3745 80156 3831 80179
rect 3913 80156 3999 80179
rect 3745 80116 3770 80156
rect 3770 80116 3810 80156
rect 3810 80116 3831 80156
rect 3913 80116 3934 80156
rect 3934 80116 3974 80156
rect 3974 80116 3999 80156
rect 3745 80093 3831 80116
rect 3913 80093 3999 80116
rect 18865 80156 18951 80179
rect 19033 80156 19119 80179
rect 18865 80116 18890 80156
rect 18890 80116 18930 80156
rect 18930 80116 18951 80156
rect 19033 80116 19054 80156
rect 19054 80116 19094 80156
rect 19094 80116 19119 80156
rect 18865 80093 18951 80116
rect 19033 80093 19119 80116
rect 4985 79400 5071 79423
rect 5153 79400 5239 79423
rect 4985 79360 5010 79400
rect 5010 79360 5050 79400
rect 5050 79360 5071 79400
rect 5153 79360 5174 79400
rect 5174 79360 5214 79400
rect 5214 79360 5239 79400
rect 4985 79337 5071 79360
rect 5153 79337 5239 79360
rect 20105 79400 20191 79423
rect 20273 79400 20359 79423
rect 20105 79360 20130 79400
rect 20130 79360 20170 79400
rect 20170 79360 20191 79400
rect 20273 79360 20294 79400
rect 20294 79360 20334 79400
rect 20334 79360 20359 79400
rect 20105 79337 20191 79360
rect 20273 79337 20359 79360
rect 3745 78644 3831 78667
rect 3913 78644 3999 78667
rect 3745 78604 3770 78644
rect 3770 78604 3810 78644
rect 3810 78604 3831 78644
rect 3913 78604 3934 78644
rect 3934 78604 3974 78644
rect 3974 78604 3999 78644
rect 3745 78581 3831 78604
rect 3913 78581 3999 78604
rect 18865 78644 18951 78667
rect 19033 78644 19119 78667
rect 18865 78604 18890 78644
rect 18890 78604 18930 78644
rect 18930 78604 18951 78644
rect 19033 78604 19054 78644
rect 19054 78604 19094 78644
rect 19094 78604 19119 78644
rect 18865 78581 18951 78604
rect 19033 78581 19119 78604
rect 4985 77888 5071 77911
rect 5153 77888 5239 77911
rect 4985 77848 5010 77888
rect 5010 77848 5050 77888
rect 5050 77848 5071 77888
rect 5153 77848 5174 77888
rect 5174 77848 5214 77888
rect 5214 77848 5239 77888
rect 4985 77825 5071 77848
rect 5153 77825 5239 77848
rect 20105 77888 20191 77911
rect 20273 77888 20359 77911
rect 20105 77848 20130 77888
rect 20130 77848 20170 77888
rect 20170 77848 20191 77888
rect 20273 77848 20294 77888
rect 20294 77848 20334 77888
rect 20334 77848 20359 77888
rect 20105 77825 20191 77848
rect 20273 77825 20359 77848
rect 3745 77132 3831 77155
rect 3913 77132 3999 77155
rect 3745 77092 3770 77132
rect 3770 77092 3810 77132
rect 3810 77092 3831 77132
rect 3913 77092 3934 77132
rect 3934 77092 3974 77132
rect 3974 77092 3999 77132
rect 3745 77069 3831 77092
rect 3913 77069 3999 77092
rect 18865 77132 18951 77155
rect 19033 77132 19119 77155
rect 18865 77092 18890 77132
rect 18890 77092 18930 77132
rect 18930 77092 18951 77132
rect 19033 77092 19054 77132
rect 19054 77092 19094 77132
rect 19094 77092 19119 77132
rect 18865 77069 18951 77092
rect 19033 77069 19119 77092
rect 4985 76376 5071 76399
rect 5153 76376 5239 76399
rect 4985 76336 5010 76376
rect 5010 76336 5050 76376
rect 5050 76336 5071 76376
rect 5153 76336 5174 76376
rect 5174 76336 5214 76376
rect 5214 76336 5239 76376
rect 4985 76313 5071 76336
rect 5153 76313 5239 76336
rect 20105 76376 20191 76399
rect 20273 76376 20359 76399
rect 20105 76336 20130 76376
rect 20130 76336 20170 76376
rect 20170 76336 20191 76376
rect 20273 76336 20294 76376
rect 20294 76336 20334 76376
rect 20334 76336 20359 76376
rect 20105 76313 20191 76336
rect 20273 76313 20359 76336
rect 3745 75620 3831 75643
rect 3913 75620 3999 75643
rect 3745 75580 3770 75620
rect 3770 75580 3810 75620
rect 3810 75580 3831 75620
rect 3913 75580 3934 75620
rect 3934 75580 3974 75620
rect 3974 75580 3999 75620
rect 3745 75557 3831 75580
rect 3913 75557 3999 75580
rect 18865 75620 18951 75643
rect 19033 75620 19119 75643
rect 18865 75580 18890 75620
rect 18890 75580 18930 75620
rect 18930 75580 18951 75620
rect 19033 75580 19054 75620
rect 19054 75580 19094 75620
rect 19094 75580 19119 75620
rect 18865 75557 18951 75580
rect 19033 75557 19119 75580
rect 4985 74864 5071 74887
rect 5153 74864 5239 74887
rect 4985 74824 5010 74864
rect 5010 74824 5050 74864
rect 5050 74824 5071 74864
rect 5153 74824 5174 74864
rect 5174 74824 5214 74864
rect 5214 74824 5239 74864
rect 4985 74801 5071 74824
rect 5153 74801 5239 74824
rect 20105 74864 20191 74887
rect 20273 74864 20359 74887
rect 20105 74824 20130 74864
rect 20130 74824 20170 74864
rect 20170 74824 20191 74864
rect 20273 74824 20294 74864
rect 20294 74824 20334 74864
rect 20334 74824 20359 74864
rect 20105 74801 20191 74824
rect 20273 74801 20359 74824
rect 3745 74108 3831 74131
rect 3913 74108 3999 74131
rect 3745 74068 3770 74108
rect 3770 74068 3810 74108
rect 3810 74068 3831 74108
rect 3913 74068 3934 74108
rect 3934 74068 3974 74108
rect 3974 74068 3999 74108
rect 3745 74045 3831 74068
rect 3913 74045 3999 74068
rect 18865 74108 18951 74131
rect 19033 74108 19119 74131
rect 18865 74068 18890 74108
rect 18890 74068 18930 74108
rect 18930 74068 18951 74108
rect 19033 74068 19054 74108
rect 19054 74068 19094 74108
rect 19094 74068 19119 74108
rect 18865 74045 18951 74068
rect 19033 74045 19119 74068
rect 4985 73352 5071 73375
rect 5153 73352 5239 73375
rect 4985 73312 5010 73352
rect 5010 73312 5050 73352
rect 5050 73312 5071 73352
rect 5153 73312 5174 73352
rect 5174 73312 5214 73352
rect 5214 73312 5239 73352
rect 4985 73289 5071 73312
rect 5153 73289 5239 73312
rect 20105 73352 20191 73375
rect 20273 73352 20359 73375
rect 20105 73312 20130 73352
rect 20130 73312 20170 73352
rect 20170 73312 20191 73352
rect 20273 73312 20294 73352
rect 20294 73312 20334 73352
rect 20334 73312 20359 73352
rect 20105 73289 20191 73312
rect 20273 73289 20359 73312
rect 15333 72701 15419 72787
rect 3745 72596 3831 72619
rect 3913 72596 3999 72619
rect 3745 72556 3770 72596
rect 3770 72556 3810 72596
rect 3810 72556 3831 72596
rect 3913 72556 3934 72596
rect 3934 72556 3974 72596
rect 3974 72556 3999 72596
rect 3745 72533 3831 72556
rect 3913 72533 3999 72556
rect 18865 72596 18951 72619
rect 19033 72596 19119 72619
rect 18865 72556 18890 72596
rect 18890 72556 18930 72596
rect 18930 72556 18951 72596
rect 19033 72556 19054 72596
rect 19054 72556 19094 72596
rect 19094 72556 19119 72596
rect 18865 72533 18951 72556
rect 19033 72533 19119 72556
rect 12141 72113 12227 72199
rect 4985 71840 5071 71863
rect 5153 71840 5239 71863
rect 4985 71800 5010 71840
rect 5010 71800 5050 71840
rect 5050 71800 5071 71840
rect 5153 71800 5174 71840
rect 5174 71800 5214 71840
rect 5214 71800 5239 71840
rect 4985 71777 5071 71800
rect 5153 71777 5239 71800
rect 20105 71840 20191 71863
rect 20273 71840 20359 71863
rect 20105 71800 20130 71840
rect 20130 71800 20170 71840
rect 20170 71800 20191 71840
rect 20273 71800 20294 71840
rect 20294 71800 20334 71840
rect 20334 71800 20359 71840
rect 20105 71777 20191 71800
rect 20273 71777 20359 71800
rect 3745 71084 3831 71107
rect 3913 71084 3999 71107
rect 3745 71044 3770 71084
rect 3770 71044 3810 71084
rect 3810 71044 3831 71084
rect 3913 71044 3934 71084
rect 3934 71044 3974 71084
rect 3974 71044 3999 71084
rect 3745 71021 3831 71044
rect 3913 71021 3999 71044
rect 18865 71084 18951 71107
rect 19033 71084 19119 71107
rect 18865 71044 18890 71084
rect 18890 71044 18930 71084
rect 18930 71044 18951 71084
rect 19033 71044 19054 71084
rect 19054 71044 19094 71084
rect 19094 71044 19119 71084
rect 18865 71021 18951 71044
rect 19033 71021 19119 71044
rect 4985 70328 5071 70351
rect 5153 70328 5239 70351
rect 4985 70288 5010 70328
rect 5010 70288 5050 70328
rect 5050 70288 5071 70328
rect 5153 70288 5174 70328
rect 5174 70288 5214 70328
rect 5214 70288 5239 70328
rect 4985 70265 5071 70288
rect 5153 70265 5239 70288
rect 20105 70328 20191 70351
rect 20273 70328 20359 70351
rect 20105 70288 20130 70328
rect 20130 70288 20170 70328
rect 20170 70288 20191 70328
rect 20273 70288 20294 70328
rect 20294 70288 20334 70328
rect 20334 70288 20359 70328
rect 20105 70265 20191 70288
rect 20273 70265 20359 70288
rect 3745 69572 3831 69595
rect 3913 69572 3999 69595
rect 3745 69532 3770 69572
rect 3770 69532 3810 69572
rect 3810 69532 3831 69572
rect 3913 69532 3934 69572
rect 3934 69532 3974 69572
rect 3974 69532 3999 69572
rect 3745 69509 3831 69532
rect 3913 69509 3999 69532
rect 18865 69572 18951 69595
rect 19033 69572 19119 69595
rect 18865 69532 18890 69572
rect 18890 69532 18930 69572
rect 18930 69532 18951 69572
rect 19033 69532 19054 69572
rect 19054 69532 19094 69572
rect 19094 69532 19119 69572
rect 18865 69509 18951 69532
rect 19033 69509 19119 69532
rect 11229 69257 11315 69343
rect 4985 68816 5071 68839
rect 5153 68816 5239 68839
rect 4985 68776 5010 68816
rect 5010 68776 5050 68816
rect 5050 68776 5071 68816
rect 5153 68776 5174 68816
rect 5174 68776 5214 68816
rect 5214 68776 5239 68816
rect 4985 68753 5071 68776
rect 5153 68753 5239 68776
rect 20105 68816 20191 68839
rect 20273 68816 20359 68839
rect 20105 68776 20130 68816
rect 20130 68776 20170 68816
rect 20170 68776 20191 68816
rect 20273 68776 20294 68816
rect 20294 68776 20334 68816
rect 20334 68776 20359 68816
rect 20105 68753 20191 68776
rect 20273 68753 20359 68776
rect 3745 68060 3831 68083
rect 3913 68060 3999 68083
rect 3745 68020 3770 68060
rect 3770 68020 3810 68060
rect 3810 68020 3831 68060
rect 3913 68020 3934 68060
rect 3934 68020 3974 68060
rect 3974 68020 3999 68060
rect 3745 67997 3831 68020
rect 3913 67997 3999 68020
rect 18865 68060 18951 68083
rect 19033 68060 19119 68083
rect 18865 68020 18890 68060
rect 18890 68020 18930 68060
rect 18930 68020 18951 68060
rect 19033 68020 19054 68060
rect 19054 68020 19094 68060
rect 19094 68020 19119 68060
rect 18865 67997 18951 68020
rect 19033 67997 19119 68020
rect 4985 67304 5071 67327
rect 5153 67304 5239 67327
rect 4985 67264 5010 67304
rect 5010 67264 5050 67304
rect 5050 67264 5071 67304
rect 5153 67264 5174 67304
rect 5174 67264 5214 67304
rect 5214 67264 5239 67304
rect 4985 67241 5071 67264
rect 5153 67241 5239 67264
rect 20105 67304 20191 67327
rect 20273 67304 20359 67327
rect 20105 67264 20130 67304
rect 20130 67264 20170 67304
rect 20170 67264 20191 67304
rect 20273 67264 20294 67304
rect 20294 67264 20334 67304
rect 20334 67264 20359 67304
rect 20105 67241 20191 67264
rect 20273 67241 20359 67264
rect 3745 66548 3831 66571
rect 3913 66548 3999 66571
rect 3745 66508 3770 66548
rect 3770 66508 3810 66548
rect 3810 66508 3831 66548
rect 3913 66508 3934 66548
rect 3934 66508 3974 66548
rect 3974 66508 3999 66548
rect 3745 66485 3831 66508
rect 3913 66485 3999 66508
rect 18865 66548 18951 66571
rect 19033 66548 19119 66571
rect 18865 66508 18890 66548
rect 18890 66508 18930 66548
rect 18930 66508 18951 66548
rect 19033 66508 19054 66548
rect 19054 66508 19094 66548
rect 19094 66508 19119 66548
rect 18865 66485 18951 66508
rect 19033 66485 19119 66508
rect 4985 65792 5071 65815
rect 5153 65792 5239 65815
rect 4985 65752 5010 65792
rect 5010 65752 5050 65792
rect 5050 65752 5071 65792
rect 5153 65752 5174 65792
rect 5174 65752 5214 65792
rect 5214 65752 5239 65792
rect 4985 65729 5071 65752
rect 5153 65729 5239 65752
rect 20105 65792 20191 65815
rect 20273 65792 20359 65815
rect 20105 65752 20130 65792
rect 20130 65752 20170 65792
rect 20170 65752 20191 65792
rect 20273 65752 20294 65792
rect 20294 65752 20334 65792
rect 20334 65752 20359 65792
rect 20105 65729 20191 65752
rect 20273 65729 20359 65752
rect 3745 65036 3831 65059
rect 3913 65036 3999 65059
rect 3745 64996 3770 65036
rect 3770 64996 3810 65036
rect 3810 64996 3831 65036
rect 3913 64996 3934 65036
rect 3934 64996 3974 65036
rect 3974 64996 3999 65036
rect 3745 64973 3831 64996
rect 3913 64973 3999 64996
rect 18865 65036 18951 65059
rect 19033 65036 19119 65059
rect 18865 64996 18890 65036
rect 18890 64996 18930 65036
rect 18930 64996 18951 65036
rect 19033 64996 19054 65036
rect 19054 64996 19094 65036
rect 19094 64996 19119 65036
rect 18865 64973 18951 64996
rect 19033 64973 19119 64996
rect 1197 64385 1283 64471
rect 4985 64280 5071 64303
rect 5153 64280 5239 64303
rect 4985 64240 5010 64280
rect 5010 64240 5050 64280
rect 5050 64240 5071 64280
rect 5153 64240 5174 64280
rect 5174 64240 5214 64280
rect 5214 64240 5239 64280
rect 4985 64217 5071 64240
rect 5153 64217 5239 64240
rect 20105 64280 20191 64303
rect 20273 64280 20359 64303
rect 20105 64240 20130 64280
rect 20130 64240 20170 64280
rect 20170 64240 20191 64280
rect 20273 64240 20294 64280
rect 20294 64240 20334 64280
rect 20334 64240 20359 64280
rect 20105 64217 20191 64240
rect 20273 64217 20359 64240
rect 3745 63524 3831 63547
rect 3913 63524 3999 63547
rect 3745 63484 3770 63524
rect 3770 63484 3810 63524
rect 3810 63484 3831 63524
rect 3913 63484 3934 63524
rect 3934 63484 3974 63524
rect 3974 63484 3999 63524
rect 3745 63461 3831 63484
rect 3913 63461 3999 63484
rect 18865 63524 18951 63547
rect 19033 63524 19119 63547
rect 18865 63484 18890 63524
rect 18890 63484 18930 63524
rect 18930 63484 18951 63524
rect 19033 63484 19054 63524
rect 19054 63484 19094 63524
rect 19094 63484 19119 63524
rect 18865 63461 18951 63484
rect 19033 63461 19119 63484
rect 9861 62957 9947 63043
rect 4985 62768 5071 62791
rect 5153 62768 5239 62791
rect 4985 62728 5010 62768
rect 5010 62728 5050 62768
rect 5050 62728 5071 62768
rect 5153 62728 5174 62768
rect 5174 62728 5214 62768
rect 5214 62728 5239 62768
rect 4985 62705 5071 62728
rect 5153 62705 5239 62728
rect 20105 62768 20191 62791
rect 20273 62768 20359 62791
rect 20105 62728 20130 62768
rect 20130 62728 20170 62768
rect 20170 62728 20191 62768
rect 20273 62728 20294 62768
rect 20294 62728 20334 62768
rect 20334 62728 20359 62768
rect 20105 62705 20191 62728
rect 20273 62705 20359 62728
rect 3745 62012 3831 62035
rect 3913 62012 3999 62035
rect 3745 61972 3770 62012
rect 3770 61972 3810 62012
rect 3810 61972 3831 62012
rect 3913 61972 3934 62012
rect 3934 61972 3974 62012
rect 3974 61972 3999 62012
rect 3745 61949 3831 61972
rect 3913 61949 3999 61972
rect 18865 62012 18951 62035
rect 19033 62012 19119 62035
rect 18865 61972 18890 62012
rect 18890 61972 18930 62012
rect 18930 61972 18951 62012
rect 19033 61972 19054 62012
rect 19054 61972 19094 62012
rect 19094 61972 19119 62012
rect 18865 61949 18951 61972
rect 19033 61949 19119 61972
rect 4985 61256 5071 61279
rect 5153 61256 5239 61279
rect 4985 61216 5010 61256
rect 5010 61216 5050 61256
rect 5050 61216 5071 61256
rect 5153 61216 5174 61256
rect 5174 61216 5214 61256
rect 5214 61216 5239 61256
rect 4985 61193 5071 61216
rect 5153 61193 5239 61216
rect 20105 61256 20191 61279
rect 20273 61256 20359 61279
rect 20105 61216 20130 61256
rect 20130 61216 20170 61256
rect 20170 61216 20191 61256
rect 20273 61216 20294 61256
rect 20294 61216 20334 61256
rect 20334 61216 20359 61256
rect 20105 61193 20191 61216
rect 20273 61193 20359 61216
rect 3745 60500 3831 60523
rect 3913 60500 3999 60523
rect 3745 60460 3770 60500
rect 3770 60460 3810 60500
rect 3810 60460 3831 60500
rect 3913 60460 3934 60500
rect 3934 60460 3974 60500
rect 3974 60460 3999 60500
rect 3745 60437 3831 60460
rect 3913 60437 3999 60460
rect 18865 60500 18951 60523
rect 19033 60500 19119 60523
rect 18865 60460 18890 60500
rect 18890 60460 18930 60500
rect 18930 60460 18951 60500
rect 19033 60460 19054 60500
rect 19054 60460 19094 60500
rect 19094 60460 19119 60500
rect 18865 60437 18951 60460
rect 19033 60437 19119 60460
rect 4985 59744 5071 59767
rect 5153 59744 5239 59767
rect 4985 59704 5010 59744
rect 5010 59704 5050 59744
rect 5050 59704 5071 59744
rect 5153 59704 5174 59744
rect 5174 59704 5214 59744
rect 5214 59704 5239 59744
rect 4985 59681 5071 59704
rect 5153 59681 5239 59704
rect 20105 59744 20191 59767
rect 20273 59744 20359 59767
rect 20105 59704 20130 59744
rect 20130 59704 20170 59744
rect 20170 59704 20191 59744
rect 20273 59704 20294 59744
rect 20294 59704 20334 59744
rect 20334 59704 20359 59744
rect 20105 59681 20191 59704
rect 20273 59681 20359 59704
rect 3745 58988 3831 59011
rect 3913 58988 3999 59011
rect 3745 58948 3770 58988
rect 3770 58948 3810 58988
rect 3810 58948 3831 58988
rect 3913 58948 3934 58988
rect 3934 58948 3974 58988
rect 3974 58948 3999 58988
rect 3745 58925 3831 58948
rect 3913 58925 3999 58948
rect 18865 58988 18951 59011
rect 19033 58988 19119 59011
rect 18865 58948 18890 58988
rect 18890 58948 18930 58988
rect 18930 58948 18951 58988
rect 19033 58948 19054 58988
rect 19054 58948 19094 58988
rect 19094 58948 19119 58988
rect 18865 58925 18951 58948
rect 19033 58925 19119 58948
rect 4985 58232 5071 58255
rect 5153 58232 5239 58255
rect 4985 58192 5010 58232
rect 5010 58192 5050 58232
rect 5050 58192 5071 58232
rect 5153 58192 5174 58232
rect 5174 58192 5214 58232
rect 5214 58192 5239 58232
rect 4985 58169 5071 58192
rect 5153 58169 5239 58192
rect 20105 58232 20191 58255
rect 20273 58232 20359 58255
rect 20105 58192 20130 58232
rect 20130 58192 20170 58232
rect 20170 58192 20191 58232
rect 20273 58192 20294 58232
rect 20294 58192 20334 58232
rect 20334 58192 20359 58232
rect 20105 58169 20191 58192
rect 20273 58169 20359 58192
rect 3745 57476 3831 57499
rect 3913 57476 3999 57499
rect 3745 57436 3770 57476
rect 3770 57436 3810 57476
rect 3810 57436 3831 57476
rect 3913 57436 3934 57476
rect 3934 57436 3974 57476
rect 3974 57436 3999 57476
rect 3745 57413 3831 57436
rect 3913 57413 3999 57436
rect 18865 57476 18951 57499
rect 19033 57476 19119 57499
rect 18865 57436 18890 57476
rect 18890 57436 18930 57476
rect 18930 57436 18951 57476
rect 19033 57436 19054 57476
rect 19054 57436 19094 57476
rect 19094 57436 19119 57476
rect 18865 57413 18951 57436
rect 19033 57413 19119 57436
rect 4985 56720 5071 56743
rect 5153 56720 5239 56743
rect 4985 56680 5010 56720
rect 5010 56680 5050 56720
rect 5050 56680 5071 56720
rect 5153 56680 5174 56720
rect 5174 56680 5214 56720
rect 5214 56680 5239 56720
rect 4985 56657 5071 56680
rect 5153 56657 5239 56680
rect 20105 56720 20191 56743
rect 20273 56720 20359 56743
rect 20105 56680 20130 56720
rect 20130 56680 20170 56720
rect 20170 56680 20191 56720
rect 20273 56680 20294 56720
rect 20294 56680 20334 56720
rect 20334 56680 20359 56720
rect 20105 56657 20191 56680
rect 20273 56657 20359 56680
rect 3745 55964 3831 55987
rect 3913 55964 3999 55987
rect 3745 55924 3770 55964
rect 3770 55924 3810 55964
rect 3810 55924 3831 55964
rect 3913 55924 3934 55964
rect 3934 55924 3974 55964
rect 3974 55924 3999 55964
rect 3745 55901 3831 55924
rect 3913 55901 3999 55924
rect 18865 55964 18951 55987
rect 19033 55964 19119 55987
rect 18865 55924 18890 55964
rect 18890 55924 18930 55964
rect 18930 55924 18951 55964
rect 19033 55924 19054 55964
rect 19054 55924 19094 55964
rect 19094 55924 19119 55964
rect 18865 55901 18951 55924
rect 19033 55901 19119 55924
rect 4985 55208 5071 55231
rect 5153 55208 5239 55231
rect 4985 55168 5010 55208
rect 5010 55168 5050 55208
rect 5050 55168 5071 55208
rect 5153 55168 5174 55208
rect 5174 55168 5214 55208
rect 5214 55168 5239 55208
rect 4985 55145 5071 55168
rect 5153 55145 5239 55168
rect 20105 55208 20191 55231
rect 20273 55208 20359 55231
rect 20105 55168 20130 55208
rect 20130 55168 20170 55208
rect 20170 55168 20191 55208
rect 20273 55168 20294 55208
rect 20294 55168 20334 55208
rect 20334 55168 20359 55208
rect 20105 55145 20191 55168
rect 20273 55145 20359 55168
rect 3745 54452 3831 54475
rect 3913 54452 3999 54475
rect 3745 54412 3770 54452
rect 3770 54412 3810 54452
rect 3810 54412 3831 54452
rect 3913 54412 3934 54452
rect 3934 54412 3974 54452
rect 3974 54412 3999 54452
rect 3745 54389 3831 54412
rect 3913 54389 3999 54412
rect 18865 54452 18951 54475
rect 19033 54452 19119 54475
rect 18865 54412 18890 54452
rect 18890 54412 18930 54452
rect 18930 54412 18951 54452
rect 19033 54412 19054 54452
rect 19054 54412 19094 54452
rect 19094 54412 19119 54452
rect 18865 54389 18951 54412
rect 19033 54389 19119 54412
rect 4985 53696 5071 53719
rect 5153 53696 5239 53719
rect 4985 53656 5010 53696
rect 5010 53656 5050 53696
rect 5050 53656 5071 53696
rect 5153 53656 5174 53696
rect 5174 53656 5214 53696
rect 5214 53656 5239 53696
rect 4985 53633 5071 53656
rect 5153 53633 5239 53656
rect 20105 53696 20191 53719
rect 20273 53696 20359 53719
rect 20105 53656 20130 53696
rect 20130 53656 20170 53696
rect 20170 53656 20191 53696
rect 20273 53656 20294 53696
rect 20294 53656 20334 53696
rect 20334 53656 20359 53696
rect 20105 53633 20191 53656
rect 20273 53633 20359 53656
rect 3745 52940 3831 52963
rect 3913 52940 3999 52963
rect 3745 52900 3770 52940
rect 3770 52900 3810 52940
rect 3810 52900 3831 52940
rect 3913 52900 3934 52940
rect 3934 52900 3974 52940
rect 3974 52900 3999 52940
rect 3745 52877 3831 52900
rect 3913 52877 3999 52900
rect 18865 52940 18951 52963
rect 19033 52940 19119 52963
rect 18865 52900 18890 52940
rect 18890 52900 18930 52940
rect 18930 52900 18951 52940
rect 19033 52900 19054 52940
rect 19054 52900 19094 52940
rect 19094 52900 19119 52940
rect 18865 52877 18951 52900
rect 19033 52877 19119 52900
rect 4985 52184 5071 52207
rect 5153 52184 5239 52207
rect 4985 52144 5010 52184
rect 5010 52144 5050 52184
rect 5050 52144 5071 52184
rect 5153 52144 5174 52184
rect 5174 52144 5214 52184
rect 5214 52144 5239 52184
rect 4985 52121 5071 52144
rect 5153 52121 5239 52144
rect 20105 52184 20191 52207
rect 20273 52184 20359 52207
rect 20105 52144 20130 52184
rect 20130 52144 20170 52184
rect 20170 52144 20191 52184
rect 20273 52144 20294 52184
rect 20294 52144 20334 52184
rect 20334 52144 20359 52184
rect 20105 52121 20191 52144
rect 20273 52121 20359 52144
rect 3745 51428 3831 51451
rect 3913 51428 3999 51451
rect 3745 51388 3770 51428
rect 3770 51388 3810 51428
rect 3810 51388 3831 51428
rect 3913 51388 3934 51428
rect 3934 51388 3974 51428
rect 3974 51388 3999 51428
rect 3745 51365 3831 51388
rect 3913 51365 3999 51388
rect 18865 51428 18951 51451
rect 19033 51428 19119 51451
rect 18865 51388 18890 51428
rect 18890 51388 18930 51428
rect 18930 51388 18951 51428
rect 19033 51388 19054 51428
rect 19054 51388 19094 51428
rect 19094 51388 19119 51428
rect 18865 51365 18951 51388
rect 19033 51365 19119 51388
rect 4985 50672 5071 50695
rect 5153 50672 5239 50695
rect 4985 50632 5010 50672
rect 5010 50632 5050 50672
rect 5050 50632 5071 50672
rect 5153 50632 5174 50672
rect 5174 50632 5214 50672
rect 5214 50632 5239 50672
rect 4985 50609 5071 50632
rect 5153 50609 5239 50632
rect 20105 50672 20191 50695
rect 20273 50672 20359 50695
rect 20105 50632 20130 50672
rect 20130 50632 20170 50672
rect 20170 50632 20191 50672
rect 20273 50632 20294 50672
rect 20294 50632 20334 50672
rect 20334 50632 20359 50672
rect 20105 50609 20191 50632
rect 20273 50609 20359 50632
rect 3745 49916 3831 49939
rect 3913 49916 3999 49939
rect 3745 49876 3770 49916
rect 3770 49876 3810 49916
rect 3810 49876 3831 49916
rect 3913 49876 3934 49916
rect 3934 49876 3974 49916
rect 3974 49876 3999 49916
rect 3745 49853 3831 49876
rect 3913 49853 3999 49876
rect 18865 49916 18951 49939
rect 19033 49916 19119 49939
rect 18865 49876 18890 49916
rect 18890 49876 18930 49916
rect 18930 49876 18951 49916
rect 19033 49876 19054 49916
rect 19054 49876 19094 49916
rect 19094 49876 19119 49916
rect 18865 49853 18951 49876
rect 19033 49853 19119 49876
rect 4985 49160 5071 49183
rect 5153 49160 5239 49183
rect 4985 49120 5010 49160
rect 5010 49120 5050 49160
rect 5050 49120 5071 49160
rect 5153 49120 5174 49160
rect 5174 49120 5214 49160
rect 5214 49120 5239 49160
rect 4985 49097 5071 49120
rect 5153 49097 5239 49120
rect 20105 49160 20191 49183
rect 20273 49160 20359 49183
rect 20105 49120 20130 49160
rect 20130 49120 20170 49160
rect 20170 49120 20191 49160
rect 20273 49120 20294 49160
rect 20294 49120 20334 49160
rect 20334 49120 20359 49160
rect 20105 49097 20191 49120
rect 20273 49097 20359 49120
rect 3745 48404 3831 48427
rect 3913 48404 3999 48427
rect 3745 48364 3770 48404
rect 3770 48364 3810 48404
rect 3810 48364 3831 48404
rect 3913 48364 3934 48404
rect 3934 48364 3974 48404
rect 3974 48364 3999 48404
rect 3745 48341 3831 48364
rect 3913 48341 3999 48364
rect 18865 48404 18951 48427
rect 19033 48404 19119 48427
rect 18865 48364 18890 48404
rect 18890 48364 18930 48404
rect 18930 48364 18951 48404
rect 19033 48364 19054 48404
rect 19054 48364 19094 48404
rect 19094 48364 19119 48404
rect 18865 48341 18951 48364
rect 19033 48341 19119 48364
rect 4985 47648 5071 47671
rect 5153 47648 5239 47671
rect 4985 47608 5010 47648
rect 5010 47608 5050 47648
rect 5050 47608 5071 47648
rect 5153 47608 5174 47648
rect 5174 47608 5214 47648
rect 5214 47608 5239 47648
rect 4985 47585 5071 47608
rect 5153 47585 5239 47608
rect 20105 47648 20191 47671
rect 20273 47648 20359 47671
rect 20105 47608 20130 47648
rect 20130 47608 20170 47648
rect 20170 47608 20191 47648
rect 20273 47608 20294 47648
rect 20294 47608 20334 47648
rect 20334 47608 20359 47648
rect 20105 47585 20191 47608
rect 20273 47585 20359 47608
rect 3745 46892 3831 46915
rect 3913 46892 3999 46915
rect 3745 46852 3770 46892
rect 3770 46852 3810 46892
rect 3810 46852 3831 46892
rect 3913 46852 3934 46892
rect 3934 46852 3974 46892
rect 3974 46852 3999 46892
rect 3745 46829 3831 46852
rect 3913 46829 3999 46852
rect 18865 46892 18951 46915
rect 19033 46892 19119 46915
rect 18865 46852 18890 46892
rect 18890 46852 18930 46892
rect 18930 46852 18951 46892
rect 19033 46852 19054 46892
rect 19054 46852 19094 46892
rect 19094 46852 19119 46892
rect 18865 46829 18951 46852
rect 19033 46829 19119 46852
rect 4985 46136 5071 46159
rect 5153 46136 5239 46159
rect 4985 46096 5010 46136
rect 5010 46096 5050 46136
rect 5050 46096 5071 46136
rect 5153 46096 5174 46136
rect 5174 46096 5214 46136
rect 5214 46096 5239 46136
rect 4985 46073 5071 46096
rect 5153 46073 5239 46096
rect 20105 46136 20191 46159
rect 20273 46136 20359 46159
rect 20105 46096 20130 46136
rect 20130 46096 20170 46136
rect 20170 46096 20191 46136
rect 20273 46096 20294 46136
rect 20294 46096 20334 46136
rect 20334 46096 20359 46136
rect 20105 46073 20191 46096
rect 20273 46073 20359 46096
rect 3745 45380 3831 45403
rect 3913 45380 3999 45403
rect 3745 45340 3770 45380
rect 3770 45340 3810 45380
rect 3810 45340 3831 45380
rect 3913 45340 3934 45380
rect 3934 45340 3974 45380
rect 3974 45340 3999 45380
rect 3745 45317 3831 45340
rect 3913 45317 3999 45340
rect 18865 45380 18951 45403
rect 19033 45380 19119 45403
rect 18865 45340 18890 45380
rect 18890 45340 18930 45380
rect 18930 45340 18951 45380
rect 19033 45340 19054 45380
rect 19054 45340 19094 45380
rect 19094 45340 19119 45380
rect 18865 45317 18951 45340
rect 19033 45317 19119 45340
rect 4985 44624 5071 44647
rect 5153 44624 5239 44647
rect 4985 44584 5010 44624
rect 5010 44584 5050 44624
rect 5050 44584 5071 44624
rect 5153 44584 5174 44624
rect 5174 44584 5214 44624
rect 5214 44584 5239 44624
rect 4985 44561 5071 44584
rect 5153 44561 5239 44584
rect 20105 44624 20191 44647
rect 20273 44624 20359 44647
rect 20105 44584 20130 44624
rect 20130 44584 20170 44624
rect 20170 44584 20191 44624
rect 20273 44584 20294 44624
rect 20294 44584 20334 44624
rect 20334 44584 20359 44624
rect 20105 44561 20191 44584
rect 20273 44561 20359 44584
rect 3745 43868 3831 43891
rect 3913 43868 3999 43891
rect 3745 43828 3770 43868
rect 3770 43828 3810 43868
rect 3810 43828 3831 43868
rect 3913 43828 3934 43868
rect 3934 43828 3974 43868
rect 3974 43828 3999 43868
rect 3745 43805 3831 43828
rect 3913 43805 3999 43828
rect 18865 43868 18951 43891
rect 19033 43868 19119 43891
rect 18865 43828 18890 43868
rect 18890 43828 18930 43868
rect 18930 43828 18951 43868
rect 19033 43828 19054 43868
rect 19054 43828 19094 43868
rect 19094 43828 19119 43868
rect 18865 43805 18951 43828
rect 19033 43805 19119 43828
rect 4985 43112 5071 43135
rect 5153 43112 5239 43135
rect 4985 43072 5010 43112
rect 5010 43072 5050 43112
rect 5050 43072 5071 43112
rect 5153 43072 5174 43112
rect 5174 43072 5214 43112
rect 5214 43072 5239 43112
rect 4985 43049 5071 43072
rect 5153 43049 5239 43072
rect 20105 43112 20191 43135
rect 20273 43112 20359 43135
rect 20105 43072 20130 43112
rect 20130 43072 20170 43112
rect 20170 43072 20191 43112
rect 20273 43072 20294 43112
rect 20294 43072 20334 43112
rect 20334 43072 20359 43112
rect 20105 43049 20191 43072
rect 20273 43049 20359 43072
rect 3745 42356 3831 42379
rect 3913 42356 3999 42379
rect 3745 42316 3770 42356
rect 3770 42316 3810 42356
rect 3810 42316 3831 42356
rect 3913 42316 3934 42356
rect 3934 42316 3974 42356
rect 3974 42316 3999 42356
rect 3745 42293 3831 42316
rect 3913 42293 3999 42316
rect 18865 42356 18951 42379
rect 19033 42356 19119 42379
rect 18865 42316 18890 42356
rect 18890 42316 18930 42356
rect 18930 42316 18951 42356
rect 19033 42316 19054 42356
rect 19054 42316 19094 42356
rect 19094 42316 19119 42356
rect 18865 42293 18951 42316
rect 19033 42293 19119 42316
rect 4985 41600 5071 41623
rect 5153 41600 5239 41623
rect 4985 41560 5010 41600
rect 5010 41560 5050 41600
rect 5050 41560 5071 41600
rect 5153 41560 5174 41600
rect 5174 41560 5214 41600
rect 5214 41560 5239 41600
rect 4985 41537 5071 41560
rect 5153 41537 5239 41560
rect 20105 41600 20191 41623
rect 20273 41600 20359 41623
rect 20105 41560 20130 41600
rect 20130 41560 20170 41600
rect 20170 41560 20191 41600
rect 20273 41560 20294 41600
rect 20294 41560 20334 41600
rect 20334 41560 20359 41600
rect 20105 41537 20191 41560
rect 20273 41537 20359 41560
rect 3745 40844 3831 40867
rect 3913 40844 3999 40867
rect 3745 40804 3770 40844
rect 3770 40804 3810 40844
rect 3810 40804 3831 40844
rect 3913 40804 3934 40844
rect 3934 40804 3974 40844
rect 3974 40804 3999 40844
rect 3745 40781 3831 40804
rect 3913 40781 3999 40804
rect 18865 40844 18951 40867
rect 19033 40844 19119 40867
rect 18865 40804 18890 40844
rect 18890 40804 18930 40844
rect 18930 40804 18951 40844
rect 19033 40804 19054 40844
rect 19054 40804 19094 40844
rect 19094 40804 19119 40844
rect 18865 40781 18951 40804
rect 19033 40781 19119 40804
rect 4985 40088 5071 40111
rect 5153 40088 5239 40111
rect 4985 40048 5010 40088
rect 5010 40048 5050 40088
rect 5050 40048 5071 40088
rect 5153 40048 5174 40088
rect 5174 40048 5214 40088
rect 5214 40048 5239 40088
rect 4985 40025 5071 40048
rect 5153 40025 5239 40048
rect 20105 40088 20191 40111
rect 20273 40088 20359 40111
rect 20105 40048 20130 40088
rect 20130 40048 20170 40088
rect 20170 40048 20191 40088
rect 20273 40048 20294 40088
rect 20294 40048 20334 40088
rect 20334 40048 20359 40088
rect 20105 40025 20191 40048
rect 20273 40025 20359 40048
rect 3745 39332 3831 39355
rect 3913 39332 3999 39355
rect 3745 39292 3770 39332
rect 3770 39292 3810 39332
rect 3810 39292 3831 39332
rect 3913 39292 3934 39332
rect 3934 39292 3974 39332
rect 3974 39292 3999 39332
rect 3745 39269 3831 39292
rect 3913 39269 3999 39292
rect 18865 39332 18951 39355
rect 19033 39332 19119 39355
rect 18865 39292 18890 39332
rect 18890 39292 18930 39332
rect 18930 39292 18951 39332
rect 19033 39292 19054 39332
rect 19054 39292 19094 39332
rect 19094 39292 19119 39332
rect 18865 39269 18951 39292
rect 19033 39269 19119 39292
rect 4985 38576 5071 38599
rect 5153 38576 5239 38599
rect 4985 38536 5010 38576
rect 5010 38536 5050 38576
rect 5050 38536 5071 38576
rect 5153 38536 5174 38576
rect 5174 38536 5214 38576
rect 5214 38536 5239 38576
rect 4985 38513 5071 38536
rect 5153 38513 5239 38536
rect 20105 38576 20191 38599
rect 20273 38576 20359 38599
rect 20105 38536 20130 38576
rect 20130 38536 20170 38576
rect 20170 38536 20191 38576
rect 20273 38536 20294 38576
rect 20294 38536 20334 38576
rect 20334 38536 20359 38576
rect 20105 38513 20191 38536
rect 20273 38513 20359 38536
rect 3745 37820 3831 37843
rect 3913 37820 3999 37843
rect 3745 37780 3770 37820
rect 3770 37780 3810 37820
rect 3810 37780 3831 37820
rect 3913 37780 3934 37820
rect 3934 37780 3974 37820
rect 3974 37780 3999 37820
rect 3745 37757 3831 37780
rect 3913 37757 3999 37780
rect 18865 37820 18951 37843
rect 19033 37820 19119 37843
rect 18865 37780 18890 37820
rect 18890 37780 18930 37820
rect 18930 37780 18951 37820
rect 19033 37780 19054 37820
rect 19054 37780 19094 37820
rect 19094 37780 19119 37820
rect 18865 37757 18951 37780
rect 19033 37757 19119 37780
rect 4985 37064 5071 37087
rect 5153 37064 5239 37087
rect 4985 37024 5010 37064
rect 5010 37024 5050 37064
rect 5050 37024 5071 37064
rect 5153 37024 5174 37064
rect 5174 37024 5214 37064
rect 5214 37024 5239 37064
rect 4985 37001 5071 37024
rect 5153 37001 5239 37024
rect 20105 37064 20191 37087
rect 20273 37064 20359 37087
rect 20105 37024 20130 37064
rect 20130 37024 20170 37064
rect 20170 37024 20191 37064
rect 20273 37024 20294 37064
rect 20294 37024 20334 37064
rect 20334 37024 20359 37064
rect 20105 37001 20191 37024
rect 20273 37001 20359 37024
rect 3745 36308 3831 36331
rect 3913 36308 3999 36331
rect 3745 36268 3770 36308
rect 3770 36268 3810 36308
rect 3810 36268 3831 36308
rect 3913 36268 3934 36308
rect 3934 36268 3974 36308
rect 3974 36268 3999 36308
rect 3745 36245 3831 36268
rect 3913 36245 3999 36268
rect 18865 36308 18951 36331
rect 19033 36308 19119 36331
rect 18865 36268 18890 36308
rect 18890 36268 18930 36308
rect 18930 36268 18951 36308
rect 19033 36268 19054 36308
rect 19054 36268 19094 36308
rect 19094 36268 19119 36308
rect 18865 36245 18951 36268
rect 19033 36245 19119 36268
rect 4985 35552 5071 35575
rect 5153 35552 5239 35575
rect 4985 35512 5010 35552
rect 5010 35512 5050 35552
rect 5050 35512 5071 35552
rect 5153 35512 5174 35552
rect 5174 35512 5214 35552
rect 5214 35512 5239 35552
rect 4985 35489 5071 35512
rect 5153 35489 5239 35512
rect 20105 35552 20191 35575
rect 20273 35552 20359 35575
rect 20105 35512 20130 35552
rect 20130 35512 20170 35552
rect 20170 35512 20191 35552
rect 20273 35512 20294 35552
rect 20294 35512 20334 35552
rect 20334 35512 20359 35552
rect 20105 35489 20191 35512
rect 20273 35489 20359 35512
rect 3745 34796 3831 34819
rect 3913 34796 3999 34819
rect 3745 34756 3770 34796
rect 3770 34756 3810 34796
rect 3810 34756 3831 34796
rect 3913 34756 3934 34796
rect 3934 34756 3974 34796
rect 3974 34756 3999 34796
rect 3745 34733 3831 34756
rect 3913 34733 3999 34756
rect 18865 34796 18951 34819
rect 19033 34796 19119 34819
rect 18865 34756 18890 34796
rect 18890 34756 18930 34796
rect 18930 34756 18951 34796
rect 19033 34756 19054 34796
rect 19054 34756 19094 34796
rect 19094 34756 19119 34796
rect 18865 34733 18951 34756
rect 19033 34733 19119 34756
rect 4985 34040 5071 34063
rect 5153 34040 5239 34063
rect 4985 34000 5010 34040
rect 5010 34000 5050 34040
rect 5050 34000 5071 34040
rect 5153 34000 5174 34040
rect 5174 34000 5214 34040
rect 5214 34000 5239 34040
rect 4985 33977 5071 34000
rect 5153 33977 5239 34000
rect 20105 34040 20191 34063
rect 20273 34040 20359 34063
rect 20105 34000 20130 34040
rect 20130 34000 20170 34040
rect 20170 34000 20191 34040
rect 20273 34000 20294 34040
rect 20294 34000 20334 34040
rect 20334 34000 20359 34040
rect 20105 33977 20191 34000
rect 20273 33977 20359 34000
rect 3745 33284 3831 33307
rect 3913 33284 3999 33307
rect 3745 33244 3770 33284
rect 3770 33244 3810 33284
rect 3810 33244 3831 33284
rect 3913 33244 3934 33284
rect 3934 33244 3974 33284
rect 3974 33244 3999 33284
rect 3745 33221 3831 33244
rect 3913 33221 3999 33244
rect 18865 33284 18951 33307
rect 19033 33284 19119 33307
rect 18865 33244 18890 33284
rect 18890 33244 18930 33284
rect 18930 33244 18951 33284
rect 19033 33244 19054 33284
rect 19054 33244 19094 33284
rect 19094 33244 19119 33284
rect 18865 33221 18951 33244
rect 19033 33221 19119 33244
rect 4985 32528 5071 32551
rect 5153 32528 5239 32551
rect 4985 32488 5010 32528
rect 5010 32488 5050 32528
rect 5050 32488 5071 32528
rect 5153 32488 5174 32528
rect 5174 32488 5214 32528
rect 5214 32488 5239 32528
rect 4985 32465 5071 32488
rect 5153 32465 5239 32488
rect 20105 32528 20191 32551
rect 20273 32528 20359 32551
rect 20105 32488 20130 32528
rect 20130 32488 20170 32528
rect 20170 32488 20191 32528
rect 20273 32488 20294 32528
rect 20294 32488 20334 32528
rect 20334 32488 20359 32528
rect 20105 32465 20191 32488
rect 20273 32465 20359 32488
rect 3745 31772 3831 31795
rect 3913 31772 3999 31795
rect 3745 31732 3770 31772
rect 3770 31732 3810 31772
rect 3810 31732 3831 31772
rect 3913 31732 3934 31772
rect 3934 31732 3974 31772
rect 3974 31732 3999 31772
rect 3745 31709 3831 31732
rect 3913 31709 3999 31732
rect 18865 31772 18951 31795
rect 19033 31772 19119 31795
rect 18865 31732 18890 31772
rect 18890 31732 18930 31772
rect 18930 31732 18951 31772
rect 19033 31732 19054 31772
rect 19054 31732 19094 31772
rect 19094 31732 19119 31772
rect 18865 31709 18951 31732
rect 19033 31709 19119 31732
rect 4985 31016 5071 31039
rect 5153 31016 5239 31039
rect 4985 30976 5010 31016
rect 5010 30976 5050 31016
rect 5050 30976 5071 31016
rect 5153 30976 5174 31016
rect 5174 30976 5214 31016
rect 5214 30976 5239 31016
rect 4985 30953 5071 30976
rect 5153 30953 5239 30976
rect 20105 31016 20191 31039
rect 20273 31016 20359 31039
rect 20105 30976 20130 31016
rect 20130 30976 20170 31016
rect 20170 30976 20191 31016
rect 20273 30976 20294 31016
rect 20294 30976 20334 31016
rect 20334 30976 20359 31016
rect 20105 30953 20191 30976
rect 20273 30953 20359 30976
rect 12141 30617 12227 30703
rect 3745 30260 3831 30283
rect 3913 30260 3999 30283
rect 3745 30220 3770 30260
rect 3770 30220 3810 30260
rect 3810 30220 3831 30260
rect 3913 30220 3934 30260
rect 3934 30220 3974 30260
rect 3974 30220 3999 30260
rect 3745 30197 3831 30220
rect 3913 30197 3999 30220
rect 18865 30260 18951 30283
rect 19033 30260 19119 30283
rect 18865 30220 18890 30260
rect 18890 30220 18930 30260
rect 18930 30220 18951 30260
rect 19033 30220 19054 30260
rect 19054 30220 19094 30260
rect 19094 30220 19119 30260
rect 18865 30197 18951 30220
rect 19033 30197 19119 30220
rect 4985 29504 5071 29527
rect 5153 29504 5239 29527
rect 4985 29464 5010 29504
rect 5010 29464 5050 29504
rect 5050 29464 5071 29504
rect 5153 29464 5174 29504
rect 5174 29464 5214 29504
rect 5214 29464 5239 29504
rect 4985 29441 5071 29464
rect 5153 29441 5239 29464
rect 20105 29504 20191 29527
rect 20273 29504 20359 29527
rect 20105 29464 20130 29504
rect 20130 29464 20170 29504
rect 20170 29464 20191 29504
rect 20273 29464 20294 29504
rect 20294 29464 20334 29504
rect 20334 29464 20359 29504
rect 20105 29441 20191 29464
rect 20273 29441 20359 29464
rect 3745 28748 3831 28771
rect 3913 28748 3999 28771
rect 3745 28708 3770 28748
rect 3770 28708 3810 28748
rect 3810 28708 3831 28748
rect 3913 28708 3934 28748
rect 3934 28708 3974 28748
rect 3974 28708 3999 28748
rect 3745 28685 3831 28708
rect 3913 28685 3999 28708
rect 18865 28748 18951 28771
rect 19033 28748 19119 28771
rect 18865 28708 18890 28748
rect 18890 28708 18930 28748
rect 18930 28708 18951 28748
rect 19033 28708 19054 28748
rect 19054 28708 19094 28748
rect 19094 28708 19119 28748
rect 18865 28685 18951 28708
rect 19033 28685 19119 28708
rect 4985 27992 5071 28015
rect 5153 27992 5239 28015
rect 4985 27952 5010 27992
rect 5010 27952 5050 27992
rect 5050 27952 5071 27992
rect 5153 27952 5174 27992
rect 5174 27952 5214 27992
rect 5214 27952 5239 27992
rect 4985 27929 5071 27952
rect 5153 27929 5239 27952
rect 20105 27992 20191 28015
rect 20273 27992 20359 28015
rect 20105 27952 20130 27992
rect 20130 27952 20170 27992
rect 20170 27952 20191 27992
rect 20273 27952 20294 27992
rect 20294 27952 20334 27992
rect 20334 27952 20359 27992
rect 20105 27929 20191 27952
rect 20273 27929 20359 27952
rect 3745 27236 3831 27259
rect 3913 27236 3999 27259
rect 3745 27196 3770 27236
rect 3770 27196 3810 27236
rect 3810 27196 3831 27236
rect 3913 27196 3934 27236
rect 3934 27196 3974 27236
rect 3974 27196 3999 27236
rect 3745 27173 3831 27196
rect 3913 27173 3999 27196
rect 18865 27236 18951 27259
rect 19033 27236 19119 27259
rect 18865 27196 18890 27236
rect 18890 27196 18930 27236
rect 18930 27196 18951 27236
rect 19033 27196 19054 27236
rect 19054 27196 19094 27236
rect 19094 27196 19119 27236
rect 18865 27173 18951 27196
rect 19033 27173 19119 27196
rect 4985 26480 5071 26503
rect 5153 26480 5239 26503
rect 4985 26440 5010 26480
rect 5010 26440 5050 26480
rect 5050 26440 5071 26480
rect 5153 26440 5174 26480
rect 5174 26440 5214 26480
rect 5214 26440 5239 26480
rect 4985 26417 5071 26440
rect 5153 26417 5239 26440
rect 9861 26417 9947 26503
rect 20105 26480 20191 26503
rect 20273 26480 20359 26503
rect 20105 26440 20130 26480
rect 20130 26440 20170 26480
rect 20170 26440 20191 26480
rect 20273 26440 20294 26480
rect 20294 26440 20334 26480
rect 20334 26440 20359 26480
rect 20105 26417 20191 26440
rect 20273 26417 20359 26440
rect 8037 26249 8123 26335
rect 3745 25724 3831 25747
rect 3913 25724 3999 25747
rect 3745 25684 3770 25724
rect 3770 25684 3810 25724
rect 3810 25684 3831 25724
rect 3913 25684 3934 25724
rect 3934 25684 3974 25724
rect 3974 25684 3999 25724
rect 3745 25661 3831 25684
rect 3913 25661 3999 25684
rect 18865 25724 18951 25747
rect 19033 25724 19119 25747
rect 18865 25684 18890 25724
rect 18890 25684 18930 25724
rect 18930 25684 18951 25724
rect 19033 25684 19054 25724
rect 19054 25684 19094 25724
rect 19094 25684 19119 25724
rect 18865 25661 18951 25684
rect 19033 25661 19119 25684
rect 4985 24968 5071 24991
rect 5153 24968 5239 24991
rect 4985 24928 5010 24968
rect 5010 24928 5050 24968
rect 5050 24928 5071 24968
rect 5153 24928 5174 24968
rect 5174 24928 5214 24968
rect 5214 24928 5239 24968
rect 4985 24905 5071 24928
rect 5153 24905 5239 24928
rect 20105 24968 20191 24991
rect 20273 24968 20359 24991
rect 20105 24928 20130 24968
rect 20130 24928 20170 24968
rect 20170 24928 20191 24968
rect 20273 24928 20294 24968
rect 20294 24928 20334 24968
rect 20334 24928 20359 24968
rect 20105 24905 20191 24928
rect 20273 24905 20359 24928
rect 3745 24212 3831 24235
rect 3913 24212 3999 24235
rect 3745 24172 3770 24212
rect 3770 24172 3810 24212
rect 3810 24172 3831 24212
rect 3913 24172 3934 24212
rect 3934 24172 3974 24212
rect 3974 24172 3999 24212
rect 3745 24149 3831 24172
rect 3913 24149 3999 24172
rect 18865 24212 18951 24235
rect 19033 24212 19119 24235
rect 18865 24172 18890 24212
rect 18890 24172 18930 24212
rect 18930 24172 18951 24212
rect 19033 24172 19054 24212
rect 19054 24172 19094 24212
rect 19094 24172 19119 24212
rect 18865 24149 18951 24172
rect 19033 24149 19119 24172
rect 4985 23456 5071 23479
rect 5153 23456 5239 23479
rect 4985 23416 5010 23456
rect 5010 23416 5050 23456
rect 5050 23416 5071 23456
rect 5153 23416 5174 23456
rect 5174 23416 5214 23456
rect 5214 23416 5239 23456
rect 4985 23393 5071 23416
rect 5153 23393 5239 23416
rect 20105 23456 20191 23479
rect 20273 23456 20359 23479
rect 20105 23416 20130 23456
rect 20130 23416 20170 23456
rect 20170 23416 20191 23456
rect 20273 23416 20294 23456
rect 20294 23416 20334 23456
rect 20334 23416 20359 23456
rect 20105 23393 20191 23416
rect 20273 23393 20359 23416
rect 3745 22700 3831 22723
rect 3913 22700 3999 22723
rect 3745 22660 3770 22700
rect 3770 22660 3810 22700
rect 3810 22660 3831 22700
rect 3913 22660 3934 22700
rect 3934 22660 3974 22700
rect 3974 22660 3999 22700
rect 3745 22637 3831 22660
rect 3913 22637 3999 22660
rect 18865 22700 18951 22723
rect 19033 22700 19119 22723
rect 18865 22660 18890 22700
rect 18890 22660 18930 22700
rect 18930 22660 18951 22700
rect 19033 22660 19054 22700
rect 19054 22660 19094 22700
rect 19094 22660 19119 22700
rect 18865 22637 18951 22660
rect 19033 22637 19119 22660
rect 4985 21944 5071 21967
rect 5153 21944 5239 21967
rect 4985 21904 5010 21944
rect 5010 21904 5050 21944
rect 5050 21904 5071 21944
rect 5153 21904 5174 21944
rect 5174 21904 5214 21944
rect 5214 21904 5239 21944
rect 4985 21881 5071 21904
rect 5153 21881 5239 21904
rect 20105 21944 20191 21967
rect 20273 21944 20359 21967
rect 20105 21904 20130 21944
rect 20130 21904 20170 21944
rect 20170 21904 20191 21944
rect 20273 21904 20294 21944
rect 20294 21904 20334 21944
rect 20334 21904 20359 21944
rect 20105 21881 20191 21904
rect 20273 21881 20359 21904
rect 3745 21188 3831 21211
rect 3913 21188 3999 21211
rect 3745 21148 3770 21188
rect 3770 21148 3810 21188
rect 3810 21148 3831 21188
rect 3913 21148 3934 21188
rect 3934 21148 3974 21188
rect 3974 21148 3999 21188
rect 3745 21125 3831 21148
rect 3913 21125 3999 21148
rect 18865 21188 18951 21211
rect 19033 21188 19119 21211
rect 18865 21148 18890 21188
rect 18890 21148 18930 21188
rect 18930 21148 18951 21188
rect 19033 21148 19054 21188
rect 19054 21148 19094 21188
rect 19094 21148 19119 21188
rect 18865 21125 18951 21148
rect 19033 21125 19119 21148
rect 4985 20432 5071 20455
rect 5153 20432 5239 20455
rect 4985 20392 5010 20432
rect 5010 20392 5050 20432
rect 5050 20392 5071 20432
rect 5153 20392 5174 20432
rect 5174 20392 5214 20432
rect 5214 20392 5239 20432
rect 4985 20369 5071 20392
rect 5153 20369 5239 20392
rect 20105 20432 20191 20455
rect 20273 20432 20359 20455
rect 20105 20392 20130 20432
rect 20130 20392 20170 20432
rect 20170 20392 20191 20432
rect 20273 20392 20294 20432
rect 20294 20392 20334 20432
rect 20334 20392 20359 20432
rect 20105 20369 20191 20392
rect 20273 20369 20359 20392
rect 3745 19676 3831 19699
rect 3913 19676 3999 19699
rect 3745 19636 3770 19676
rect 3770 19636 3810 19676
rect 3810 19636 3831 19676
rect 3913 19636 3934 19676
rect 3934 19636 3974 19676
rect 3974 19636 3999 19676
rect 3745 19613 3831 19636
rect 3913 19613 3999 19636
rect 18865 19676 18951 19699
rect 19033 19676 19119 19699
rect 18865 19636 18890 19676
rect 18890 19636 18930 19676
rect 18930 19636 18951 19676
rect 19033 19636 19054 19676
rect 19054 19636 19094 19676
rect 19094 19636 19119 19676
rect 18865 19613 18951 19636
rect 19033 19613 19119 19636
rect 4985 18920 5071 18943
rect 5153 18920 5239 18943
rect 4985 18880 5010 18920
rect 5010 18880 5050 18920
rect 5050 18880 5071 18920
rect 5153 18880 5174 18920
rect 5174 18880 5214 18920
rect 5214 18880 5239 18920
rect 4985 18857 5071 18880
rect 5153 18857 5239 18880
rect 20105 18920 20191 18943
rect 20273 18920 20359 18943
rect 20105 18880 20130 18920
rect 20130 18880 20170 18920
rect 20170 18880 20191 18920
rect 20273 18880 20294 18920
rect 20294 18880 20334 18920
rect 20334 18880 20359 18920
rect 20105 18857 20191 18880
rect 20273 18857 20359 18880
rect 3745 18164 3831 18187
rect 3913 18164 3999 18187
rect 3745 18124 3770 18164
rect 3770 18124 3810 18164
rect 3810 18124 3831 18164
rect 3913 18124 3934 18164
rect 3934 18124 3974 18164
rect 3974 18124 3999 18164
rect 3745 18101 3831 18124
rect 3913 18101 3999 18124
rect 18865 18164 18951 18187
rect 19033 18164 19119 18187
rect 18865 18124 18890 18164
rect 18890 18124 18930 18164
rect 18930 18124 18951 18164
rect 19033 18124 19054 18164
rect 19054 18124 19094 18164
rect 19094 18124 19119 18164
rect 18865 18101 18951 18124
rect 19033 18101 19119 18124
rect 15333 17597 15419 17683
rect 4985 17408 5071 17431
rect 5153 17408 5239 17431
rect 4985 17368 5010 17408
rect 5010 17368 5050 17408
rect 5050 17368 5071 17408
rect 5153 17368 5174 17408
rect 5174 17368 5214 17408
rect 5214 17368 5239 17408
rect 4985 17345 5071 17368
rect 5153 17345 5239 17368
rect 20105 17408 20191 17431
rect 20273 17408 20359 17431
rect 20105 17368 20130 17408
rect 20130 17368 20170 17408
rect 20170 17368 20191 17408
rect 20273 17368 20294 17408
rect 20294 17368 20334 17408
rect 20334 17368 20359 17408
rect 20105 17345 20191 17368
rect 20273 17345 20359 17368
rect 3745 16652 3831 16675
rect 3913 16652 3999 16675
rect 3745 16612 3770 16652
rect 3770 16612 3810 16652
rect 3810 16612 3831 16652
rect 3913 16612 3934 16652
rect 3934 16612 3974 16652
rect 3974 16612 3999 16652
rect 3745 16589 3831 16612
rect 3913 16589 3999 16612
rect 18865 16652 18951 16675
rect 19033 16652 19119 16675
rect 18865 16612 18890 16652
rect 18890 16612 18930 16652
rect 18930 16612 18951 16652
rect 19033 16612 19054 16652
rect 19054 16612 19094 16652
rect 19094 16612 19119 16652
rect 18865 16589 18951 16612
rect 19033 16589 19119 16612
rect 4985 15896 5071 15919
rect 5153 15896 5239 15919
rect 4985 15856 5010 15896
rect 5010 15856 5050 15896
rect 5050 15856 5071 15896
rect 5153 15856 5174 15896
rect 5174 15856 5214 15896
rect 5214 15856 5239 15896
rect 4985 15833 5071 15856
rect 5153 15833 5239 15856
rect 20105 15896 20191 15919
rect 20273 15896 20359 15919
rect 20105 15856 20130 15896
rect 20130 15856 20170 15896
rect 20170 15856 20191 15896
rect 20273 15856 20294 15896
rect 20294 15856 20334 15896
rect 20334 15856 20359 15896
rect 20105 15833 20191 15856
rect 20273 15833 20359 15856
rect 3745 15140 3831 15163
rect 3913 15140 3999 15163
rect 3745 15100 3770 15140
rect 3770 15100 3810 15140
rect 3810 15100 3831 15140
rect 3913 15100 3934 15140
rect 3934 15100 3974 15140
rect 3974 15100 3999 15140
rect 3745 15077 3831 15100
rect 3913 15077 3999 15100
rect 18865 15140 18951 15163
rect 19033 15140 19119 15163
rect 18865 15100 18890 15140
rect 18890 15100 18930 15140
rect 18930 15100 18951 15140
rect 19033 15100 19054 15140
rect 19054 15100 19094 15140
rect 19094 15100 19119 15140
rect 18865 15077 18951 15100
rect 19033 15077 19119 15100
rect 4985 14384 5071 14407
rect 5153 14384 5239 14407
rect 4985 14344 5010 14384
rect 5010 14344 5050 14384
rect 5050 14344 5071 14384
rect 5153 14344 5174 14384
rect 5174 14344 5214 14384
rect 5214 14344 5239 14384
rect 4985 14321 5071 14344
rect 5153 14321 5239 14344
rect 20105 14384 20191 14407
rect 20273 14384 20359 14407
rect 20105 14344 20130 14384
rect 20130 14344 20170 14384
rect 20170 14344 20191 14384
rect 20273 14344 20294 14384
rect 20294 14344 20334 14384
rect 20334 14344 20359 14384
rect 20105 14321 20191 14344
rect 20273 14321 20359 14344
rect 3745 13628 3831 13651
rect 3913 13628 3999 13651
rect 3745 13588 3770 13628
rect 3770 13588 3810 13628
rect 3810 13588 3831 13628
rect 3913 13588 3934 13628
rect 3934 13588 3974 13628
rect 3974 13588 3999 13628
rect 3745 13565 3831 13588
rect 3913 13565 3999 13588
rect 18865 13628 18951 13651
rect 19033 13628 19119 13651
rect 18865 13588 18890 13628
rect 18890 13588 18930 13628
rect 18930 13588 18951 13628
rect 19033 13588 19054 13628
rect 19054 13588 19094 13628
rect 19094 13588 19119 13628
rect 18865 13565 18951 13588
rect 19033 13565 19119 13588
rect 4985 12872 5071 12895
rect 5153 12872 5239 12895
rect 4985 12832 5010 12872
rect 5010 12832 5050 12872
rect 5050 12832 5071 12872
rect 5153 12832 5174 12872
rect 5174 12832 5214 12872
rect 5214 12832 5239 12872
rect 4985 12809 5071 12832
rect 5153 12809 5239 12832
rect 20105 12872 20191 12895
rect 20273 12872 20359 12895
rect 20105 12832 20130 12872
rect 20130 12832 20170 12872
rect 20170 12832 20191 12872
rect 20273 12832 20294 12872
rect 20294 12832 20334 12872
rect 20334 12832 20359 12872
rect 20105 12809 20191 12832
rect 20273 12809 20359 12832
rect 3745 12116 3831 12139
rect 3913 12116 3999 12139
rect 3745 12076 3770 12116
rect 3770 12076 3810 12116
rect 3810 12076 3831 12116
rect 3913 12076 3934 12116
rect 3934 12076 3974 12116
rect 3974 12076 3999 12116
rect 3745 12053 3831 12076
rect 3913 12053 3999 12076
rect 18865 12116 18951 12139
rect 19033 12116 19119 12139
rect 18865 12076 18890 12116
rect 18890 12076 18930 12116
rect 18930 12076 18951 12116
rect 19033 12076 19054 12116
rect 19054 12076 19094 12116
rect 19094 12076 19119 12116
rect 18865 12053 18951 12076
rect 19033 12053 19119 12076
rect 4985 11360 5071 11383
rect 5153 11360 5239 11383
rect 4985 11320 5010 11360
rect 5010 11320 5050 11360
rect 5050 11320 5071 11360
rect 5153 11320 5174 11360
rect 5174 11320 5214 11360
rect 5214 11320 5239 11360
rect 4985 11297 5071 11320
rect 5153 11297 5239 11320
rect 20105 11360 20191 11383
rect 20273 11360 20359 11383
rect 20105 11320 20130 11360
rect 20130 11320 20170 11360
rect 20170 11320 20191 11360
rect 20273 11320 20294 11360
rect 20294 11320 20334 11360
rect 20334 11320 20359 11360
rect 20105 11297 20191 11320
rect 20273 11297 20359 11320
rect 3745 10604 3831 10627
rect 3913 10604 3999 10627
rect 3745 10564 3770 10604
rect 3770 10564 3810 10604
rect 3810 10564 3831 10604
rect 3913 10564 3934 10604
rect 3934 10564 3974 10604
rect 3974 10564 3999 10604
rect 3745 10541 3831 10564
rect 3913 10541 3999 10564
rect 18865 10604 18951 10627
rect 19033 10604 19119 10627
rect 18865 10564 18890 10604
rect 18890 10564 18930 10604
rect 18930 10564 18951 10604
rect 19033 10564 19054 10604
rect 19054 10564 19094 10604
rect 19094 10564 19119 10604
rect 18865 10541 18951 10564
rect 19033 10541 19119 10564
rect 4985 9848 5071 9871
rect 5153 9848 5239 9871
rect 4985 9808 5010 9848
rect 5010 9808 5050 9848
rect 5050 9808 5071 9848
rect 5153 9808 5174 9848
rect 5174 9808 5214 9848
rect 5214 9808 5239 9848
rect 4985 9785 5071 9808
rect 5153 9785 5239 9808
rect 20105 9848 20191 9871
rect 20273 9848 20359 9871
rect 20105 9808 20130 9848
rect 20130 9808 20170 9848
rect 20170 9808 20191 9848
rect 20273 9808 20294 9848
rect 20294 9808 20334 9848
rect 20334 9808 20359 9848
rect 20105 9785 20191 9808
rect 20273 9785 20359 9808
rect 3745 9092 3831 9115
rect 3913 9092 3999 9115
rect 3745 9052 3770 9092
rect 3770 9052 3810 9092
rect 3810 9052 3831 9092
rect 3913 9052 3934 9092
rect 3934 9052 3974 9092
rect 3974 9052 3999 9092
rect 3745 9029 3831 9052
rect 3913 9029 3999 9052
rect 18865 9092 18951 9115
rect 19033 9092 19119 9115
rect 18865 9052 18890 9092
rect 18890 9052 18930 9092
rect 18930 9052 18951 9092
rect 19033 9052 19054 9092
rect 19054 9052 19094 9092
rect 19094 9052 19119 9092
rect 18865 9029 18951 9052
rect 19033 9029 19119 9052
rect 4985 8336 5071 8359
rect 5153 8336 5239 8359
rect 4985 8296 5010 8336
rect 5010 8296 5050 8336
rect 5050 8296 5071 8336
rect 5153 8296 5174 8336
rect 5174 8296 5214 8336
rect 5214 8296 5239 8336
rect 4985 8273 5071 8296
rect 5153 8273 5239 8296
rect 20105 8336 20191 8359
rect 20273 8336 20359 8359
rect 20105 8296 20130 8336
rect 20130 8296 20170 8336
rect 20170 8296 20191 8336
rect 20273 8296 20294 8336
rect 20294 8296 20334 8336
rect 20334 8296 20359 8336
rect 20105 8273 20191 8296
rect 20273 8273 20359 8296
rect 3745 7580 3831 7603
rect 3913 7580 3999 7603
rect 3745 7540 3770 7580
rect 3770 7540 3810 7580
rect 3810 7540 3831 7580
rect 3913 7540 3934 7580
rect 3934 7540 3974 7580
rect 3974 7540 3999 7580
rect 3745 7517 3831 7540
rect 3913 7517 3999 7540
rect 18865 7580 18951 7603
rect 19033 7580 19119 7603
rect 18865 7540 18890 7580
rect 18890 7540 18930 7580
rect 18930 7540 18951 7580
rect 19033 7540 19054 7580
rect 19054 7540 19094 7580
rect 19094 7540 19119 7580
rect 18865 7517 18951 7540
rect 19033 7517 19119 7540
rect 4985 6824 5071 6847
rect 5153 6824 5239 6847
rect 4985 6784 5010 6824
rect 5010 6784 5050 6824
rect 5050 6784 5071 6824
rect 5153 6784 5174 6824
rect 5174 6784 5214 6824
rect 5214 6784 5239 6824
rect 4985 6761 5071 6784
rect 5153 6761 5239 6784
rect 20105 6824 20191 6847
rect 20273 6824 20359 6847
rect 20105 6784 20130 6824
rect 20130 6784 20170 6824
rect 20170 6784 20191 6824
rect 20273 6784 20294 6824
rect 20294 6784 20334 6824
rect 20334 6784 20359 6824
rect 20105 6761 20191 6784
rect 20273 6761 20359 6784
rect 17157 6257 17243 6343
rect 3745 6068 3831 6091
rect 3913 6068 3999 6091
rect 3745 6028 3770 6068
rect 3770 6028 3810 6068
rect 3810 6028 3831 6068
rect 3913 6028 3934 6068
rect 3934 6028 3974 6068
rect 3974 6028 3999 6068
rect 3745 6005 3831 6028
rect 3913 6005 3999 6028
rect 18865 6068 18951 6091
rect 19033 6068 19119 6091
rect 18865 6028 18890 6068
rect 18890 6028 18930 6068
rect 18930 6028 18951 6068
rect 19033 6028 19054 6068
rect 19054 6028 19094 6068
rect 19094 6028 19119 6068
rect 18865 6005 18951 6028
rect 19033 6005 19119 6028
rect 4985 5312 5071 5335
rect 5153 5312 5239 5335
rect 4985 5272 5010 5312
rect 5010 5272 5050 5312
rect 5050 5272 5071 5312
rect 5153 5272 5174 5312
rect 5174 5272 5214 5312
rect 5214 5272 5239 5312
rect 4985 5249 5071 5272
rect 5153 5249 5239 5272
rect 20105 5312 20191 5335
rect 20273 5312 20359 5335
rect 20105 5272 20130 5312
rect 20130 5272 20170 5312
rect 20170 5272 20191 5312
rect 20273 5272 20294 5312
rect 20294 5272 20334 5312
rect 20334 5272 20359 5312
rect 20105 5249 20191 5272
rect 20273 5249 20359 5272
rect 3745 4556 3831 4579
rect 3913 4556 3999 4579
rect 3745 4516 3770 4556
rect 3770 4516 3810 4556
rect 3810 4516 3831 4556
rect 3913 4516 3934 4556
rect 3934 4516 3974 4556
rect 3974 4516 3999 4556
rect 3745 4493 3831 4516
rect 3913 4493 3999 4516
rect 18865 4556 18951 4579
rect 19033 4556 19119 4579
rect 18865 4516 18890 4556
rect 18890 4516 18930 4556
rect 18930 4516 18951 4556
rect 19033 4516 19054 4556
rect 19054 4516 19094 4556
rect 19094 4516 19119 4556
rect 18865 4493 18951 4516
rect 19033 4493 19119 4516
rect 4985 3800 5071 3823
rect 5153 3800 5239 3823
rect 4985 3760 5010 3800
rect 5010 3760 5050 3800
rect 5050 3760 5071 3800
rect 5153 3760 5174 3800
rect 5174 3760 5214 3800
rect 5214 3760 5239 3800
rect 4985 3737 5071 3760
rect 5153 3737 5239 3760
rect 20105 3800 20191 3823
rect 20273 3800 20359 3823
rect 20105 3760 20130 3800
rect 20130 3760 20170 3800
rect 20170 3760 20191 3800
rect 20273 3760 20294 3800
rect 20294 3760 20334 3800
rect 20334 3760 20359 3800
rect 20105 3737 20191 3760
rect 20273 3737 20359 3760
rect 11229 3401 11315 3487
rect 3745 3044 3831 3067
rect 3913 3044 3999 3067
rect 3745 3004 3770 3044
rect 3770 3004 3810 3044
rect 3810 3004 3831 3044
rect 3913 3004 3934 3044
rect 3934 3004 3974 3044
rect 3974 3004 3999 3044
rect 3745 2981 3831 3004
rect 3913 2981 3999 3004
rect 18865 3044 18951 3067
rect 19033 3044 19119 3067
rect 18865 3004 18890 3044
rect 18890 3004 18930 3044
rect 18930 3004 18951 3044
rect 19033 3004 19054 3044
rect 19054 3004 19094 3044
rect 19094 3004 19119 3044
rect 18865 2981 18951 3004
rect 19033 2981 19119 3004
rect 4985 2288 5071 2311
rect 5153 2288 5239 2311
rect 4985 2248 5010 2288
rect 5010 2248 5050 2288
rect 5050 2248 5071 2288
rect 5153 2248 5174 2288
rect 5174 2248 5214 2288
rect 5214 2248 5239 2288
rect 4985 2225 5071 2248
rect 5153 2225 5239 2248
rect 20105 2288 20191 2311
rect 20273 2288 20359 2311
rect 20105 2248 20130 2288
rect 20130 2248 20170 2288
rect 20170 2248 20191 2288
rect 20273 2248 20294 2288
rect 20294 2248 20334 2288
rect 20334 2248 20359 2288
rect 20105 2225 20191 2248
rect 20273 2225 20359 2248
rect 3745 1532 3831 1555
rect 3913 1532 3999 1555
rect 3745 1492 3770 1532
rect 3770 1492 3810 1532
rect 3810 1492 3831 1532
rect 3913 1492 3934 1532
rect 3934 1492 3974 1532
rect 3974 1492 3999 1532
rect 3745 1469 3831 1492
rect 3913 1469 3999 1492
rect 18865 1532 18951 1555
rect 19033 1532 19119 1555
rect 18865 1492 18890 1532
rect 18890 1492 18930 1532
rect 18930 1492 18951 1532
rect 19033 1492 19054 1532
rect 19054 1492 19094 1532
rect 19094 1492 19119 1532
rect 18865 1469 18951 1492
rect 19033 1469 19119 1492
rect 1197 1217 1283 1303
rect 13509 1049 13595 1135
rect 4985 776 5071 799
rect 5153 776 5239 799
rect 4985 736 5010 776
rect 5010 736 5050 776
rect 5050 736 5071 776
rect 5153 736 5174 776
rect 5174 736 5214 776
rect 5214 736 5239 776
rect 4985 713 5071 736
rect 5153 713 5239 736
rect 20105 776 20191 799
rect 20273 776 20359 799
rect 20105 736 20130 776
rect 20130 736 20170 776
rect 20170 736 20191 776
rect 20273 736 20294 776
rect 20294 736 20334 776
rect 20334 736 20359 776
rect 20105 713 20191 736
rect 20273 713 20359 736
rect 12141 209 12227 295
<< metal6 >>
rect 3652 84715 4092 86016
rect 3652 84629 3745 84715
rect 3831 84629 3913 84715
rect 3999 84629 4092 84715
rect 3652 83203 4092 84629
rect 3652 83117 3745 83203
rect 3831 83117 3913 83203
rect 3999 83117 4092 83203
rect 3652 81691 4092 83117
rect 3652 81605 3745 81691
rect 3831 81605 3913 81691
rect 3999 81605 4092 81691
rect 3652 80179 4092 81605
rect 3652 80093 3745 80179
rect 3831 80093 3913 80179
rect 3999 80093 4092 80179
rect 3652 78667 4092 80093
rect 3652 78581 3745 78667
rect 3831 78581 3913 78667
rect 3999 78581 4092 78667
rect 3652 77155 4092 78581
rect 3652 77069 3745 77155
rect 3831 77069 3913 77155
rect 3999 77069 4092 77155
rect 3652 75643 4092 77069
rect 3652 75557 3745 75643
rect 3831 75557 3913 75643
rect 3999 75557 4092 75643
rect 3652 74131 4092 75557
rect 3652 74045 3745 74131
rect 3831 74045 3913 74131
rect 3999 74045 4092 74131
rect 3652 72619 4092 74045
rect 3652 72533 3745 72619
rect 3831 72533 3913 72619
rect 3999 72533 4092 72619
rect 3652 71107 4092 72533
rect 3652 71021 3745 71107
rect 3831 71021 3913 71107
rect 3999 71021 4092 71107
rect 3652 69595 4092 71021
rect 3652 69509 3745 69595
rect 3831 69509 3913 69595
rect 3999 69509 4092 69595
rect 3652 68083 4092 69509
rect 3652 67997 3745 68083
rect 3831 67997 3913 68083
rect 3999 67997 4092 68083
rect 3652 66571 4092 67997
rect 3652 66485 3745 66571
rect 3831 66485 3913 66571
rect 3999 66485 4092 66571
rect 3652 65059 4092 66485
rect 3652 64973 3745 65059
rect 3831 64973 3913 65059
rect 3999 64973 4092 65059
rect 1076 64471 1404 64592
rect 1076 64385 1197 64471
rect 1283 64385 1404 64471
rect 1076 1303 1404 64385
rect 1076 1217 1197 1303
rect 1283 1217 1404 1303
rect 1076 1096 1404 1217
rect 3652 63547 4092 64973
rect 3652 63461 3745 63547
rect 3831 63461 3913 63547
rect 3999 63461 4092 63547
rect 3652 62035 4092 63461
rect 3652 61949 3745 62035
rect 3831 61949 3913 62035
rect 3999 61949 4092 62035
rect 3652 60523 4092 61949
rect 3652 60437 3745 60523
rect 3831 60437 3913 60523
rect 3999 60437 4092 60523
rect 3652 59011 4092 60437
rect 3652 58925 3745 59011
rect 3831 58925 3913 59011
rect 3999 58925 4092 59011
rect 3652 57499 4092 58925
rect 3652 57413 3745 57499
rect 3831 57413 3913 57499
rect 3999 57413 4092 57499
rect 3652 55987 4092 57413
rect 3652 55901 3745 55987
rect 3831 55901 3913 55987
rect 3999 55901 4092 55987
rect 3652 54475 4092 55901
rect 3652 54389 3745 54475
rect 3831 54389 3913 54475
rect 3999 54389 4092 54475
rect 3652 52963 4092 54389
rect 3652 52877 3745 52963
rect 3831 52877 3913 52963
rect 3999 52877 4092 52963
rect 3652 51451 4092 52877
rect 3652 51365 3745 51451
rect 3831 51365 3913 51451
rect 3999 51365 4092 51451
rect 3652 49939 4092 51365
rect 3652 49853 3745 49939
rect 3831 49853 3913 49939
rect 3999 49853 4092 49939
rect 3652 48427 4092 49853
rect 3652 48341 3745 48427
rect 3831 48341 3913 48427
rect 3999 48341 4092 48427
rect 3652 46915 4092 48341
rect 3652 46829 3745 46915
rect 3831 46829 3913 46915
rect 3999 46829 4092 46915
rect 3652 45403 4092 46829
rect 3652 45317 3745 45403
rect 3831 45317 3913 45403
rect 3999 45317 4092 45403
rect 3652 43891 4092 45317
rect 3652 43805 3745 43891
rect 3831 43805 3913 43891
rect 3999 43805 4092 43891
rect 3652 42379 4092 43805
rect 3652 42293 3745 42379
rect 3831 42293 3913 42379
rect 3999 42293 4092 42379
rect 3652 40867 4092 42293
rect 3652 40781 3745 40867
rect 3831 40781 3913 40867
rect 3999 40781 4092 40867
rect 3652 39355 4092 40781
rect 3652 39269 3745 39355
rect 3831 39269 3913 39355
rect 3999 39269 4092 39355
rect 3652 37843 4092 39269
rect 3652 37757 3745 37843
rect 3831 37757 3913 37843
rect 3999 37757 4092 37843
rect 3652 36331 4092 37757
rect 3652 36245 3745 36331
rect 3831 36245 3913 36331
rect 3999 36245 4092 36331
rect 3652 34819 4092 36245
rect 3652 34733 3745 34819
rect 3831 34733 3913 34819
rect 3999 34733 4092 34819
rect 3652 33307 4092 34733
rect 3652 33221 3745 33307
rect 3831 33221 3913 33307
rect 3999 33221 4092 33307
rect 3652 31795 4092 33221
rect 3652 31709 3745 31795
rect 3831 31709 3913 31795
rect 3999 31709 4092 31795
rect 3652 30283 4092 31709
rect 3652 30197 3745 30283
rect 3831 30197 3913 30283
rect 3999 30197 4092 30283
rect 3652 28771 4092 30197
rect 3652 28685 3745 28771
rect 3831 28685 3913 28771
rect 3999 28685 4092 28771
rect 3652 27259 4092 28685
rect 3652 27173 3745 27259
rect 3831 27173 3913 27259
rect 3999 27173 4092 27259
rect 3652 25747 4092 27173
rect 3652 25661 3745 25747
rect 3831 25661 3913 25747
rect 3999 25661 4092 25747
rect 3652 24235 4092 25661
rect 3652 24149 3745 24235
rect 3831 24149 3913 24235
rect 3999 24149 4092 24235
rect 3652 22723 4092 24149
rect 3652 22637 3745 22723
rect 3831 22637 3913 22723
rect 3999 22637 4092 22723
rect 3652 21211 4092 22637
rect 3652 21125 3745 21211
rect 3831 21125 3913 21211
rect 3999 21125 4092 21211
rect 3652 19699 4092 21125
rect 3652 19613 3745 19699
rect 3831 19613 3913 19699
rect 3999 19613 4092 19699
rect 3652 18187 4092 19613
rect 3652 18101 3745 18187
rect 3831 18101 3913 18187
rect 3999 18101 4092 18187
rect 3652 16675 4092 18101
rect 3652 16589 3745 16675
rect 3831 16589 3913 16675
rect 3999 16589 4092 16675
rect 3652 15163 4092 16589
rect 3652 15077 3745 15163
rect 3831 15077 3913 15163
rect 3999 15077 4092 15163
rect 3652 13651 4092 15077
rect 3652 13565 3745 13651
rect 3831 13565 3913 13651
rect 3999 13565 4092 13651
rect 3652 12139 4092 13565
rect 3652 12053 3745 12139
rect 3831 12053 3913 12139
rect 3999 12053 4092 12139
rect 3652 10627 4092 12053
rect 3652 10541 3745 10627
rect 3831 10541 3913 10627
rect 3999 10541 4092 10627
rect 3652 9115 4092 10541
rect 3652 9029 3745 9115
rect 3831 9029 3913 9115
rect 3999 9029 4092 9115
rect 3652 7603 4092 9029
rect 3652 7517 3745 7603
rect 3831 7517 3913 7603
rect 3999 7517 4092 7603
rect 3652 6091 4092 7517
rect 3652 6005 3745 6091
rect 3831 6005 3913 6091
rect 3999 6005 4092 6091
rect 3652 4579 4092 6005
rect 3652 4493 3745 4579
rect 3831 4493 3913 4579
rect 3999 4493 4092 4579
rect 3652 3067 4092 4493
rect 3652 2981 3745 3067
rect 3831 2981 3913 3067
rect 3999 2981 4092 3067
rect 3652 1555 4092 2981
rect 3652 1469 3745 1555
rect 3831 1469 3913 1555
rect 3999 1469 4092 1555
rect 3652 0 4092 1469
rect 4892 83959 5332 86016
rect 4892 83873 4985 83959
rect 5071 83873 5153 83959
rect 5239 83873 5332 83959
rect 4892 82447 5332 83873
rect 18772 84715 19212 86016
rect 18772 84629 18865 84715
rect 18951 84629 19033 84715
rect 19119 84629 19212 84715
rect 4892 82361 4985 82447
rect 5071 82361 5153 82447
rect 5239 82361 5332 82447
rect 4892 80935 5332 82361
rect 4892 80849 4985 80935
rect 5071 80849 5153 80935
rect 5239 80849 5332 80935
rect 4892 79423 5332 80849
rect 4892 79337 4985 79423
rect 5071 79337 5153 79423
rect 5239 79337 5332 79423
rect 4892 77911 5332 79337
rect 4892 77825 4985 77911
rect 5071 77825 5153 77911
rect 5239 77825 5332 77911
rect 4892 76399 5332 77825
rect 4892 76313 4985 76399
rect 5071 76313 5153 76399
rect 5239 76313 5332 76399
rect 4892 74887 5332 76313
rect 4892 74801 4985 74887
rect 5071 74801 5153 74887
rect 5239 74801 5332 74887
rect 4892 73375 5332 74801
rect 4892 73289 4985 73375
rect 5071 73289 5153 73375
rect 5239 73289 5332 73375
rect 4892 71863 5332 73289
rect 4892 71777 4985 71863
rect 5071 71777 5153 71863
rect 5239 71777 5332 71863
rect 4892 70351 5332 71777
rect 4892 70265 4985 70351
rect 5071 70265 5153 70351
rect 5239 70265 5332 70351
rect 4892 68839 5332 70265
rect 4892 68753 4985 68839
rect 5071 68753 5153 68839
rect 5239 68753 5332 68839
rect 4892 67327 5332 68753
rect 4892 67241 4985 67327
rect 5071 67241 5153 67327
rect 5239 67241 5332 67327
rect 4892 65815 5332 67241
rect 4892 65729 4985 65815
rect 5071 65729 5153 65815
rect 5239 65729 5332 65815
rect 4892 64303 5332 65729
rect 4892 64217 4985 64303
rect 5071 64217 5153 64303
rect 5239 64217 5332 64303
rect 4892 62791 5332 64217
rect 4892 62705 4985 62791
rect 5071 62705 5153 62791
rect 5239 62705 5332 62791
rect 4892 61279 5332 62705
rect 4892 61193 4985 61279
rect 5071 61193 5153 61279
rect 5239 61193 5332 61279
rect 4892 59767 5332 61193
rect 4892 59681 4985 59767
rect 5071 59681 5153 59767
rect 5239 59681 5332 59767
rect 4892 58255 5332 59681
rect 4892 58169 4985 58255
rect 5071 58169 5153 58255
rect 5239 58169 5332 58255
rect 4892 56743 5332 58169
rect 4892 56657 4985 56743
rect 5071 56657 5153 56743
rect 5239 56657 5332 56743
rect 4892 55231 5332 56657
rect 4892 55145 4985 55231
rect 5071 55145 5153 55231
rect 5239 55145 5332 55231
rect 4892 53719 5332 55145
rect 4892 53633 4985 53719
rect 5071 53633 5153 53719
rect 5239 53633 5332 53719
rect 4892 52207 5332 53633
rect 4892 52121 4985 52207
rect 5071 52121 5153 52207
rect 5239 52121 5332 52207
rect 4892 50695 5332 52121
rect 4892 50609 4985 50695
rect 5071 50609 5153 50695
rect 5239 50609 5332 50695
rect 4892 49183 5332 50609
rect 4892 49097 4985 49183
rect 5071 49097 5153 49183
rect 5239 49097 5332 49183
rect 4892 47671 5332 49097
rect 4892 47585 4985 47671
rect 5071 47585 5153 47671
rect 5239 47585 5332 47671
rect 4892 46159 5332 47585
rect 4892 46073 4985 46159
rect 5071 46073 5153 46159
rect 5239 46073 5332 46159
rect 4892 44647 5332 46073
rect 4892 44561 4985 44647
rect 5071 44561 5153 44647
rect 5239 44561 5332 44647
rect 4892 43135 5332 44561
rect 4892 43049 4985 43135
rect 5071 43049 5153 43135
rect 5239 43049 5332 43135
rect 4892 41623 5332 43049
rect 4892 41537 4985 41623
rect 5071 41537 5153 41623
rect 5239 41537 5332 41623
rect 4892 40111 5332 41537
rect 4892 40025 4985 40111
rect 5071 40025 5153 40111
rect 5239 40025 5332 40111
rect 4892 38599 5332 40025
rect 4892 38513 4985 38599
rect 5071 38513 5153 38599
rect 5239 38513 5332 38599
rect 4892 37087 5332 38513
rect 4892 37001 4985 37087
rect 5071 37001 5153 37087
rect 5239 37001 5332 37087
rect 4892 35575 5332 37001
rect 4892 35489 4985 35575
rect 5071 35489 5153 35575
rect 5239 35489 5332 35575
rect 4892 34063 5332 35489
rect 4892 33977 4985 34063
rect 5071 33977 5153 34063
rect 5239 33977 5332 34063
rect 4892 32551 5332 33977
rect 4892 32465 4985 32551
rect 5071 32465 5153 32551
rect 5239 32465 5332 32551
rect 4892 31039 5332 32465
rect 4892 30953 4985 31039
rect 5071 30953 5153 31039
rect 5239 30953 5332 31039
rect 4892 29527 5332 30953
rect 4892 29441 4985 29527
rect 5071 29441 5153 29527
rect 5239 29441 5332 29527
rect 4892 28015 5332 29441
rect 4892 27929 4985 28015
rect 5071 27929 5153 28015
rect 5239 27929 5332 28015
rect 4892 26503 5332 27929
rect 4892 26417 4985 26503
rect 5071 26417 5153 26503
rect 5239 26417 5332 26503
rect 4892 24991 5332 26417
rect 7916 83539 8244 83660
rect 7916 83453 8037 83539
rect 8123 83453 8244 83539
rect 17036 83539 17364 83660
rect 7916 26335 8244 83453
rect 13388 83371 13716 83492
rect 13388 83285 13509 83371
rect 13595 83285 13716 83371
rect 12020 72199 12348 72320
rect 12020 72113 12141 72199
rect 12227 72113 12348 72199
rect 11108 69343 11436 69464
rect 11108 69257 11229 69343
rect 11315 69257 11436 69343
rect 7916 26249 8037 26335
rect 8123 26249 8244 26335
rect 9740 63043 10068 63164
rect 9740 62957 9861 63043
rect 9947 62957 10068 63043
rect 9740 26503 10068 62957
rect 9740 26417 9861 26503
rect 9947 26417 10068 26503
rect 9740 26296 10068 26417
rect 7916 26128 8244 26249
rect 4892 24905 4985 24991
rect 5071 24905 5153 24991
rect 5239 24905 5332 24991
rect 4892 23479 5332 24905
rect 4892 23393 4985 23479
rect 5071 23393 5153 23479
rect 5239 23393 5332 23479
rect 4892 21967 5332 23393
rect 4892 21881 4985 21967
rect 5071 21881 5153 21967
rect 5239 21881 5332 21967
rect 4892 20455 5332 21881
rect 4892 20369 4985 20455
rect 5071 20369 5153 20455
rect 5239 20369 5332 20455
rect 4892 18943 5332 20369
rect 4892 18857 4985 18943
rect 5071 18857 5153 18943
rect 5239 18857 5332 18943
rect 4892 17431 5332 18857
rect 4892 17345 4985 17431
rect 5071 17345 5153 17431
rect 5239 17345 5332 17431
rect 4892 15919 5332 17345
rect 4892 15833 4985 15919
rect 5071 15833 5153 15919
rect 5239 15833 5332 15919
rect 4892 14407 5332 15833
rect 4892 14321 4985 14407
rect 5071 14321 5153 14407
rect 5239 14321 5332 14407
rect 4892 12895 5332 14321
rect 4892 12809 4985 12895
rect 5071 12809 5153 12895
rect 5239 12809 5332 12895
rect 4892 11383 5332 12809
rect 4892 11297 4985 11383
rect 5071 11297 5153 11383
rect 5239 11297 5332 11383
rect 4892 9871 5332 11297
rect 4892 9785 4985 9871
rect 5071 9785 5153 9871
rect 5239 9785 5332 9871
rect 4892 8359 5332 9785
rect 4892 8273 4985 8359
rect 5071 8273 5153 8359
rect 5239 8273 5332 8359
rect 4892 6847 5332 8273
rect 4892 6761 4985 6847
rect 5071 6761 5153 6847
rect 5239 6761 5332 6847
rect 4892 5335 5332 6761
rect 4892 5249 4985 5335
rect 5071 5249 5153 5335
rect 5239 5249 5332 5335
rect 4892 3823 5332 5249
rect 4892 3737 4985 3823
rect 5071 3737 5153 3823
rect 5239 3737 5332 3823
rect 4892 2311 5332 3737
rect 11108 3487 11436 69257
rect 11108 3401 11229 3487
rect 11315 3401 11436 3487
rect 11108 3280 11436 3401
rect 12020 30703 12348 72113
rect 12020 30617 12141 30703
rect 12227 30617 12348 30703
rect 4892 2225 4985 2311
rect 5071 2225 5153 2311
rect 5239 2225 5332 2311
rect 4892 799 5332 2225
rect 4892 713 4985 799
rect 5071 713 5153 799
rect 5239 713 5332 799
rect 4892 0 5332 713
rect 12020 295 12348 30617
rect 13388 1135 13716 83285
rect 17036 83453 17157 83539
rect 17243 83453 17364 83539
rect 15212 72787 15540 72908
rect 15212 72701 15333 72787
rect 15419 72701 15540 72787
rect 15212 17683 15540 72701
rect 15212 17597 15333 17683
rect 15419 17597 15540 17683
rect 15212 17476 15540 17597
rect 17036 6343 17364 83453
rect 17036 6257 17157 6343
rect 17243 6257 17364 6343
rect 17036 6136 17364 6257
rect 18772 83203 19212 84629
rect 18772 83117 18865 83203
rect 18951 83117 19033 83203
rect 19119 83117 19212 83203
rect 18772 81691 19212 83117
rect 18772 81605 18865 81691
rect 18951 81605 19033 81691
rect 19119 81605 19212 81691
rect 18772 80179 19212 81605
rect 18772 80093 18865 80179
rect 18951 80093 19033 80179
rect 19119 80093 19212 80179
rect 18772 78667 19212 80093
rect 18772 78581 18865 78667
rect 18951 78581 19033 78667
rect 19119 78581 19212 78667
rect 18772 77155 19212 78581
rect 18772 77069 18865 77155
rect 18951 77069 19033 77155
rect 19119 77069 19212 77155
rect 18772 75643 19212 77069
rect 18772 75557 18865 75643
rect 18951 75557 19033 75643
rect 19119 75557 19212 75643
rect 18772 74131 19212 75557
rect 18772 74045 18865 74131
rect 18951 74045 19033 74131
rect 19119 74045 19212 74131
rect 18772 72619 19212 74045
rect 18772 72533 18865 72619
rect 18951 72533 19033 72619
rect 19119 72533 19212 72619
rect 18772 71107 19212 72533
rect 18772 71021 18865 71107
rect 18951 71021 19033 71107
rect 19119 71021 19212 71107
rect 18772 69595 19212 71021
rect 18772 69509 18865 69595
rect 18951 69509 19033 69595
rect 19119 69509 19212 69595
rect 18772 68083 19212 69509
rect 18772 67997 18865 68083
rect 18951 67997 19033 68083
rect 19119 67997 19212 68083
rect 18772 66571 19212 67997
rect 18772 66485 18865 66571
rect 18951 66485 19033 66571
rect 19119 66485 19212 66571
rect 18772 65059 19212 66485
rect 18772 64973 18865 65059
rect 18951 64973 19033 65059
rect 19119 64973 19212 65059
rect 18772 63547 19212 64973
rect 18772 63461 18865 63547
rect 18951 63461 19033 63547
rect 19119 63461 19212 63547
rect 18772 62035 19212 63461
rect 18772 61949 18865 62035
rect 18951 61949 19033 62035
rect 19119 61949 19212 62035
rect 18772 60523 19212 61949
rect 18772 60437 18865 60523
rect 18951 60437 19033 60523
rect 19119 60437 19212 60523
rect 18772 59011 19212 60437
rect 18772 58925 18865 59011
rect 18951 58925 19033 59011
rect 19119 58925 19212 59011
rect 18772 57499 19212 58925
rect 18772 57413 18865 57499
rect 18951 57413 19033 57499
rect 19119 57413 19212 57499
rect 18772 55987 19212 57413
rect 18772 55901 18865 55987
rect 18951 55901 19033 55987
rect 19119 55901 19212 55987
rect 18772 54475 19212 55901
rect 18772 54389 18865 54475
rect 18951 54389 19033 54475
rect 19119 54389 19212 54475
rect 18772 52963 19212 54389
rect 18772 52877 18865 52963
rect 18951 52877 19033 52963
rect 19119 52877 19212 52963
rect 18772 51451 19212 52877
rect 18772 51365 18865 51451
rect 18951 51365 19033 51451
rect 19119 51365 19212 51451
rect 18772 49939 19212 51365
rect 18772 49853 18865 49939
rect 18951 49853 19033 49939
rect 19119 49853 19212 49939
rect 18772 48427 19212 49853
rect 18772 48341 18865 48427
rect 18951 48341 19033 48427
rect 19119 48341 19212 48427
rect 18772 46915 19212 48341
rect 18772 46829 18865 46915
rect 18951 46829 19033 46915
rect 19119 46829 19212 46915
rect 18772 45403 19212 46829
rect 18772 45317 18865 45403
rect 18951 45317 19033 45403
rect 19119 45317 19212 45403
rect 18772 43891 19212 45317
rect 18772 43805 18865 43891
rect 18951 43805 19033 43891
rect 19119 43805 19212 43891
rect 18772 42379 19212 43805
rect 18772 42293 18865 42379
rect 18951 42293 19033 42379
rect 19119 42293 19212 42379
rect 18772 40867 19212 42293
rect 18772 40781 18865 40867
rect 18951 40781 19033 40867
rect 19119 40781 19212 40867
rect 18772 39355 19212 40781
rect 18772 39269 18865 39355
rect 18951 39269 19033 39355
rect 19119 39269 19212 39355
rect 18772 37843 19212 39269
rect 18772 37757 18865 37843
rect 18951 37757 19033 37843
rect 19119 37757 19212 37843
rect 18772 36331 19212 37757
rect 18772 36245 18865 36331
rect 18951 36245 19033 36331
rect 19119 36245 19212 36331
rect 18772 34819 19212 36245
rect 18772 34733 18865 34819
rect 18951 34733 19033 34819
rect 19119 34733 19212 34819
rect 18772 33307 19212 34733
rect 18772 33221 18865 33307
rect 18951 33221 19033 33307
rect 19119 33221 19212 33307
rect 18772 31795 19212 33221
rect 18772 31709 18865 31795
rect 18951 31709 19033 31795
rect 19119 31709 19212 31795
rect 18772 30283 19212 31709
rect 18772 30197 18865 30283
rect 18951 30197 19033 30283
rect 19119 30197 19212 30283
rect 18772 28771 19212 30197
rect 18772 28685 18865 28771
rect 18951 28685 19033 28771
rect 19119 28685 19212 28771
rect 18772 27259 19212 28685
rect 18772 27173 18865 27259
rect 18951 27173 19033 27259
rect 19119 27173 19212 27259
rect 18772 25747 19212 27173
rect 18772 25661 18865 25747
rect 18951 25661 19033 25747
rect 19119 25661 19212 25747
rect 18772 24235 19212 25661
rect 18772 24149 18865 24235
rect 18951 24149 19033 24235
rect 19119 24149 19212 24235
rect 18772 22723 19212 24149
rect 18772 22637 18865 22723
rect 18951 22637 19033 22723
rect 19119 22637 19212 22723
rect 18772 21211 19212 22637
rect 18772 21125 18865 21211
rect 18951 21125 19033 21211
rect 19119 21125 19212 21211
rect 18772 19699 19212 21125
rect 18772 19613 18865 19699
rect 18951 19613 19033 19699
rect 19119 19613 19212 19699
rect 18772 18187 19212 19613
rect 18772 18101 18865 18187
rect 18951 18101 19033 18187
rect 19119 18101 19212 18187
rect 18772 16675 19212 18101
rect 18772 16589 18865 16675
rect 18951 16589 19033 16675
rect 19119 16589 19212 16675
rect 18772 15163 19212 16589
rect 18772 15077 18865 15163
rect 18951 15077 19033 15163
rect 19119 15077 19212 15163
rect 18772 13651 19212 15077
rect 18772 13565 18865 13651
rect 18951 13565 19033 13651
rect 19119 13565 19212 13651
rect 18772 12139 19212 13565
rect 18772 12053 18865 12139
rect 18951 12053 19033 12139
rect 19119 12053 19212 12139
rect 18772 10627 19212 12053
rect 18772 10541 18865 10627
rect 18951 10541 19033 10627
rect 19119 10541 19212 10627
rect 18772 9115 19212 10541
rect 18772 9029 18865 9115
rect 18951 9029 19033 9115
rect 19119 9029 19212 9115
rect 18772 7603 19212 9029
rect 18772 7517 18865 7603
rect 18951 7517 19033 7603
rect 19119 7517 19212 7603
rect 13388 1049 13509 1135
rect 13595 1049 13716 1135
rect 13388 928 13716 1049
rect 18772 6091 19212 7517
rect 18772 6005 18865 6091
rect 18951 6005 19033 6091
rect 19119 6005 19212 6091
rect 18772 4579 19212 6005
rect 18772 4493 18865 4579
rect 18951 4493 19033 4579
rect 19119 4493 19212 4579
rect 18772 3067 19212 4493
rect 18772 2981 18865 3067
rect 18951 2981 19033 3067
rect 19119 2981 19212 3067
rect 18772 1555 19212 2981
rect 18772 1469 18865 1555
rect 18951 1469 19033 1555
rect 19119 1469 19212 1555
rect 12020 209 12141 295
rect 12227 209 12348 295
rect 12020 88 12348 209
rect 18772 0 19212 1469
rect 20012 83959 20452 86016
rect 20012 83873 20105 83959
rect 20191 83873 20273 83959
rect 20359 83873 20452 83959
rect 20012 82447 20452 83873
rect 20012 82361 20105 82447
rect 20191 82361 20273 82447
rect 20359 82361 20452 82447
rect 20012 80935 20452 82361
rect 20012 80849 20105 80935
rect 20191 80849 20273 80935
rect 20359 80849 20452 80935
rect 20012 79423 20452 80849
rect 20012 79337 20105 79423
rect 20191 79337 20273 79423
rect 20359 79337 20452 79423
rect 20012 77911 20452 79337
rect 20012 77825 20105 77911
rect 20191 77825 20273 77911
rect 20359 77825 20452 77911
rect 20012 76399 20452 77825
rect 20012 76313 20105 76399
rect 20191 76313 20273 76399
rect 20359 76313 20452 76399
rect 20012 74887 20452 76313
rect 20012 74801 20105 74887
rect 20191 74801 20273 74887
rect 20359 74801 20452 74887
rect 20012 73375 20452 74801
rect 20012 73289 20105 73375
rect 20191 73289 20273 73375
rect 20359 73289 20452 73375
rect 20012 71863 20452 73289
rect 20012 71777 20105 71863
rect 20191 71777 20273 71863
rect 20359 71777 20452 71863
rect 20012 70351 20452 71777
rect 20012 70265 20105 70351
rect 20191 70265 20273 70351
rect 20359 70265 20452 70351
rect 20012 68839 20452 70265
rect 20012 68753 20105 68839
rect 20191 68753 20273 68839
rect 20359 68753 20452 68839
rect 20012 67327 20452 68753
rect 20012 67241 20105 67327
rect 20191 67241 20273 67327
rect 20359 67241 20452 67327
rect 20012 65815 20452 67241
rect 20012 65729 20105 65815
rect 20191 65729 20273 65815
rect 20359 65729 20452 65815
rect 20012 64303 20452 65729
rect 20012 64217 20105 64303
rect 20191 64217 20273 64303
rect 20359 64217 20452 64303
rect 20012 62791 20452 64217
rect 20012 62705 20105 62791
rect 20191 62705 20273 62791
rect 20359 62705 20452 62791
rect 20012 61279 20452 62705
rect 20012 61193 20105 61279
rect 20191 61193 20273 61279
rect 20359 61193 20452 61279
rect 20012 59767 20452 61193
rect 20012 59681 20105 59767
rect 20191 59681 20273 59767
rect 20359 59681 20452 59767
rect 20012 58255 20452 59681
rect 20012 58169 20105 58255
rect 20191 58169 20273 58255
rect 20359 58169 20452 58255
rect 20012 56743 20452 58169
rect 20012 56657 20105 56743
rect 20191 56657 20273 56743
rect 20359 56657 20452 56743
rect 20012 55231 20452 56657
rect 20012 55145 20105 55231
rect 20191 55145 20273 55231
rect 20359 55145 20452 55231
rect 20012 53719 20452 55145
rect 20012 53633 20105 53719
rect 20191 53633 20273 53719
rect 20359 53633 20452 53719
rect 20012 52207 20452 53633
rect 20012 52121 20105 52207
rect 20191 52121 20273 52207
rect 20359 52121 20452 52207
rect 20012 50695 20452 52121
rect 20012 50609 20105 50695
rect 20191 50609 20273 50695
rect 20359 50609 20452 50695
rect 20012 49183 20452 50609
rect 20012 49097 20105 49183
rect 20191 49097 20273 49183
rect 20359 49097 20452 49183
rect 20012 47671 20452 49097
rect 20012 47585 20105 47671
rect 20191 47585 20273 47671
rect 20359 47585 20452 47671
rect 20012 46159 20452 47585
rect 20012 46073 20105 46159
rect 20191 46073 20273 46159
rect 20359 46073 20452 46159
rect 20012 44647 20452 46073
rect 20012 44561 20105 44647
rect 20191 44561 20273 44647
rect 20359 44561 20452 44647
rect 20012 43135 20452 44561
rect 20012 43049 20105 43135
rect 20191 43049 20273 43135
rect 20359 43049 20452 43135
rect 20012 41623 20452 43049
rect 20012 41537 20105 41623
rect 20191 41537 20273 41623
rect 20359 41537 20452 41623
rect 20012 40111 20452 41537
rect 20012 40025 20105 40111
rect 20191 40025 20273 40111
rect 20359 40025 20452 40111
rect 20012 38599 20452 40025
rect 20012 38513 20105 38599
rect 20191 38513 20273 38599
rect 20359 38513 20452 38599
rect 20012 37087 20452 38513
rect 20012 37001 20105 37087
rect 20191 37001 20273 37087
rect 20359 37001 20452 37087
rect 20012 35575 20452 37001
rect 20012 35489 20105 35575
rect 20191 35489 20273 35575
rect 20359 35489 20452 35575
rect 20012 34063 20452 35489
rect 20012 33977 20105 34063
rect 20191 33977 20273 34063
rect 20359 33977 20452 34063
rect 20012 32551 20452 33977
rect 20012 32465 20105 32551
rect 20191 32465 20273 32551
rect 20359 32465 20452 32551
rect 20012 31039 20452 32465
rect 20012 30953 20105 31039
rect 20191 30953 20273 31039
rect 20359 30953 20452 31039
rect 20012 29527 20452 30953
rect 20012 29441 20105 29527
rect 20191 29441 20273 29527
rect 20359 29441 20452 29527
rect 20012 28015 20452 29441
rect 20012 27929 20105 28015
rect 20191 27929 20273 28015
rect 20359 27929 20452 28015
rect 20012 26503 20452 27929
rect 20012 26417 20105 26503
rect 20191 26417 20273 26503
rect 20359 26417 20452 26503
rect 20012 24991 20452 26417
rect 20012 24905 20105 24991
rect 20191 24905 20273 24991
rect 20359 24905 20452 24991
rect 20012 23479 20452 24905
rect 20012 23393 20105 23479
rect 20191 23393 20273 23479
rect 20359 23393 20452 23479
rect 20012 21967 20452 23393
rect 20012 21881 20105 21967
rect 20191 21881 20273 21967
rect 20359 21881 20452 21967
rect 20012 20455 20452 21881
rect 20012 20369 20105 20455
rect 20191 20369 20273 20455
rect 20359 20369 20452 20455
rect 20012 18943 20452 20369
rect 20012 18857 20105 18943
rect 20191 18857 20273 18943
rect 20359 18857 20452 18943
rect 20012 17431 20452 18857
rect 20012 17345 20105 17431
rect 20191 17345 20273 17431
rect 20359 17345 20452 17431
rect 20012 15919 20452 17345
rect 20012 15833 20105 15919
rect 20191 15833 20273 15919
rect 20359 15833 20452 15919
rect 20012 14407 20452 15833
rect 20012 14321 20105 14407
rect 20191 14321 20273 14407
rect 20359 14321 20452 14407
rect 20012 12895 20452 14321
rect 20012 12809 20105 12895
rect 20191 12809 20273 12895
rect 20359 12809 20452 12895
rect 20012 11383 20452 12809
rect 20012 11297 20105 11383
rect 20191 11297 20273 11383
rect 20359 11297 20452 11383
rect 20012 9871 20452 11297
rect 20012 9785 20105 9871
rect 20191 9785 20273 9871
rect 20359 9785 20452 9871
rect 20012 8359 20452 9785
rect 20012 8273 20105 8359
rect 20191 8273 20273 8359
rect 20359 8273 20452 8359
rect 20012 6847 20452 8273
rect 20012 6761 20105 6847
rect 20191 6761 20273 6847
rect 20359 6761 20452 6847
rect 20012 5335 20452 6761
rect 20012 5249 20105 5335
rect 20191 5249 20273 5335
rect 20359 5249 20452 5335
rect 20012 3823 20452 5249
rect 20012 3737 20105 3823
rect 20191 3737 20273 3823
rect 20359 3737 20452 3823
rect 20012 2311 20452 3737
rect 20012 2225 20105 2311
rect 20191 2225 20273 2311
rect 20359 2225 20452 2311
rect 20012 799 20452 2225
rect 20012 713 20105 799
rect 20191 713 20273 799
rect 20359 713 20452 799
rect 20012 0 20452 713
use sg13g2_inv_1  _0357_
timestamp 1676382929
transform 1 0 11808 0 1 59724
box -48 -56 336 834
use sg13g2_inv_1  _0358_
timestamp 1676382929
transform 1 0 17760 0 1 64260
box -48 -56 336 834
use sg13g2_inv_1  _0359_
timestamp 1676382929
transform 1 0 5376 0 -1 74844
box -48 -56 336 834
use sg13g2_inv_1  _0360_
timestamp 1676382929
transform 1 0 4992 0 -1 61236
box -48 -56 336 834
use sg13g2_inv_1  _0361_
timestamp 1676382929
transform 1 0 6528 0 -1 68796
box -48 -56 336 834
use sg13g2_inv_1  _0362_
timestamp 1676382929
transform 1 0 12672 0 1 65772
box -48 -56 336 834
use sg13g2_inv_1  _0363_
timestamp 1676382929
transform 1 0 15936 0 1 65772
box -48 -56 336 834
use sg13g2_inv_1  _0364_
timestamp 1676382929
transform -1 0 6912 0 1 71820
box -48 -56 336 834
use sg13g2_inv_1  _0365_
timestamp 1676382929
transform 1 0 14208 0 -1 37044
box -48 -56 336 834
use sg13g2_inv_1  _0366_
timestamp 1676382929
transform 1 0 12864 0 -1 37044
box -48 -56 336 834
use sg13g2_inv_1  _0367_
timestamp 1676382929
transform 1 0 7872 0 -1 38556
box -48 -56 336 834
use sg13g2_inv_1  _0368_
timestamp 1676382929
transform 1 0 15552 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  _0369_
timestamp 1676382929
transform 1 0 14304 0 -1 20412
box -48 -56 336 834
use sg13g2_inv_1  _0370_
timestamp 1676382929
transform 1 0 1536 0 -1 30996
box -48 -56 336 834
use sg13g2_inv_1  _0371_
timestamp 1676382929
transform -1 0 9120 0 -1 23436
box -48 -56 336 834
use sg13g2_inv_1  _0372_
timestamp 1676382929
transform 1 0 16896 0 1 21924
box -48 -56 336 834
use sg13g2_inv_1  _0373_
timestamp 1676382929
transform -1 0 18240 0 -1 29484
box -48 -56 336 834
use sg13g2_inv_1  _0374_
timestamp 1676382929
transform 1 0 9024 0 1 30996
box -48 -56 336 834
use sg13g2_inv_1  _0375_
timestamp 1676382929
transform -1 0 13920 0 1 32508
box -48 -56 336 834
use sg13g2_inv_1  _0376_
timestamp 1676382929
transform -1 0 13920 0 -1 32508
box -48 -56 336 834
use sg13g2_inv_1  _0377_
timestamp 1676382929
transform -1 0 14304 0 -1 38556
box -48 -56 336 834
use sg13g2_nand2b_1  _0378_
timestamp 1676567195
transform 1 0 13440 0 1 58212
box -48 -56 528 834
use sg13g2_nor3_1  _0379_
timestamp 1676639442
transform -1 0 13152 0 -1 61236
box -48 -56 528 834
use sg13g2_a221oi_1  _0380_
timestamp 1685197497
transform -1 0 13440 0 1 58212
box -48 -56 816 834
use sg13g2_mux4_1  _0381_
timestamp 1677257233
transform 1 0 12096 0 1 59724
box -48 -56 2064 834
use sg13g2_nand2b_1  _0382_
timestamp 1676567195
transform 1 0 15072 0 1 17388
box -48 -56 528 834
use sg13g2_nor3_1  _0383_
timestamp 1676639442
transform 1 0 14400 0 1 15876
box -48 -56 528 834
use sg13g2_a221oi_1  _0384_
timestamp 1685197497
transform 1 0 15360 0 -1 18900
box -48 -56 816 834
use sg13g2_mux4_1  _0385_
timestamp 1677257233
transform 1 0 13344 0 -1 21924
box -48 -56 2064 834
use sg13g2_mux4_1  _0386_
timestamp 1677257233
transform 1 0 13056 0 -1 49140
box -48 -56 2064 834
use sg13g2_mux4_1  _0387_
timestamp 1677257233
transform 1 0 11808 0 -1 62748
box -48 -56 2064 834
use sg13g2_nand2b_1  _0388_
timestamp 1676567195
transform -1 0 18432 0 -1 64260
box -48 -56 528 834
use sg13g2_nor3_1  _0389_
timestamp 1676639442
transform -1 0 18528 0 1 62748
box -48 -56 528 834
use sg13g2_a221oi_1  _0390_
timestamp 1685197497
transform -1 0 17952 0 -1 64260
box -48 -56 816 834
use sg13g2_mux4_1  _0391_
timestamp 1677257233
transform 1 0 16032 0 -1 65772
box -48 -56 2064 834
use sg13g2_nand2b_1  _0392_
timestamp 1676567195
transform 1 0 17376 0 -1 29484
box -48 -56 528 834
use sg13g2_nor3_1  _0393_
timestamp 1676639442
transform 1 0 16128 0 -1 29484
box -48 -56 528 834
use sg13g2_a221oi_1  _0394_
timestamp 1685197497
transform 1 0 16608 0 -1 29484
box -48 -56 816 834
use sg13g2_mux4_1  _0395_
timestamp 1677257233
transform 1 0 15936 0 1 30996
box -48 -56 2064 834
use sg13g2_mux4_1  _0396_
timestamp 1677257233
transform 1 0 16608 0 1 56700
box -48 -56 2064 834
use sg13g2_mux4_1  _0397_
timestamp 1677257233
transform 1 0 15552 0 1 71820
box -48 -56 2064 834
use sg13g2_nand2b_1  _0398_
timestamp 1676567195
transform -1 0 7776 0 -1 74844
box -48 -56 528 834
use sg13g2_nor3_1  _0399_
timestamp 1676639442
transform 1 0 6240 0 -1 73332
box -48 -56 528 834
use sg13g2_a221oi_1  _0400_
timestamp 1685197497
transform 1 0 6720 0 1 73332
box -48 -56 816 834
use sg13g2_mux4_1  _0401_
timestamp 1677257233
transform 1 0 4608 0 1 73332
box -48 -56 2064 834
use sg13g2_nand2b_1  _0402_
timestamp 1676567195
transform -1 0 7872 0 -1 38556
box -48 -56 528 834
use sg13g2_nor3_1  _0403_
timestamp 1676639442
transform 1 0 5856 0 -1 40068
box -48 -56 528 834
use sg13g2_a221oi_1  _0404_
timestamp 1685197497
transform 1 0 6336 0 -1 40068
box -48 -56 816 834
use sg13g2_mux4_1  _0405_
timestamp 1677257233
transform 1 0 5280 0 -1 38556
box -48 -56 2064 834
use sg13g2_mux4_1  _0406_
timestamp 1677257233
transform 1 0 7968 0 -1 76356
box -48 -56 2064 834
use sg13g2_mux4_1  _0407_
timestamp 1677257233
transform 1 0 4128 0 1 74844
box -48 -56 2064 834
use sg13g2_mux4_1  _0408_
timestamp 1677257233
transform 1 0 1440 0 -1 65772
box -48 -56 2064 834
use sg13g2_mux2_1  _0409_
timestamp 1677247768
transform 1 0 3264 0 1 26460
box -48 -56 1008 834
use sg13g2_nor2_1  _0410_
timestamp 1676627187
transform -1 0 5760 0 -1 27972
box -48 -56 432 834
use sg13g2_nand2b_1  _0411_
timestamp 1676567195
transform 1 0 3072 0 1 27972
box -48 -56 528 834
use sg13g2_nand2_1  _0412_
timestamp 1676557249
transform -1 0 4320 0 -1 29484
box -48 -56 432 834
use sg13g2_nand3_1  _0413_
timestamp 1683988354
transform 1 0 3552 0 1 27972
box -48 -56 528 834
use sg13g2_nand2b_1  _0414_
timestamp 1676567195
transform -1 0 4896 0 -1 27972
box -48 -56 528 834
use sg13g2_nor2b_1  _0415_
timestamp 1685181386
transform 1 0 4896 0 -1 27972
box -54 -56 528 834
use sg13g2_mux4_1  _0416_
timestamp 1677257233
transform 1 0 1248 0 1 26460
box -48 -56 2064 834
use sg13g2_mux4_1  _0417_
timestamp 1677257233
transform 1 0 2688 0 -1 77868
box -48 -56 2064 834
use sg13g2_mux4_1  _0418_
timestamp 1677257233
transform 1 0 1344 0 -1 76356
box -48 -56 2064 834
use sg13g2_mux4_1  _0419_
timestamp 1677257233
transform 1 0 2208 0 1 67284
box -48 -56 2064 834
use sg13g2_mux2_1  _0420_
timestamp 1677247768
transform 1 0 9696 0 1 2268
box -48 -56 1008 834
use sg13g2_nor2_1  _0421_
timestamp 1676627187
transform -1 0 11040 0 1 2268
box -48 -56 432 834
use sg13g2_nand2b_1  _0422_
timestamp 1676567195
transform 1 0 9312 0 -1 2268
box -48 -56 528 834
use sg13g2_nand2_1  _0423_
timestamp 1676557249
transform -1 0 11040 0 -1 3780
box -48 -56 432 834
use sg13g2_nand3_1  _0424_
timestamp 1683988354
transform 1 0 9792 0 -1 2268
box -48 -56 528 834
use sg13g2_nand2b_1  _0425_
timestamp 1676567195
transform -1 0 10560 0 1 3780
box -48 -56 528 834
use sg13g2_nor2b_1  _0426_
timestamp 1685181386
transform 1 0 10176 0 -1 3780
box -54 -56 528 834
use sg13g2_mux4_1  _0427_
timestamp 1677257233
transform 1 0 9120 0 -1 24948
box -48 -56 2064 834
use sg13g2_mux4_1  _0428_
timestamp 1677257233
transform 1 0 9792 0 1 68796
box -48 -56 2064 834
use sg13g2_mux4_1  _0429_
timestamp 1677257233
transform 1 0 1728 0 1 68796
box -48 -56 2064 834
use sg13g2_mux4_1  _0430_
timestamp 1677257233
transform 1 0 9408 0 1 67284
box -48 -56 2064 834
use sg13g2_mux2_1  _0431_
timestamp 1677247768
transform 1 0 11904 0 -1 30996
box -48 -56 1008 834
use sg13g2_nor2_1  _0432_
timestamp 1676627187
transform -1 0 13440 0 1 30996
box -48 -56 432 834
use sg13g2_nand2b_1  _0433_
timestamp 1676567195
transform -1 0 11424 0 1 30996
box -48 -56 528 834
use sg13g2_nand2_1  _0434_
timestamp 1676557249
transform 1 0 12192 0 1 32508
box -48 -56 432 834
use sg13g2_nand3_1  _0435_
timestamp 1683988354
transform 1 0 12768 0 -1 32508
box -48 -56 528 834
use sg13g2_nand2b_1  _0436_
timestamp 1676567195
transform 1 0 12864 0 -1 30996
box -48 -56 528 834
use sg13g2_nor2b_1  _0437_
timestamp 1685181386
transform -1 0 13056 0 1 29484
box -54 -56 528 834
use sg13g2_mux4_1  _0438_
timestamp 1677257233
transform 1 0 11712 0 -1 29484
box -48 -56 2064 834
use sg13g2_mux4_1  _0439_
timestamp 1677257233
transform 1 0 11712 0 1 71820
box -48 -56 2064 834
use sg13g2_mux4_1  _0440_
timestamp 1677257233
transform 1 0 8448 0 -1 68796
box -48 -56 2064 834
use sg13g2_mux4_1  _0441_
timestamp 1677257233
transform 1 0 1824 0 1 71820
box -48 -56 2064 834
use sg13g2_mux2_1  _0442_
timestamp 1677247768
transform -1 0 4320 0 -1 35532
box -48 -56 1008 834
use sg13g2_nor2_1  _0443_
timestamp 1676627187
transform 1 0 2976 0 -1 35532
box -48 -56 432 834
use sg13g2_nand2b_1  _0444_
timestamp 1676567195
transform 1 0 4416 0 1 35532
box -48 -56 528 834
use sg13g2_nand2_1  _0445_
timestamp 1676557249
transform -1 0 5280 0 -1 37044
box -48 -56 432 834
use sg13g2_nand3_1  _0446_
timestamp 1683988354
transform -1 0 4896 0 -1 37044
box -48 -56 528 834
use sg13g2_nand2b_1  _0447_
timestamp 1676567195
transform 1 0 4032 0 1 34020
box -48 -56 528 834
use sg13g2_nor2b_1  _0448_
timestamp 1685181386
transform -1 0 3936 0 -1 34020
box -54 -56 528 834
use sg13g2_mux4_1  _0449_
timestamp 1677257233
transform 1 0 2016 0 1 34020
box -48 -56 2064 834
use sg13g2_mux4_1  _0450_
timestamp 1677257233
transform 1 0 3456 0 1 79380
box -48 -56 2064 834
use sg13g2_mux4_1  _0451_
timestamp 1677257233
transform 1 0 1632 0 1 73332
box -48 -56 2064 834
use sg13g2_mux4_1  _0452_
timestamp 1677257233
transform 1 0 2592 0 1 62748
box -48 -56 2064 834
use sg13g2_mux4_1  _0453_
timestamp 1677257233
transform 1 0 3840 0 -1 40068
box -48 -56 2064 834
use sg13g2_mux4_1  _0454_
timestamp 1677257233
transform 1 0 1824 0 -1 40068
box -48 -56 2064 834
use sg13g2_mux4_1  _0455_
timestamp 1677257233
transform 1 0 4800 0 -1 43092
box -48 -56 2064 834
use sg13g2_mux4_1  _0456_
timestamp 1677257233
transform 1 0 2112 0 -1 64260
box -48 -56 2064 834
use sg13g2_mux4_1  _0457_
timestamp 1677257233
transform 1 0 2400 0 -1 59724
box -48 -56 2064 834
use sg13g2_mux4_1  _0458_
timestamp 1677257233
transform 1 0 9216 0 1 40068
box -48 -56 2064 834
use sg13g2_mux4_1  _0459_
timestamp 1677257233
transform 1 0 9312 0 -1 26460
box -48 -56 2064 834
use sg13g2_mux4_1  _0460_
timestamp 1677257233
transform 1 0 10656 0 1 74844
box -48 -56 2064 834
use sg13g2_mux4_1  _0461_
timestamp 1677257233
transform 1 0 2304 0 1 70308
box -48 -56 2064 834
use sg13g2_mux4_1  _0462_
timestamp 1677257233
transform 1 0 9024 0 1 59724
box -48 -56 2064 834
use sg13g2_mux4_1  _0463_
timestamp 1677257233
transform 1 0 10272 0 -1 41580
box -48 -56 2064 834
use sg13g2_mux4_1  _0464_
timestamp 1677257233
transform 1 0 10656 0 -1 20412
box -48 -56 2064 834
use sg13g2_mux4_1  _0465_
timestamp 1677257233
transform 1 0 11424 0 -1 70308
box -48 -56 2064 834
use sg13g2_mux4_1  _0466_
timestamp 1677257233
transform 1 0 9024 0 -1 61236
box -48 -56 2064 834
use sg13g2_mux4_1  _0467_
timestamp 1677257233
transform 1 0 2688 0 -1 61236
box -48 -56 2064 834
use sg13g2_mux4_1  _0468_
timestamp 1677257233
transform 1 0 5184 0 -1 41580
box -48 -56 2064 834
use sg13g2_mux4_1  _0469_
timestamp 1677257233
transform 1 0 2208 0 1 37044
box -48 -56 2064 834
use sg13g2_mux4_1  _0470_
timestamp 1677257233
transform 1 0 5280 0 -1 80892
box -48 -56 2064 834
use sg13g2_mux4_1  _0471_
timestamp 1677257233
transform 1 0 2016 0 1 61236
box -48 -56 2064 834
use sg13g2_nand2b_1  _0472_
timestamp 1676567195
transform 1 0 6912 0 1 59724
box -48 -56 528 834
use sg13g2_nor3_1  _0473_
timestamp 1676639442
transform 1 0 6912 0 -1 61236
box -48 -56 528 834
use sg13g2_a221oi_1  _0474_
timestamp 1685197497
transform 1 0 8352 0 -1 59724
box -48 -56 816 834
use sg13g2_mux4_1  _0475_
timestamp 1677257233
transform 1 0 5472 0 1 61236
box -48 -56 2064 834
use sg13g2_nand2b_1  _0476_
timestamp 1676567195
transform 1 0 3552 0 1 30996
box -48 -56 528 834
use sg13g2_nor3_1  _0477_
timestamp 1676639442
transform 1 0 1824 0 -1 30996
box -48 -56 528 834
use sg13g2_a221oi_1  _0478_
timestamp 1685197497
transform 1 0 2784 0 1 30996
box -48 -56 816 834
use sg13g2_mux4_1  _0479_
timestamp 1677257233
transform 1 0 4320 0 1 30996
box -48 -56 2064 834
use sg13g2_mux4_1  _0480_
timestamp 1677257233
transform 1 0 7776 0 1 43092
box -48 -56 2064 834
use sg13g2_mux4_1  _0481_
timestamp 1677257233
transform 1 0 12384 0 1 46116
box -48 -56 2064 834
use sg13g2_mux4_1  _0482_
timestamp 1677257233
transform 1 0 15552 0 -1 44604
box -48 -56 2064 834
use sg13g2_mux4_1  _0483_
timestamp 1677257233
transform 1 0 8640 0 -1 49140
box -48 -56 2064 834
use sg13g2_mux4_1  _0484_
timestamp 1677257233
transform 1 0 5376 0 -1 44604
box -48 -56 2064 834
use sg13g2_mux4_1  _0485_
timestamp 1677257233
transform 1 0 17760 0 1 46116
box -48 -56 2064 834
use sg13g2_mux4_1  _0486_
timestamp 1677257233
transform 1 0 9696 0 1 46116
box -48 -56 2064 834
use sg13g2_mux4_1  _0487_
timestamp 1677257233
transform -1 0 4128 0 -1 55188
box -48 -56 2064 834
use sg13g2_mux4_1  _0488_
timestamp 1677257233
transform -1 0 4224 0 1 41580
box -48 -56 2064 834
use sg13g2_mux4_1  _0489_
timestamp 1677257233
transform 1 0 14976 0 -1 46116
box -48 -56 2064 834
use sg13g2_mux4_1  _0490_
timestamp 1677257233
transform 1 0 11616 0 -1 44604
box -48 -56 2064 834
use sg13g2_mux4_1  _0491_
timestamp 1677257233
transform -1 0 4320 0 1 44604
box -48 -56 2064 834
use sg13g2_mux4_1  _0492_
timestamp 1677257233
transform 1 0 5472 0 1 44604
box -48 -56 2064 834
use sg13g2_mux4_1  _0493_
timestamp 1677257233
transform 1 0 17760 0 1 44604
box -48 -56 2064 834
use sg13g2_mux4_1  _0494_
timestamp 1677257233
transform 1 0 9312 0 -1 46116
box -48 -56 2064 834
use sg13g2_mux4_1  _0495_
timestamp 1677257233
transform 1 0 2112 0 -1 47628
box -48 -56 2064 834
use sg13g2_mux4_1  _0496_
timestamp 1677257233
transform -1 0 4416 0 1 43092
box -48 -56 2064 834
use sg13g2_mux4_1  _0497_
timestamp 1677257233
transform 1 0 14880 0 -1 47628
box -48 -56 2064 834
use sg13g2_mux4_1  _0498_
timestamp 1677257233
transform 1 0 11520 0 1 43092
box -48 -56 2064 834
use sg13g2_mux4_1  _0499_
timestamp 1677257233
transform -1 0 4224 0 1 49140
box -48 -56 2064 834
use sg13g2_mux4_1  _0500_
timestamp 1677257233
transform -1 0 6624 0 -1 50652
box -48 -56 2064 834
use sg13g2_mux4_1  _0501_
timestamp 1677257233
transform 1 0 18144 0 -1 52164
box -48 -56 2064 834
use sg13g2_mux4_1  _0502_
timestamp 1677257233
transform 1 0 11424 0 1 49140
box -48 -56 2064 834
use sg13g2_mux4_1  _0503_
timestamp 1677257233
transform 1 0 7296 0 -1 56700
box -48 -56 2064 834
use sg13g2_mux4_1  _0504_
timestamp 1677257233
transform 1 0 4992 0 1 55188
box -48 -56 2064 834
use sg13g2_mux4_1  _0505_
timestamp 1677257233
transform 1 0 8256 0 1 76356
box -48 -56 2064 834
use sg13g2_mux4_1  _0506_
timestamp 1677257233
transform -1 0 7200 0 1 47628
box -48 -56 2064 834
use sg13g2_mux4_1  _0507_
timestamp 1677257233
transform 1 0 17280 0 -1 56700
box -48 -56 2064 834
use sg13g2_mux4_1  _0508_
timestamp 1677257233
transform 1 0 15168 0 1 49140
box -48 -56 2064 834
use sg13g2_mux4_1  _0509_
timestamp 1677257233
transform 1 0 13056 0 1 50652
box -48 -56 2064 834
use sg13g2_mux4_1  _0510_
timestamp 1677257233
transform 1 0 10272 0 1 50652
box -48 -56 2064 834
use sg13g2_mux4_1  _0511_
timestamp 1677257233
transform 1 0 7392 0 -1 53676
box -48 -56 2064 834
use sg13g2_mux4_1  _0512_
timestamp 1677257233
transform -1 0 4320 0 -1 52164
box -48 -56 2064 834
use sg13g2_mux4_1  _0513_
timestamp 1677257233
transform 1 0 7584 0 -1 77868
box -48 -56 2064 834
use sg13g2_mux4_1  _0514_
timestamp 1677257233
transform -1 0 9696 0 1 47628
box -48 -56 2064 834
use sg13g2_mux4_1  _0515_
timestamp 1677257233
transform 1 0 17376 0 1 59724
box -48 -56 2064 834
use sg13g2_mux4_1  _0516_
timestamp 1677257233
transform 1 0 17856 0 -1 49140
box -48 -56 2064 834
use sg13g2_mux4_1  _0517_
timestamp 1677257233
transform 1 0 12480 0 1 52164
box -48 -56 2064 834
use sg13g2_mux4_1  _0518_
timestamp 1677257233
transform 1 0 10176 0 1 52164
box -48 -56 2064 834
use sg13g2_mux4_1  _0519_
timestamp 1677257233
transform 1 0 6720 0 1 52164
box -48 -56 2064 834
use sg13g2_mux4_1  _0520_
timestamp 1677257233
transform -1 0 5088 0 -1 53676
box -48 -56 2064 834
use sg13g2_mux4_1  _0521_
timestamp 1677257233
transform 1 0 8256 0 1 77868
box -48 -56 2064 834
use sg13g2_mux4_1  _0522_
timestamp 1677257233
transform 1 0 5184 0 1 50652
box -48 -56 2064 834
use sg13g2_mux4_1  _0523_
timestamp 1677257233
transform 1 0 17376 0 -1 59724
box -48 -56 2064 834
use sg13g2_mux4_1  _0524_
timestamp 1677257233
transform 1 0 15552 0 -1 52164
box -48 -56 2064 834
use sg13g2_mux4_1  _0525_
timestamp 1677257233
transform 1 0 12864 0 -1 55188
box -48 -56 2064 834
use sg13g2_mux4_1  _0526_
timestamp 1677257233
transform 1 0 17184 0 -1 55188
box -48 -56 2064 834
use sg13g2_mux4_1  _0527_
timestamp 1677257233
transform 1 0 7008 0 1 56700
box -48 -56 2064 834
use sg13g2_mux4_1  _0528_
timestamp 1677257233
transform -1 0 4992 0 -1 56700
box -48 -56 2064 834
use sg13g2_mux4_1  _0529_
timestamp 1677257233
transform 1 0 7776 0 1 55188
box -48 -56 2064 834
use sg13g2_mux4_1  _0530_
timestamp 1677257233
transform 1 0 14880 0 -1 55188
box -48 -56 2064 834
use sg13g2_mux4_1  _0531_
timestamp 1677257233
transform 1 0 13632 0 1 56700
box -48 -56 2064 834
use sg13g2_mux4_1  _0532_
timestamp 1677257233
transform 1 0 8256 0 -1 58212
box -48 -56 2064 834
use sg13g2_mux4_1  _0533_
timestamp 1677257233
transform 1 0 4800 0 -1 47628
box -48 -56 2064 834
use sg13g2_mux4_1  _0534_
timestamp 1677257233
transform 1 0 17376 0 -1 50652
box -48 -56 2064 834
use sg13g2_mux4_1  _0535_
timestamp 1677257233
transform 1 0 10560 0 1 55188
box -48 -56 2064 834
use sg13g2_mux4_1  _0536_
timestamp 1677257233
transform 1 0 3168 0 1 53676
box -48 -56 2064 834
use sg13g2_mux4_1  _0537_
timestamp 1677257233
transform 1 0 7392 0 1 50652
box -48 -56 2064 834
use sg13g2_mux4_1  _0538_
timestamp 1677257233
transform 1 0 14976 0 -1 53676
box -48 -56 2064 834
use sg13g2_mux4_1  _0539_
timestamp 1677257233
transform 1 0 11424 0 1 56700
box -48 -56 2064 834
use sg13g2_mux4_1  _0540_
timestamp 1677257233
transform 1 0 3456 0 -1 58212
box -48 -56 2064 834
use sg13g2_nand2b_1  _0541_
timestamp 1676567195
transform -1 0 6336 0 -1 65772
box -48 -56 528 834
use sg13g2_o21ai_1  _0542_
timestamp 1685175443
transform -1 0 4320 0 1 65772
box -48 -56 538 834
use sg13g2_o21ai_1  _0543_
timestamp 1685175443
transform -1 0 3840 0 1 65772
box -48 -56 538 834
use sg13g2_mux2_1  _0544_
timestamp 1677247768
transform 1 0 6336 0 1 65772
box -48 -56 1008 834
use sg13g2_a21oi_1  _0545_
timestamp 1683973020
transform 1 0 6336 0 -1 65772
box -48 -56 528 834
use sg13g2_mux4_1  _0546_
timestamp 1677257233
transform 1 0 4320 0 1 65772
box -48 -56 2064 834
use sg13g2_nor2_1  _0547_
timestamp 1676627187
transform 1 0 5088 0 1 64260
box -48 -56 432 834
use sg13g2_nor2_1  _0548_
timestamp 1676627187
transform -1 0 9888 0 -1 67284
box -48 -56 432 834
use sg13g2_nand2b_1  _0549_
timestamp 1676567195
transform 1 0 12480 0 1 62748
box -48 -56 528 834
use sg13g2_o21ai_1  _0550_
timestamp 1685175443
transform 1 0 13152 0 1 64260
box -48 -56 538 834
use sg13g2_o21ai_1  _0551_
timestamp 1685175443
transform 1 0 12672 0 -1 65772
box -48 -56 538 834
use sg13g2_mux2_1  _0552_
timestamp 1677247768
transform 1 0 12384 0 -1 64260
box -48 -56 1008 834
use sg13g2_a21oi_1  _0553_
timestamp 1683973020
transform 1 0 13152 0 -1 65772
box -48 -56 528 834
use sg13g2_mux4_1  _0554_
timestamp 1677257233
transform 1 0 11136 0 1 64260
box -48 -56 2064 834
use sg13g2_nor2_1  _0555_
timestamp 1676627187
transform -1 0 14016 0 1 64260
box -48 -56 432 834
use sg13g2_nor2_1  _0556_
timestamp 1676627187
transform -1 0 12672 0 1 65772
box -48 -56 432 834
use sg13g2_nand2b_1  _0557_
timestamp 1676567195
transform -1 0 17280 0 -1 70308
box -48 -56 528 834
use sg13g2_o21ai_1  _0558_
timestamp 1685175443
transform -1 0 16800 0 -1 70308
box -48 -56 538 834
use sg13g2_o21ai_1  _0559_
timestamp 1685175443
transform 1 0 15168 0 1 70308
box -48 -56 538 834
use sg13g2_mux2_1  _0560_
timestamp 1677247768
transform -1 0 16224 0 1 68796
box -48 -56 1008 834
use sg13g2_a21oi_1  _0561_
timestamp 1683973020
transform -1 0 15168 0 1 70308
box -48 -56 528 834
use sg13g2_mux4_1  _0562_
timestamp 1677257233
transform 1 0 14304 0 -1 70308
box -48 -56 2064 834
use sg13g2_nor2_1  _0563_
timestamp 1676627187
transform 1 0 15456 0 -1 71820
box -48 -56 432 834
use sg13g2_nor2_1  _0564_
timestamp 1676627187
transform -1 0 16032 0 1 70308
box -48 -56 432 834
use sg13g2_nand2b_1  _0565_
timestamp 1676567195
transform 1 0 5952 0 1 76356
box -48 -56 528 834
use sg13g2_o21ai_1  _0566_
timestamp 1685175443
transform 1 0 6816 0 -1 76356
box -48 -56 538 834
use sg13g2_o21ai_1  _0567_
timestamp 1685175443
transform 1 0 7296 0 -1 76356
box -48 -56 538 834
use sg13g2_mux2_1  _0568_
timestamp 1677247768
transform 1 0 4992 0 -1 77868
box -48 -56 1008 834
use sg13g2_a21oi_1  _0569_
timestamp 1683973020
transform 1 0 7776 0 -1 79380
box -48 -56 528 834
use sg13g2_mux4_1  _0570_
timestamp 1677257233
transform 1 0 4800 0 -1 76356
box -48 -56 2064 834
use sg13g2_nor2_1  _0571_
timestamp 1676627187
transform 1 0 5760 0 -1 79380
box -48 -56 432 834
use sg13g2_nor2_1  _0572_
timestamp 1676627187
transform -1 0 7488 0 1 79380
box -48 -56 432 834
use sg13g2_nand2b_1  _0573_
timestamp 1676567195
transform 1 0 8832 0 1 64260
box -48 -56 528 834
use sg13g2_o21ai_1  _0574_
timestamp 1685175443
transform 1 0 9504 0 -1 62748
box -48 -56 538 834
use sg13g2_o21ai_1  _0575_
timestamp 1685175443
transform 1 0 10176 0 1 62748
box -48 -56 538 834
use sg13g2_inv_1  _0576_
timestamp 1676382929
transform 1 0 11040 0 1 62748
box -48 -56 336 834
use sg13g2_nand2b_1  _0577_
timestamp 1676567195
transform 1 0 7776 0 -1 64260
box -48 -56 528 834
use sg13g2_and2_1  _0578_
timestamp 1676901763
transform 1 0 8256 0 -1 64260
box -48 -56 528 834
use sg13g2_o21ai_1  _0579_
timestamp 1685175443
transform 1 0 9024 0 -1 62748
box -48 -56 538 834
use sg13g2_mux4_1  _0580_
timestamp 1677257233
transform 1 0 7488 0 1 62748
box -48 -56 2064 834
use sg13g2_nor2_1  _0581_
timestamp 1676627187
transform -1 0 11040 0 1 62748
box -48 -56 432 834
use sg13g2_a21oi_1  _0582_
timestamp 1683973020
transform -1 0 10176 0 1 62748
box -48 -56 528 834
use sg13g2_nand2b_1  _0583_
timestamp 1676567195
transform 1 0 14688 0 1 61236
box -48 -56 528 834
use sg13g2_o21ai_1  _0584_
timestamp 1685175443
transform -1 0 15648 0 -1 62748
box -48 -56 538 834
use sg13g2_o21ai_1  _0585_
timestamp 1685175443
transform 1 0 15168 0 1 61236
box -48 -56 538 834
use sg13g2_inv_1  _0586_
timestamp 1676382929
transform 1 0 17472 0 -1 58212
box -48 -56 336 834
use sg13g2_nand2b_1  _0587_
timestamp 1676567195
transform -1 0 16224 0 1 58212
box -48 -56 528 834
use sg13g2_and2_1  _0588_
timestamp 1676901763
transform 1 0 15648 0 -1 62748
box -48 -56 528 834
use sg13g2_o21ai_1  _0589_
timestamp 1685175443
transform 1 0 16224 0 1 58212
box -48 -56 538 834
use sg13g2_mux4_1  _0590_
timestamp 1677257233
transform 1 0 13728 0 -1 61236
box -48 -56 2064 834
use sg13g2_nor2_1  _0591_
timestamp 1676627187
transform 1 0 14304 0 1 61236
box -48 -56 432 834
use sg13g2_a21oi_1  _0592_
timestamp 1683973020
transform 1 0 15744 0 -1 61236
box -48 -56 528 834
use sg13g2_nand2b_1  _0593_
timestamp 1676567195
transform 1 0 19584 0 1 68796
box -48 -56 528 834
use sg13g2_o21ai_1  _0594_
timestamp 1685175443
transform 1 0 18144 0 1 68796
box -48 -56 538 834
use sg13g2_o21ai_1  _0595_
timestamp 1685175443
transform 1 0 18624 0 1 68796
box -48 -56 538 834
use sg13g2_inv_1  _0596_
timestamp 1676382929
transform 1 0 19296 0 -1 71820
box -48 -56 336 834
use sg13g2_nand2b_1  _0597_
timestamp 1676567195
transform 1 0 19104 0 1 68796
box -48 -56 528 834
use sg13g2_and2_1  _0598_
timestamp 1676901763
transform 1 0 19680 0 1 70308
box -48 -56 528 834
use sg13g2_o21ai_1  _0599_
timestamp 1685175443
transform 1 0 19200 0 1 70308
box -48 -56 538 834
use sg13g2_mux4_1  _0600_
timestamp 1677257233
transform 1 0 17472 0 -1 70308
box -48 -56 2064 834
use sg13g2_nor2_1  _0601_
timestamp 1676627187
transform -1 0 20352 0 -1 70308
box -48 -56 432 834
use sg13g2_a21oi_1  _0602_
timestamp 1683973020
transform -1 0 19968 0 -1 70308
box -48 -56 528 834
use sg13g2_nand2b_1  _0603_
timestamp 1676567195
transform 1 0 8544 0 -1 74844
box -48 -56 528 834
use sg13g2_o21ai_1  _0604_
timestamp 1685175443
transform 1 0 9024 0 -1 74844
box -48 -56 538 834
use sg13g2_o21ai_1  _0605_
timestamp 1685175443
transform 1 0 9984 0 1 73332
box -48 -56 538 834
use sg13g2_inv_1  _0606_
timestamp 1676382929
transform 1 0 10464 0 1 73332
box -48 -56 336 834
use sg13g2_nand2b_1  _0607_
timestamp 1676567195
transform 1 0 7680 0 1 73332
box -48 -56 528 834
use sg13g2_and2_1  _0608_
timestamp 1676901763
transform 1 0 9504 0 -1 74844
box -48 -56 528 834
use sg13g2_o21ai_1  _0609_
timestamp 1685175443
transform 1 0 9984 0 -1 74844
box -48 -56 538 834
use sg13g2_mux4_1  _0610_
timestamp 1677257233
transform 1 0 8352 0 -1 73332
box -48 -56 2064 834
use sg13g2_nor2_1  _0611_
timestamp 1676627187
transform -1 0 10656 0 -1 76356
box -48 -56 432 834
use sg13g2_a21oi_1  _0612_
timestamp 1683973020
transform -1 0 10848 0 -1 73332
box -48 -56 528 834
use sg13g2_mux4_1  _0613_
timestamp 1677257233
transform 1 0 6048 0 1 26460
box -48 -56 2064 834
use sg13g2_mux4_1  _0614_
timestamp 1677257233
transform 1 0 14976 0 1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _0615_
timestamp 1677257233
transform 1 0 16512 0 1 15876
box -48 -56 2064 834
use sg13g2_mux4_1  _0616_
timestamp 1677257233
transform 1 0 8352 0 -1 38556
box -48 -56 2064 834
use sg13g2_a21oi_1  _0617_
timestamp 1683973020
transform -1 0 4512 0 -1 68796
box -48 -56 528 834
use sg13g2_o21ai_1  _0618_
timestamp 1685175443
transform 1 0 6048 0 -1 70308
box -48 -56 538 834
use sg13g2_mux4_1  _0619_
timestamp 1677257233
transform 1 0 4512 0 -1 68796
box -48 -56 2064 834
use sg13g2_nor2_1  _0620_
timestamp 1676627187
transform -1 0 7104 0 -1 70308
box -48 -56 432 834
use sg13g2_a21oi_1  _0621_
timestamp 1683973020
transform -1 0 7488 0 1 68796
box -48 -56 528 834
use sg13g2_a21oi_1  _0622_
timestamp 1683973020
transform -1 0 13920 0 1 65772
box -48 -56 528 834
use sg13g2_o21ai_1  _0623_
timestamp 1685175443
transform 1 0 12960 0 1 65772
box -48 -56 538 834
use sg13g2_mux4_1  _0624_
timestamp 1677257233
transform 1 0 11904 0 -1 67284
box -48 -56 2064 834
use sg13g2_nor2_1  _0625_
timestamp 1676627187
transform -1 0 14400 0 1 67284
box -48 -56 432 834
use sg13g2_a21oi_1  _0626_
timestamp 1683973020
transform -1 0 14592 0 1 65772
box -48 -56 528 834
use sg13g2_a21oi_1  _0627_
timestamp 1683973020
transform 1 0 16704 0 1 67284
box -48 -56 528 834
use sg13g2_o21ai_1  _0628_
timestamp 1685175443
transform 1 0 16224 0 1 65772
box -48 -56 538 834
use sg13g2_mux4_1  _0629_
timestamp 1677257233
transform 1 0 14688 0 1 67284
box -48 -56 2064 834
use sg13g2_nor2_1  _0630_
timestamp 1676627187
transform -1 0 17088 0 1 65772
box -48 -56 432 834
use sg13g2_a21oi_1  _0631_
timestamp 1683973020
transform -1 0 17664 0 -1 67284
box -48 -56 528 834
use sg13g2_a21oi_1  _0632_
timestamp 1683973020
transform -1 0 5856 0 -1 71820
box -48 -56 528 834
use sg13g2_o21ai_1  _0633_
timestamp 1685175443
transform 1 0 6144 0 1 71820
box -48 -56 538 834
use sg13g2_mux4_1  _0634_
timestamp 1677257233
transform 1 0 4896 0 1 70308
box -48 -56 2064 834
use sg13g2_nor2_1  _0635_
timestamp 1676627187
transform -1 0 7776 0 1 70308
box -48 -56 432 834
use sg13g2_a21oi_1  _0636_
timestamp 1683973020
transform -1 0 7392 0 1 70308
box -48 -56 528 834
use sg13g2_nor2b_1  _0637_
timestamp 1685181386
transform -1 0 7392 0 -1 65772
box -54 -56 528 834
use sg13g2_o21ai_1  _0638_
timestamp 1685175443
transform 1 0 8544 0 -1 67284
box -48 -56 538 834
use sg13g2_mux4_1  _0639_
timestamp 1677257233
transform 1 0 7392 0 -1 65772
box -48 -56 2064 834
use sg13g2_nor2b_1  _0640_
timestamp 1685181386
transform 1 0 9312 0 1 65772
box -54 -56 528 834
use sg13g2_nor3_1  _0641_
timestamp 1676639442
transform 1 0 9024 0 -1 67284
box -48 -56 528 834
use sg13g2_or2_1  _0642_
timestamp 1684236171
transform 1 0 9792 0 1 65772
box -48 -56 528 834
use sg13g2_nor2b_1  _0643_
timestamp 1685181386
transform 1 0 15648 0 -1 64260
box -54 -56 528 834
use sg13g2_o21ai_1  _0644_
timestamp 1685175443
transform 1 0 14688 0 -1 62748
box -48 -56 538 834
use sg13g2_mux4_1  _0645_
timestamp 1677257233
transform 1 0 13632 0 -1 64260
box -48 -56 2064 834
use sg13g2_nor2b_1  _0646_
timestamp 1685181386
transform 1 0 15648 0 1 64260
box -54 -56 528 834
use sg13g2_nor3_1  _0647_
timestamp 1676639442
transform 1 0 16128 0 -1 64260
box -48 -56 528 834
use sg13g2_or2_1  _0648_
timestamp 1684236171
transform 1 0 16608 0 -1 64260
box -48 -56 528 834
use sg13g2_nor2b_1  _0649_
timestamp 1685181386
transform -1 0 19008 0 -1 68796
box -54 -56 528 834
use sg13g2_o21ai_1  _0650_
timestamp 1685175443
transform 1 0 19392 0 1 67284
box -48 -56 538 834
use sg13g2_mux4_1  _0651_
timestamp 1677257233
transform 1 0 17376 0 1 67284
box -48 -56 2064 834
use sg13g2_nor2b_1  _0652_
timestamp 1685181386
transform -1 0 20352 0 1 67284
box -54 -56 528 834
use sg13g2_nor3_1  _0653_
timestamp 1676639442
transform 1 0 19008 0 -1 68796
box -48 -56 528 834
use sg13g2_or2_1  _0654_
timestamp 1684236171
transform 1 0 19584 0 -1 67284
box -48 -56 528 834
use sg13g2_nor2b_1  _0655_
timestamp 1685181386
transform 1 0 8544 0 1 71820
box -54 -56 528 834
use sg13g2_o21ai_1  _0656_
timestamp 1685175443
transform 1 0 9024 0 1 71820
box -48 -56 538 834
use sg13g2_mux4_1  _0657_
timestamp 1677257233
transform 1 0 7872 0 1 70308
box -48 -56 2064 834
use sg13g2_nor2b_1  _0658_
timestamp 1685181386
transform 1 0 9984 0 1 71820
box -54 -56 528 834
use sg13g2_nor3_1  _0659_
timestamp 1676639442
transform 1 0 9504 0 1 71820
box -48 -56 528 834
use sg13g2_or2_1  _0660_
timestamp 1684236171
transform 1 0 10176 0 1 70308
box -48 -56 528 834
use sg13g2_mux4_1  _0661_
timestamp 1677257233
transform 1 0 5280 0 -1 64260
box -48 -56 2064 834
use sg13g2_mux4_1  _0662_
timestamp 1677257233
transform 1 0 3936 0 -1 30996
box -48 -56 2064 834
use sg13g2_mux4_1  _0663_
timestamp 1677257233
transform 1 0 13344 0 1 18900
box -48 -56 2064 834
use sg13g2_mux4_1  _0664_
timestamp 1677257233
transform 1 0 14304 0 1 27972
box -48 -56 2064 834
use sg13g2_mux4_1  _0665_
timestamp 1677257233
transform 1 0 5856 0 1 37044
box -48 -56 2064 834
use sg13g2_mux4_1  _0666_
timestamp 1677257233
transform 1 0 1344 0 1 20412
box -48 -56 2064 834
use sg13g2_mux4_1  _0667_
timestamp 1677257233
transform 1 0 9120 0 -1 21924
box -48 -56 2064 834
use sg13g2_mux4_1  _0668_
timestamp 1677257233
transform 1 0 11616 0 1 26460
box -48 -56 2064 834
use sg13g2_mux4_1  _0669_
timestamp 1677257233
transform 1 0 2496 0 1 32508
box -48 -56 2064 834
use sg13g2_mux4_1  _0670_
timestamp 1677257233
transform 1 0 7104 0 1 20412
box -48 -56 2064 834
use sg13g2_mux4_1  _0671_
timestamp 1677257233
transform 1 0 9216 0 -1 17388
box -48 -56 2064 834
use sg13g2_mux4_1  _0672_
timestamp 1677257233
transform 1 0 10848 0 -1 18900
box -48 -56 2064 834
use sg13g2_mux4_1  _0673_
timestamp 1677257233
transform 1 0 8448 0 1 18900
box -48 -56 2064 834
use sg13g2_mux4_1  _0674_
timestamp 1677257233
transform 1 0 6816 0 -1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _0675_
timestamp 1677257233
transform 1 0 12672 0 -1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _0676_
timestamp 1677257233
transform 1 0 16992 0 1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _0677_
timestamp 1677257233
transform 1 0 6336 0 1 5292
box -48 -56 2064 834
use sg13g2_nand2b_1  _0678_
timestamp 1676567195
transform 1 0 2784 0 -1 18900
box -48 -56 528 834
use sg13g2_nor3_1  _0679_
timestamp 1676639442
transform 1 0 1248 0 1 17388
box -48 -56 528 834
use sg13g2_a221oi_1  _0680_
timestamp 1685197497
transform 1 0 2784 0 -1 17388
box -48 -56 816 834
use sg13g2_nand2b_1  _0681_
timestamp 1676567195
transform 1 0 5568 0 -1 2268
box -48 -56 528 834
use sg13g2_nor3_1  _0682_
timestamp 1676639442
transform -1 0 5568 0 1 756
box -48 -56 528 834
use sg13g2_a221oi_1  _0683_
timestamp 1685197497
transform 1 0 5088 0 1 2268
box -48 -56 816 834
use sg13g2_nand2b_1  _0684_
timestamp 1676567195
transform 1 0 9984 0 -1 5292
box -48 -56 528 834
use sg13g2_nor3_1  _0685_
timestamp 1676639442
transform 1 0 9504 0 1 3780
box -48 -56 528 834
use sg13g2_a221oi_1  _0686_
timestamp 1685197497
transform 1 0 10080 0 1 5292
box -48 -56 816 834
use sg13g2_nand2b_1  _0687_
timestamp 1676567195
transform -1 0 2880 0 1 8316
box -48 -56 528 834
use sg13g2_nor3_1  _0688_
timestamp 1676639442
transform -1 0 3168 0 -1 9828
box -48 -56 528 834
use sg13g2_a221oi_1  _0689_
timestamp 1685197497
transform 1 0 2880 0 1 8316
box -48 -56 816 834
use sg13g2_nand2b_1  _0690_
timestamp 1676567195
transform 1 0 3360 0 1 14364
box -48 -56 528 834
use sg13g2_nor3_1  _0691_
timestamp 1676639442
transform -1 0 3648 0 1 15876
box -48 -56 528 834
use sg13g2_a221oi_1  _0692_
timestamp 1685197497
transform 1 0 3360 0 -1 15876
box -48 -56 816 834
use sg13g2_nand2b_1  _0693_
timestamp 1676567195
transform -1 0 9120 0 -1 6804
box -48 -56 528 834
use sg13g2_nor3_1  _0694_
timestamp 1676639442
transform -1 0 11232 0 1 6804
box -48 -56 528 834
use sg13g2_a221oi_1  _0695_
timestamp 1685197497
transform 1 0 10752 0 -1 6804
box -48 -56 816 834
use sg13g2_nand2b_1  _0696_
timestamp 1676567195
transform 1 0 7968 0 -1 3780
box -48 -56 528 834
use sg13g2_nor3_1  _0697_
timestamp 1676639442
transform 1 0 7296 0 -1 2268
box -48 -56 528 834
use sg13g2_a221oi_1  _0698_
timestamp 1685197497
transform 1 0 7296 0 1 3780
box -48 -56 816 834
use sg13g2_nand2b_1  _0699_
timestamp 1676567195
transform 1 0 3552 0 -1 12852
box -48 -56 528 834
use sg13g2_nor3_1  _0700_
timestamp 1676639442
transform 1 0 2016 0 -1 14364
box -48 -56 528 834
use sg13g2_a221oi_1  _0701_
timestamp 1685197497
transform 1 0 2784 0 -1 12852
box -48 -56 816 834
use sg13g2_nand2b_1  _0702_
timestamp 1676567195
transform -1 0 3264 0 1 3780
box -48 -56 528 834
use sg13g2_nor3_1  _0703_
timestamp 1676639442
transform 1 0 2016 0 -1 6804
box -48 -56 528 834
use sg13g2_a221oi_1  _0704_
timestamp 1685197497
transform 1 0 2496 0 -1 6804
box -48 -56 816 834
use sg13g2_nand2b_1  _0705_
timestamp 1676567195
transform -1 0 5952 0 1 3780
box -48 -56 528 834
use sg13g2_nor3_1  _0706_
timestamp 1676639442
transform -1 0 5568 0 -1 2268
box -48 -56 528 834
use sg13g2_a221oi_1  _0707_
timestamp 1685197497
transform 1 0 5184 0 -1 3780
box -48 -56 816 834
use sg13g2_nand2b_1  _0708_
timestamp 1676567195
transform 1 0 10272 0 -1 11340
box -48 -56 528 834
use sg13g2_nor3_1  _0709_
timestamp 1676639442
transform 1 0 7872 0 -1 9828
box -48 -56 528 834
use sg13g2_a221oi_1  _0710_
timestamp 1685197497
transform 1 0 9888 0 1 8316
box -48 -56 816 834
use sg13g2_nand2b_1  _0711_
timestamp 1676567195
transform 1 0 4128 0 1 9828
box -48 -56 528 834
use sg13g2_nor3_1  _0712_
timestamp 1676639442
transform 1 0 3168 0 -1 9828
box -48 -56 528 834
use sg13g2_a221oi_1  _0713_
timestamp 1685197497
transform 1 0 3360 0 1 9828
box -48 -56 816 834
use sg13g2_nand2b_1  _0714_
timestamp 1676567195
transform 1 0 5088 0 1 6804
box -48 -56 528 834
use sg13g2_nor3_1  _0715_
timestamp 1676639442
transform 1 0 4032 0 -1 9828
box -48 -56 528 834
use sg13g2_a221oi_1  _0716_
timestamp 1685197497
transform 1 0 4512 0 -1 9828
box -48 -56 816 834
use sg13g2_nand2b_1  _0717_
timestamp 1676567195
transform -1 0 12672 0 -1 5292
box -48 -56 528 834
use sg13g2_nor3_1  _0718_
timestamp 1676639442
transform -1 0 13152 0 -1 5292
box -48 -56 528 834
use sg13g2_a221oi_1  _0719_
timestamp 1685197497
transform -1 0 12288 0 -1 6804
box -48 -56 816 834
use sg13g2_nand2b_1  _0720_
timestamp 1676567195
transform 1 0 6432 0 -1 6804
box -48 -56 528 834
use sg13g2_nor3_1  _0721_
timestamp 1676639442
transform 1 0 6816 0 1 3780
box -48 -56 528 834
use sg13g2_a221oi_1  _0722_
timestamp 1685197497
transform 1 0 7296 0 -1 5292
box -48 -56 816 834
use sg13g2_nand2b_1  _0723_
timestamp 1676567195
transform 1 0 4992 0 -1 5292
box -48 -56 528 834
use sg13g2_nor3_1  _0724_
timestamp 1676639442
transform 1 0 3552 0 -1 6804
box -48 -56 528 834
use sg13g2_a221oi_1  _0725_
timestamp 1685197497
transform 1 0 4032 0 -1 6804
box -48 -56 816 834
use sg13g2_mux4_1  _0726_
timestamp 1677257233
transform 1 0 3360 0 1 17388
box -48 -56 2064 834
use sg13g2_mux4_1  _0727_
timestamp 1677257233
transform 1 0 17280 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _0728_
timestamp 1677257233
transform 1 0 12384 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _0729_
timestamp 1677257233
transform -1 0 7680 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _0730_
timestamp 1677257233
transform 1 0 8160 0 1 35532
box -48 -56 2064 834
use sg13g2_mux4_1  _0731_
timestamp 1677257233
transform 1 0 9120 0 1 15876
box -48 -56 2064 834
use sg13g2_mux4_1  _0732_
timestamp 1677257233
transform 1 0 16896 0 1 14364
box -48 -56 2064 834
use sg13g2_mux4_1  _0733_
timestamp 1677257233
transform 1 0 12960 0 1 11340
box -48 -56 2064 834
use sg13g2_mux4_1  _0734_
timestamp 1677257233
transform 1 0 14880 0 -1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _0735_
timestamp 1677257233
transform 1 0 10656 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _0736_
timestamp 1677257233
transform 1 0 5664 0 1 27972
box -48 -56 2064 834
use sg13g2_mux4_1  _0737_
timestamp 1677257233
transform 1 0 4416 0 1 12852
box -48 -56 2064 834
use sg13g2_mux4_1  _0738_
timestamp 1677257233
transform 1 0 8448 0 1 38556
box -48 -56 2064 834
use sg13g2_mux4_1  _0739_
timestamp 1677257233
transform 1 0 8160 0 1 11340
box -48 -56 2064 834
use sg13g2_mux4_1  _0740_
timestamp 1677257233
transform 1 0 16800 0 -1 18900
box -48 -56 2064 834
use sg13g2_mux4_1  _0741_
timestamp 1677257233
transform -1 0 19680 0 -1 11340
box -48 -56 2064 834
use sg13g2_mux4_1  _0742_
timestamp 1677257233
transform 1 0 15168 0 1 9828
box -48 -56 2064 834
use sg13g2_mux4_1  _0743_
timestamp 1677257233
transform -1 0 12672 0 1 9828
box -48 -56 2064 834
use sg13g2_mux4_1  _0744_
timestamp 1677257233
transform 1 0 6048 0 1 24948
box -48 -56 2064 834
use sg13g2_mux4_1  _0745_
timestamp 1677257233
transform 1 0 5856 0 -1 11340
box -48 -56 2064 834
use sg13g2_mux4_1  _0746_
timestamp 1677257233
transform 1 0 8256 0 1 34020
box -48 -56 2064 834
use sg13g2_mux4_1  _0747_
timestamp 1677257233
transform 1 0 9216 0 -1 14364
box -48 -56 2064 834
use sg13g2_mux4_1  _0748_
timestamp 1677257233
transform 1 0 16800 0 -1 17388
box -48 -56 2064 834
use sg13g2_mux4_1  _0749_
timestamp 1677257233
transform 1 0 13152 0 1 12852
box -48 -56 2064 834
use sg13g2_mux4_1  _0750_
timestamp 1677257233
transform 1 0 14496 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _0751_
timestamp 1677257233
transform 1 0 12672 0 -1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _0752_
timestamp 1677257233
transform 1 0 5760 0 1 18900
box -48 -56 2064 834
use sg13g2_mux4_1  _0753_
timestamp 1677257233
transform 1 0 3744 0 1 11340
box -48 -56 2064 834
use sg13g2_mux4_1  _0754_
timestamp 1677257233
transform 1 0 5856 0 -1 18900
box -48 -56 2064 834
use sg13g2_mux4_1  _0755_
timestamp 1677257233
transform 1 0 15744 0 1 11340
box -48 -56 2064 834
use sg13g2_mux4_1  _0756_
timestamp 1677257233
transform 1 0 12192 0 -1 15876
box -48 -56 2064 834
use sg13g2_mux4_1  _0757_
timestamp 1677257233
transform 1 0 6720 0 -1 29484
box -48 -56 2064 834
use sg13g2_mux4_1  _0758_
timestamp 1677257233
transform 1 0 5664 0 1 15876
box -48 -56 2064 834
use sg13g2_mux4_1  _0759_
timestamp 1677257233
transform 1 0 13344 0 1 14364
box -48 -56 2064 834
use sg13g2_mux4_1  _0760_
timestamp 1677257233
transform 1 0 11040 0 -1 12852
box -48 -56 2064 834
use sg13g2_mux4_1  _0761_
timestamp 1677257233
transform 1 0 3936 0 1 14364
box -48 -56 2064 834
use sg13g2_mux4_1  _0762_
timestamp 1677257233
transform 1 0 6816 0 -1 15876
box -48 -56 2064 834
use sg13g2_mux4_1  _0763_
timestamp 1677257233
transform 1 0 15456 0 -1 14364
box -48 -56 2064 834
use sg13g2_mux4_1  _0764_
timestamp 1677257233
transform 1 0 13056 0 1 9828
box -48 -56 2064 834
use sg13g2_mux4_1  _0765_
timestamp 1677257233
transform -1 0 8736 0 1 12852
box -48 -56 2064 834
use sg13g2_mux2_1  _0766_
timestamp 1677247768
transform -1 0 5760 0 -1 20412
box -48 -56 1008 834
use sg13g2_nand2b_1  _0767_
timestamp 1676567195
transform 1 0 4992 0 1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  _0768_
timestamp 1685175443
transform 1 0 6624 0 -1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  _0769_
timestamp 1683973020
transform -1 0 4800 0 -1 20412
box -48 -56 528 834
use sg13g2_nor2b_1  _0770_
timestamp 1685181386
transform -1 0 6624 0 -1 21924
box -54 -56 528 834
use sg13g2_mux4_1  _0771_
timestamp 1677257233
transform 1 0 3456 0 -1 21924
box -48 -56 2064 834
use sg13g2_nor2_1  _0772_
timestamp 1676627187
transform -1 0 7488 0 -1 21924
box -48 -56 432 834
use sg13g2_a21oi_1  _0773_
timestamp 1683973020
transform -1 0 6144 0 -1 21924
box -48 -56 528 834
use sg13g2_mux2_1  _0774_
timestamp 1677247768
transform 1 0 12000 0 1 21924
box -48 -56 1008 834
use sg13g2_nand2b_1  _0775_
timestamp 1676567195
transform -1 0 13248 0 1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  _0776_
timestamp 1685175443
transform -1 0 12000 0 1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  _0777_
timestamp 1683973020
transform 1 0 12960 0 1 21924
box -48 -56 528 834
use sg13g2_nor2b_1  _0778_
timestamp 1685181386
transform 1 0 11808 0 1 23436
box -54 -56 528 834
use sg13g2_mux4_1  _0779_
timestamp 1677257233
transform -1 0 13632 0 -1 23436
box -48 -56 2064 834
use sg13g2_nor2_1  _0780_
timestamp 1676627187
transform 1 0 11424 0 1 23436
box -48 -56 432 834
use sg13g2_a21oi_1  _0781_
timestamp 1683973020
transform 1 0 12288 0 1 23436
box -48 -56 528 834
use sg13g2_mux2_1  _0782_
timestamp 1677247768
transform 1 0 14784 0 1 29484
box -48 -56 1008 834
use sg13g2_nand2b_1  _0783_
timestamp 1676567195
transform 1 0 15744 0 1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  _0784_
timestamp 1685175443
transform 1 0 15552 0 -1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  _0785_
timestamp 1683973020
transform -1 0 14784 0 -1 32508
box -48 -56 528 834
use sg13g2_nor2b_1  _0786_
timestamp 1685181386
transform -1 0 15264 0 -1 32508
box -54 -56 528 834
use sg13g2_mux4_1  _0787_
timestamp 1677257233
transform 1 0 13536 0 -1 30996
box -48 -56 2064 834
use sg13g2_nor2_1  _0788_
timestamp 1676627187
transform -1 0 15936 0 1 30996
box -48 -56 432 834
use sg13g2_a21oi_1  _0789_
timestamp 1683973020
transform -1 0 15552 0 1 30996
box -48 -56 528 834
use sg13g2_mux2_1  _0790_
timestamp 1677247768
transform 1 0 6432 0 -1 34020
box -48 -56 1008 834
use sg13g2_nand2b_1  _0791_
timestamp 1676567195
transform 1 0 7392 0 -1 34020
box -48 -56 528 834
use sg13g2_o21ai_1  _0792_
timestamp 1685175443
transform -1 0 5376 0 1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  _0793_
timestamp 1683973020
transform -1 0 6432 0 -1 34020
box -48 -56 528 834
use sg13g2_nor2b_1  _0794_
timestamp 1685181386
transform -1 0 7872 0 1 34020
box -54 -56 528 834
use sg13g2_mux4_1  _0795_
timestamp 1677257233
transform 1 0 5376 0 1 34020
box -48 -56 2064 834
use sg13g2_nor2_1  _0796_
timestamp 1676627187
transform -1 0 8256 0 1 34020
box -48 -56 432 834
use sg13g2_a21oi_1  _0797_
timestamp 1683973020
transform -1 0 6816 0 -1 35532
box -48 -56 528 834
use sg13g2_mux2_1  _0798_
timestamp 1677247768
transform 1 0 6528 0 -1 24948
box -48 -56 1008 834
use sg13g2_nand2b_1  _0799_
timestamp 1676567195
transform 1 0 8064 0 1 24948
box -48 -56 528 834
use sg13g2_mux2_1  _0800_
timestamp 1677247768
transform 1 0 7584 0 1 23436
box -48 -56 1008 834
use sg13g2_a21oi_1  _0801_
timestamp 1683973020
transform -1 0 8448 0 1 21924
box -48 -56 528 834
use sg13g2_mux4_1  _0802_
timestamp 1677257233
transform 1 0 5568 0 1 23436
box -48 -56 2064 834
use sg13g2_nor2_1  _0803_
timestamp 1676627187
transform -1 0 9408 0 1 23436
box -48 -56 432 834
use sg13g2_a21oi_1  _0804_
timestamp 1683973020
transform -1 0 9024 0 1 23436
box -48 -56 528 834
use sg13g2_mux2_1  _0805_
timestamp 1677247768
transform 1 0 16032 0 1 20412
box -48 -56 1008 834
use sg13g2_nand2b_1  _0806_
timestamp 1676567195
transform 1 0 17952 0 1 20412
box -48 -56 528 834
use sg13g2_mux2_1  _0807_
timestamp 1677247768
transform 1 0 16992 0 1 20412
box -48 -56 1008 834
use sg13g2_a21oi_1  _0808_
timestamp 1683973020
transform 1 0 17664 0 -1 20412
box -48 -56 528 834
use sg13g2_mux4_1  _0809_
timestamp 1677257233
transform 1 0 15456 0 -1 21924
box -48 -56 2064 834
use sg13g2_nor2_1  _0810_
timestamp 1676627187
transform -1 0 18816 0 1 20412
box -48 -56 432 834
use sg13g2_a21oi_1  _0811_
timestamp 1683973020
transform 1 0 17184 0 -1 20412
box -48 -56 528 834
use sg13g2_mux2_1  _0812_
timestamp 1677247768
transform 1 0 19392 0 1 29484
box -48 -56 1008 834
use sg13g2_nand2b_1  _0813_
timestamp 1676567195
transform -1 0 20160 0 -1 30996
box -48 -56 528 834
use sg13g2_mux2_1  _0814_
timestamp 1677247768
transform 1 0 18240 0 -1 30996
box -48 -56 1008 834
use sg13g2_a21oi_1  _0815_
timestamp 1683973020
transform 1 0 19872 0 -1 29484
box -48 -56 528 834
use sg13g2_mux4_1  _0816_
timestamp 1677257233
transform 1 0 17376 0 1 29484
box -48 -56 2064 834
use sg13g2_nor2_1  _0817_
timestamp 1676627187
transform -1 0 20160 0 1 30996
box -48 -56 432 834
use sg13g2_a21oi_1  _0818_
timestamp 1683973020
transform 1 0 19200 0 -1 30996
box -48 -56 528 834
use sg13g2_mux2_1  _0819_
timestamp 1677247768
transform 1 0 10656 0 -1 30996
box -48 -56 1008 834
use sg13g2_nand2b_1  _0820_
timestamp 1676567195
transform -1 0 11136 0 -1 32508
box -48 -56 528 834
use sg13g2_mux2_1  _0821_
timestamp 1677247768
transform 1 0 9312 0 1 29484
box -48 -56 1008 834
use sg13g2_a21oi_1  _0822_
timestamp 1683973020
transform 1 0 10560 0 -1 29484
box -48 -56 528 834
use sg13g2_mux4_1  _0823_
timestamp 1677257233
transform 1 0 8640 0 -1 30996
box -48 -56 2064 834
use sg13g2_nor2_1  _0824_
timestamp 1676627187
transform 1 0 8928 0 1 29484
box -48 -56 432 834
use sg13g2_a21oi_1  _0825_
timestamp 1683973020
transform 1 0 10368 0 1 29484
box -48 -56 528 834
use sg13g2_nor2_1  _0826_
timestamp 1676627187
transform 1 0 6528 0 1 21924
box -48 -56 432 834
use sg13g2_nor2b_1  _0827_
timestamp 1685181386
transform 1 0 1344 0 -1 23436
box -54 -56 528 834
use sg13g2_mux4_1  _0828_
timestamp 1677257233
transform 1 0 1824 0 -1 23436
box -48 -56 2064 834
use sg13g2_nor3_1  _0829_
timestamp 1676639442
transform -1 0 6528 0 1 21924
box -48 -56 528 834
use sg13g2_mux2_1  _0830_
timestamp 1677247768
transform 1 0 2976 0 1 23436
box -48 -56 1008 834
use sg13g2_mux2_1  _0831_
timestamp 1677247768
transform 1 0 15552 0 -1 23436
box -48 -56 1008 834
use sg13g2_nand3b_1  _0832_
timestamp 1676573470
transform 1 0 15744 0 1 24948
box -48 -56 720 834
use sg13g2_mux4_1  _0833_
timestamp 1677257233
transform 1 0 13344 0 1 23436
box -48 -56 2064 834
use sg13g2_inv_1  _0834_
timestamp 1676382929
transform 1 0 15456 0 1 23436
box -48 -56 336 834
use sg13g2_o21ai_1  _0835_
timestamp 1685175443
transform 1 0 16896 0 -1 24948
box -48 -56 538 834
use sg13g2_nor2b_1  _0836_
timestamp 1685181386
transform 1 0 15264 0 1 24948
box -54 -56 528 834
use sg13g2_nor2_1  _0837_
timestamp 1676627187
transform 1 0 14880 0 1 24948
box -48 -56 432 834
use sg13g2_mux4_1  _0838_
timestamp 1677257233
transform 1 0 13920 0 -1 26460
box -48 -56 2064 834
use sg13g2_nor3_1  _0839_
timestamp 1676639442
transform 1 0 15744 0 1 26460
box -48 -56 528 834
use sg13g2_mux2_1  _0840_
timestamp 1677247768
transform 1 0 16512 0 1 24948
box -48 -56 1008 834
use sg13g2_nor2_1  _0841_
timestamp 1676627187
transform 1 0 6432 0 1 30996
box -48 -56 432 834
use sg13g2_nor2b_1  _0842_
timestamp 1685181386
transform 1 0 8160 0 1 32508
box -54 -56 528 834
use sg13g2_mux4_1  _0843_
timestamp 1677257233
transform 1 0 5664 0 -1 32508
box -48 -56 2064 834
use sg13g2_nor3_1  _0844_
timestamp 1676639442
transform 1 0 7680 0 1 32508
box -48 -56 528 834
use sg13g2_mux2_1  _0845_
timestamp 1677247768
transform 1 0 7872 0 -1 32508
box -48 -56 1008 834
use sg13g2_mux4_1  _0846_
timestamp 1677257233
transform 1 0 2592 0 1 24948
box -48 -56 2064 834
use sg13g2_nand2b_1  _0847_
timestamp 1676567195
transform 1 0 5088 0 -1 26460
box -48 -56 528 834
use sg13g2_nand2b_1  _0848_
timestamp 1676567195
transform -1 0 2592 0 1 24948
box -48 -56 528 834
use sg13g2_nand2b_1  _0849_
timestamp 1676567195
transform -1 0 6048 0 1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  _0850_
timestamp 1685175443
transform -1 0 5568 0 1 24948
box -48 -56 538 834
use sg13g2_o21ai_1  _0851_
timestamp 1685175443
transform 1 0 4608 0 1 24948
box -48 -56 538 834
use sg13g2_mux4_1  _0852_
timestamp 1677257233
transform 1 0 15744 0 1 23436
box -48 -56 2064 834
use sg13g2_nand2b_1  _0853_
timestamp 1676567195
transform 1 0 19680 0 1 23436
box -48 -56 528 834
use sg13g2_nand2b_1  _0854_
timestamp 1676567195
transform 1 0 19104 0 -1 23436
box -48 -56 528 834
use sg13g2_nand2b_1  _0855_
timestamp 1676567195
transform 1 0 17376 0 1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  _0856_
timestamp 1685175443
transform 1 0 18336 0 -1 23436
box -48 -56 538 834
use sg13g2_o21ai_1  _0857_
timestamp 1685175443
transform 1 0 19584 0 -1 23436
box -48 -56 538 834
use sg13g2_nand2b_1  _0858_
timestamp 1676567195
transform 1 0 19680 0 1 26460
box -48 -56 528 834
use sg13g2_nand2b_1  _0859_
timestamp 1676567195
transform 1 0 19680 0 -1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  _0860_
timestamp 1685175443
transform 1 0 19200 0 1 26460
box -48 -56 538 834
use sg13g2_mux4_1  _0861_
timestamp 1677257233
transform 1 0 17184 0 1 26460
box -48 -56 2064 834
use sg13g2_nand2b_1  _0862_
timestamp 1676567195
transform -1 0 19680 0 -1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  _0863_
timestamp 1685175443
transform 1 0 19776 0 1 27972
box -48 -56 538 834
use sg13g2_mux4_1  _0864_
timestamp 1677257233
transform 1 0 8448 0 -1 27972
box -48 -56 2064 834
use sg13g2_nand2b_1  _0865_
timestamp 1676567195
transform 1 0 11040 0 -1 29484
box -48 -56 528 834
use sg13g2_nand2b_1  _0866_
timestamp 1676567195
transform 1 0 10464 0 1 26460
box -48 -56 528 834
use sg13g2_nand2b_1  _0867_
timestamp 1676567195
transform 1 0 10944 0 1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  _0868_
timestamp 1685175443
transform 1 0 9984 0 1 26460
box -48 -56 538 834
use sg13g2_o21ai_1  _0869_
timestamp 1685175443
transform 1 0 11424 0 1 27972
box -48 -56 538 834
use sg13g2_nor2b_1  _0870_
timestamp 1685181386
transform 1 0 10752 0 -1 35532
box -54 -56 528 834
use sg13g2_nor2_1  _0871_
timestamp 1676627187
transform -1 0 14496 0 1 34020
box -48 -56 432 834
use sg13g2_a21oi_1  _0872_
timestamp 1683973020
transform 1 0 11520 0 -1 34020
box -48 -56 528 834
use sg13g2_mux2_1  _0873_
timestamp 1677247768
transform 1 0 12384 0 1 34020
box -48 -56 1008 834
use sg13g2_nor3_1  _0874_
timestamp 1676639442
transform 1 0 12576 0 -1 34020
box -48 -56 528 834
use sg13g2_mux4_1  _0875_
timestamp 1677257233
transform 1 0 10368 0 1 34020
box -48 -56 2064 834
use sg13g2_inv_1  _0876_
timestamp 1676382929
transform 1 0 12288 0 -1 34020
box -48 -56 336 834
use sg13g2_a221oi_1  _0877_
timestamp 1685197497
transform 1 0 13344 0 1 34020
box -48 -56 816 834
use sg13g2_nor3_1  _0878_
timestamp 1676639442
transform -1 0 13632 0 1 35532
box -48 -56 528 834
use sg13g2_mux2_1  _0879_
timestamp 1677247768
transform 1 0 11232 0 -1 35532
box -48 -56 1008 834
use sg13g2_o21ai_1  _0880_
timestamp 1685175443
transform 1 0 12864 0 -1 35532
box -48 -56 538 834
use sg13g2_nand2b_1  _0881_
timestamp 1676567195
transform 1 0 13344 0 -1 35532
box -48 -56 528 834
use sg13g2_a22oi_1  _0882_
timestamp 1685173987
transform 1 0 13056 0 -1 34020
box -48 -56 624 834
use sg13g2_nor3_1  _0883_
timestamp 1676639442
transform 1 0 13632 0 -1 34020
box -48 -56 528 834
use sg13g2_nor3_1  _0884_
timestamp 1676639442
transform 1 0 13152 0 1 32508
box -48 -56 528 834
use sg13g2_nor2b_1  _0885_
timestamp 1685181386
transform -1 0 14592 0 -1 34020
box -54 -56 528 834
use sg13g2_o21ai_1  _0886_
timestamp 1685175443
transform 1 0 13632 0 1 35532
box -48 -56 538 834
use sg13g2_o21ai_1  _0887_
timestamp 1685175443
transform 1 0 14112 0 1 35532
box -48 -56 538 834
use sg13g2_inv_1  _0888_
timestamp 1676382929
transform 1 0 19680 0 1 34020
box -48 -56 336 834
use sg13g2_nor2b_1  _0889_
timestamp 1685181386
transform -1 0 12672 0 1 35532
box -54 -56 528 834
use sg13g2_nor2b_1  _0890_
timestamp 1685181386
transform -1 0 12960 0 1 37044
box -54 -56 528 834
use sg13g2_nor2b_1  _0891_
timestamp 1685181386
transform 1 0 11232 0 1 35532
box -54 -56 528 834
use sg13g2_nand2_1  _0892_
timestamp 1676557249
transform 1 0 10368 0 -1 35532
box -48 -56 432 834
use sg13g2_nand3_1  _0893_
timestamp 1683988354
transform 1 0 11712 0 1 35532
box -48 -56 528 834
use sg13g2_mux2_1  _0894_
timestamp 1677247768
transform 1 0 11136 0 -1 37044
box -48 -56 1008 834
use sg13g2_nor3_1  _0895_
timestamp 1676639442
transform 1 0 11520 0 1 37044
box -48 -56 528 834
use sg13g2_nor2b_1  _0896_
timestamp 1685181386
transform 1 0 10656 0 1 35532
box -54 -56 528 834
use sg13g2_a21oi_1  _0897_
timestamp 1683973020
transform 1 0 11040 0 1 37044
box -48 -56 528 834
use sg13g2_nor2b_1  _0898_
timestamp 1685181386
transform 1 0 10176 0 1 35532
box -54 -56 528 834
use sg13g2_a21oi_1  _0899_
timestamp 1683973020
transform -1 0 10656 0 -1 37044
box -48 -56 528 834
use sg13g2_a221oi_1  _0900_
timestamp 1685197497
transform 1 0 12096 0 -1 37044
box -48 -56 816 834
use sg13g2_o21ai_1  _0901_
timestamp 1685175443
transform 1 0 12192 0 -1 35532
box -48 -56 538 834
use sg13g2_nand2b_1  _0902_
timestamp 1676567195
transform 1 0 12672 0 1 35532
box -48 -56 528 834
use sg13g2_nor3_1  _0903_
timestamp 1676639442
transform 1 0 10656 0 -1 37044
box -48 -56 528 834
use sg13g2_a21oi_1  _0904_
timestamp 1683973020
transform 1 0 12000 0 1 37044
box -48 -56 528 834
use sg13g2_nand3_1  _0905_
timestamp 1683988354
transform 1 0 12960 0 1 37044
box -48 -56 528 834
use sg13g2_nor3_1  _0906_
timestamp 1676639442
transform 1 0 12576 0 -1 40068
box -48 -56 528 834
use sg13g2_o21ai_1  _0907_
timestamp 1685175443
transform -1 0 14208 0 -1 37044
box -48 -56 538 834
use sg13g2_nor2b_1  _0908_
timestamp 1685181386
transform 1 0 13056 0 1 38556
box -54 -56 528 834
use sg13g2_nor3_1  _0909_
timestamp 1676639442
transform 1 0 13056 0 -1 38556
box -48 -56 528 834
use sg13g2_a21oi_1  _0910_
timestamp 1683973020
transform -1 0 14016 0 -1 38556
box -48 -56 528 834
use sg13g2_a22oi_1  _0911_
timestamp 1685173987
transform -1 0 13728 0 -1 37044
box -48 -56 624 834
use sg13g2_dlhq_1  _0912_
timestamp 1678805552
transform 1 0 5664 0 -1 74844
box -50 -56 1692 834
use sg13g2_dlhq_1  _0913_
timestamp 1678805552
transform 1 0 6144 0 1 74844
box -50 -56 1692 834
use sg13g2_dlhq_1  _0914_
timestamp 1678805552
transform 1 0 16416 0 1 62748
box -50 -56 1692 834
use sg13g2_dlhq_1  _0915_
timestamp 1678805552
transform 1 0 16416 0 -1 62748
box -50 -56 1692 834
use sg13g2_dlhq_1  _0916_
timestamp 1678805552
transform 1 0 11232 0 -1 59724
box -50 -56 1692 834
use sg13g2_dlhq_1  _0917_
timestamp 1678805552
transform 1 0 11040 0 1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _0918_
timestamp 1678805552
transform 1 0 5280 0 -1 61236
box -50 -56 1692 834
use sg13g2_dlhq_1  _0919_
timestamp 1678805552
transform 1 0 5280 0 1 59724
box -50 -56 1692 834
use sg13g2_dlhq_1  _0920_
timestamp 1678805552
transform 1 0 4032 0 1 82404
box -50 -56 1692 834
use sg13g2_dlhq_1  _0921_
timestamp 1678805552
transform 1 0 6048 0 1 80892
box -50 -56 1692 834
use sg13g2_dlhq_1  _0922_
timestamp 1678805552
transform 1 0 10656 0 1 70308
box -50 -56 1692 834
use sg13g2_dlhq_1  _0923_
timestamp 1678805552
transform 1 0 11904 0 1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _0924_
timestamp 1678805552
transform 1 0 9024 0 1 74844
box -50 -56 1692 834
use sg13g2_dlhq_1  _0925_
timestamp 1678805552
transform 1 0 11232 0 -1 74844
box -50 -56 1692 834
use sg13g2_dlhq_1  _0926_
timestamp 1678805552
transform 1 0 3168 0 -1 43092
box -50 -56 1692 834
use sg13g2_dlhq_1  _0927_
timestamp 1678805552
transform 1 0 5184 0 1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _0928_
timestamp 1678805552
transform 1 0 1824 0 1 82404
box -50 -56 1692 834
use sg13g2_dlhq_1  _0929_
timestamp 1678805552
transform 1 0 3648 0 -1 82404
box -50 -56 1692 834
use sg13g2_dlhq_1  _0930_
timestamp 1678805552
transform 1 0 10848 0 -1 73332
box -50 -56 1692 834
use sg13g2_dlhq_1  _0931_
timestamp 1678805552
transform 1 0 12096 0 -1 71820
box -50 -56 1692 834
use sg13g2_dlhq_1  _0932_
timestamp 1678805552
transform 1 0 8160 0 -1 70308
box -50 -56 1692 834
use sg13g2_dlhq_1  _0933_
timestamp 1678805552
transform 1 0 9792 0 -1 70308
box -50 -56 1692 834
use sg13g2_dlhq_1  _0934_
timestamp 1678805552
transform 1 0 1152 0 -1 82404
box -50 -56 1692 834
use sg13g2_dlhq_1  _0935_
timestamp 1678805552
transform 1 0 2784 0 1 80892
box -50 -56 1692 834
use sg13g2_dlhq_1  _0936_
timestamp 1678805552
transform -1 0 12576 0 -1 76356
box -50 -56 1692 834
use sg13g2_dlhq_1  _0937_
timestamp 1678805552
transform 1 0 6624 0 1 76356
box -50 -56 1692 834
use sg13g2_dlhq_1  _0938_
timestamp 1678805552
transform 1 0 16704 0 1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _0939_
timestamp 1678805552
transform 1 0 15168 0 -1 56700
box -50 -56 1692 834
use sg13g2_dlhq_1  _0940_
timestamp 1678805552
transform 1 0 13440 0 1 49140
box -50 -56 1692 834
use sg13g2_dlhq_1  _0941_
timestamp 1678805552
transform 1 0 11424 0 -1 49140
box -50 -56 1692 834
use sg13g2_dlhq_1  _0942_
timestamp 1678805552
transform 1 0 5664 0 -1 56700
box -50 -56 1692 834
use sg13g2_dlhq_1  _0943_
timestamp 1678805552
transform 1 0 5376 0 1 56700
box -50 -56 1692 834
use sg13g2_dlhq_1  _0944_
timestamp 1678805552
transform -1 0 11904 0 1 76356
box -50 -56 1692 834
use sg13g2_dlhq_1  _0945_
timestamp 1678805552
transform 1 0 5952 0 -1 77868
box -50 -56 1692 834
use sg13g2_dlhq_1  _0946_
timestamp 1678805552
transform -1 0 20256 0 1 56700
box -50 -56 1692 834
use sg13g2_dlhq_1  _0947_
timestamp 1678805552
transform 1 0 15840 0 -1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _0948_
timestamp 1678805552
transform 1 0 13440 0 -1 52164
box -50 -56 1692 834
use sg13g2_dlhq_1  _0949_
timestamp 1678805552
transform 1 0 11808 0 -1 52164
box -50 -56 1692 834
use sg13g2_dlhq_1  _0950_
timestamp 1678805552
transform 1 0 8256 0 1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _0951_
timestamp 1678805552
transform 1 0 5760 0 -1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _0952_
timestamp 1678805552
transform 1 0 7872 0 1 79380
box -50 -56 1692 834
use sg13g2_dlhq_1  _0953_
timestamp 1678805552
transform 1 0 6144 0 -1 79380
box -50 -56 1692 834
use sg13g2_dlhq_1  _0954_
timestamp 1678805552
transform 1 0 18144 0 -1 61236
box -50 -56 1692 834
use sg13g2_dlhq_1  _0955_
timestamp 1678805552
transform 1 0 16320 0 -1 61236
box -50 -56 1692 834
use sg13g2_dlhq_1  _0956_
timestamp 1678805552
transform 1 0 12672 0 -1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _0957_
timestamp 1678805552
transform 1 0 11040 0 -1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _0958_
timestamp 1678805552
transform 1 0 6624 0 1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _0959_
timestamp 1678805552
transform 1 0 5376 0 -1 55188
box -50 -56 1692 834
use sg13g2_dlhq_1  _0960_
timestamp 1678805552
transform 1 0 8832 0 -1 79380
box -50 -56 1692 834
use sg13g2_dlhq_1  _0961_
timestamp 1678805552
transform 1 0 6624 0 1 77868
box -50 -56 1692 834
use sg13g2_dlhq_1  _0962_
timestamp 1678805552
transform 1 0 18336 0 1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _0963_
timestamp 1678805552
transform 1 0 15744 0 1 59724
box -50 -56 1692 834
use sg13g2_dlhq_1  _0964_
timestamp 1678805552
transform 1 0 13056 0 1 55188
box -50 -56 1692 834
use sg13g2_dlhq_1  _0965_
timestamp 1678805552
transform 1 0 11232 0 -1 55188
box -50 -56 1692 834
use sg13g2_dlhq_1  _0966_
timestamp 1678805552
transform 1 0 7296 0 1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _0967_
timestamp 1678805552
transform 1 0 5088 0 -1 59724
box -50 -56 1692 834
use sg13g2_dlhq_1  _0968_
timestamp 1678805552
transform 1 0 7680 0 -1 71820
box -50 -56 1692 834
use sg13g2_dlhq_1  _0969_
timestamp 1678805552
transform -1 0 10944 0 -1 71820
box -50 -56 1692 834
use sg13g2_dlhq_1  _0970_
timestamp 1678805552
transform 1 0 6912 0 1 71820
box -50 -56 1692 834
use sg13g2_dlhq_1  _0971_
timestamp 1678805552
transform 1 0 17952 0 -1 67284
box -50 -56 1692 834
use sg13g2_dlhq_1  _0972_
timestamp 1678805552
transform 1 0 18336 0 1 65772
box -50 -56 1692 834
use sg13g2_dlhq_1  _0973_
timestamp 1678805552
transform 1 0 16896 0 -1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _0974_
timestamp 1678805552
transform 1 0 14016 0 1 64260
box -50 -56 1692 834
use sg13g2_dlhq_1  _0975_
timestamp 1678805552
transform -1 0 16416 0 1 62748
box -50 -56 1692 834
use sg13g2_dlhq_1  _0976_
timestamp 1678805552
transform 1 0 13152 0 1 62748
box -50 -56 1692 834
use sg13g2_dlhq_1  _0977_
timestamp 1678805552
transform 1 0 7584 0 1 65772
box -50 -56 1692 834
use sg13g2_dlhq_1  _0978_
timestamp 1678805552
transform -1 0 11040 0 -1 65772
box -50 -56 1692 834
use sg13g2_dlhq_1  _0979_
timestamp 1678805552
transform 1 0 6720 0 -1 67284
box -50 -56 1692 834
use sg13g2_dlhq_1  _0980_
timestamp 1678805552
transform 1 0 4512 0 1 71820
box -50 -56 1692 834
use sg13g2_dlhq_1  _0981_
timestamp 1678805552
transform 1 0 5856 0 -1 71820
box -50 -56 1692 834
use sg13g2_dlhq_1  _0982_
timestamp 1678805552
transform 1 0 4416 0 -1 73332
box -50 -56 1692 834
use sg13g2_dlhq_1  _0983_
timestamp 1678805552
transform 1 0 15264 0 -1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _0984_
timestamp 1678805552
transform 1 0 15552 0 -1 67284
box -50 -56 1692 834
use sg13g2_dlhq_1  _0985_
timestamp 1678805552
transform 1 0 13632 0 -1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _0986_
timestamp 1678805552
transform 1 0 12000 0 1 67284
box -50 -56 1692 834
use sg13g2_dlhq_1  _0987_
timestamp 1678805552
transform -1 0 15552 0 -1 67284
box -50 -56 1692 834
use sg13g2_dlhq_1  _0988_
timestamp 1678805552
transform 1 0 11424 0 -1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _0989_
timestamp 1678805552
transform -1 0 6048 0 -1 70308
box -50 -56 1692 834
use sg13g2_dlhq_1  _0990_
timestamp 1678805552
transform 1 0 5856 0 1 67284
box -50 -56 1692 834
use sg13g2_dlhq_1  _0991_
timestamp 1678805552
transform -1 0 7008 0 1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _0992_
timestamp 1678805552
transform 1 0 1632 0 -1 62748
box -50 -56 1692 834
use sg13g2_dlhq_1  _0993_
timestamp 1678805552
transform 1 0 3648 0 1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _0994_
timestamp 1678805552
transform 1 0 9792 0 1 56700
box -50 -56 1692 834
use sg13g2_dlhq_1  _0995_
timestamp 1678805552
transform 1 0 11616 0 -1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _0996_
timestamp 1678805552
transform 1 0 13728 0 1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _0997_
timestamp 1678805552
transform 1 0 15456 0 1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _0998_
timestamp 1678805552
transform 1 0 5760 0 1 49140
box -50 -56 1692 834
use sg13g2_dlhq_1  _0999_
timestamp 1678805552
transform 1 0 7488 0 -1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _1000_
timestamp 1678805552
transform 1 0 3360 0 1 55188
box -50 -56 1692 834
use sg13g2_dlhq_1  _1001_
timestamp 1678805552
transform 1 0 1344 0 -1 56700
box -50 -56 1692 834
use sg13g2_dlhq_1  _1002_
timestamp 1678805552
transform 1 0 10656 0 -1 56700
box -50 -56 1692 834
use sg13g2_dlhq_1  _1003_
timestamp 1678805552
transform 1 0 9504 0 -1 55188
box -50 -56 1692 834
use sg13g2_dlhq_1  _1004_
timestamp 1678805552
transform -1 0 18816 0 1 49140
box -50 -56 1692 834
use sg13g2_dlhq_1  _1005_
timestamp 1678805552
transform 1 0 17856 0 1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _1006_
timestamp 1678805552
transform 1 0 3360 0 -1 49140
box -50 -56 1692 834
use sg13g2_dlhq_1  _1007_
timestamp 1678805552
transform 1 0 4992 0 -1 49140
box -50 -56 1692 834
use sg13g2_dlhq_1  _1008_
timestamp 1678805552
transform 1 0 8928 0 1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _1009_
timestamp 1678805552
transform 1 0 6720 0 -1 59724
box -50 -56 1692 834
use sg13g2_dlhq_1  _1010_
timestamp 1678805552
transform 1 0 14016 0 1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _1011_
timestamp 1678805552
transform -1 0 14880 0 -1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _1012_
timestamp 1678805552
transform 1 0 14976 0 1 55188
box -50 -56 1692 834
use sg13g2_dlhq_1  _1013_
timestamp 1678805552
transform 1 0 13152 0 -1 56700
box -50 -56 1692 834
use sg13g2_dlhq_1  _1014_
timestamp 1678805552
transform 1 0 7872 0 -1 55188
box -50 -56 1692 834
use sg13g2_dlhq_1  _1015_
timestamp 1678805552
transform 1 0 6240 0 -1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _1016_
timestamp 1678805552
transform 1 0 2112 0 1 56700
box -50 -56 1692 834
use sg13g2_dlhq_1  _1017_
timestamp 1678805552
transform 1 0 1344 0 1 59724
box -50 -56 1692 834
use sg13g2_dlhq_1  _1018_
timestamp 1678805552
transform 1 0 17760 0 1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _1019_
timestamp 1678805552
transform -1 0 18240 0 1 55188
box -50 -56 1692 834
use sg13g2_dlhq_1  _1020_
timestamp 1678805552
transform 1 0 16128 0 1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _1021_
timestamp 1678805552
transform 1 0 14496 0 1 52164
box -50 -56 1692 834
use sg13g2_dlhq_1  _1022_
timestamp 1678805552
transform 1 0 5856 0 -1 52164
box -50 -56 1692 834
use sg13g2_dlhq_1  _1023_
timestamp 1678805552
transform 1 0 3744 0 1 52164
box -50 -56 1692 834
use sg13g2_dlhq_1  _1024_
timestamp 1678805552
transform 1 0 1440 0 -1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _1025_
timestamp 1678805552
transform 1 0 1344 0 1 55188
box -50 -56 1692 834
use sg13g2_dlhq_1  _1026_
timestamp 1678805552
transform 1 0 10272 0 1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _1027_
timestamp 1678805552
transform 1 0 9408 0 -1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _1028_
timestamp 1678805552
transform 1 0 18144 0 1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _1029_
timestamp 1678805552
transform 1 0 16512 0 1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _1030_
timestamp 1678805552
transform -1 0 9600 0 -1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _1031_
timestamp 1678805552
transform 1 0 6720 0 -1 49140
box -50 -56 1692 834
use sg13g2_dlhq_1  _1032_
timestamp 1678805552
transform -1 0 3744 0 1 52164
box -50 -56 1692 834
use sg13g2_dlhq_1  _1033_
timestamp 1678805552
transform 1 0 1152 0 1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _1034_
timestamp 1678805552
transform 1 0 10176 0 -1 52164
box -50 -56 1692 834
use sg13g2_dlhq_1  _1035_
timestamp 1678805552
transform 1 0 8544 0 -1 52164
box -50 -56 1692 834
use sg13g2_dlhq_1  _1036_
timestamp 1678805552
transform 1 0 15552 0 -1 49140
box -50 -56 1692 834
use sg13g2_dlhq_1  _1037_
timestamp 1678805552
transform 1 0 13920 0 -1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _1038_
timestamp 1678805552
transform 1 0 4416 0 1 46116
box -50 -56 1692 834
use sg13g2_dlhq_1  _1039_
timestamp 1678805552
transform 1 0 3552 0 1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _1040_
timestamp 1678805552
transform 1 0 5280 0 1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _1041_
timestamp 1678805552
transform 1 0 3744 0 1 56700
box -50 -56 1692 834
use sg13g2_dlhq_1  _1042_
timestamp 1678805552
transform 1 0 11520 0 -1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _1043_
timestamp 1678805552
transform 1 0 9792 0 1 49140
box -50 -56 1692 834
use sg13g2_dlhq_1  _1044_
timestamp 1678805552
transform 1 0 18432 0 -1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _1045_
timestamp 1678805552
transform 1 0 17376 0 1 52164
box -50 -56 1692 834
use sg13g2_dlhq_1  _1046_
timestamp 1678805552
transform 1 0 2976 0 -1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _1047_
timestamp 1678805552
transform 1 0 3264 0 1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _1048_
timestamp 1678805552
transform 1 0 1344 0 -1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _1049_
timestamp 1678805552
transform 1 0 1152 0 1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _1050_
timestamp 1678805552
transform 1 0 12000 0 1 44604
box -50 -56 1692 834
use sg13g2_dlhq_1  _1051_
timestamp 1678805552
transform 1 0 9984 0 -1 44604
box -50 -56 1692 834
use sg13g2_dlhq_1  _1052_
timestamp 1678805552
transform 1 0 15168 0 1 46116
box -50 -56 1692 834
use sg13g2_dlhq_1  _1053_
timestamp 1678805552
transform 1 0 13536 0 1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _1054_
timestamp 1678805552
transform -1 0 3744 0 -1 44604
box -50 -56 1692 834
use sg13g2_dlhq_1  _1055_
timestamp 1678805552
transform 1 0 1152 0 -1 43092
box -50 -56 1692 834
use sg13g2_dlhq_1  _1056_
timestamp 1678805552
transform 1 0 1920 0 1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _1057_
timestamp 1678805552
transform 1 0 1152 0 -1 49140
box -50 -56 1692 834
use sg13g2_dlhq_1  _1058_
timestamp 1678805552
transform 1 0 9504 0 1 44604
box -50 -56 1692 834
use sg13g2_dlhq_1  _1059_
timestamp 1678805552
transform 1 0 7872 0 1 44604
box -50 -56 1692 834
use sg13g2_dlhq_1  _1060_
timestamp 1678805552
transform 1 0 18048 0 -1 44604
box -50 -56 1692 834
use sg13g2_dlhq_1  _1061_
timestamp 1678805552
transform 1 0 16992 0 -1 46116
box -50 -56 1692 834
use sg13g2_dlhq_1  _1062_
timestamp 1678805552
transform 1 0 6240 0 -1 46116
box -50 -56 1692 834
use sg13g2_dlhq_1  _1063_
timestamp 1678805552
transform 1 0 4032 0 -1 46116
box -50 -56 1692 834
use sg13g2_dlhq_1  _1064_
timestamp 1678805552
transform -1 0 4032 0 -1 46116
box -50 -56 1692 834
use sg13g2_dlhq_1  _1065_
timestamp 1678805552
transform 1 0 1152 0 1 46116
box -50 -56 1692 834
use sg13g2_dlhq_1  _1066_
timestamp 1678805552
transform 1 0 12288 0 -1 43092
box -50 -56 1692 834
use sg13g2_dlhq_1  _1067_
timestamp 1678805552
transform 1 0 9888 0 1 43092
box -50 -56 1692 834
use sg13g2_dlhq_1  _1068_
timestamp 1678805552
transform 1 0 15168 0 1 44604
box -50 -56 1692 834
use sg13g2_dlhq_1  _1069_
timestamp 1678805552
transform 1 0 13344 0 -1 46116
box -50 -56 1692 834
use sg13g2_dlhq_1  _1070_
timestamp 1678805552
transform 1 0 1824 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1071_
timestamp 1678805552
transform 1 0 1152 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1072_
timestamp 1678805552
transform -1 0 3456 0 -1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _1073_
timestamp 1678805552
transform 1 0 1152 0 1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _1074_
timestamp 1678805552
transform 1 0 10176 0 1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _1075_
timestamp 1678805552
transform 1 0 8064 0 1 46116
box -50 -56 1692 834
use sg13g2_dlhq_1  _1076_
timestamp 1678805552
transform 1 0 18528 0 -1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _1077_
timestamp 1678805552
transform 1 0 16896 0 -1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _1078_
timestamp 1678805552
transform 1 0 6048 0 1 46116
box -50 -56 1692 834
use sg13g2_dlhq_1  _1079_
timestamp 1678805552
transform 1 0 3744 0 -1 44604
box -50 -56 1692 834
use sg13g2_dlhq_1  _1080_
timestamp 1678805552
transform 1 0 7392 0 1 49140
box -50 -56 1692 834
use sg13g2_dlhq_1  _1081_
timestamp 1678805552
transform 1 0 9120 0 -1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _1082_
timestamp 1678805552
transform 1 0 13920 0 -1 44604
box -50 -56 1692 834
use sg13g2_dlhq_1  _1083_
timestamp 1678805552
transform 1 0 15744 0 1 43092
box -50 -56 1692 834
use sg13g2_dlhq_1  _1084_
timestamp 1678805552
transform 1 0 11040 0 -1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _1085_
timestamp 1678805552
transform 1 0 12672 0 -1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _1086_
timestamp 1678805552
transform 1 0 6144 0 1 43092
box -50 -56 1692 834
use sg13g2_dlhq_1  _1087_
timestamp 1678805552
transform 1 0 8064 0 -1 43092
box -50 -56 1692 834
use sg13g2_dlhq_1  _1088_
timestamp 1678805552
transform 1 0 8160 0 1 73332
box -50 -56 1692 834
use sg13g2_dlhq_1  _1089_
timestamp 1678805552
transform -1 0 12384 0 1 73332
box -50 -56 1692 834
use sg13g2_dlhq_1  _1090_
timestamp 1678805552
transform 1 0 6720 0 -1 73332
box -50 -56 1692 834
use sg13g2_dlhq_1  _1091_
timestamp 1678805552
transform 1 0 17472 0 -1 71820
box -50 -56 1692 834
use sg13g2_dlhq_1  _1092_
timestamp 1678805552
transform 1 0 17568 0 1 70308
box -50 -56 1692 834
use sg13g2_dlhq_1  _1093_
timestamp 1678805552
transform 1 0 16320 0 1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _1094_
timestamp 1678805552
transform -1 0 17280 0 1 61236
box -50 -56 1692 834
use sg13g2_dlhq_1  _1095_
timestamp 1678805552
transform -1 0 16128 0 -1 59724
box -50 -56 1692 834
use sg13g2_dlhq_1  _1096_
timestamp 1678805552
transform -1 0 15744 0 1 59724
box -50 -56 1692 834
use sg13g2_dlhq_1  _1097_
timestamp 1678805552
transform 1 0 7392 0 -1 62748
box -50 -56 1692 834
use sg13g2_dlhq_1  _1098_
timestamp 1678805552
transform 1 0 8736 0 -1 64260
box -50 -56 1692 834
use sg13g2_dlhq_1  _1099_
timestamp 1678805552
transform 1 0 5856 0 1 62748
box -50 -56 1692 834
use sg13g2_dlhq_1  _1100_
timestamp 1678805552
transform 1 0 3456 0 1 64260
box -50 -56 1692 834
use sg13g2_dlhq_1  _1101_
timestamp 1678805552
transform 1 0 1152 0 1 65772
box -50 -56 1692 834
use sg13g2_dlhq_1  _1102_
timestamp 1678805552
transform 1 0 9408 0 -1 59724
box -50 -56 1692 834
use sg13g2_dlhq_1  _1103_
timestamp 1678805552
transform 1 0 7392 0 1 59724
box -50 -56 1692 834
use sg13g2_dlhq_1  _1104_
timestamp 1678805552
transform 1 0 2976 0 1 59724
box -50 -56 1692 834
use sg13g2_dlhq_1  _1105_
timestamp 1678805552
transform 1 0 1152 0 1 64260
box -50 -56 1692 834
use sg13g2_dlhq_1  _1106_
timestamp 1678805552
transform 1 0 1152 0 -1 70308
box -50 -56 1692 834
use sg13g2_dlhq_1  _1107_
timestamp 1678805552
transform 1 0 3456 0 -1 67284
box -50 -56 1692 834
use sg13g2_dlhq_1  _1108_
timestamp 1678805552
transform 1 0 2016 0 1 76356
box -50 -56 1692 834
use sg13g2_dlhq_1  _1109_
timestamp 1678805552
transform 1 0 1152 0 1 77868
box -50 -56 1692 834
use sg13g2_dlhq_1  _1110_
timestamp 1678805552
transform 1 0 10176 0 -1 67284
box -50 -56 1692 834
use sg13g2_dlhq_1  _1111_
timestamp 1678805552
transform 1 0 7776 0 1 67284
box -50 -56 1692 834
use sg13g2_dlhq_1  _1112_
timestamp 1678805552
transform 1 0 2784 0 -1 71820
box -50 -56 1692 834
use sg13g2_dlhq_1  _1113_
timestamp 1678805552
transform 1 0 1152 0 -1 73332
box -50 -56 1692 834
use sg13g2_dlhq_1  _1114_
timestamp 1678805552
transform -1 0 4416 0 -1 70308
box -50 -56 1692 834
use sg13g2_dlhq_1  _1115_
timestamp 1678805552
transform 1 0 1152 0 -1 71820
box -50 -56 1692 834
use sg13g2_dlhq_1  _1116_
timestamp 1678805552
transform 1 0 4320 0 1 76356
box -50 -56 1692 834
use sg13g2_dlhq_1  _1117_
timestamp 1678805552
transform 1 0 3264 0 1 77868
box -50 -56 1692 834
use sg13g2_dlhq_1  _1118_
timestamp 1678805552
transform 1 0 16128 0 1 64260
box -50 -56 1692 834
use sg13g2_dlhq_1  _1119_
timestamp 1678805552
transform 1 0 14400 0 -1 65772
box -50 -56 1692 834
use sg13g2_dlhq_1  _1120_
timestamp 1678805552
transform 1 0 12864 0 -1 59724
box -50 -56 1692 834
use sg13g2_dlhq_1  _1121_
timestamp 1678805552
transform 1 0 11040 0 -1 61236
box -50 -56 1692 834
use sg13g2_dlhq_1  _1122_
timestamp 1678805552
transform 1 0 4128 0 -1 62748
box -50 -56 1692 834
use sg13g2_dlhq_1  _1123_
timestamp 1678805552
transform 1 0 5760 0 -1 62748
box -50 -56 1692 834
use sg13g2_dlhq_1  _1124_
timestamp 1678805552
transform 1 0 4416 0 1 80892
box -50 -56 1692 834
use sg13g2_dlhq_1  _1125_
timestamp 1678805552
transform 1 0 5472 0 1 79380
box -50 -56 1692 834
use sg13g2_dlhq_1  _1126_
timestamp 1678805552
transform 1 0 3648 0 -1 80892
box -50 -56 1692 834
use sg13g2_dlhq_1  _1127_
timestamp 1678805552
transform 1 0 13632 0 1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _1128_
timestamp 1678805552
transform 1 0 13728 0 -1 71820
box -50 -56 1692 834
use sg13g2_dlhq_1  _1129_
timestamp 1678805552
transform 1 0 12960 0 1 70308
box -50 -56 1692 834
use sg13g2_dlhq_1  _1130_
timestamp 1678805552
transform 1 0 10752 0 -1 64260
box -50 -56 1692 834
use sg13g2_dlhq_1  _1131_
timestamp 1678805552
transform 1 0 11040 0 -1 65772
box -50 -56 1692 834
use sg13g2_dlhq_1  _1132_
timestamp 1678805552
transform 1 0 9504 0 1 64260
box -50 -56 1692 834
use sg13g2_dlhq_1  _1133_
timestamp 1678805552
transform -1 0 5856 0 1 67284
box -50 -56 1692 834
use sg13g2_dlhq_1  _1134_
timestamp 1678805552
transform -1 0 6720 0 -1 67284
box -50 -56 1692 834
use sg13g2_dlhq_1  _1135_
timestamp 1678805552
transform -1 0 5376 0 1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _1136_
timestamp 1678805552
transform 1 0 1632 0 -1 67284
box -50 -56 1692 834
use sg13g2_dlhq_1  _1137_
timestamp 1678805552
transform -1 0 9120 0 1 61236
box -50 -56 1692 834
use sg13g2_dlhq_1  _1138_
timestamp 1678805552
transform 1 0 9600 0 1 61236
box -50 -56 1692 834
use sg13g2_dlhq_1  _1139_
timestamp 1678805552
transform 1 0 7392 0 -1 61236
box -50 -56 1692 834
use sg13g2_dlhq_1  _1140_
timestamp 1678805552
transform 1 0 2784 0 -1 74844
box -50 -56 1692 834
use sg13g2_dlhq_1  _1141_
timestamp 1678805552
transform 1 0 1152 0 1 74844
box -50 -56 1692 834
use sg13g2_dlhq_1  _1142_
timestamp 1678805552
transform 1 0 2304 0 -1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _1143_
timestamp 1678805552
transform -1 0 8736 0 1 64260
box -50 -56 1692 834
use sg13g2_dlhq_1  _1144_
timestamp 1678805552
transform 1 0 1824 0 -1 79380
box -50 -56 1692 834
use sg13g2_dlhq_1  _1145_
timestamp 1678805552
transform -1 0 2784 0 1 79380
box -50 -56 1692 834
use sg13g2_dlhq_1  _1146_
timestamp 1678805552
transform 1 0 8160 0 1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _1147_
timestamp 1678805552
transform 1 0 6816 0 -1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _1148_
timestamp 1678805552
transform -1 0 4416 0 -1 73332
box -50 -56 1692 834
use sg13g2_dlhq_1  _1149_
timestamp 1678805552
transform -1 0 2784 0 -1 74844
box -50 -56 1692 834
use sg13g2_dlhq_1  _1150_
timestamp 1678805552
transform 1 0 1536 0 -1 80892
box -50 -56 1692 834
use sg13g2_dlhq_1  _1151_
timestamp 1678805552
transform -1 0 2784 0 1 80892
box -50 -56 1692 834
use sg13g2_dlhq_1  _1152_
timestamp 1678805552
transform 1 0 4128 0 -1 79380
box -50 -56 1692 834
use sg13g2_dlhq_1  _1153_
timestamp 1678805552
transform -1 0 6528 0 1 77868
box -50 -56 1692 834
use sg13g2_dlhq_1  _1154_
timestamp 1678805552
transform 1 0 15840 0 -1 71820
box -50 -56 1692 834
use sg13g2_dlhq_1  _1155_
timestamp 1678805552
transform 1 0 13920 0 1 71820
box -50 -56 1692 834
use sg13g2_dlhq_1  _1156_
timestamp 1678805552
transform 1 0 12096 0 1 61236
box -50 -56 1692 834
use sg13g2_dlhq_1  _1157_
timestamp 1678805552
transform 1 0 10176 0 -1 62748
box -50 -56 1692 834
use sg13g2_dlhq_1  _1158_
timestamp 1678805552
transform 1 0 4224 0 -1 65772
box -50 -56 1692 834
use sg13g2_dlhq_1  _1159_
timestamp 1678805552
transform 1 0 5472 0 1 64260
box -50 -56 1692 834
use sg13g2_dlhq_1  _1160_
timestamp 1678805552
transform 1 0 5184 0 1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1161_
timestamp 1678805552
transform -1 0 9120 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1162_
timestamp 1678805552
transform -1 0 17952 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1163_
timestamp 1678805552
transform 1 0 15840 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1164_
timestamp 1678805552
transform 1 0 13440 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1165_
timestamp 1678805552
transform 1 0 13536 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1166_
timestamp 1678805552
transform 1 0 1152 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1167_
timestamp 1678805552
transform 1 0 1152 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1168_
timestamp 1678805552
transform 1 0 5856 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1169_
timestamp 1678805552
transform 1 0 3552 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1170_
timestamp 1678805552
transform 1 0 10752 0 1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1171_
timestamp 1678805552
transform 1 0 7584 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1172_
timestamp 1678805552
transform 1 0 9120 0 1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1173_
timestamp 1678805552
transform 1 0 7488 0 1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1174_
timestamp 1678805552
transform 1 0 3840 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1175_
timestamp 1678805552
transform 1 0 1920 0 1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1176_
timestamp 1678805552
transform 1 0 2784 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1177_
timestamp 1678805552
transform 1 0 1344 0 -1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1178_
timestamp 1678805552
transform 1 0 11424 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1179_
timestamp 1678805552
transform -1 0 12768 0 -1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1180_
timestamp 1678805552
transform 1 0 8544 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _1181_
timestamp 1678805552
transform 1 0 8064 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _1182_
timestamp 1678805552
transform 1 0 2784 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1183_
timestamp 1678805552
transform 1 0 1440 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1184_
timestamp 1678805552
transform 1 0 8928 0 1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1185_
timestamp 1678805552
transform 1 0 7392 0 -1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1186_
timestamp 1678805552
transform 1 0 16512 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1187_
timestamp 1678805552
transform 1 0 14880 0 1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1188_
timestamp 1678805552
transform 1 0 15360 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _1189_
timestamp 1678805552
transform 1 0 13728 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _1190_
timestamp 1678805552
transform -1 0 9696 0 1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1191_
timestamp 1678805552
transform 1 0 4416 0 1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1192_
timestamp 1678805552
transform 1 0 8448 0 -1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1193_
timestamp 1678805552
transform 1 0 6528 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1194_
timestamp 1678805552
transform 1 0 17664 0 -1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1195_
timestamp 1678805552
transform 1 0 15840 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1196_
timestamp 1678805552
transform 1 0 15360 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1197_
timestamp 1678805552
transform -1 0 16320 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1198_
timestamp 1678805552
transform 1 0 5856 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1199_
timestamp 1678805552
transform 1 0 4032 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1200_
timestamp 1678805552
transform 1 0 7584 0 -1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1201_
timestamp 1678805552
transform 1 0 6816 0 1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1202_
timestamp 1678805552
transform 1 0 17376 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1203_
timestamp 1678805552
transform 1 0 15552 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1204_
timestamp 1678805552
transform 1 0 15744 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1205_
timestamp 1678805552
transform 1 0 14112 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1206_
timestamp 1678805552
transform 1 0 6048 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1207_
timestamp 1678805552
transform 1 0 4800 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1208_
timestamp 1678805552
transform 1 0 8256 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1209_
timestamp 1678805552
transform 1 0 6816 0 -1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1210_
timestamp 1678805552
transform 1 0 17568 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1211_
timestamp 1678805552
transform 1 0 15168 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1212_
timestamp 1678805552
transform 1 0 14784 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _1213_
timestamp 1678805552
transform 1 0 12864 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _1214_
timestamp 1678805552
transform 1 0 5760 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1215_
timestamp 1678805552
transform 1 0 4128 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1216_
timestamp 1678805552
transform 1 0 13536 0 1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1217_
timestamp 1678805552
transform 1 0 11424 0 1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1218_
timestamp 1678805552
transform 1 0 11424 0 -1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1219_
timestamp 1678805552
transform -1 0 12000 0 -1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1220_
timestamp 1678805552
transform -1 0 16224 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1221_
timestamp 1678805552
transform -1 0 16128 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1222_
timestamp 1678805552
transform -1 0 15648 0 -1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1223_
timestamp 1678805552
transform 1 0 9888 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1224_
timestamp 1678805552
transform 1 0 9792 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1225_
timestamp 1678805552
transform 1 0 7968 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1226_
timestamp 1678805552
transform 1 0 8928 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1227_
timestamp 1678805552
transform 1 0 18144 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1228_
timestamp 1678805552
transform -1 0 19200 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1229_
timestamp 1678805552
transform 1 0 18048 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1230_
timestamp 1678805552
transform 1 0 18048 0 1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1231_
timestamp 1678805552
transform -1 0 19584 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1232_
timestamp 1678805552
transform 1 0 16704 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1233_
timestamp 1678805552
transform -1 0 4512 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1234_
timestamp 1678805552
transform 1 0 1152 0 1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1235_
timestamp 1678805552
transform 1 0 3456 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1236_
timestamp 1678805552
transform 1 0 6816 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1237_
timestamp 1678805552
transform 1 0 6048 0 1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1238_
timestamp 1678805552
transform 1 0 4032 0 -1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1239_
timestamp 1678805552
transform -1 0 17568 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1240_
timestamp 1678805552
transform 1 0 14112 0 1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1241_
timestamp 1678805552
transform 1 0 13056 0 1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1242_
timestamp 1678805552
transform 1 0 15264 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1243_
timestamp 1678805552
transform 1 0 13920 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1244_
timestamp 1678805552
transform 1 0 13056 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1245_
timestamp 1678805552
transform -1 0 4416 0 1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1246_
timestamp 1678805552
transform 1 0 1632 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1247_
timestamp 1678805552
transform 1 0 3840 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1248_
timestamp 1678805552
transform 1 0 5760 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1249_
timestamp 1678805552
transform 1 0 6144 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1250_
timestamp 1678805552
transform 1 0 11904 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1251_
timestamp 1678805552
transform 1 0 13536 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1252_
timestamp 1678805552
transform 1 0 13824 0 -1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1253_
timestamp 1678805552
transform 1 0 15936 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1254_
timestamp 1678805552
transform 1 0 5184 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1255_
timestamp 1678805552
transform 1 0 7296 0 -1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1256_
timestamp 1678805552
transform 1 0 2496 0 -1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1257_
timestamp 1678805552
transform 1 0 4128 0 -1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1258_
timestamp 1678805552
transform 1 0 9408 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1259_
timestamp 1678805552
transform 1 0 11136 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1260_
timestamp 1678805552
transform 1 0 11712 0 1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1261_
timestamp 1678805552
transform 1 0 14208 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1262_
timestamp 1678805552
transform 1 0 4032 0 1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1263_
timestamp 1678805552
transform 1 0 5952 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1264_
timestamp 1678805552
transform 1 0 7008 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1265_
timestamp 1678805552
transform 1 0 5088 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1266_
timestamp 1678805552
transform 1 0 12384 0 1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1267_
timestamp 1678805552
transform 1 0 10560 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1268_
timestamp 1678805552
transform -1 0 19392 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1269_
timestamp 1678805552
transform 1 0 14976 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1270_
timestamp 1678805552
transform 1 0 5568 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1271_
timestamp 1678805552
transform 1 0 4224 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1272_
timestamp 1678805552
transform 1 0 2112 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1273_
timestamp 1678805552
transform 1 0 4224 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1274_
timestamp 1678805552
transform 1 0 13056 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1275_
timestamp 1678805552
transform 1 0 11424 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1276_
timestamp 1678805552
transform 1 0 11808 0 -1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1277_
timestamp 1678805552
transform 1 0 13632 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1278_
timestamp 1678805552
transform 1 0 9696 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1279_
timestamp 1678805552
transform 1 0 7776 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1280_
timestamp 1678805552
transform 1 0 4608 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1281_
timestamp 1678805552
transform 1 0 6240 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1282_
timestamp 1678805552
transform -1 0 11904 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1283_
timestamp 1678805552
transform 1 0 9024 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1284_
timestamp 1678805552
transform 1 0 17184 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1285_
timestamp 1678805552
transform -1 0 19680 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1286_
timestamp 1678805552
transform 1 0 8640 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1287_
timestamp 1678805552
transform 1 0 7008 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1288_
timestamp 1678805552
transform 1 0 2784 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1289_
timestamp 1678805552
transform 1 0 4512 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1290_
timestamp 1678805552
transform 1 0 10944 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1291_
timestamp 1678805552
transform 1 0 9120 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1292_
timestamp 1678805552
transform 1 0 11616 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1293_
timestamp 1678805552
transform 1 0 13344 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1294_
timestamp 1678805552
transform 1 0 9696 0 1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1295_
timestamp 1678805552
transform 1 0 7968 0 1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1296_
timestamp 1678805552
transform 1 0 4032 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1297_
timestamp 1678805552
transform 1 0 5184 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1298_
timestamp 1678805552
transform 1 0 12864 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _1299_
timestamp 1678805552
transform 1 0 11232 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _1300_
timestamp 1678805552
transform -1 0 18528 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1301_
timestamp 1678805552
transform 1 0 17664 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1302_
timestamp 1678805552
transform 1 0 3648 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1303_
timestamp 1678805552
transform 1 0 1728 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1304_
timestamp 1678805552
transform 1 0 3072 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _1305_
timestamp 1678805552
transform 1 0 3360 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _1306_
timestamp 1678805552
transform 1 0 5664 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _1307_
timestamp 1678805552
transform 1 0 4704 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _1308_
timestamp 1678805552
transform 1 0 10560 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _1309_
timestamp 1678805552
transform 1 0 10656 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _1310_
timestamp 1678805552
transform 1 0 3456 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1311_
timestamp 1678805552
transform 1 0 3552 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1312_
timestamp 1678805552
transform 1 0 1728 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1313_
timestamp 1678805552
transform 1 0 2016 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1314_
timestamp 1678805552
transform -1 0 9888 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1315_
timestamp 1678805552
transform -1 0 9984 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1316_
timestamp 1678805552
transform 1 0 3456 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _1317_
timestamp 1678805552
transform 1 0 3552 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _1318_
timestamp 1678805552
transform 1 0 1344 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _1319_
timestamp 1678805552
transform 1 0 1344 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _1320_
timestamp 1678805552
transform 1 0 1152 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1321_
timestamp 1678805552
transform 1 0 1152 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1322_
timestamp 1678805552
transform 1 0 6240 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _1323_
timestamp 1678805552
transform 1 0 6336 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _1324_
timestamp 1678805552
transform 1 0 9120 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1325_
timestamp 1678805552
transform -1 0 10752 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1326_
timestamp 1678805552
transform 1 0 1728 0 1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1327_
timestamp 1678805552
transform 1 0 1728 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1328_
timestamp 1678805552
transform 1 0 1440 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1329_
timestamp 1678805552
transform 1 0 1536 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1330_
timestamp 1678805552
transform 1 0 8352 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _1331_
timestamp 1678805552
transform 1 0 8448 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _1332_
timestamp 1678805552
transform 1 0 3456 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _1333_
timestamp 1678805552
transform 1 0 3552 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _1334_
timestamp 1678805552
transform 1 0 1152 0 1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1335_
timestamp 1678805552
transform 1 0 1152 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1336_
timestamp 1678805552
transform 1 0 4800 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1337_
timestamp 1678805552
transform 1 0 6912 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1338_
timestamp 1678805552
transform 1 0 15456 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _1339_
timestamp 1678805552
transform 1 0 17088 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1340_
timestamp 1678805552
transform 1 0 11040 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _1341_
timestamp 1678805552
transform 1 0 12864 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _1342_
timestamp 1678805552
transform 1 0 5664 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1343_
timestamp 1678805552
transform 1 0 7296 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1344_
timestamp 1678805552
transform -1 0 10656 0 -1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1345_
timestamp 1678805552
transform 1 0 9312 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1346_
timestamp 1678805552
transform 1 0 7008 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1347_
timestamp 1678805552
transform 1 0 18240 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1348_
timestamp 1678805552
transform 1 0 18144 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1349_
timestamp 1678805552
transform 1 0 16416 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1350_
timestamp 1678805552
transform 1 0 15552 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1351_
timestamp 1678805552
transform -1 0 19104 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1352_
timestamp 1678805552
transform 1 0 14304 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1353_
timestamp 1678805552
transform 1 0 7200 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1354_
timestamp 1678805552
transform 1 0 5568 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1355_
timestamp 1678805552
transform 1 0 3936 0 1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1356_
timestamp 1678805552
transform 1 0 7200 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1357_
timestamp 1678805552
transform 1 0 8832 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1358_
timestamp 1678805552
transform 1 0 9216 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1359_
timestamp 1678805552
transform 1 0 11424 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1360_
timestamp 1678805552
transform 1 0 7584 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1361_
timestamp 1678805552
transform -1 0 12864 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1362_
timestamp 1678805552
transform 1 0 5472 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1363_
timestamp 1678805552
transform 1 0 7392 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1364_
timestamp 1678805552
transform 1 0 2400 0 -1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1365_
timestamp 1678805552
transform 1 0 1152 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1366_
timestamp 1678805552
transform 1 0 11904 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1367_
timestamp 1678805552
transform 1 0 10848 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1368_
timestamp 1678805552
transform 1 0 9504 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1369_
timestamp 1678805552
transform 1 0 7488 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1370_
timestamp 1678805552
transform 1 0 1248 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1371_
timestamp 1678805552
transform 1 0 1152 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1372_
timestamp 1678805552
transform 1 0 5760 0 -1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1373_
timestamp 1678805552
transform 1 0 4224 0 1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1374_
timestamp 1678805552
transform 1 0 14400 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1375_
timestamp 1678805552
transform 1 0 12960 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1376_
timestamp 1678805552
transform 1 0 13728 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1377_
timestamp 1678805552
transform 1 0 12672 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1378_
timestamp 1678805552
transform 1 0 2880 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1379_
timestamp 1678805552
transform 1 0 2304 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1380_
timestamp 1678805552
transform 1 0 4896 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1381_
timestamp 1678805552
transform 1 0 4128 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1382_
timestamp 1678805552
transform 1 0 4416 0 -1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1383_
timestamp 1678805552
transform 1 0 13920 0 1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1384_
timestamp 1678805552
transform 1 0 13152 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1385_
timestamp 1678805552
transform 1 0 13440 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1386_
timestamp 1678805552
transform -1 0 12768 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1387_
timestamp 1678805552
transform 1 0 9984 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1388_
timestamp 1678805552
transform 1 0 11328 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1389_
timestamp 1678805552
transform 1 0 4416 0 1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1390_
timestamp 1678805552
transform 1 0 2400 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1391_
timestamp 1678805552
transform 1 0 3360 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1392_
timestamp 1678805552
transform 1 0 2784 0 -1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1393_
timestamp 1678805552
transform 1 0 1152 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1394_
timestamp 1678805552
transform 1 0 11136 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1395_
timestamp 1678805552
transform 1 0 9024 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1396_
timestamp 1678805552
transform 1 0 9696 0 1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1397_
timestamp 1678805552
transform 1 0 7680 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1398_
timestamp 1678805552
transform 1 0 1536 0 -1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1399_
timestamp 1678805552
transform 1 0 1152 0 -1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1400_
timestamp 1678805552
transform 1 0 1632 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1401_
timestamp 1678805552
transform 1 0 1152 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1402_
timestamp 1678805552
transform 1 0 12000 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1403_
timestamp 1678805552
transform 1 0 10848 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1404_
timestamp 1678805552
transform 1 0 9408 0 1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1405_
timestamp 1678805552
transform 1 0 7488 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1406_
timestamp 1678805552
transform 1 0 1248 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1407_
timestamp 1678805552
transform -1 0 2784 0 1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1408_
timestamp 1678805552
transform 1 0 3552 0 1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1409_
timestamp 1678805552
transform 1 0 3648 0 -1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1410_
timestamp 1678805552
transform 1 0 15264 0 -1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1411_
timestamp 1678805552
transform 1 0 16128 0 1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1412_
timestamp 1678805552
transform 1 0 12192 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1413_
timestamp 1678805552
transform 1 0 13632 0 1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1414_
timestamp 1678805552
transform 1 0 2304 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1415_
timestamp 1678805552
transform 1 0 4512 0 1 29484
box -50 -56 1692 834
use sg13g2_buf_1  _1416_
timestamp 1676381911
transform 1 0 16320 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  _1417_
timestamp 1676381911
transform 1 0 18912 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1418_
timestamp 1676381911
transform 1 0 18912 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1419_
timestamp 1676381911
transform 1 0 18528 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1420_
timestamp 1676381911
transform 1 0 19296 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1421_
timestamp 1676381911
transform 1 0 18912 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1422_
timestamp 1676381911
transform 1 0 19968 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1423_
timestamp 1676381911
transform 1 0 19584 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1424_
timestamp 1676381911
transform 1 0 19584 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1425_
timestamp 1676381911
transform 1 0 19680 0 -1 43092
box -48 -56 432 834
use sg13g2_buf_1  _1426_
timestamp 1676381911
transform 1 0 19296 0 1 43092
box -48 -56 432 834
use sg13g2_buf_1  _1427_
timestamp 1676381911
transform 1 0 17760 0 1 43092
box -48 -56 432 834
use sg13g2_buf_1  _1428_
timestamp 1676381911
transform 1 0 19680 0 -1 44604
box -48 -56 432 834
use sg13g2_buf_1  _1429_
timestamp 1676381911
transform 1 0 19776 0 1 44604
box -48 -56 432 834
use sg13g2_buf_1  _1430_
timestamp 1676381911
transform 1 0 19488 0 -1 46116
box -48 -56 432 834
use sg13g2_buf_1  _1431_
timestamp 1676381911
transform 1 0 11808 0 1 46116
box -48 -56 432 834
use sg13g2_buf_1  _1432_
timestamp 1676381911
transform 1 0 19776 0 1 46116
box -48 -56 432 834
use sg13g2_buf_1  _1433_
timestamp 1676381911
transform 1 0 19776 0 1 47628
box -48 -56 432 834
use sg13g2_buf_1  _1434_
timestamp 1676381911
transform 1 0 19872 0 -1 49140
box -48 -56 432 834
use sg13g2_buf_1  _1435_
timestamp 1676381911
transform 1 0 19296 0 1 49140
box -48 -56 432 834
use sg13g2_buf_1  _1436_
timestamp 1676381911
transform 1 0 19680 0 1 49140
box -48 -56 432 834
use sg13g2_buf_1  _1437_
timestamp 1676381911
transform 1 0 19392 0 -1 50652
box -48 -56 432 834
use sg13g2_buf_1  _1438_
timestamp 1676381911
transform 1 0 19776 0 -1 50652
box -48 -56 432 834
use sg13g2_buf_1  _1439_
timestamp 1676381911
transform 1 0 19872 0 1 50652
box -48 -56 432 834
use sg13g2_buf_1  _1440_
timestamp 1676381911
transform 1 0 19680 0 1 52164
box -48 -56 432 834
use sg13g2_buf_1  _1441_
timestamp 1676381911
transform 1 0 19392 0 1 53676
box -48 -56 432 834
use sg13g2_buf_1  _1442_
timestamp 1676381911
transform 1 0 9888 0 1 53676
box -48 -56 432 834
use sg13g2_buf_1  _1443_
timestamp 1676381911
transform 1 0 19776 0 1 53676
box -48 -56 432 834
use sg13g2_buf_1  _1444_
timestamp 1676381911
transform 1 0 19584 0 -1 55188
box -48 -56 432 834
use sg13g2_buf_1  _1445_
timestamp 1676381911
transform 1 0 19968 0 -1 55188
box -48 -56 432 834
use sg13g2_buf_1  _1446_
timestamp 1676381911
transform 1 0 19296 0 1 55188
box -48 -56 432 834
use sg13g2_buf_1  _1447_
timestamp 1676381911
transform 1 0 10272 0 -1 56700
box -48 -56 432 834
use sg13g2_buf_1  _1448_
timestamp 1676381911
transform 1 0 19296 0 -1 56700
box -48 -56 432 834
use sg13g2_buf_1  _1449_
timestamp 1676381911
transform 1 0 15552 0 1 80892
box -48 -56 432 834
use sg13g2_buf_1  _1450_
timestamp 1676381911
transform 1 0 15744 0 1 79380
box -48 -56 432 834
use sg13g2_buf_1  _1451_
timestamp 1676381911
transform 1 0 15936 0 -1 73332
box -48 -56 432 834
use sg13g2_buf_1  _1452_
timestamp 1676381911
transform -1 0 16608 0 1 56700
box -48 -56 432 834
use sg13g2_buf_1  _1453_
timestamp 1676381911
transform -1 0 17184 0 -1 56700
box -48 -56 432 834
use sg13g2_buf_1  _1454_
timestamp 1676381911
transform 1 0 16512 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1455_
timestamp 1676381911
transform 1 0 16704 0 -1 79380
box -48 -56 432 834
use sg13g2_buf_1  _1456_
timestamp 1676381911
transform 1 0 16896 0 1 76356
box -48 -56 432 834
use sg13g2_buf_1  _1457_
timestamp 1676381911
transform -1 0 17664 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1458_
timestamp 1676381911
transform -1 0 18048 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1459_
timestamp 1676381911
transform -1 0 18432 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1460_
timestamp 1676381911
transform -1 0 18816 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1461_
timestamp 1676381911
transform 1 0 17952 0 1 82404
box -48 -56 432 834
use sg13g2_buf_1  _1462_
timestamp 1676381911
transform -1 0 19200 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1463_
timestamp 1676381911
transform 1 0 18336 0 1 82404
box -48 -56 432 834
use sg13g2_buf_1  _1464_
timestamp 1676381911
transform -1 0 19584 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1465_
timestamp 1676381911
transform 1 0 18720 0 1 82404
box -48 -56 432 834
use sg13g2_buf_1  _1466_
timestamp 1676381911
transform -1 0 19968 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1467_
timestamp 1676381911
transform 1 0 19104 0 1 82404
box -48 -56 432 834
use sg13g2_buf_1  _1468_
timestamp 1676381911
transform -1 0 20352 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1469_
timestamp 1676381911
transform -1 0 6720 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1470_
timestamp 1676381911
transform 1 0 1632 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1471_
timestamp 1676381911
transform -1 0 17280 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1472_
timestamp 1676381911
transform -1 0 5856 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1473_
timestamp 1676381911
transform 1 0 2016 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1474_
timestamp 1676381911
transform -1 0 3360 0 1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1475_
timestamp 1676381911
transform -1 0 3744 0 1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1476_
timestamp 1676381911
transform 1 0 2400 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1477_
timestamp 1676381911
transform -1 0 3936 0 1 82404
box -48 -56 432 834
use sg13g2_buf_1  _1478_
timestamp 1676381911
transform 1 0 3168 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1479_
timestamp 1676381911
transform -1 0 10368 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1480_
timestamp 1676381911
transform 1 0 3552 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1481_
timestamp 1676381911
transform 1 0 2784 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1482_
timestamp 1676381911
transform -1 0 9888 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1483_
timestamp 1676381911
transform -1 0 5088 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1484_
timestamp 1676381911
transform 1 0 3936 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1485_
timestamp 1676381911
transform 1 0 4320 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1486_
timestamp 1676381911
transform -1 0 10752 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1487_
timestamp 1676381911
transform -1 0 11616 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1488_
timestamp 1676381911
transform 1 0 5088 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1489_
timestamp 1676381911
transform -1 0 6240 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1490_
timestamp 1676381911
transform -1 0 6624 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1491_
timestamp 1676381911
transform -1 0 7008 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1492_
timestamp 1676381911
transform -1 0 6528 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1493_
timestamp 1676381911
transform -1 0 6912 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1494_
timestamp 1676381911
transform -1 0 7680 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1495_
timestamp 1676381911
transform -1 0 7296 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1496_
timestamp 1676381911
transform -1 0 8064 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1497_
timestamp 1676381911
transform 1 0 5952 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1498_
timestamp 1676381911
transform -1 0 7872 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1499_
timestamp 1676381911
transform -1 0 8256 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1500_
timestamp 1676381911
transform 1 0 6720 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1501_
timestamp 1676381911
transform 1 0 7200 0 1 82404
box -48 -56 432 834
use sg13g2_buf_1  _1502_
timestamp 1676381911
transform -1 0 8736 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1503_
timestamp 1676381911
transform -1 0 9120 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1504_
timestamp 1676381911
transform 1 0 7104 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1505_
timestamp 1676381911
transform -1 0 16032 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1506_
timestamp 1676381911
transform -1 0 9312 0 -1 44604
box -48 -56 432 834
use sg13g2_buf_1  _1507_
timestamp 1676381911
transform -1 0 14208 0 1 43092
box -48 -56 432 834
use sg13g2_buf_1  _1508_
timestamp 1676381911
transform -1 0 17760 0 1 43092
box -48 -56 432 834
use sg13g2_buf_1  _1509_
timestamp 1676381911
transform -1 0 9984 0 -1 44604
box -48 -56 432 834
use sg13g2_buf_1  _1510_
timestamp 1676381911
transform -1 0 2208 0 1 44604
box -48 -56 432 834
use sg13g2_buf_1  _1511_
timestamp 1676381911
transform -1 0 19104 0 -1 46116
box -48 -56 432 834
use sg13g2_buf_1  _1512_
timestamp 1676381911
transform -1 0 11712 0 -1 46116
box -48 -56 432 834
use sg13g2_buf_1  _1513_
timestamp 1676381911
transform -1 0 1824 0 1 44604
box -48 -56 432 834
use sg13g2_buf_1  _1514_
timestamp 1676381911
transform -1 0 2208 0 1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1515_
timestamp 1676381911
transform -1 0 17184 0 1 44604
box -48 -56 432 834
use sg13g2_buf_1  _1516_
timestamp 1676381911
transform -1 0 14016 0 1 44604
box -48 -56 432 834
use sg13g2_buf_1  _1517_
timestamp 1676381911
transform -1 0 1824 0 -1 46116
box -48 -56 432 834
use sg13g2_buf_1  _1518_
timestamp 1676381911
transform -1 0 2208 0 -1 46116
box -48 -56 432 834
use sg13g2_buf_1  _1519_
timestamp 1676381911
transform -1 0 19488 0 -1 46116
box -48 -56 432 834
use sg13g2_buf_1  _1520_
timestamp 1676381911
transform -1 0 10944 0 -1 47628
box -48 -56 432 834
use sg13g2_buf_1  _1521_
timestamp 1676381911
transform -1 0 2112 0 -1 47628
box -48 -56 432 834
use sg13g2_buf_1  _1522_
timestamp 1676381911
transform -1 0 2112 0 -1 44604
box -48 -56 432 834
use sg13g2_buf_1  _1523_
timestamp 1676381911
transform -1 0 16512 0 1 47628
box -48 -56 432 834
use sg13g2_buf_1  _1524_
timestamp 1676381911
transform -1 0 13248 0 -1 46116
box -48 -56 432 834
use sg13g2_buf_1  _1525_
timestamp 1676381911
transform -1 0 1824 0 1 49140
box -48 -56 432 834
use sg13g2_buf_1  _1526_
timestamp 1676381911
transform -1 0 10176 0 1 55188
box -48 -56 432 834
use sg13g2_buf_1  _1527_
timestamp 1676381911
transform -1 0 16128 0 1 56700
box -48 -56 432 834
use sg13g2_buf_1  _1528_
timestamp 1676381911
transform -1 0 15168 0 -1 56700
box -48 -56 432 834
use sg13g2_buf_1  _1529_
timestamp 1676381911
transform -1 0 9792 0 1 56700
box -48 -56 432 834
use sg13g2_buf_1  _1530_
timestamp 1676381911
transform -1 0 1920 0 1 47628
box -48 -56 432 834
use sg13g2_buf_1  _1531_
timestamp 1676381911
transform -1 0 19872 0 1 50652
box -48 -56 432 834
use sg13g2_buf_1  _1532_
timestamp 1676381911
transform -1 0 12672 0 -1 56700
box -48 -56 432 834
use sg13g2_buf_1  _1533_
timestamp 1676381911
transform -1 0 2112 0 1 56700
box -48 -56 432 834
use sg13g2_buf_1  _1534_
timestamp 1676381911
transform -1 0 3168 0 1 50652
box -48 -56 432 834
use sg13g2_buf_1  _1535_
timestamp 1676381911
transform -1 0 17472 0 1 53676
box -48 -56 432 834
use sg13g2_buf_1  _1536_
timestamp 1676381911
transform -1 0 11616 0 -1 58212
box -48 -56 432 834
use sg13g2_buf_1  _1537_
timestamp 1676381911
transform -1 0 2208 0 -1 59724
box -48 -56 432 834
use sg13g2_buf_1  _1538_
timestamp 1676381911
transform -1 0 2208 0 -1 52164
box -48 -56 432 834
use sg13g2_buf_1  _1539_
timestamp 1676381911
transform -1 0 19680 0 1 52164
box -48 -56 432 834
use sg13g2_buf_1  _1540_
timestamp 1676381911
transform -1 0 13536 0 -1 50652
box -48 -56 432 834
use sg13g2_buf_1  _1541_
timestamp 1676381911
transform -1 0 1824 0 -1 52164
box -48 -56 432 834
use sg13g2_buf_1  _1542_
timestamp 1676381911
transform -1 0 3168 0 -1 49140
box -48 -56 432 834
use sg13g2_buf_1  _1543_
timestamp 1676381911
transform -1 0 16128 0 -1 50652
box -48 -56 432 834
use sg13g2_buf_1  _1544_
timestamp 1676381911
transform -1 0 12672 0 1 50652
box -48 -56 432 834
use sg13g2_buf_1  _1545_
timestamp 1676381911
transform -1 0 1728 0 1 52164
box -48 -56 432 834
use sg13g2_buf_1  _1546_
timestamp 1676381911
transform -1 0 2208 0 1 49140
box -48 -56 432 834
use sg13g2_buf_1  _1547_
timestamp 1676381911
transform -1 0 19296 0 1 49140
box -48 -56 432 834
use sg13g2_buf_1  _1548_
timestamp 1676381911
transform -1 0 12288 0 1 53676
box -48 -56 432 834
use sg13g2_buf_1  _1549_
timestamp 1676381911
transform -1 0 2112 0 -1 55188
box -48 -56 432 834
use sg13g2_buf_1  _1550_
timestamp 1676381911
transform -1 0 2112 0 1 52164
box -48 -56 432 834
use sg13g2_buf_1  _1551_
timestamp 1676381911
transform -1 0 17376 0 -1 53676
box -48 -56 432 834
use sg13g2_buf_1  _1552_
timestamp 1676381911
transform -1 0 19584 0 -1 55188
box -48 -56 432 834
use sg13g2_buf_1  _1553_
timestamp 1676381911
transform -1 0 3360 0 1 55188
box -48 -56 432 834
use sg13g2_buf_1  _1554_
timestamp 1676381911
transform 1 0 19296 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  _1555_
timestamp 1676381911
transform 1 0 19680 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  _1556_
timestamp 1676381911
transform 1 0 18912 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  _1557_
timestamp 1676381911
transform 1 0 18912 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  _1558_
timestamp 1676381911
transform 1 0 19296 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1559_
timestamp 1676381911
transform 1 0 19680 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1560_
timestamp 1676381911
transform 1 0 12960 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1561_
timestamp 1676381911
transform 1 0 14400 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1562_
timestamp 1676381911
transform 1 0 19296 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  _1563_
timestamp 1676381911
transform 1 0 19296 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  _1564_
timestamp 1676381911
transform 1 0 14304 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1565_
timestamp 1676381911
transform 1 0 15264 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1566_
timestamp 1676381911
transform 1 0 19296 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1567_
timestamp 1676381911
transform 1 0 19680 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1568_
timestamp 1676381911
transform 1 0 19296 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1569_
timestamp 1676381911
transform 1 0 19296 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1570_
timestamp 1676381911
transform 1 0 18816 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1571_
timestamp 1676381911
transform 1 0 12672 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1572_
timestamp 1676381911
transform 1 0 19296 0 -1 43092
box -48 -56 432 834
use sg13g2_buf_1  _1573_
timestamp 1676381911
transform 1 0 16896 0 1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1574_
timestamp 1676381911
transform 1 0 19776 0 1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1575_
timestamp 1676381911
transform 1 0 18624 0 1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1576_
timestamp 1676381911
transform 1 0 19200 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1577_
timestamp 1676381911
transform 1 0 19392 0 1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1578_
timestamp 1676381911
transform 1 0 19200 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1579_
timestamp 1676381911
transform 1 0 18816 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1580_
timestamp 1676381911
transform 1 0 18240 0 1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1581_
timestamp 1676381911
transform 1 0 19008 0 1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1582_
timestamp 1676381911
transform 1 0 18528 0 -1 43092
box -48 -56 432 834
use sg13g2_buf_1  _1583_
timestamp 1676381911
transform 1 0 18912 0 -1 43092
box -48 -56 432 834
use sg13g2_buf_1  _1584_
timestamp 1676381911
transform 1 0 18912 0 1 43092
box -48 -56 432 834
use sg13g2_buf_1  _1585_
timestamp 1676381911
transform 1 0 14784 0 1 43092
box -48 -56 432 834
use sg13g2_buf_1  _1586_
timestamp 1676381911
transform 1 0 7776 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1587_
timestamp 1676381911
transform -1 0 15360 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1588_
timestamp 1676381911
transform -1 0 16128 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1589_
timestamp 1676381911
transform 1 0 8160 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1590_
timestamp 1676381911
transform 1 0 3072 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1591_
timestamp 1676381911
transform 1 0 9312 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1592_
timestamp 1676381911
transform -1 0 13056 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1593_
timestamp 1676381911
transform 1 0 8928 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1594_
timestamp 1676381911
transform 1 0 8544 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1595_
timestamp 1676381911
transform 1 0 10080 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1596_
timestamp 1676381911
transform -1 0 12000 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1597_
timestamp 1676381911
transform 1 0 9696 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1598_
timestamp 1676381911
transform -1 0 11424 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1599_
timestamp 1676381911
transform 1 0 8928 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1600_
timestamp 1676381911
transform -1 0 12384 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1601_
timestamp 1676381911
transform 1 0 10464 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1602_
timestamp 1676381911
transform 1 0 10848 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1603_
timestamp 1676381911
transform 1 0 10464 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1604_
timestamp 1676381911
transform 1 0 10848 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1605_
timestamp 1676381911
transform 1 0 11232 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1606_
timestamp 1676381911
transform -1 0 13440 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1607_
timestamp 1676381911
transform -1 0 13824 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1608_
timestamp 1676381911
transform -1 0 14208 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1609_
timestamp 1676381911
transform -1 0 14592 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1610_
timestamp 1676381911
transform -1 0 14976 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1611_
timestamp 1676381911
transform -1 0 14496 0 1 82404
box -48 -56 432 834
use sg13g2_buf_1  _1612_
timestamp 1676381911
transform -1 0 15360 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1613_
timestamp 1676381911
transform -1 0 14880 0 1 82404
box -48 -56 432 834
use sg13g2_buf_1  _1614_
timestamp 1676381911
transform 1 0 13152 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1615_
timestamp 1676381911
transform -1 0 15744 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1616_
timestamp 1676381911
transform -1 0 15264 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1617_
timestamp 1676381911
transform 1 0 13824 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1618_
timestamp 1676381911
transform 1 0 14208 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1619_
timestamp 1676381911
transform -1 0 16128 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1620_
timestamp 1676381911
transform -1 0 16512 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1621_
timestamp 1676381911
transform 1 0 14592 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1622_
timestamp 1676381911
transform -1 0 2208 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1623_
timestamp 1676381911
transform -1 0 2976 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1624_
timestamp 1676381911
transform -1 0 2592 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1625_
timestamp 1676381911
transform -1 0 1824 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1626_
timestamp 1676381911
transform -1 0 2592 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1627_
timestamp 1676381911
transform -1 0 1824 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1628_
timestamp 1676381911
transform -1 0 2208 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1629_
timestamp 1676381911
transform -1 0 2688 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1630_
timestamp 1676381911
transform -1 0 3360 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _1631_
timestamp 1676381911
transform -1 0 2208 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1632_
timestamp 1676381911
transform -1 0 1824 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1633_
timestamp 1676381911
transform -1 0 2976 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _1634_
timestamp 1676381911
transform -1 0 2592 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _1635_
timestamp 1676381911
transform -1 0 1824 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _1636_
timestamp 1676381911
transform -1 0 2208 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _1637_
timestamp 1676381911
transform -1 0 3360 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _1638_
timestamp 1676381911
transform -1 0 2208 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _1639_
timestamp 1676381911
transform -1 0 2592 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _1640_
timestamp 1676381911
transform -1 0 1824 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _1641_
timestamp 1676381911
transform -1 0 3456 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _1642_
timestamp 1676381911
transform -1 0 7776 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  _1643_
timestamp 1676381911
transform -1 0 17952 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  _1644_
timestamp 1676381911
transform -1 0 2016 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  _1645_
timestamp 1676381911
transform -1 0 2208 0 -1 29484
box -48 -56 432 834
use sg13g2_buf_1  _1646_
timestamp 1676381911
transform -1 0 1728 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  _1647_
timestamp 1676381911
transform -1 0 4512 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  _1648_
timestamp 1676381911
transform -1 0 2112 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  _1649_
timestamp 1676381911
transform -1 0 3168 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  _1650_
timestamp 1676381911
transform -1 0 7968 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  _1651_
timestamp 1676381911
transform -1 0 1632 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  _1652_
timestamp 1676381911
transform -1 0 1728 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  _1653_
timestamp 1676381911
transform -1 0 1728 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  _1654_
timestamp 1676381911
transform -1 0 2016 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _1655_
timestamp 1676381911
transform -1 0 18912 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _1656_
timestamp 1676381911
transform -1 0 1632 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _1657_
timestamp 1676381911
transform -1 0 3552 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _1658_
timestamp 1676381911
transform -1 0 1824 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _1659_
timestamp 1676381911
transform -1 0 2208 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _1660_
timestamp 1676381911
transform -1 0 1536 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _1661_
timestamp 1676381911
transform -1 0 1824 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _1662_
timestamp 1676381911
transform -1 0 1632 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  _1663_
timestamp 1676381911
transform -1 0 2208 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _1664_
timestamp 1676381911
transform -1 0 2592 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _1665_
timestamp 1676381911
transform -1 0 8256 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  _1666_
timestamp 1676381911
transform -1 0 10848 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  _1667_
timestamp 1676381911
transform -1 0 1728 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  _1668_
timestamp 1676381911
transform -1 0 4032 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _1669_
timestamp 1676381911
transform -1 0 2016 0 -1 11340
box -48 -56 432 834
use sg13g2_antennanp  ANTENNA_1
timestamp 1679999689
transform -1 0 5088 0 1 41580
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_2
timestamp 1679999689
transform 1 0 18048 0 1 83916
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_3
timestamp 1679999689
transform 1 0 18432 0 1 83916
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_4
timestamp 1679999689
transform 1 0 17952 0 -1 82404
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_5
timestamp 1679999689
transform 1 0 18816 0 1 83916
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_6
timestamp 1679999689
transform 1 0 18336 0 -1 82404
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_7
timestamp 1679999689
transform 1 0 19200 0 1 83916
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_8
timestamp 1679999689
transform 1 0 18720 0 -1 82404
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_9
timestamp 1679999689
transform 1 0 19584 0 1 82404
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_10
timestamp 1679999689
transform 1 0 19104 0 -1 82404
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_11
timestamp 1679999689
transform 1 0 17280 0 1 82404
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_12
timestamp 1679999689
transform 1 0 17664 0 1 82404
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_13
timestamp 1679999689
transform 1 0 9216 0 -1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_14
timestamp 1679999689
transform 1 0 10656 0 -1 74844
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_15
timestamp 1679999689
transform 1 0 9216 0 -1 41580
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_16
timestamp 1679999689
transform -1 0 10944 0 -1 76356
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_17
timestamp 1679999689
transform 1 0 19968 0 1 82404
box -48 -56 336 834
use sg13g2_buf_8  clkbuf_0_Tile_X0Y1_UserCLK
timestamp 1676451365
transform 1 0 16128 0 -1 59724
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_1_0__f_Tile_X0Y1_UserCLK
timestamp 1676451365
transform -1 0 17376 0 -1 50652
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_1_1__f_Tile_X0Y1_UserCLK
timestamp 1676451365
transform -1 0 17280 0 1 70308
box -48 -56 1296 834
use sg13g2_fill_2  FILLER_0_0
timestamp 1677580104
transform 1 0 1152 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_2
timestamp 1677579658
transform 1 0 1344 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_15
timestamp 1679581782
transform 1 0 2592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_22
timestamp 1679581782
transform 1 0 3264 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_29
timestamp 1679581782
transform 1 0 3936 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_36
timestamp 1679577901
transform 1 0 4608 0 1 756
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_40
timestamp 1677579658
transform 1 0 4992 0 1 756
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_46
timestamp 1677580104
transform 1 0 5568 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_48
timestamp 1677579658
transform 1 0 5760 0 1 756
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_61
timestamp 1677580104
transform 1 0 7008 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_63
timestamp 1677579658
transform 1 0 7200 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_72
timestamp 1679581782
transform 1 0 8064 0 1 756
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_79
timestamp 1677580104
transform 1 0 8736 0 1 756
box -48 -56 240 834
use sg13g2_decap_8  FILLER_0_105
timestamp 1679581782
transform 1 0 11232 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_112
timestamp 1679581782
transform 1 0 11904 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_119
timestamp 1679581782
transform 1 0 12576 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_126
timestamp 1679581782
transform 1 0 13248 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_133
timestamp 1679581782
transform 1 0 13920 0 1 756
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_140
timestamp 1677580104
transform 1 0 14592 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_142
timestamp 1677579658
transform 1 0 14784 0 1 756
box -48 -56 144 834
use sg13g2_decap_4  FILLER_0_147
timestamp 1679577901
transform 1 0 15264 0 1 756
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_151
timestamp 1677579658
transform 1 0 15648 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_156
timestamp 1679581782
transform 1 0 16128 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_163
timestamp 1679581782
transform 1 0 16800 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_170
timestamp 1679581782
transform 1 0 17472 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_177
timestamp 1679581782
transform 1 0 18144 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_184
timestamp 1679581782
transform 1 0 18816 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_191
timestamp 1679581782
transform 1 0 19488 0 1 756
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_198
timestamp 1677580104
transform 1 0 20160 0 1 756
box -48 -56 240 834
use sg13g2_fill_2  FILLER_1_0
timestamp 1677580104
transform 1 0 1152 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_2
timestamp 1677579658
transform 1 0 1344 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_19
timestamp 1677579658
transform 1 0 2976 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_51
timestamp 1677579658
transform 1 0 6048 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_95
timestamp 1677580104
transform 1 0 10272 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_1_117
timestamp 1677580104
transform 1 0 12384 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_119
timestamp 1677579658
transform 1 0 12576 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_124
timestamp 1677579658
transform 1 0 13056 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_129
timestamp 1677580104
transform 1 0 13536 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_131
timestamp 1677579658
transform 1 0 13728 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_160
timestamp 1679581782
transform 1 0 16512 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_167
timestamp 1679581782
transform 1 0 17184 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_174
timestamp 1679581782
transform 1 0 17856 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_181
timestamp 1679581782
transform 1 0 18528 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_188
timestamp 1679581782
transform 1 0 19200 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_195
timestamp 1679577901
transform 1 0 19872 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_199
timestamp 1677579658
transform 1 0 20256 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_0
timestamp 1677580104
transform 1 0 1152 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_2
timestamp 1677579658
transform 1 0 1344 0 1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_11
timestamp 1677579658
transform 1 0 2208 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_16
timestamp 1679581782
transform 1 0 2688 0 1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_23
timestamp 1677579658
transform 1 0 3360 0 1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_49
timestamp 1679577901
transform 1 0 5856 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_70
timestamp 1677580104
transform 1 0 7872 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_107
timestamp 1679581782
transform 1 0 11424 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_114
timestamp 1679581782
transform 1 0 12096 0 1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_121
timestamp 1677579658
transform 1 0 12768 0 1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_139
timestamp 1677580104
transform 1 0 14496 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_141
timestamp 1677579658
transform 1 0 14688 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_159
timestamp 1679581782
transform 1 0 16416 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_166
timestamp 1679581782
transform 1 0 17088 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_173
timestamp 1679581782
transform 1 0 17760 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_180
timestamp 1679581782
transform 1 0 18432 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_187
timestamp 1679581782
transform 1 0 19104 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_194
timestamp 1679577901
transform 1 0 19776 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_198
timestamp 1677580104
transform 1 0 20160 0 1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_0
timestamp 1677580104
transform 1 0 1152 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_2
timestamp 1677579658
transform 1 0 1344 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_23
timestamp 1677580104
transform 1 0 3360 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_4  FILLER_3_50
timestamp 1679577901
transform 1 0 5952 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_76
timestamp 1677579658
transform 1 0 8448 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_141
timestamp 1679581782
transform 1 0 14688 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_165
timestamp 1679581782
transform 1 0 16992 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_172
timestamp 1679581782
transform 1 0 17664 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_179
timestamp 1679581782
transform 1 0 18336 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_186
timestamp 1679581782
transform 1 0 19008 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_193
timestamp 1679581782
transform 1 0 19680 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_0
timestamp 1677580104
transform 1 0 1152 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_2
timestamp 1677579658
transform 1 0 1344 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_15
timestamp 1677580104
transform 1 0 2592 0 1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_22
timestamp 1677580104
transform 1 0 3264 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_24
timestamp 1677579658
transform 1 0 3456 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_42
timestamp 1677580104
transform 1 0 5184 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_44
timestamp 1677579658
transform 1 0 5376 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_50
timestamp 1679581782
transform 1 0 5952 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_57
timestamp 1677580104
transform 1 0 6624 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_72
timestamp 1679581782
transform 1 0 8064 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_79
timestamp 1679581782
transform 1 0 8736 0 1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_86
timestamp 1677579658
transform 1 0 9408 0 1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_92
timestamp 1677579658
transform 1 0 9984 0 1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_98
timestamp 1677579658
transform 1 0 10560 0 1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_4_116
timestamp 1679577901
transform 1 0 12288 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_120
timestamp 1677580104
transform 1 0 12672 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_160
timestamp 1679581782
transform 1 0 16512 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_167
timestamp 1679581782
transform 1 0 17184 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_174
timestamp 1679581782
transform 1 0 17856 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_181
timestamp 1679581782
transform 1 0 18528 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_188
timestamp 1679581782
transform 1 0 19200 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_195
timestamp 1679577901
transform 1 0 19872 0 1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_199
timestamp 1677579658
transform 1 0 20256 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_0
timestamp 1677580104
transform 1 0 1152 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_2  FILLER_5_45
timestamp 1677580104
transform 1 0 5472 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_2  FILLER_5_72
timestamp 1677580104
transform 1 0 8064 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_74
timestamp 1677579658
transform 1 0 8256 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_97
timestamp 1677579658
transform 1 0 10464 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_5_125
timestamp 1679577901
transform 1 0 13152 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_129
timestamp 1677580104
transform 1 0 13536 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_148
timestamp 1677579658
transform 1 0 15360 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_166
timestamp 1679581782
transform 1 0 17088 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_173
timestamp 1679581782
transform 1 0 17760 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_180
timestamp 1679581782
transform 1 0 18432 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_187
timestamp 1679581782
transform 1 0 19104 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_194
timestamp 1679577901
transform 1 0 19776 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_198
timestamp 1677580104
transform 1 0 20160 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_2  FILLER_6_0
timestamp 1677580104
transform 1 0 1152 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_19
timestamp 1677579658
transform 1 0 2976 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_75
timestamp 1677579658
transform 1 0 8352 0 1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_6_101
timestamp 1679577901
transform 1 0 10848 0 1 5292
box -48 -56 432 834
use sg13g2_decap_4  FILLER_6_139
timestamp 1679577901
transform 1 0 14496 0 1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_143
timestamp 1677579658
transform 1 0 14880 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_186
timestamp 1679581782
transform 1 0 19008 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_193
timestamp 1679581782
transform 1 0 19680 0 1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_0
timestamp 1677579658
transform 1 0 1152 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_22
timestamp 1677580104
transform 1 0 3264 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_24
timestamp 1677579658
transform 1 0 3456 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_77
timestamp 1677579658
transform 1 0 8544 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_116
timestamp 1677579658
transform 1 0 12288 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_138
timestamp 1679581782
transform 1 0 14400 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_145
timestamp 1677580104
transform 1 0 15072 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_147
timestamp 1677579658
transform 1 0 15264 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_165
timestamp 1677579658
transform 1 0 16992 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_183
timestamp 1679581782
transform 1 0 18720 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_190
timestamp 1679581782
transform 1 0 19392 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_197
timestamp 1677580104
transform 1 0 20064 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_199
timestamp 1677579658
transform 1 0 20256 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_0
timestamp 1677580104
transform 1 0 1152 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_2
timestamp 1677579658
transform 1 0 1344 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_46
timestamp 1677579658
transform 1 0 5568 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_81
timestamp 1677580104
transform 1 0 8928 0 1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_105
timestamp 1677580104
transform 1 0 11232 0 1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_158
timestamp 1679581782
transform 1 0 16320 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_165
timestamp 1679581782
transform 1 0 16992 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_172
timestamp 1679581782
transform 1 0 17664 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_179
timestamp 1679581782
transform 1 0 18336 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_186
timestamp 1679581782
transform 1 0 19008 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_193
timestamp 1679581782
transform 1 0 19680 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_80
timestamp 1677580104
transform 1 0 8832 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_82
timestamp 1677579658
transform 1 0 9024 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_100
timestamp 1677580104
transform 1 0 10752 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_119
timestamp 1677579658
transform 1 0 12576 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_141
timestamp 1677580104
transform 1 0 14688 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_185
timestamp 1679581782
transform 1 0 18912 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_192
timestamp 1679581782
transform 1 0 19584 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_199
timestamp 1677579658
transform 1 0 20256 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_0
timestamp 1677580104
transform 1 0 1152 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_2
timestamp 1677579658
transform 1 0 1344 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_11
timestamp 1677580104
transform 1 0 2208 0 1 8316
box -48 -56 240 834
use sg13g2_decap_4  FILLER_10_68
timestamp 1679577901
transform 1 0 7680 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_72
timestamp 1677580104
transform 1 0 8064 0 1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_120
timestamp 1679581782
transform 1 0 12672 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_127
timestamp 1679581782
transform 1 0 13344 0 1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_134
timestamp 1677579658
transform 1 0 14016 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_152
timestamp 1679581782
transform 1 0 15744 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_159
timestamp 1679581782
transform 1 0 16416 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_166
timestamp 1677580104
transform 1 0 17088 0 1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_189
timestamp 1679581782
transform 1 0 19296 0 1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_196
timestamp 1679577901
transform 1 0 19968 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_0
timestamp 1677580104
transform 1 0 1152 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_2
timestamp 1677579658
transform 1 0 1344 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_15
timestamp 1677579658
transform 1 0 2592 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_11_26
timestamp 1679577901
transform 1 0 3648 0 -1 9828
box -48 -56 432 834
use sg13g2_decap_8  FILLER_11_43
timestamp 1679581782
transform 1 0 5280 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_50
timestamp 1677580104
transform 1 0 5952 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_52
timestamp 1677579658
transform 1 0 6144 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_92
timestamp 1677580104
transform 1 0 9984 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_94
timestamp 1677579658
transform 1 0 10176 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_11_146
timestamp 1679577901
transform 1 0 15168 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_150
timestamp 1677580104
transform 1 0 15552 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_169
timestamp 1677580104
transform 1 0 17376 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_171
timestamp 1677579658
transform 1 0 17568 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_189
timestamp 1679581782
transform 1 0 19296 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_196
timestamp 1679577901
transform 1 0 19968 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_12_0
timestamp 1677580104
transform 1 0 1152 0 1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_12_53
timestamp 1679581782
transform 1 0 6240 0 1 9828
box -48 -56 720 834
use sg13g2_fill_1  FILLER_12_60
timestamp 1677579658
transform 1 0 6912 0 1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_12_78
timestamp 1679577901
transform 1 0 8640 0 1 9828
box -48 -56 432 834
use sg13g2_decap_4  FILLER_12_120
timestamp 1679577901
transform 1 0 12672 0 1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_12_145
timestamp 1677579658
transform 1 0 15072 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_184
timestamp 1679581782
transform 1 0 18816 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_191
timestamp 1679581782
transform 1 0 19488 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_198
timestamp 1677580104
transform 1 0 20160 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_0
timestamp 1677579658
transform 1 0 1152 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_4  FILLER_13_26
timestamp 1679577901
transform 1 0 3648 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_13_30
timestamp 1677580104
transform 1 0 4032 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_4  FILLER_13_74
timestamp 1679577901
transform 1 0 8256 0 -1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_13_100
timestamp 1679581782
transform 1 0 10752 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_13_107
timestamp 1677580104
transform 1 0 11424 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_126
timestamp 1677579658
transform 1 0 13248 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_161
timestamp 1679581782
transform 1 0 16608 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_168
timestamp 1679577901
transform 1 0 17280 0 -1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_13_193
timestamp 1679581782
transform 1 0 19680 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_14_0
timestamp 1677580104
transform 1 0 1152 0 1 11340
box -48 -56 240 834
use sg13g2_decap_4  FILLER_14_69
timestamp 1679577901
transform 1 0 7776 0 1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_14_94
timestamp 1677580104
transform 1 0 10176 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_96
timestamp 1677579658
transform 1 0 10368 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_101
timestamp 1677580104
transform 1 0 10848 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_103
timestamp 1677579658
transform 1 0 11040 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_121
timestamp 1677580104
transform 1 0 12768 0 1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_14_144
timestamp 1679581782
transform 1 0 14976 0 1 11340
box -48 -56 720 834
use sg13g2_fill_1  FILLER_14_151
timestamp 1677579658
transform 1 0 15648 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_190
timestamp 1679581782
transform 1 0 19392 0 1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_14_197
timestamp 1677580104
transform 1 0 20064 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_199
timestamp 1677579658
transform 1 0 20256 0 1 11340
box -48 -56 144 834
use sg13g2_decap_4  FILLER_15_30
timestamp 1679577901
transform 1 0 4032 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_15_34
timestamp 1677579658
transform 1 0 4416 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_15_124
timestamp 1679577901
transform 1 0 13056 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_15_128
timestamp 1677580104
transform 1 0 13440 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_15_147
timestamp 1679581782
transform 1 0 15264 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_15_175
timestamp 1677579658
transform 1 0 17952 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_193
timestamp 1679581782
transform 1 0 19680 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_16_55
timestamp 1677580104
transform 1 0 6432 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_57
timestamp 1677579658
transform 1 0 6624 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_79
timestamp 1679581782
transform 1 0 8736 0 1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_16_86
timestamp 1677580104
transform 1 0 9408 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_88
timestamp 1677579658
transform 1 0 9600 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_106
timestamp 1679581782
transform 1 0 11328 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_113
timestamp 1679581782
transform 1 0 12000 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_120
timestamp 1679577901
transform 1 0 12672 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_124
timestamp 1677579658
transform 1 0 13056 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_146
timestamp 1679581782
transform 1 0 15168 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_170
timestamp 1679581782
transform 1 0 17472 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_177
timestamp 1679581782
transform 1 0 18144 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_184
timestamp 1679581782
transform 1 0 18816 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_191
timestamp 1679581782
transform 1 0 19488 0 1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_16_198
timestamp 1677580104
transform 1 0 20160 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_0
timestamp 1677579658
transform 1 0 1152 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_48
timestamp 1679581782
transform 1 0 5760 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_55
timestamp 1679581782
transform 1 0 6432 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_62
timestamp 1677580104
transform 1 0 7104 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_17_81
timestamp 1677580104
transform 1 0 8928 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_83
timestamp 1677579658
transform 1 0 9120 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_4  FILLER_17_105
timestamp 1679577901
transform 1 0 11232 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_17_109
timestamp 1677580104
transform 1 0 11616 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_4  FILLER_17_128
timestamp 1679577901
transform 1 0 13440 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_17_170
timestamp 1677580104
transform 1 0 17472 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_17_189
timestamp 1679581782
transform 1 0 19296 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_17_196
timestamp 1679577901
transform 1 0 19968 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_18_0
timestamp 1677580104
transform 1 0 1152 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_28
timestamp 1677579658
transform 1 0 3840 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_50
timestamp 1679581782
transform 1 0 5952 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_57
timestamp 1679581782
transform 1 0 6624 0 1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_64
timestamp 1677580104
transform 1 0 7296 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_66
timestamp 1677579658
transform 1 0 7488 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_88
timestamp 1677579658
transform 1 0 9600 0 1 14364
box -48 -56 144 834
use sg13g2_decap_4  FILLER_18_106
timestamp 1679577901
transform 1 0 11328 0 1 14364
box -48 -56 432 834
use sg13g2_decap_8  FILLER_18_148
timestamp 1679581782
transform 1 0 15360 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_155
timestamp 1679581782
transform 1 0 16032 0 1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_162
timestamp 1677580104
transform 1 0 16704 0 1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_18_185
timestamp 1679581782
transform 1 0 18912 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_192
timestamp 1679581782
transform 1 0 19584 0 1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_18_199
timestamp 1677579658
transform 1 0 20256 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_0
timestamp 1677580104
transform 1 0 1152 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_19_35
timestamp 1679581782
transform 1 0 4512 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_80
timestamp 1679581782
transform 1 0 8832 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_87
timestamp 1679581782
transform 1 0 9504 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_19_94
timestamp 1679577901
transform 1 0 10176 0 -1 15876
box -48 -56 432 834
use sg13g2_decap_8  FILLER_19_153
timestamp 1679581782
transform 1 0 15840 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_177
timestamp 1679581782
transform 1 0 18144 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_184
timestamp 1679581782
transform 1 0 18816 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_191
timestamp 1679581782
transform 1 0 19488 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_198
timestamp 1677580104
transform 1 0 20160 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_4  FILLER_20_26
timestamp 1679577901
transform 1 0 3648 0 1 15876
box -48 -56 432 834
use sg13g2_decap_8  FILLER_20_68
timestamp 1679581782
transform 1 0 7680 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_75
timestamp 1679581782
transform 1 0 8352 0 1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_20_82
timestamp 1677579658
transform 1 0 9024 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_104
timestamp 1679581782
transform 1 0 11136 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_111
timestamp 1679577901
transform 1 0 11808 0 1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_20_115
timestamp 1677580104
transform 1 0 12192 0 1 15876
box -48 -56 240 834
use sg13g2_decap_4  FILLER_20_134
timestamp 1679577901
transform 1 0 14016 0 1 15876
box -48 -56 432 834
use sg13g2_decap_8  FILLER_20_181
timestamp 1679581782
transform 1 0 18528 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_188
timestamp 1679581782
transform 1 0 19200 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_195
timestamp 1679577901
transform 1 0 19872 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_199
timestamp 1677579658
transform 1 0 20256 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_21_25
timestamp 1677579658
transform 1 0 3552 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_43
timestamp 1679581782
transform 1 0 5280 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_122
timestamp 1679581782
transform 1 0 12864 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_184
timestamp 1679581782
transform 1 0 18816 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_191
timestamp 1679581782
transform 1 0 19488 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_21_198
timestamp 1677580104
transform 1 0 20160 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_0
timestamp 1677579658
transform 1 0 1152 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_44
timestamp 1677580104
transform 1 0 5376 0 1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_22_97
timestamp 1679581782
transform 1 0 10464 0 1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_22_104
timestamp 1677580104
transform 1 0 11136 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_106
timestamp 1677579658
transform 1 0 11328 0 1 17388
box -48 -56 144 834
use sg13g2_decap_4  FILLER_22_124
timestamp 1679577901
transform 1 0 13056 0 1 17388
box -48 -56 432 834
use sg13g2_decap_4  FILLER_22_167
timestamp 1679577901
transform 1 0 17184 0 1 17388
box -48 -56 432 834
use sg13g2_decap_8  FILLER_22_188
timestamp 1679581782
transform 1 0 19200 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_195
timestamp 1679577901
transform 1 0 19872 0 1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_22_199
timestamp 1677579658
transform 1 0 20256 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_22
timestamp 1679581782
transform 1 0 3264 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_23_29
timestamp 1677580104
transform 1 0 3936 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_31
timestamp 1677579658
transform 1 0 4128 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_70
timestamp 1679581782
transform 1 0 7872 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_77
timestamp 1679581782
transform 1 0 8544 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_122
timestamp 1679581782
transform 1 0 12864 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_23_129
timestamp 1677580104
transform 1 0 13536 0 -1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_23_156
timestamp 1679581782
transform 1 0 16128 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_184
timestamp 1679581782
transform 1 0 18816 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_191
timestamp 1679581782
transform 1 0 19488 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_23_198
timestamp 1677580104
transform 1 0 20160 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_0
timestamp 1677579658
transform 1 0 1152 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_18
timestamp 1679581782
transform 1 0 2880 0 1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_24_25
timestamp 1679577901
transform 1 0 3552 0 1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_24_29
timestamp 1677580104
transform 1 0 3936 0 1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_24_69
timestamp 1679581782
transform 1 0 7776 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_97
timestamp 1679581782
transform 1 0 10464 0 1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_24_121
timestamp 1679577901
transform 1 0 12768 0 1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_24_125
timestamp 1677580104
transform 1 0 13152 0 1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_24_148
timestamp 1679581782
transform 1 0 15360 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_155
timestamp 1679581782
transform 1 0 16032 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_162
timestamp 1679581782
transform 1 0 16704 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_186
timestamp 1679581782
transform 1 0 19008 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_193
timestamp 1679581782
transform 1 0 19680 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_0
timestamp 1679581782
transform 1 0 1152 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_7
timestamp 1679577901
transform 1 0 1824 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_25_11
timestamp 1677580104
transform 1 0 2208 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_2  FILLER_25_30
timestamp 1677580104
transform 1 0 4032 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_32
timestamp 1677579658
transform 1 0 4224 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_140
timestamp 1679581782
transform 1 0 14592 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_147
timestamp 1677580104
transform 1 0 15264 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_149
timestamp 1677579658
transform 1 0 15456 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_177
timestamp 1679581782
transform 1 0 18144 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_184
timestamp 1679581782
transform 1 0 18816 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_191
timestamp 1679581782
transform 1 0 19488 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_198
timestamp 1677580104
transform 1 0 20160 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_2  FILLER_26_0
timestamp 1677580104
transform 1 0 1152 0 1 20412
box -48 -56 240 834
use sg13g2_decap_4  FILLER_26_83
timestamp 1679577901
transform 1 0 9120 0 1 20412
box -48 -56 432 834
use sg13g2_decap_8  FILLER_26_104
timestamp 1679581782
transform 1 0 11136 0 1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_26_111
timestamp 1679577901
transform 1 0 11808 0 1 20412
box -48 -56 432 834
use sg13g2_decap_4  FILLER_26_132
timestamp 1679577901
transform 1 0 13824 0 1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_26_136
timestamp 1677579658
transform 1 0 14208 0 1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_26_154
timestamp 1677579658
transform 1 0 15936 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_184
timestamp 1679581782
transform 1 0 18816 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_191
timestamp 1679581782
transform 1 0 19488 0 1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_26_198
timestamp 1677580104
transform 1 0 20160 0 1 20412
box -48 -56 240 834
use sg13g2_decap_4  FILLER_27_0
timestamp 1679577901
transform 1 0 1152 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_27_4
timestamp 1677579658
transform 1 0 1536 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_27_22
timestamp 1677580104
transform 1 0 3264 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_27_45
timestamp 1677580104
transform 1 0 5472 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_27_104
timestamp 1677580104
transform 1 0 11136 0 -1 21924
box -48 -56 240 834
use sg13g2_decap_4  FILLER_27_123
timestamp 1679577901
transform 1 0 12960 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_27_148
timestamp 1677579658
transform 1 0 15360 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_187
timestamp 1679581782
transform 1 0 19104 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_194
timestamp 1679577901
transform 1 0 19776 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_27_198
timestamp 1677580104
transform 1 0 20160 0 -1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_28_60
timestamp 1679581782
transform 1 0 6912 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_67
timestamp 1679577901
transform 1 0 7584 0 1 21924
box -48 -56 432 834
use sg13g2_decap_8  FILLER_28_76
timestamp 1679581782
transform 1 0 8448 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_83
timestamp 1679581782
transform 1 0 9120 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_90
timestamp 1679581782
transform 1 0 9792 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_97
timestamp 1679581782
transform 1 0 10464 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_104
timestamp 1679577901
transform 1 0 11136 0 1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_28_128
timestamp 1677580104
transform 1 0 13440 0 1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_28_147
timestamp 1679581782
transform 1 0 15264 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_154
timestamp 1679581782
transform 1 0 15936 0 1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_28_161
timestamp 1677580104
transform 1 0 16608 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_163
timestamp 1677579658
transform 1 0 16800 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_167
timestamp 1677580104
transform 1 0 17184 0 1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_28_174
timestamp 1679581782
transform 1 0 17856 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_181
timestamp 1679581782
transform 1 0 18528 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_188
timestamp 1679581782
transform 1 0 19200 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_195
timestamp 1679577901
transform 1 0 19872 0 1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_28_199
timestamp 1677579658
transform 1 0 20256 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_0
timestamp 1677580104
transform 1 0 1152 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_45
timestamp 1677579658
transform 1 0 5472 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_29_83
timestamp 1679581782
transform 1 0 9120 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_29_90
timestamp 1677580104
transform 1 0 9792 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_2  FILLER_29_130
timestamp 1677580104
transform 1 0 13632 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_132
timestamp 1677579658
transform 1 0 13824 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_160
timestamp 1677580104
transform 1 0 16512 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_2  FILLER_29_184
timestamp 1677580104
transform 1 0 18816 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_186
timestamp 1677579658
transform 1 0 19008 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_197
timestamp 1677580104
transform 1 0 20064 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_199
timestamp 1677579658
transform 1 0 20256 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_17
timestamp 1677580104
transform 1 0 2784 0 1 23436
box -48 -56 240 834
use sg13g2_decap_4  FILLER_30_103
timestamp 1679577901
transform 1 0 11040 0 1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_30_126
timestamp 1677579658
transform 1 0 13248 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_148
timestamp 1677579658
transform 1 0 15360 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_173
timestamp 1677580104
transform 1 0 17760 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_175
timestamp 1677579658
transform 1 0 17952 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_198
timestamp 1677580104
transform 1 0 20160 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_0
timestamp 1677579658
transform 1 0 1152 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_31_35
timestamp 1677580104
transform 1 0 4512 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_37
timestamp 1677579658
transform 1 0 4704 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_31_55
timestamp 1677579658
transform 1 0 6432 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_31_121
timestamp 1677580104
transform 1 0 12768 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_123
timestamp 1677579658
transform 1 0 12960 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_31_141
timestamp 1679577901
transform 1 0 14688 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_145
timestamp 1677580104
transform 1 0 15072 0 -1 24948
box -48 -56 240 834
use sg13g2_decap_4  FILLER_31_169
timestamp 1679577901
transform 1 0 17376 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_173
timestamp 1677580104
transform 1 0 17760 0 -1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_31_192
timestamp 1679581782
transform 1 0 19584 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_1  FILLER_31_199
timestamp 1677579658
transform 1 0 20256 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_0
timestamp 1679581782
transform 1 0 1152 0 1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_32_7
timestamp 1677580104
transform 1 0 1824 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_9
timestamp 1677579658
transform 1 0 2016 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_77
timestamp 1679581782
transform 1 0 8544 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_84
timestamp 1679577901
transform 1 0 9216 0 1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_32_88
timestamp 1677579658
transform 1 0 9600 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_106
timestamp 1679581782
transform 1 0 11328 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_113
timestamp 1679581782
transform 1 0 12000 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_120
timestamp 1679577901
transform 1 0 12672 0 1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_32_141
timestamp 1677580104
transform 1 0 14688 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_159
timestamp 1677579658
transform 1 0 16416 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_170
timestamp 1679581782
transform 1 0 17472 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_177
timestamp 1679581782
transform 1 0 18144 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_184
timestamp 1679581782
transform 1 0 18816 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_191
timestamp 1679581782
transform 1 0 19488 0 1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_32_198
timestamp 1677580104
transform 1 0 20160 0 1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_33_0
timestamp 1677580104
transform 1 0 1152 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_2
timestamp 1677579658
transform 1 0 1344 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_4  FILLER_33_20
timestamp 1679577901
transform 1 0 3072 0 -1 26460
box -48 -56 432 834
use sg13g2_decap_4  FILLER_33_46
timestamp 1679577901
transform 1 0 5568 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_33_50
timestamp 1677579658
transform 1 0 5952 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_4  FILLER_33_106
timestamp 1679577901
transform 1 0 11328 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_33_110
timestamp 1677580104
transform 1 0 11712 0 -1 26460
box -48 -56 240 834
use sg13g2_decap_4  FILLER_33_129
timestamp 1679577901
transform 1 0 13536 0 -1 26460
box -48 -56 432 834
use sg13g2_decap_8  FILLER_33_193
timestamp 1679581782
transform 1 0 19680 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_1  FILLER_34_0
timestamp 1677579658
transform 1 0 1152 0 1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_34_32
timestamp 1677580104
transform 1 0 4224 0 1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_34_89
timestamp 1677580104
transform 1 0 9696 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_91
timestamp 1677579658
transform 1 0 9888 0 1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_34_107
timestamp 1677580104
transform 1 0 11424 0 1 26460
box -48 -56 240 834
use sg13g2_decap_4  FILLER_34_130
timestamp 1679577901
transform 1 0 13632 0 1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_34_134
timestamp 1677579658
transform 1 0 14016 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_157
timestamp 1679581782
transform 1 0 16224 0 1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_34_164
timestamp 1677580104
transform 1 0 16896 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_166
timestamp 1677579658
transform 1 0 17088 0 1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_34_198
timestamp 1677580104
transform 1 0 20160 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_48
timestamp 1677579658
transform 1 0 5760 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_66
timestamp 1679581782
transform 1 0 7488 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_35_73
timestamp 1677580104
transform 1 0 8160 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_75
timestamp 1677579658
transform 1 0 8352 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_4  FILLER_35_97
timestamp 1679577901
transform 1 0 10464 0 -1 27972
box -48 -56 432 834
use sg13g2_decap_4  FILLER_35_118
timestamp 1679577901
transform 1 0 12480 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_35_122
timestamp 1677579658
transform 1 0 12864 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_140
timestamp 1679581782
transform 1 0 14592 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_35_147
timestamp 1677580104
transform 1 0 15264 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_149
timestamp 1677579658
transform 1 0 15456 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_4  FILLER_35_170
timestamp 1679577901
transform 1 0 17472 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_35_174
timestamp 1677580104
transform 1 0 17856 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_2  FILLER_35_198
timestamp 1677580104
transform 1 0 20160 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_2  FILLER_36_17
timestamp 1677580104
transform 1 0 2784 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_19
timestamp 1677579658
transform 1 0 2976 0 1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_36_68
timestamp 1677580104
transform 1 0 7680 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_70
timestamp 1677579658
transform 1 0 7872 0 1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_36_88
timestamp 1677580104
transform 1 0 9600 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_112
timestamp 1677579658
transform 1 0 11904 0 1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_36_130
timestamp 1679581782
transform 1 0 13632 0 1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_36_175
timestamp 1677580104
transform 1 0 17952 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_199
timestamp 1677579658
transform 1 0 20256 0 1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_0
timestamp 1679581782
transform 1 0 1152 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_1  FILLER_37_11
timestamp 1677579658
transform 1 0 2208 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_33
timestamp 1679581782
transform 1 0 4320 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_1  FILLER_37_40
timestamp 1677579658
transform 1 0 4992 0 -1 29484
box -48 -56 144 834
use sg13g2_fill_2  FILLER_37_79
timestamp 1677580104
transform 1 0 8736 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_37_108
timestamp 1677580104
transform 1 0 11520 0 -1 29484
box -48 -56 240 834
use sg13g2_decap_8  FILLER_37_131
timestamp 1679581782
transform 1 0 13728 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_1  FILLER_37_155
timestamp 1677579658
transform 1 0 16032 0 -1 29484
box -48 -56 144 834
use sg13g2_fill_1  FILLER_37_174
timestamp 1677579658
transform 1 0 17856 0 -1 29484
box -48 -56 144 834
use sg13g2_fill_1  FILLER_38_17
timestamp 1677579658
transform 1 0 2784 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_52
timestamp 1679581782
transform 1 0 6144 0 1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_38_59
timestamp 1677580104
transform 1 0 6816 0 1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_38_78
timestamp 1677580104
transform 1 0 8640 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_80
timestamp 1677579658
transform 1 0 8832 0 1 29484
box -48 -56 144 834
use sg13g2_fill_1  FILLER_38_95
timestamp 1677579658
transform 1 0 10272 0 1 29484
box -48 -56 144 834
use sg13g2_fill_1  FILLER_38_118
timestamp 1677579658
transform 1 0 12480 0 1 29484
box -48 -56 144 834
use sg13g2_fill_1  FILLER_38_124
timestamp 1677579658
transform 1 0 13056 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_157
timestamp 1679581782
transform 1 0 16224 0 1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_38_164
timestamp 1679577901
transform 1 0 16896 0 1 29484
box -48 -56 432 834
use sg13g2_fill_1  FILLER_38_168
timestamp 1677579658
transform 1 0 17280 0 1 29484
box -48 -56 144 834
use sg13g2_decap_4  FILLER_39_0
timestamp 1679577901
transform 1 0 1152 0 -1 30996
box -48 -56 432 834
use sg13g2_decap_8  FILLER_39_50
timestamp 1679581782
transform 1 0 5952 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_39_57
timestamp 1679577901
transform 1 0 6624 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_39_109
timestamp 1677580104
transform 1 0 11616 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_111
timestamp 1677579658
transform 1 0 11808 0 -1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_39_127
timestamp 1677580104
transform 1 0 13344 0 -1 30996
box -48 -56 240 834
use sg13g2_decap_4  FILLER_39_155
timestamp 1679577901
transform 1 0 16032 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_39_176
timestamp 1677580104
transform 1 0 18048 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_2  FILLER_39_198
timestamp 1677580104
transform 1 0 20160 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_2  FILLER_40_30
timestamp 1677580104
transform 1 0 4032 0 1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_40_32
timestamp 1677579658
transform 1 0 4224 0 1 30996
box -48 -56 144 834
use sg13g2_fill_1  FILLER_40_54
timestamp 1677579658
transform 1 0 6336 0 1 30996
box -48 -56 144 834
use sg13g2_decap_4  FILLER_40_76
timestamp 1679577901
transform 1 0 8448 0 1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_40_80
timestamp 1677580104
transform 1 0 8832 0 1 30996
box -48 -56 240 834
use sg13g2_fill_2  FILLER_40_175
timestamp 1677580104
transform 1 0 17952 0 1 30996
box -48 -56 240 834
use sg13g2_fill_2  FILLER_40_198
timestamp 1677580104
transform 1 0 20160 0 1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_41_0
timestamp 1679581782
transform 1 0 1152 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_41_7
timestamp 1679577901
transform 1 0 1824 0 -1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_41_11
timestamp 1677580104
transform 1 0 2208 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_2  FILLER_41_68
timestamp 1677580104
transform 1 0 7680 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_2  FILLER_41_80
timestamp 1677580104
transform 1 0 8832 0 -1 32508
box -48 -56 240 834
use sg13g2_decap_4  FILLER_41_126
timestamp 1679577901
transform 1 0 13248 0 -1 32508
box -48 -56 432 834
use sg13g2_decap_4  FILLER_41_133
timestamp 1679577901
transform 1 0 13920 0 -1 32508
box -48 -56 432 834
use sg13g2_decap_8  FILLER_41_164
timestamp 1679581782
transform 1 0 16896 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_171
timestamp 1679581782
transform 1 0 17568 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_178
timestamp 1679581782
transform 1 0 18240 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_185
timestamp 1679581782
transform 1 0 18912 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_192
timestamp 1679581782
transform 1 0 19584 0 -1 32508
box -48 -56 720 834
use sg13g2_fill_1  FILLER_41_199
timestamp 1677579658
transform 1 0 20256 0 -1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_0
timestamp 1679581782
transform 1 0 1152 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_7
timestamp 1679581782
transform 1 0 1824 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_35
timestamp 1679581782
transform 1 0 4512 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_42
timestamp 1679581782
transform 1 0 5184 0 1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_42_49
timestamp 1677580104
transform 1 0 5856 0 1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_42_78
timestamp 1679581782
transform 1 0 8640 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_85
timestamp 1679581782
transform 1 0 9312 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_92
timestamp 1679581782
transform 1 0 9984 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_99
timestamp 1679581782
transform 1 0 10656 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_106
timestamp 1679581782
transform 1 0 11328 0 1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_42_113
timestamp 1677580104
transform 1 0 12000 0 1 32508
box -48 -56 240 834
use sg13g2_decap_4  FILLER_42_119
timestamp 1679577901
transform 1 0 12576 0 1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_42_123
timestamp 1677580104
transform 1 0 12960 0 1 32508
box -48 -56 240 834
use sg13g2_decap_4  FILLER_42_150
timestamp 1679577901
transform 1 0 15552 0 1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_42_154
timestamp 1677580104
transform 1 0 15936 0 1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_42_173
timestamp 1679581782
transform 1 0 17760 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_180
timestamp 1679581782
transform 1 0 18432 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_187
timestamp 1679581782
transform 1 0 19104 0 1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_42_194
timestamp 1679577901
transform 1 0 19776 0 1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_42_198
timestamp 1677580104
transform 1 0 20160 0 1 32508
box -48 -56 240 834
use sg13g2_decap_4  FILLER_43_0
timestamp 1679577901
transform 1 0 1152 0 -1 34020
box -48 -56 432 834
use sg13g2_fill_1  FILLER_43_4
timestamp 1677579658
transform 1 0 1536 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_43_22
timestamp 1677580104
transform 1 0 3264 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_2  FILLER_43_29
timestamp 1677580104
transform 1 0 3936 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_2  FILLER_43_48
timestamp 1677580104
transform 1 0 5760 0 -1 34020
box -48 -56 240 834
use sg13g2_decap_4  FILLER_43_70
timestamp 1679577901
transform 1 0 7872 0 -1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_43_113
timestamp 1677580104
transform 1 0 12000 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_43_115
timestamp 1677579658
transform 1 0 12192 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_157
timestamp 1679581782
transform 1 0 16224 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_164
timestamp 1679581782
transform 1 0 16896 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_171
timestamp 1679581782
transform 1 0 17568 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_178
timestamp 1679581782
transform 1 0 18240 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_185
timestamp 1679581782
transform 1 0 18912 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_192
timestamp 1679581782
transform 1 0 19584 0 -1 34020
box -48 -56 720 834
use sg13g2_fill_1  FILLER_43_199
timestamp 1677579658
transform 1 0 20256 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_44_0
timestamp 1679581782
transform 1 0 1152 0 1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_44_7
timestamp 1677580104
transform 1 0 1824 0 1 34020
box -48 -56 240 834
use sg13g2_decap_4  FILLER_44_35
timestamp 1679577901
transform 1 0 4512 0 1 34020
box -48 -56 432 834
use sg13g2_fill_1  FILLER_44_95
timestamp 1677579658
transform 1 0 10272 0 1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_44_156
timestamp 1679581782
transform 1 0 16128 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_163
timestamp 1679581782
transform 1 0 16800 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_170
timestamp 1679581782
transform 1 0 17472 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_177
timestamp 1679581782
transform 1 0 18144 0 1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_44_184
timestamp 1679577901
transform 1 0 18816 0 1 34020
box -48 -56 432 834
use sg13g2_fill_1  FILLER_44_188
timestamp 1677579658
transform 1 0 19200 0 1 34020
box -48 -56 144 834
use sg13g2_decap_4  FILLER_44_196
timestamp 1679577901
transform 1 0 19968 0 1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_45_0
timestamp 1677580104
transform 1 0 1152 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_45_33
timestamp 1677579658
transform 1 0 4320 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_45_51
timestamp 1677580104
transform 1 0 6048 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_45_53
timestamp 1677579658
transform 1 0 6240 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_45_93
timestamp 1677580104
transform 1 0 10080 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_45_95
timestamp 1677579658
transform 1 0 10272 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_45_120
timestamp 1677580104
transform 1 0 12672 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_2  FILLER_45_132
timestamp 1677580104
transform 1 0 13824 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_45_151
timestamp 1679581782
transform 1 0 15648 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_162
timestamp 1679581782
transform 1 0 16704 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_169
timestamp 1679581782
transform 1 0 17376 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_176
timestamp 1679581782
transform 1 0 18048 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_45_183
timestamp 1677580104
transform 1 0 18720 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_45_193
timestamp 1679581782
transform 1 0 19680 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_46_104
timestamp 1677579658
transform 1 0 11136 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_140
timestamp 1679581782
transform 1 0 14592 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_147
timestamp 1679581782
transform 1 0 15264 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_154
timestamp 1679581782
transform 1 0 15936 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_161
timestamp 1679581782
transform 1 0 16608 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_168
timestamp 1679581782
transform 1 0 17280 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_175
timestamp 1679581782
transform 1 0 17952 0 1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_46_182
timestamp 1677580104
transform 1 0 18624 0 1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_46_184
timestamp 1677579658
transform 1 0 18816 0 1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_46_197
timestamp 1677580104
transform 1 0 20064 0 1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_46_199
timestamp 1677579658
transform 1 0 20256 0 1 35532
box -48 -56 144 834
use sg13g2_decap_4  FILLER_47_43
timestamp 1679577901
transform 1 0 5280 0 -1 37044
box -48 -56 432 834
use sg13g2_fill_1  FILLER_47_47
timestamp 1677579658
transform 1 0 5664 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_47_82
timestamp 1679581782
transform 1 0 9024 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_47_89
timestamp 1679577901
transform 1 0 9696 0 -1 37044
box -48 -56 432 834
use sg13g2_fill_1  FILLER_47_93
timestamp 1677579658
transform 1 0 10080 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_47_139
timestamp 1679581782
transform 1 0 14496 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_146
timestamp 1679581782
transform 1 0 15168 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_153
timestamp 1679581782
transform 1 0 15840 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_160
timestamp 1679581782
transform 1 0 16512 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_167
timestamp 1679581782
transform 1 0 17184 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_174
timestamp 1679581782
transform 1 0 17856 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_47_181
timestamp 1679577901
transform 1 0 18528 0 -1 37044
box -48 -56 432 834
use sg13g2_decap_8  FILLER_47_193
timestamp 1679581782
transform 1 0 19680 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_0
timestamp 1679581782
transform 1 0 1152 0 1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_48_7
timestamp 1679577901
transform 1 0 1824 0 1 37044
box -48 -56 432 834
use sg13g2_decap_8  FILLER_48_70
timestamp 1679581782
transform 1 0 7872 0 1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_48_77
timestamp 1679577901
transform 1 0 8544 0 1 37044
box -48 -56 432 834
use sg13g2_decap_4  FILLER_48_98
timestamp 1679577901
transform 1 0 10560 0 1 37044
box -48 -56 432 834
use sg13g2_fill_1  FILLER_48_102
timestamp 1677579658
transform 1 0 10944 0 1 37044
box -48 -56 144 834
use sg13g2_fill_1  FILLER_48_128
timestamp 1677579658
transform 1 0 13440 0 1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_48_146
timestamp 1679581782
transform 1 0 15168 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_153
timestamp 1679581782
transform 1 0 15840 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_160
timestamp 1679581782
transform 1 0 16512 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_167
timestamp 1679581782
transform 1 0 17184 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_174
timestamp 1679581782
transform 1 0 17856 0 1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_48_181
timestamp 1679577901
transform 1 0 18528 0 1 37044
box -48 -56 432 834
use sg13g2_fill_2  FILLER_48_197
timestamp 1677580104
transform 1 0 20064 0 1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_48_199
timestamp 1677579658
transform 1 0 20256 0 1 37044
box -48 -56 144 834
use sg13g2_decap_4  FILLER_49_0
timestamp 1679577901
transform 1 0 1152 0 -1 38556
box -48 -56 432 834
use sg13g2_decap_4  FILLER_49_21
timestamp 1679577901
transform 1 0 3168 0 -1 38556
box -48 -56 432 834
use sg13g2_fill_1  FILLER_49_25
timestamp 1677579658
transform 1 0 3552 0 -1 38556
box -48 -56 144 834
use sg13g2_fill_1  FILLER_49_64
timestamp 1677579658
transform 1 0 7296 0 -1 38556
box -48 -56 144 834
use sg13g2_fill_2  FILLER_49_73
timestamp 1677580104
transform 1 0 8160 0 -1 38556
box -48 -56 240 834
use sg13g2_decap_8  FILLER_49_96
timestamp 1679581782
transform 1 0 10368 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_4  FILLER_49_103
timestamp 1679577901
transform 1 0 11040 0 -1 38556
box -48 -56 432 834
use sg13g2_decap_4  FILLER_49_141
timestamp 1679577901
transform 1 0 14688 0 -1 38556
box -48 -56 432 834
use sg13g2_fill_2  FILLER_49_145
timestamp 1677580104
transform 1 0 15072 0 -1 38556
box -48 -56 240 834
use sg13g2_decap_8  FILLER_49_151
timestamp 1679581782
transform 1 0 15648 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_158
timestamp 1679581782
transform 1 0 16320 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_165
timestamp 1679581782
transform 1 0 16992 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_172
timestamp 1679581782
transform 1 0 17664 0 -1 38556
box -48 -56 720 834
use sg13g2_fill_2  FILLER_49_179
timestamp 1677580104
transform 1 0 18336 0 -1 38556
box -48 -56 240 834
use sg13g2_decap_4  FILLER_49_185
timestamp 1679577901
transform 1 0 18912 0 -1 38556
box -48 -56 432 834
use sg13g2_decap_8  FILLER_49_193
timestamp 1679581782
transform 1 0 19680 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_0
timestamp 1679581782
transform 1 0 1152 0 1 38556
box -48 -56 720 834
use sg13g2_fill_1  FILLER_50_7
timestamp 1677579658
transform 1 0 1824 0 1 38556
box -48 -56 144 834
use sg13g2_decap_8  FILLER_50_97
timestamp 1679581782
transform 1 0 10464 0 1 38556
box -48 -56 720 834
use sg13g2_fill_2  FILLER_50_104
timestamp 1677580104
transform 1 0 11136 0 1 38556
box -48 -56 240 834
use sg13g2_fill_1  FILLER_50_106
timestamp 1677579658
transform 1 0 11328 0 1 38556
box -48 -56 144 834
use sg13g2_decap_8  FILLER_50_129
timestamp 1679581782
transform 1 0 13536 0 1 38556
box -48 -56 720 834
use sg13g2_fill_2  FILLER_50_136
timestamp 1677580104
transform 1 0 14208 0 1 38556
box -48 -56 240 834
use sg13g2_decap_8  FILLER_50_142
timestamp 1679581782
transform 1 0 14784 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_149
timestamp 1679581782
transform 1 0 15456 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_156
timestamp 1679581782
transform 1 0 16128 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_163
timestamp 1679581782
transform 1 0 16800 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_170
timestamp 1679581782
transform 1 0 17472 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_177
timestamp 1679581782
transform 1 0 18144 0 1 38556
box -48 -56 720 834
use sg13g2_decap_4  FILLER_50_184
timestamp 1679577901
transform 1 0 18816 0 1 38556
box -48 -56 432 834
use sg13g2_fill_1  FILLER_50_188
timestamp 1677579658
transform 1 0 19200 0 1 38556
box -48 -56 144 834
use sg13g2_decap_8  FILLER_50_193
timestamp 1679581782
transform 1 0 19680 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_0
timestamp 1679581782
transform 1 0 1152 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_4  FILLER_51_62
timestamp 1679577901
transform 1 0 7104 0 -1 40068
box -48 -56 432 834
use sg13g2_fill_1  FILLER_51_66
timestamp 1677579658
transform 1 0 7488 0 -1 40068
box -48 -56 144 834
use sg13g2_decap_8  FILLER_51_87
timestamp 1679581782
transform 1 0 9504 0 -1 40068
box -48 -56 720 834
use sg13g2_fill_2  FILLER_51_94
timestamp 1677580104
transform 1 0 10176 0 -1 40068
box -48 -56 240 834
use sg13g2_decap_4  FILLER_51_113
timestamp 1679577901
transform 1 0 12000 0 -1 40068
box -48 -56 432 834
use sg13g2_fill_2  FILLER_51_117
timestamp 1677580104
transform 1 0 12384 0 -1 40068
box -48 -56 240 834
use sg13g2_decap_8  FILLER_51_124
timestamp 1679581782
transform 1 0 13056 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_131
timestamp 1679581782
transform 1 0 13728 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_138
timestamp 1679581782
transform 1 0 14400 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_145
timestamp 1679581782
transform 1 0 15072 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_152
timestamp 1679581782
transform 1 0 15744 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_159
timestamp 1679581782
transform 1 0 16416 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_166
timestamp 1679581782
transform 1 0 17088 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_173
timestamp 1679581782
transform 1 0 17760 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_4  FILLER_51_180
timestamp 1679577901
transform 1 0 18432 0 -1 40068
box -48 -56 432 834
use sg13g2_fill_1  FILLER_51_184
timestamp 1677579658
transform 1 0 18816 0 -1 40068
box -48 -56 144 834
use sg13g2_fill_2  FILLER_51_197
timestamp 1677580104
transform 1 0 20064 0 -1 40068
box -48 -56 240 834
use sg13g2_fill_1  FILLER_51_199
timestamp 1677579658
transform 1 0 20256 0 -1 40068
box -48 -56 144 834
use sg13g2_decap_8  FILLER_52_17
timestamp 1679581782
transform 1 0 2784 0 1 40068
box -48 -56 720 834
use sg13g2_decap_4  FILLER_52_24
timestamp 1679577901
transform 1 0 3456 0 1 40068
box -48 -56 432 834
use sg13g2_decap_4  FILLER_52_45
timestamp 1679577901
transform 1 0 5472 0 1 40068
box -48 -56 432 834
use sg13g2_fill_1  FILLER_52_83
timestamp 1677579658
transform 1 0 9120 0 1 40068
box -48 -56 144 834
use sg13g2_decap_8  FILLER_52_105
timestamp 1679581782
transform 1 0 11232 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_112
timestamp 1679581782
transform 1 0 11904 0 1 40068
box -48 -56 720 834
use sg13g2_decap_4  FILLER_52_119
timestamp 1679577901
transform 1 0 12576 0 1 40068
box -48 -56 432 834
use sg13g2_decap_8  FILLER_52_127
timestamp 1679581782
transform 1 0 13344 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_134
timestamp 1679581782
transform 1 0 14016 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_141
timestamp 1679581782
transform 1 0 14688 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_148
timestamp 1679581782
transform 1 0 15360 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_155
timestamp 1679581782
transform 1 0 16032 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_162
timestamp 1679581782
transform 1 0 16704 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_169
timestamp 1679581782
transform 1 0 17376 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_176
timestamp 1679581782
transform 1 0 18048 0 1 40068
box -48 -56 720 834
use sg13g2_fill_1  FILLER_52_183
timestamp 1677579658
transform 1 0 18720 0 1 40068
box -48 -56 144 834
use sg13g2_decap_8  FILLER_53_0
timestamp 1679581782
transform 1 0 1152 0 -1 41580
box -48 -56 720 834
use sg13g2_fill_1  FILLER_53_24
timestamp 1677579658
transform 1 0 3456 0 -1 41580
box -48 -56 144 834
use sg13g2_decap_4  FILLER_53_63
timestamp 1679577901
transform 1 0 7200 0 -1 41580
box -48 -56 432 834
use sg13g2_decap_8  FILLER_53_87
timestamp 1679581782
transform 1 0 9504 0 -1 41580
box -48 -56 720 834
use sg13g2_fill_1  FILLER_53_94
timestamp 1677579658
transform 1 0 10176 0 -1 41580
box -48 -56 144 834
use sg13g2_decap_4  FILLER_53_116
timestamp 1679577901
transform 1 0 12288 0 -1 41580
box -48 -56 432 834
use sg13g2_decap_8  FILLER_53_124
timestamp 1679581782
transform 1 0 13056 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_131
timestamp 1679581782
transform 1 0 13728 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_138
timestamp 1679581782
transform 1 0 14400 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_145
timestamp 1679581782
transform 1 0 15072 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_152
timestamp 1679581782
transform 1 0 15744 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_159
timestamp 1679581782
transform 1 0 16416 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_166
timestamp 1679581782
transform 1 0 17088 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_173
timestamp 1679581782
transform 1 0 17760 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_4  FILLER_53_180
timestamp 1679577901
transform 1 0 18432 0 -1 41580
box -48 -56 432 834
use sg13g2_decap_4  FILLER_53_196
timestamp 1679577901
transform 1 0 19968 0 -1 41580
box -48 -56 432 834
use sg13g2_decap_8  FILLER_54_0
timestamp 1679581782
transform 1 0 1152 0 1 41580
box -48 -56 720 834
use sg13g2_decap_4  FILLER_54_32
timestamp 1679577901
transform 1 0 4224 0 1 41580
box -48 -56 432 834
use sg13g2_fill_2  FILLER_54_36
timestamp 1677580104
transform 1 0 4608 0 1 41580
box -48 -56 240 834
use sg13g2_fill_1  FILLER_54_41
timestamp 1677579658
transform 1 0 5088 0 1 41580
box -48 -56 144 834
use sg13g2_decap_8  FILLER_54_59
timestamp 1679581782
transform 1 0 6816 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_117
timestamp 1679581782
transform 1 0 12384 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_124
timestamp 1679581782
transform 1 0 13056 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_131
timestamp 1679581782
transform 1 0 13728 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_138
timestamp 1679581782
transform 1 0 14400 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_145
timestamp 1679581782
transform 1 0 15072 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_152
timestamp 1679581782
transform 1 0 15744 0 1 41580
box -48 -56 720 834
use sg13g2_decap_4  FILLER_54_159
timestamp 1679577901
transform 1 0 16416 0 1 41580
box -48 -56 432 834
use sg13g2_fill_1  FILLER_54_163
timestamp 1677579658
transform 1 0 16800 0 1 41580
box -48 -56 144 834
use sg13g2_decap_8  FILLER_54_168
timestamp 1679581782
transform 1 0 17280 0 1 41580
box -48 -56 720 834
use sg13g2_fill_2  FILLER_54_175
timestamp 1677580104
transform 1 0 17952 0 1 41580
box -48 -56 240 834
use sg13g2_fill_1  FILLER_54_177
timestamp 1677579658
transform 1 0 18144 0 1 41580
box -48 -56 144 834
use sg13g2_fill_2  FILLER_54_198
timestamp 1677580104
transform 1 0 20160 0 1 41580
box -48 -56 240 834
use sg13g2_decap_4  FILLER_55_17
timestamp 1679577901
transform 1 0 2784 0 -1 43092
box -48 -56 432 834
use sg13g2_decap_8  FILLER_55_59
timestamp 1679581782
transform 1 0 6816 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_4  FILLER_55_66
timestamp 1679577901
transform 1 0 7488 0 -1 43092
box -48 -56 432 834
use sg13g2_fill_2  FILLER_55_70
timestamp 1677580104
transform 1 0 7872 0 -1 43092
box -48 -56 240 834
use sg13g2_decap_8  FILLER_55_89
timestamp 1679581782
transform 1 0 9696 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_96
timestamp 1679581782
transform 1 0 10368 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_103
timestamp 1679581782
transform 1 0 11040 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_4  FILLER_55_110
timestamp 1679577901
transform 1 0 11712 0 -1 43092
box -48 -56 432 834
use sg13g2_fill_2  FILLER_55_114
timestamp 1677580104
transform 1 0 12096 0 -1 43092
box -48 -56 240 834
use sg13g2_decap_8  FILLER_55_133
timestamp 1679581782
transform 1 0 13920 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_140
timestamp 1679581782
transform 1 0 14592 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_147
timestamp 1679581782
transform 1 0 15264 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_154
timestamp 1679581782
transform 1 0 15936 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_161
timestamp 1679581782
transform 1 0 16608 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_168
timestamp 1679581782
transform 1 0 17280 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_4  FILLER_55_175
timestamp 1679577901
transform 1 0 17952 0 -1 43092
box -48 -56 432 834
use sg13g2_fill_2  FILLER_55_179
timestamp 1677580104
transform 1 0 18336 0 -1 43092
box -48 -56 240 834
use sg13g2_fill_2  FILLER_55_197
timestamp 1677580104
transform 1 0 20064 0 -1 43092
box -48 -56 240 834
use sg13g2_fill_1  FILLER_55_199
timestamp 1677579658
transform 1 0 20256 0 -1 43092
box -48 -56 144 834
use sg13g2_decap_8  FILLER_56_0
timestamp 1679581782
transform 1 0 1152 0 1 43092
box -48 -56 720 834
use sg13g2_decap_4  FILLER_56_7
timestamp 1679577901
transform 1 0 1824 0 1 43092
box -48 -56 432 834
use sg13g2_fill_2  FILLER_56_11
timestamp 1677580104
transform 1 0 2208 0 1 43092
box -48 -56 240 834
use sg13g2_decap_8  FILLER_56_34
timestamp 1679581782
transform 1 0 4416 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_41
timestamp 1679581782
transform 1 0 5088 0 1 43092
box -48 -56 720 834
use sg13g2_decap_4  FILLER_56_48
timestamp 1679577901
transform 1 0 5760 0 1 43092
box -48 -56 432 834
use sg13g2_fill_1  FILLER_56_90
timestamp 1677579658
transform 1 0 9792 0 1 43092
box -48 -56 144 834
use sg13g2_fill_2  FILLER_56_129
timestamp 1677580104
transform 1 0 13536 0 1 43092
box -48 -56 240 834
use sg13g2_fill_1  FILLER_56_131
timestamp 1677579658
transform 1 0 13728 0 1 43092
box -48 -56 144 834
use sg13g2_decap_4  FILLER_56_136
timestamp 1679577901
transform 1 0 14208 0 1 43092
box -48 -56 432 834
use sg13g2_fill_2  FILLER_56_140
timestamp 1677580104
transform 1 0 14592 0 1 43092
box -48 -56 240 834
use sg13g2_decap_4  FILLER_56_146
timestamp 1679577901
transform 1 0 15168 0 1 43092
box -48 -56 432 834
use sg13g2_fill_2  FILLER_56_150
timestamp 1677580104
transform 1 0 15552 0 1 43092
box -48 -56 240 834
use sg13g2_decap_8  FILLER_56_177
timestamp 1679581782
transform 1 0 18144 0 1 43092
box -48 -56 720 834
use sg13g2_fill_1  FILLER_56_184
timestamp 1677579658
transform 1 0 18816 0 1 43092
box -48 -56 144 834
use sg13g2_decap_8  FILLER_56_193
timestamp 1679581782
transform 1 0 19680 0 1 43092
box -48 -56 720 834
use sg13g2_decap_4  FILLER_57_0
timestamp 1679577901
transform 1 0 1152 0 -1 44604
box -48 -56 432 834
use sg13g2_fill_2  FILLER_57_4
timestamp 1677580104
transform 1 0 1536 0 -1 44604
box -48 -56 240 834
use sg13g2_decap_8  FILLER_57_65
timestamp 1679581782
transform 1 0 7392 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_72
timestamp 1679581782
transform 1 0 8064 0 -1 44604
box -48 -56 720 834
use sg13g2_fill_2  FILLER_57_79
timestamp 1677580104
transform 1 0 8736 0 -1 44604
box -48 -56 240 834
use sg13g2_fill_2  FILLER_57_85
timestamp 1677580104
transform 1 0 9312 0 -1 44604
box -48 -56 240 834
use sg13g2_fill_1  FILLER_57_87
timestamp 1677579658
transform 1 0 9504 0 -1 44604
box -48 -56 144 834
use sg13g2_fill_2  FILLER_57_130
timestamp 1677580104
transform 1 0 13632 0 -1 44604
box -48 -56 240 834
use sg13g2_fill_1  FILLER_57_132
timestamp 1677579658
transform 1 0 13824 0 -1 44604
box -48 -56 144 834
use sg13g2_decap_4  FILLER_57_171
timestamp 1679577901
transform 1 0 17568 0 -1 44604
box -48 -56 432 834
use sg13g2_fill_1  FILLER_57_175
timestamp 1677579658
transform 1 0 17952 0 -1 44604
box -48 -56 144 834
use sg13g2_fill_2  FILLER_57_197
timestamp 1677580104
transform 1 0 20064 0 -1 44604
box -48 -56 240 834
use sg13g2_fill_1  FILLER_57_199
timestamp 1677579658
transform 1 0 20256 0 -1 44604
box -48 -56 144 834
use sg13g2_fill_2  FILLER_58_0
timestamp 1677580104
transform 1 0 1152 0 1 44604
box -48 -56 240 834
use sg13g2_fill_1  FILLER_58_2
timestamp 1677579658
transform 1 0 1344 0 1 44604
box -48 -56 144 834
use sg13g2_fill_1  FILLER_58_11
timestamp 1677579658
transform 1 0 2208 0 1 44604
box -48 -56 144 834
use sg13g2_decap_8  FILLER_58_33
timestamp 1679581782
transform 1 0 4320 0 1 44604
box -48 -56 720 834
use sg13g2_decap_4  FILLER_58_40
timestamp 1679577901
transform 1 0 4992 0 1 44604
box -48 -56 432 834
use sg13g2_fill_1  FILLER_58_44
timestamp 1677579658
transform 1 0 5376 0 1 44604
box -48 -56 144 834
use sg13g2_decap_4  FILLER_58_66
timestamp 1679577901
transform 1 0 7488 0 1 44604
box -48 -56 432 834
use sg13g2_decap_8  FILLER_58_104
timestamp 1679581782
transform 1 0 11136 0 1 44604
box -48 -56 720 834
use sg13g2_fill_2  FILLER_58_111
timestamp 1677580104
transform 1 0 11808 0 1 44604
box -48 -56 240 834
use sg13g2_decap_8  FILLER_58_134
timestamp 1679581782
transform 1 0 14016 0 1 44604
box -48 -56 720 834
use sg13g2_decap_4  FILLER_58_141
timestamp 1679577901
transform 1 0 14688 0 1 44604
box -48 -56 432 834
use sg13g2_fill_1  FILLER_58_145
timestamp 1677579658
transform 1 0 15072 0 1 44604
box -48 -56 144 834
use sg13g2_decap_4  FILLER_58_167
timestamp 1679577901
transform 1 0 17184 0 1 44604
box -48 -56 432 834
use sg13g2_fill_2  FILLER_58_171
timestamp 1677580104
transform 1 0 17568 0 1 44604
box -48 -56 240 834
use sg13g2_fill_2  FILLER_58_198
timestamp 1677580104
transform 1 0 20160 0 1 44604
box -48 -56 240 834
use sg13g2_fill_2  FILLER_59_0
timestamp 1677580104
transform 1 0 1152 0 -1 46116
box -48 -56 240 834
use sg13g2_fill_1  FILLER_59_2
timestamp 1677579658
transform 1 0 1344 0 -1 46116
box -48 -56 144 834
use sg13g2_fill_2  FILLER_59_11
timestamp 1677580104
transform 1 0 2208 0 -1 46116
box -48 -56 240 834
use sg13g2_decap_4  FILLER_59_47
timestamp 1679577901
transform 1 0 5664 0 -1 46116
box -48 -56 432 834
use sg13g2_fill_2  FILLER_59_51
timestamp 1677580104
transform 1 0 6048 0 -1 46116
box -48 -56 240 834
use sg13g2_decap_8  FILLER_59_70
timestamp 1679581782
transform 1 0 7872 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_77
timestamp 1679581782
transform 1 0 8544 0 -1 46116
box -48 -56 720 834
use sg13g2_fill_1  FILLER_59_84
timestamp 1677579658
transform 1 0 9216 0 -1 46116
box -48 -56 144 834
use sg13g2_decap_8  FILLER_59_110
timestamp 1679581782
transform 1 0 11712 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_4  FILLER_59_117
timestamp 1679577901
transform 1 0 12384 0 -1 46116
box -48 -56 432 834
use sg13g2_fill_1  FILLER_59_121
timestamp 1677579658
transform 1 0 12768 0 -1 46116
box -48 -56 144 834
use sg13g2_fill_1  FILLER_59_126
timestamp 1677579658
transform 1 0 13248 0 -1 46116
box -48 -56 144 834
use sg13g2_fill_1  FILLER_59_182
timestamp 1677579658
transform 1 0 18624 0 -1 46116
box -48 -56 144 834
use sg13g2_decap_4  FILLER_59_195
timestamp 1679577901
transform 1 0 19872 0 -1 46116
box -48 -56 432 834
use sg13g2_fill_1  FILLER_59_199
timestamp 1677579658
transform 1 0 20256 0 -1 46116
box -48 -56 144 834
use sg13g2_decap_8  FILLER_60_17
timestamp 1679581782
transform 1 0 2784 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_24
timestamp 1679581782
transform 1 0 3456 0 1 46116
box -48 -56 720 834
use sg13g2_fill_2  FILLER_60_31
timestamp 1677580104
transform 1 0 4128 0 1 46116
box -48 -56 240 834
use sg13g2_fill_1  FILLER_60_33
timestamp 1677579658
transform 1 0 4320 0 1 46116
box -48 -56 144 834
use sg13g2_decap_4  FILLER_60_68
timestamp 1679577901
transform 1 0 7680 0 1 46116
box -48 -56 432 834
use sg13g2_fill_1  FILLER_60_110
timestamp 1677579658
transform 1 0 11712 0 1 46116
box -48 -56 144 834
use sg13g2_fill_2  FILLER_60_115
timestamp 1677580104
transform 1 0 12192 0 1 46116
box -48 -56 240 834
use sg13g2_decap_8  FILLER_60_138
timestamp 1679581782
transform 1 0 14400 0 1 46116
box -48 -56 720 834
use sg13g2_fill_1  FILLER_60_145
timestamp 1677579658
transform 1 0 15072 0 1 46116
box -48 -56 144 834
use sg13g2_decap_8  FILLER_60_163
timestamp 1679581782
transform 1 0 16800 0 1 46116
box -48 -56 720 834
use sg13g2_fill_2  FILLER_60_170
timestamp 1677580104
transform 1 0 17472 0 1 46116
box -48 -56 240 834
use sg13g2_fill_1  FILLER_60_172
timestamp 1677579658
transform 1 0 17664 0 1 46116
box -48 -56 144 834
use sg13g2_fill_2  FILLER_60_198
timestamp 1677580104
transform 1 0 20160 0 1 46116
box -48 -56 240 834
use sg13g2_decap_4  FILLER_61_0
timestamp 1679577901
transform 1 0 1152 0 -1 47628
box -48 -56 432 834
use sg13g2_fill_2  FILLER_61_4
timestamp 1677580104
transform 1 0 1536 0 -1 47628
box -48 -56 240 834
use sg13g2_decap_8  FILLER_61_31
timestamp 1679581782
transform 1 0 4128 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_59
timestamp 1679581782
transform 1 0 6816 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_4  FILLER_61_66
timestamp 1679577901
transform 1 0 7488 0 -1 47628
box -48 -56 432 834
use sg13g2_fill_1  FILLER_61_70
timestamp 1677579658
transform 1 0 7872 0 -1 47628
box -48 -56 144 834
use sg13g2_decap_8  FILLER_61_88
timestamp 1679581782
transform 1 0 9600 0 -1 47628
box -48 -56 720 834
use sg13g2_fill_2  FILLER_61_95
timestamp 1677580104
transform 1 0 10272 0 -1 47628
box -48 -56 240 834
use sg13g2_fill_1  FILLER_61_97
timestamp 1677579658
transform 1 0 10464 0 -1 47628
box -48 -56 144 834
use sg13g2_fill_1  FILLER_61_102
timestamp 1677579658
transform 1 0 10944 0 -1 47628
box -48 -56 144 834
use sg13g2_decap_4  FILLER_61_137
timestamp 1679577901
transform 1 0 14304 0 -1 47628
box -48 -56 432 834
use sg13g2_fill_2  FILLER_61_141
timestamp 1677580104
transform 1 0 14688 0 -1 47628
box -48 -56 240 834
use sg13g2_fill_2  FILLER_61_198
timestamp 1677580104
transform 1 0 20160 0 -1 47628
box -48 -56 240 834
use sg13g2_decap_4  FILLER_62_0
timestamp 1679577901
transform 1 0 1152 0 1 47628
box -48 -56 432 834
use sg13g2_decap_4  FILLER_62_63
timestamp 1679577901
transform 1 0 7200 0 1 47628
box -48 -56 432 834
use sg13g2_fill_1  FILLER_62_67
timestamp 1677579658
transform 1 0 7584 0 1 47628
box -48 -56 144 834
use sg13g2_decap_4  FILLER_62_89
timestamp 1679577901
transform 1 0 9696 0 1 47628
box -48 -56 432 834
use sg13g2_fill_1  FILLER_62_93
timestamp 1677579658
transform 1 0 10080 0 1 47628
box -48 -56 144 834
use sg13g2_decap_8  FILLER_62_111
timestamp 1679581782
transform 1 0 11808 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_118
timestamp 1679581782
transform 1 0 12480 0 1 47628
box -48 -56 720 834
use sg13g2_decap_4  FILLER_62_125
timestamp 1679577901
transform 1 0 13152 0 1 47628
box -48 -56 432 834
use sg13g2_decap_8  FILLER_62_146
timestamp 1679581782
transform 1 0 15168 0 1 47628
box -48 -56 720 834
use sg13g2_fill_2  FILLER_62_153
timestamp 1677580104
transform 1 0 15840 0 1 47628
box -48 -56 240 834
use sg13g2_fill_1  FILLER_62_155
timestamp 1677579658
transform 1 0 16032 0 1 47628
box -48 -56 144 834
use sg13g2_fill_2  FILLER_62_198
timestamp 1677580104
transform 1 0 20160 0 1 47628
box -48 -56 240 834
use sg13g2_fill_2  FILLER_63_21
timestamp 1677580104
transform 1 0 3168 0 -1 49140
box -48 -56 240 834
use sg13g2_fill_1  FILLER_63_57
timestamp 1677579658
transform 1 0 6624 0 -1 49140
box -48 -56 144 834
use sg13g2_fill_2  FILLER_63_75
timestamp 1677580104
transform 1 0 8352 0 -1 49140
box -48 -56 240 834
use sg13g2_fill_1  FILLER_63_77
timestamp 1677579658
transform 1 0 8544 0 -1 49140
box -48 -56 144 834
use sg13g2_decap_8  FILLER_63_99
timestamp 1679581782
transform 1 0 10656 0 -1 49140
box -48 -56 720 834
use sg13g2_fill_1  FILLER_63_106
timestamp 1677579658
transform 1 0 11328 0 -1 49140
box -48 -56 144 834
use sg13g2_decap_4  FILLER_63_145
timestamp 1679577901
transform 1 0 15072 0 -1 49140
box -48 -56 432 834
use sg13g2_fill_1  FILLER_63_149
timestamp 1677579658
transform 1 0 15456 0 -1 49140
box -48 -56 144 834
use sg13g2_decap_8  FILLER_63_167
timestamp 1679581782
transform 1 0 17184 0 -1 49140
box -48 -56 720 834
use sg13g2_fill_1  FILLER_63_199
timestamp 1677579658
transform 1 0 20256 0 -1 49140
box -48 -56 144 834
use sg13g2_fill_2  FILLER_64_0
timestamp 1677580104
transform 1 0 1152 0 1 49140
box -48 -56 240 834
use sg13g2_fill_1  FILLER_64_2
timestamp 1677579658
transform 1 0 1344 0 1 49140
box -48 -56 144 834
use sg13g2_decap_8  FILLER_64_32
timestamp 1679581782
transform 1 0 4224 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_39
timestamp 1679581782
transform 1 0 4896 0 1 49140
box -48 -56 720 834
use sg13g2_fill_2  FILLER_64_46
timestamp 1677580104
transform 1 0 5568 0 1 49140
box -48 -56 240 834
use sg13g2_decap_8  FILLER_64_82
timestamp 1679581782
transform 1 0 9024 0 1 49140
box -48 -56 720 834
use sg13g2_fill_1  FILLER_64_89
timestamp 1677579658
transform 1 0 9696 0 1 49140
box -48 -56 144 834
use sg13g2_fill_1  FILLER_64_145
timestamp 1677579658
transform 1 0 15072 0 1 49140
box -48 -56 144 834
use sg13g2_fill_1  FILLER_64_184
timestamp 1677579658
transform 1 0 18816 0 1 49140
box -48 -56 144 834
use sg13g2_fill_2  FILLER_64_197
timestamp 1677580104
transform 1 0 20064 0 1 49140
box -48 -56 240 834
use sg13g2_fill_1  FILLER_64_199
timestamp 1677579658
transform 1 0 20256 0 1 49140
box -48 -56 144 834
use sg13g2_fill_2  FILLER_65_0
timestamp 1677580104
transform 1 0 1152 0 -1 50652
box -48 -56 240 834
use sg13g2_decap_8  FILLER_65_57
timestamp 1679581782
transform 1 0 6624 0 -1 50652
box -48 -56 720 834
use sg13g2_fill_2  FILLER_65_64
timestamp 1677580104
transform 1 0 7296 0 -1 50652
box -48 -56 240 834
use sg13g2_decap_8  FILLER_65_100
timestamp 1679581782
transform 1 0 10752 0 -1 50652
box -48 -56 720 834
use sg13g2_fill_1  FILLER_65_107
timestamp 1677579658
transform 1 0 11424 0 -1 50652
box -48 -56 144 834
use sg13g2_decap_4  FILLER_65_129
timestamp 1679577901
transform 1 0 13536 0 -1 50652
box -48 -56 432 834
use sg13g2_fill_2  FILLER_65_150
timestamp 1677580104
transform 1 0 15552 0 -1 50652
box -48 -56 240 834
use sg13g2_fill_2  FILLER_65_198
timestamp 1677580104
transform 1 0 20160 0 -1 50652
box -48 -56 240 834
use sg13g2_fill_1  FILLER_66_21
timestamp 1677579658
transform 1 0 3168 0 1 50652
box -48 -56 144 834
use sg13g2_fill_2  FILLER_66_39
timestamp 1677580104
transform 1 0 4896 0 1 50652
box -48 -56 240 834
use sg13g2_fill_1  FILLER_66_41
timestamp 1677579658
transform 1 0 5088 0 1 50652
box -48 -56 144 834
use sg13g2_fill_2  FILLER_66_63
timestamp 1677580104
transform 1 0 7200 0 1 50652
box -48 -56 240 834
use sg13g2_decap_8  FILLER_66_86
timestamp 1679581782
transform 1 0 9408 0 1 50652
box -48 -56 720 834
use sg13g2_fill_2  FILLER_66_93
timestamp 1677580104
transform 1 0 10080 0 1 50652
box -48 -56 240 834
use sg13g2_decap_4  FILLER_66_120
timestamp 1679577901
transform 1 0 12672 0 1 50652
box -48 -56 432 834
use sg13g2_decap_8  FILLER_66_145
timestamp 1679581782
transform 1 0 15072 0 1 50652
box -48 -56 720 834
use sg13g2_decap_4  FILLER_66_152
timestamp 1679577901
transform 1 0 15744 0 1 50652
box -48 -56 432 834
use sg13g2_fill_1  FILLER_66_173
timestamp 1677579658
transform 1 0 17760 0 1 50652
box -48 -56 144 834
use sg13g2_fill_1  FILLER_66_199
timestamp 1677579658
transform 1 0 20256 0 1 50652
box -48 -56 144 834
use sg13g2_fill_2  FILLER_67_0
timestamp 1677580104
transform 1 0 1152 0 -1 52164
box -48 -56 240 834
use sg13g2_fill_1  FILLER_67_2
timestamp 1677579658
transform 1 0 1344 0 -1 52164
box -48 -56 144 834
use sg13g2_fill_1  FILLER_67_11
timestamp 1677579658
transform 1 0 2208 0 -1 52164
box -48 -56 144 834
use sg13g2_decap_8  FILLER_67_33
timestamp 1679581782
transform 1 0 4320 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_40
timestamp 1679581782
transform 1 0 4992 0 -1 52164
box -48 -56 720 834
use sg13g2_fill_2  FILLER_67_47
timestamp 1677580104
transform 1 0 5664 0 -1 52164
box -48 -56 240 834
use sg13g2_decap_8  FILLER_67_66
timestamp 1679581782
transform 1 0 7488 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_4  FILLER_67_73
timestamp 1679577901
transform 1 0 8160 0 -1 52164
box -48 -56 432 834
use sg13g2_decap_4  FILLER_67_145
timestamp 1679577901
transform 1 0 15072 0 -1 52164
box -48 -56 432 834
use sg13g2_fill_1  FILLER_67_149
timestamp 1677579658
transform 1 0 15456 0 -1 52164
box -48 -56 144 834
use sg13g2_decap_4  FILLER_67_171
timestamp 1679577901
transform 1 0 17568 0 -1 52164
box -48 -56 432 834
use sg13g2_fill_2  FILLER_67_175
timestamp 1677580104
transform 1 0 17952 0 -1 52164
box -48 -56 240 834
use sg13g2_fill_2  FILLER_67_198
timestamp 1677580104
transform 1 0 20160 0 -1 52164
box -48 -56 240 834
use sg13g2_fill_2  FILLER_68_0
timestamp 1677580104
transform 1 0 1152 0 1 52164
box -48 -56 240 834
use sg13g2_decap_8  FILLER_68_44
timestamp 1679581782
transform 1 0 5376 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_51
timestamp 1679581782
transform 1 0 6048 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_79
timestamp 1679581782
transform 1 0 8736 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_86
timestamp 1679581782
transform 1 0 9408 0 1 52164
box -48 -56 720 834
use sg13g2_fill_1  FILLER_68_93
timestamp 1677579658
transform 1 0 10080 0 1 52164
box -48 -56 144 834
use sg13g2_fill_2  FILLER_68_115
timestamp 1677580104
transform 1 0 12192 0 1 52164
box -48 -56 240 834
use sg13g2_fill_1  FILLER_68_117
timestamp 1677579658
transform 1 0 12384 0 1 52164
box -48 -56 144 834
use sg13g2_decap_8  FILLER_68_156
timestamp 1679581782
transform 1 0 16128 0 1 52164
box -48 -56 720 834
use sg13g2_decap_4  FILLER_68_163
timestamp 1679577901
transform 1 0 16800 0 1 52164
box -48 -56 432 834
use sg13g2_fill_2  FILLER_68_167
timestamp 1677580104
transform 1 0 17184 0 1 52164
box -48 -56 240 834
use sg13g2_fill_2  FILLER_68_186
timestamp 1677580104
transform 1 0 19008 0 1 52164
box -48 -56 240 834
use sg13g2_fill_1  FILLER_68_188
timestamp 1677579658
transform 1 0 19200 0 1 52164
box -48 -56 144 834
use sg13g2_fill_2  FILLER_68_197
timestamp 1677580104
transform 1 0 20064 0 1 52164
box -48 -56 240 834
use sg13g2_fill_1  FILLER_68_199
timestamp 1677579658
transform 1 0 20256 0 1 52164
box -48 -56 144 834
use sg13g2_fill_2  FILLER_69_0
timestamp 1677580104
transform 1 0 1152 0 -1 53676
box -48 -56 240 834
use sg13g2_fill_1  FILLER_69_2
timestamp 1677579658
transform 1 0 1344 0 -1 53676
box -48 -56 144 834
use sg13g2_decap_8  FILLER_69_41
timestamp 1679581782
transform 1 0 5088 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_137
timestamp 1679581782
transform 1 0 14304 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_169
timestamp 1679581782
transform 1 0 17376 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_4  FILLER_69_176
timestamp 1679577901
transform 1 0 18048 0 -1 53676
box -48 -56 432 834
use sg13g2_fill_2  FILLER_69_197
timestamp 1677580104
transform 1 0 20064 0 -1 53676
box -48 -56 240 834
use sg13g2_fill_1  FILLER_69_199
timestamp 1677579658
transform 1 0 20256 0 -1 53676
box -48 -56 144 834
use sg13g2_decap_4  FILLER_70_17
timestamp 1679577901
transform 1 0 2784 0 1 53676
box -48 -56 432 834
use sg13g2_decap_8  FILLER_70_42
timestamp 1679581782
transform 1 0 5184 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_49
timestamp 1679581782
transform 1 0 5856 0 1 53676
box -48 -56 720 834
use sg13g2_fill_1  FILLER_70_56
timestamp 1677579658
transform 1 0 6528 0 1 53676
box -48 -56 144 834
use sg13g2_decap_8  FILLER_70_116
timestamp 1679581782
transform 1 0 12288 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_123
timestamp 1679581782
transform 1 0 12960 0 1 53676
box -48 -56 720 834
use sg13g2_fill_1  FILLER_70_130
timestamp 1677579658
transform 1 0 13632 0 1 53676
box -48 -56 144 834
use sg13g2_fill_1  FILLER_70_148
timestamp 1677579658
transform 1 0 15360 0 1 53676
box -48 -56 144 834
use sg13g2_fill_2  FILLER_70_170
timestamp 1677580104
transform 1 0 17472 0 1 53676
box -48 -56 240 834
use sg13g2_fill_1  FILLER_70_172
timestamp 1677579658
transform 1 0 17664 0 1 53676
box -48 -56 144 834
use sg13g2_fill_2  FILLER_70_198
timestamp 1677580104
transform 1 0 20160 0 1 53676
box -48 -56 240 834
use sg13g2_decap_4  FILLER_71_0
timestamp 1679577901
transform 1 0 1152 0 -1 55188
box -48 -56 432 834
use sg13g2_fill_2  FILLER_71_4
timestamp 1677580104
transform 1 0 1536 0 -1 55188
box -48 -56 240 834
use sg13g2_decap_8  FILLER_71_31
timestamp 1679581782
transform 1 0 4128 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_4  FILLER_71_38
timestamp 1679577901
transform 1 0 4800 0 -1 55188
box -48 -56 432 834
use sg13g2_fill_2  FILLER_71_42
timestamp 1677580104
transform 1 0 5184 0 -1 55188
box -48 -56 240 834
use sg13g2_decap_8  FILLER_71_61
timestamp 1679581782
transform 1 0 7008 0 -1 55188
box -48 -56 720 834
use sg13g2_fill_2  FILLER_71_68
timestamp 1677580104
transform 1 0 7680 0 -1 55188
box -48 -56 240 834
use sg13g2_fill_1  FILLER_71_104
timestamp 1677579658
transform 1 0 11136 0 -1 55188
box -48 -56 144 834
use sg13g2_fill_2  FILLER_71_164
timestamp 1677580104
transform 1 0 16896 0 -1 55188
box -48 -56 240 834
use sg13g2_fill_1  FILLER_71_166
timestamp 1677579658
transform 1 0 17088 0 -1 55188
box -48 -56 144 834
use sg13g2_fill_2  FILLER_72_0
timestamp 1677580104
transform 1 0 1152 0 1 55188
box -48 -56 240 834
use sg13g2_decap_8  FILLER_72_61
timestamp 1679581782
transform 1 0 7008 0 1 55188
box -48 -56 720 834
use sg13g2_fill_1  FILLER_72_68
timestamp 1677579658
transform 1 0 7680 0 1 55188
box -48 -56 144 834
use sg13g2_decap_4  FILLER_72_94
timestamp 1679577901
transform 1 0 10176 0 1 55188
box -48 -56 432 834
use sg13g2_decap_4  FILLER_72_119
timestamp 1679577901
transform 1 0 12576 0 1 55188
box -48 -56 432 834
use sg13g2_fill_1  FILLER_72_123
timestamp 1677579658
transform 1 0 12960 0 1 55188
box -48 -56 144 834
use sg13g2_fill_2  FILLER_72_141
timestamp 1677580104
transform 1 0 14688 0 1 55188
box -48 -56 240 834
use sg13g2_fill_1  FILLER_72_143
timestamp 1677579658
transform 1 0 14880 0 1 55188
box -48 -56 144 834
use sg13g2_decap_8  FILLER_72_178
timestamp 1679581782
transform 1 0 18240 0 1 55188
box -48 -56 720 834
use sg13g2_decap_4  FILLER_72_185
timestamp 1679577901
transform 1 0 18912 0 1 55188
box -48 -56 432 834
use sg13g2_decap_8  FILLER_72_193
timestamp 1679581782
transform 1 0 19680 0 1 55188
box -48 -56 720 834
use sg13g2_fill_2  FILLER_73_0
timestamp 1677580104
transform 1 0 1152 0 -1 56700
box -48 -56 240 834
use sg13g2_decap_8  FILLER_73_40
timestamp 1679581782
transform 1 0 4992 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_85
timestamp 1679581782
transform 1 0 9312 0 -1 56700
box -48 -56 720 834
use sg13g2_fill_2  FILLER_73_92
timestamp 1677580104
transform 1 0 9984 0 -1 56700
box -48 -56 240 834
use sg13g2_fill_1  FILLER_73_94
timestamp 1677579658
transform 1 0 10176 0 -1 56700
box -48 -56 144 834
use sg13g2_decap_4  FILLER_73_120
timestamp 1679577901
transform 1 0 12672 0 -1 56700
box -48 -56 432 834
use sg13g2_fill_1  FILLER_73_124
timestamp 1677579658
transform 1 0 13056 0 -1 56700
box -48 -56 144 834
use sg13g2_fill_1  FILLER_73_167
timestamp 1677579658
transform 1 0 17184 0 -1 56700
box -48 -56 144 834
use sg13g2_decap_8  FILLER_73_193
timestamp 1679581782
transform 1 0 19680 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_4  FILLER_74_0
timestamp 1679577901
transform 1 0 1152 0 1 56700
box -48 -56 432 834
use sg13g2_fill_2  FILLER_74_4
timestamp 1677580104
transform 1 0 1536 0 1 56700
box -48 -56 240 834
use sg13g2_decap_4  FILLER_74_82
timestamp 1679577901
transform 1 0 9024 0 1 56700
box -48 -56 432 834
use sg13g2_fill_2  FILLER_74_128
timestamp 1677580104
transform 1 0 13440 0 1 56700
box -48 -56 240 834
use sg13g2_fill_1  FILLER_74_151
timestamp 1677579658
transform 1 0 15648 0 1 56700
box -48 -56 144 834
use sg13g2_fill_1  FILLER_74_156
timestamp 1677579658
transform 1 0 16128 0 1 56700
box -48 -56 144 834
use sg13g2_fill_1  FILLER_74_199
timestamp 1677579658
transform 1 0 20256 0 1 56700
box -48 -56 144 834
use sg13g2_decap_8  FILLER_75_0
timestamp 1679581782
transform 1 0 1152 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_45
timestamp 1679581782
transform 1 0 5472 0 -1 58212
box -48 -56 720 834
use sg13g2_fill_1  FILLER_75_52
timestamp 1677579658
transform 1 0 6144 0 -1 58212
box -48 -56 144 834
use sg13g2_decap_4  FILLER_75_70
timestamp 1679577901
transform 1 0 7872 0 -1 58212
box -48 -56 432 834
use sg13g2_decap_8  FILLER_75_95
timestamp 1679581782
transform 1 0 10272 0 -1 58212
box -48 -56 720 834
use sg13g2_fill_2  FILLER_75_102
timestamp 1677580104
transform 1 0 10944 0 -1 58212
box -48 -56 240 834
use sg13g2_fill_1  FILLER_75_104
timestamp 1677579658
transform 1 0 11136 0 -1 58212
box -48 -56 144 834
use sg13g2_decap_8  FILLER_75_143
timestamp 1679581782
transform 1 0 14880 0 -1 58212
box -48 -56 720 834
use sg13g2_fill_2  FILLER_75_150
timestamp 1677580104
transform 1 0 15552 0 -1 58212
box -48 -56 240 834
use sg13g2_fill_1  FILLER_75_152
timestamp 1677579658
transform 1 0 15744 0 -1 58212
box -48 -56 144 834
use sg13g2_decap_8  FILLER_75_173
timestamp 1679581782
transform 1 0 17760 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_180
timestamp 1679581782
transform 1 0 18432 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_187
timestamp 1679581782
transform 1 0 19104 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_4  FILLER_75_194
timestamp 1679577901
transform 1 0 19776 0 -1 58212
box -48 -56 432 834
use sg13g2_fill_2  FILLER_75_198
timestamp 1677580104
transform 1 0 20160 0 -1 58212
box -48 -56 240 834
use sg13g2_decap_8  FILLER_76_17
timestamp 1679581782
transform 1 0 2784 0 1 58212
box -48 -56 720 834
use sg13g2_fill_2  FILLER_76_24
timestamp 1677580104
transform 1 0 3456 0 1 58212
box -48 -56 240 834
use sg13g2_decap_4  FILLER_76_60
timestamp 1679577901
transform 1 0 6912 0 1 58212
box -48 -56 432 834
use sg13g2_decap_4  FILLER_76_98
timestamp 1679577901
transform 1 0 10560 0 1 58212
box -48 -56 432 834
use sg13g2_fill_1  FILLER_76_102
timestamp 1677579658
transform 1 0 10944 0 1 58212
box -48 -56 144 834
use sg13g2_fill_1  FILLER_76_133
timestamp 1677579658
transform 1 0 13920 0 1 58212
box -48 -56 144 834
use sg13g2_fill_1  FILLER_76_151
timestamp 1677579658
transform 1 0 15648 0 1 58212
box -48 -56 144 834
use sg13g2_decap_4  FILLER_76_196
timestamp 1679577901
transform 1 0 19968 0 1 58212
box -48 -56 432 834
use sg13g2_decap_8  FILLER_77_0
timestamp 1679581782
transform 1 0 1152 0 -1 59724
box -48 -56 720 834
use sg13g2_fill_2  FILLER_77_11
timestamp 1677580104
transform 1 0 2208 0 -1 59724
box -48 -56 240 834
use sg13g2_decap_8  FILLER_77_34
timestamp 1679581782
transform 1 0 4416 0 -1 59724
box -48 -56 720 834
use sg13g2_fill_2  FILLER_77_83
timestamp 1677580104
transform 1 0 9120 0 -1 59724
box -48 -56 240 834
use sg13g2_fill_1  FILLER_77_85
timestamp 1677579658
transform 1 0 9312 0 -1 59724
box -48 -56 144 834
use sg13g2_fill_2  FILLER_77_103
timestamp 1677580104
transform 1 0 11040 0 -1 59724
box -48 -56 240 834
use sg13g2_decap_8  FILLER_77_190
timestamp 1679581782
transform 1 0 19392 0 -1 59724
box -48 -56 720 834
use sg13g2_fill_2  FILLER_77_197
timestamp 1677580104
transform 1 0 20064 0 -1 59724
box -48 -56 240 834
use sg13g2_fill_1  FILLER_77_199
timestamp 1677579658
transform 1 0 20256 0 -1 59724
box -48 -56 144 834
use sg13g2_fill_2  FILLER_78_0
timestamp 1677580104
transform 1 0 1152 0 1 59724
box -48 -56 240 834
use sg13g2_decap_8  FILLER_78_36
timestamp 1679581782
transform 1 0 4608 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_103
timestamp 1679581782
transform 1 0 11040 0 1 59724
box -48 -56 720 834
use sg13g2_fill_1  FILLER_78_110
timestamp 1677579658
transform 1 0 11712 0 1 59724
box -48 -56 144 834
use sg13g2_decap_8  FILLER_78_190
timestamp 1679581782
transform 1 0 19392 0 1 59724
box -48 -56 720 834
use sg13g2_fill_2  FILLER_78_197
timestamp 1677580104
transform 1 0 20064 0 1 59724
box -48 -56 240 834
use sg13g2_fill_1  FILLER_78_199
timestamp 1677579658
transform 1 0 20256 0 1 59724
box -48 -56 144 834
use sg13g2_decap_8  FILLER_79_0
timestamp 1679581782
transform 1 0 1152 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_7
timestamp 1679581782
transform 1 0 1824 0 -1 61236
box -48 -56 720 834
use sg13g2_fill_2  FILLER_79_14
timestamp 1677580104
transform 1 0 2496 0 -1 61236
box -48 -56 240 834
use sg13g2_fill_2  FILLER_79_37
timestamp 1677580104
transform 1 0 4704 0 -1 61236
box -48 -56 240 834
use sg13g2_fill_1  FILLER_79_39
timestamp 1677579658
transform 1 0 4896 0 -1 61236
box -48 -56 144 834
use sg13g2_decap_4  FILLER_79_125
timestamp 1679577901
transform 1 0 13152 0 -1 61236
box -48 -56 432 834
use sg13g2_fill_2  FILLER_79_129
timestamp 1677580104
transform 1 0 13536 0 -1 61236
box -48 -56 240 834
use sg13g2_fill_1  FILLER_79_157
timestamp 1677579658
transform 1 0 16224 0 -1 61236
box -48 -56 144 834
use sg13g2_fill_2  FILLER_79_175
timestamp 1677580104
transform 1 0 17952 0 -1 61236
box -48 -56 240 834
use sg13g2_decap_4  FILLER_79_194
timestamp 1679577901
transform 1 0 19776 0 -1 61236
box -48 -56 432 834
use sg13g2_fill_2  FILLER_79_198
timestamp 1677580104
transform 1 0 20160 0 -1 61236
box -48 -56 240 834
use sg13g2_decap_8  FILLER_80_0
timestamp 1679581782
transform 1 0 1152 0 1 61236
box -48 -56 720 834
use sg13g2_fill_2  FILLER_80_7
timestamp 1677580104
transform 1 0 1824 0 1 61236
box -48 -56 240 834
use sg13g2_decap_8  FILLER_80_30
timestamp 1679581782
transform 1 0 4032 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_37
timestamp 1679581782
transform 1 0 4704 0 1 61236
box -48 -56 720 834
use sg13g2_fill_1  FILLER_80_44
timestamp 1677579658
transform 1 0 5376 0 1 61236
box -48 -56 144 834
use sg13g2_decap_4  FILLER_80_83
timestamp 1679577901
transform 1 0 9120 0 1 61236
box -48 -56 432 834
use sg13g2_fill_1  FILLER_80_87
timestamp 1677579658
transform 1 0 9504 0 1 61236
box -48 -56 144 834
use sg13g2_decap_8  FILLER_80_105
timestamp 1679581782
transform 1 0 11232 0 1 61236
box -48 -56 720 834
use sg13g2_fill_2  FILLER_80_112
timestamp 1677580104
transform 1 0 11904 0 1 61236
box -48 -56 240 834
use sg13g2_decap_4  FILLER_80_131
timestamp 1679577901
transform 1 0 13728 0 1 61236
box -48 -56 432 834
use sg13g2_fill_2  FILLER_80_135
timestamp 1677580104
transform 1 0 14112 0 1 61236
box -48 -56 240 834
use sg13g2_decap_8  FILLER_80_168
timestamp 1679581782
transform 1 0 17280 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_175
timestamp 1679581782
transform 1 0 17952 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_182
timestamp 1679581782
transform 1 0 18624 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_189
timestamp 1679581782
transform 1 0 19296 0 1 61236
box -48 -56 720 834
use sg13g2_decap_4  FILLER_80_196
timestamp 1679577901
transform 1 0 19968 0 1 61236
box -48 -56 432 834
use sg13g2_decap_4  FILLER_81_0
timestamp 1679577901
transform 1 0 1152 0 -1 62748
box -48 -56 432 834
use sg13g2_fill_1  FILLER_81_4
timestamp 1677579658
transform 1 0 1536 0 -1 62748
box -48 -56 144 834
use sg13g2_decap_8  FILLER_81_22
timestamp 1679581782
transform 1 0 3264 0 -1 62748
box -48 -56 720 834
use sg13g2_fill_2  FILLER_81_29
timestamp 1677580104
transform 1 0 3936 0 -1 62748
box -48 -56 240 834
use sg13g2_fill_2  FILLER_81_92
timestamp 1677580104
transform 1 0 9984 0 -1 62748
box -48 -56 240 834
use sg13g2_decap_8  FILLER_81_132
timestamp 1679581782
transform 1 0 13824 0 -1 62748
box -48 -56 720 834
use sg13g2_fill_2  FILLER_81_139
timestamp 1677580104
transform 1 0 14496 0 -1 62748
box -48 -56 240 834
use sg13g2_fill_2  FILLER_81_156
timestamp 1677580104
transform 1 0 16128 0 -1 62748
box -48 -56 240 834
use sg13g2_fill_1  FILLER_81_158
timestamp 1677579658
transform 1 0 16320 0 -1 62748
box -48 -56 144 834
use sg13g2_decap_8  FILLER_81_176
timestamp 1679581782
transform 1 0 18048 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_183
timestamp 1679581782
transform 1 0 18720 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_190
timestamp 1679581782
transform 1 0 19392 0 -1 62748
box -48 -56 720 834
use sg13g2_fill_2  FILLER_81_197
timestamp 1677580104
transform 1 0 20064 0 -1 62748
box -48 -56 240 834
use sg13g2_fill_1  FILLER_81_199
timestamp 1677579658
transform 1 0 20256 0 -1 62748
box -48 -56 144 834
use sg13g2_decap_8  FILLER_82_0
timestamp 1679581782
transform 1 0 1152 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_7
timestamp 1679581782
transform 1 0 1824 0 1 62748
box -48 -56 720 834
use sg13g2_fill_1  FILLER_82_14
timestamp 1677579658
transform 1 0 2496 0 1 62748
box -48 -56 144 834
use sg13g2_decap_8  FILLER_82_36
timestamp 1679581782
transform 1 0 4608 0 1 62748
box -48 -56 720 834
use sg13g2_decap_4  FILLER_82_43
timestamp 1679577901
transform 1 0 5280 0 1 62748
box -48 -56 432 834
use sg13g2_fill_2  FILLER_82_47
timestamp 1677580104
transform 1 0 5664 0 1 62748
box -48 -56 240 834
use sg13g2_fill_2  FILLER_82_87
timestamp 1677580104
transform 1 0 9504 0 1 62748
box -48 -56 240 834
use sg13g2_decap_8  FILLER_82_106
timestamp 1679581782
transform 1 0 11328 0 1 62748
box -48 -56 720 834
use sg13g2_decap_4  FILLER_82_113
timestamp 1679577901
transform 1 0 12000 0 1 62748
box -48 -56 432 834
use sg13g2_fill_1  FILLER_82_117
timestamp 1677579658
transform 1 0 12384 0 1 62748
box -48 -56 144 834
use sg13g2_fill_2  FILLER_82_123
timestamp 1677580104
transform 1 0 12960 0 1 62748
box -48 -56 240 834
use sg13g2_decap_8  FILLER_82_181
timestamp 1679581782
transform 1 0 18528 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_188
timestamp 1679581782
transform 1 0 19200 0 1 62748
box -48 -56 720 834
use sg13g2_decap_4  FILLER_82_195
timestamp 1679577901
transform 1 0 19872 0 1 62748
box -48 -56 432 834
use sg13g2_fill_1  FILLER_82_199
timestamp 1677579658
transform 1 0 20256 0 1 62748
box -48 -56 144 834
use sg13g2_decap_8  FILLER_83_0
timestamp 1679581782
transform 1 0 1152 0 -1 64260
box -48 -56 720 834
use sg13g2_fill_2  FILLER_83_7
timestamp 1677580104
transform 1 0 1824 0 -1 64260
box -48 -56 240 834
use sg13g2_fill_1  FILLER_83_9
timestamp 1677579658
transform 1 0 2016 0 -1 64260
box -48 -56 144 834
use sg13g2_decap_8  FILLER_83_31
timestamp 1679581782
transform 1 0 4128 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_4  FILLER_83_38
timestamp 1679577901
transform 1 0 4800 0 -1 64260
box -48 -56 432 834
use sg13g2_fill_1  FILLER_83_42
timestamp 1677579658
transform 1 0 5184 0 -1 64260
box -48 -56 144 834
use sg13g2_decap_4  FILLER_83_64
timestamp 1679577901
transform 1 0 7296 0 -1 64260
box -48 -56 432 834
use sg13g2_fill_1  FILLER_83_68
timestamp 1677579658
transform 1 0 7680 0 -1 64260
box -48 -56 144 834
use sg13g2_decap_4  FILLER_83_96
timestamp 1679577901
transform 1 0 10368 0 -1 64260
box -48 -56 432 834
use sg13g2_fill_2  FILLER_83_127
timestamp 1677580104
transform 1 0 13344 0 -1 64260
box -48 -56 240 834
use sg13g2_fill_1  FILLER_83_129
timestamp 1677579658
transform 1 0 13536 0 -1 64260
box -48 -56 144 834
use sg13g2_fill_1  FILLER_83_166
timestamp 1677579658
transform 1 0 17088 0 -1 64260
box -48 -56 144 834
use sg13g2_decap_8  FILLER_83_180
timestamp 1679581782
transform 1 0 18432 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_187
timestamp 1679581782
transform 1 0 19104 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_4  FILLER_83_194
timestamp 1679577901
transform 1 0 19776 0 -1 64260
box -48 -56 432 834
use sg13g2_fill_2  FILLER_83_198
timestamp 1677580104
transform 1 0 20160 0 -1 64260
box -48 -56 240 834
use sg13g2_decap_8  FILLER_84_17
timestamp 1679581782
transform 1 0 2784 0 1 64260
box -48 -56 720 834
use sg13g2_fill_1  FILLER_84_79
timestamp 1677579658
transform 1 0 8736 0 1 64260
box -48 -56 144 834
use sg13g2_fill_2  FILLER_84_85
timestamp 1677580104
transform 1 0 9312 0 1 64260
box -48 -56 240 834
use sg13g2_decap_8  FILLER_84_176
timestamp 1679581782
transform 1 0 18048 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_183
timestamp 1679581782
transform 1 0 18720 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_190
timestamp 1679581782
transform 1 0 19392 0 1 64260
box -48 -56 720 834
use sg13g2_fill_2  FILLER_84_197
timestamp 1677580104
transform 1 0 20064 0 1 64260
box -48 -56 240 834
use sg13g2_fill_1  FILLER_84_199
timestamp 1677579658
transform 1 0 20256 0 1 64260
box -48 -56 144 834
use sg13g2_fill_2  FILLER_85_0
timestamp 1677580104
transform 1 0 1152 0 -1 65772
box -48 -56 240 834
use sg13g2_fill_1  FILLER_85_2
timestamp 1677579658
transform 1 0 1344 0 -1 65772
box -48 -56 144 834
use sg13g2_decap_8  FILLER_85_24
timestamp 1679581782
transform 1 0 3456 0 -1 65772
box -48 -56 720 834
use sg13g2_fill_1  FILLER_85_31
timestamp 1677579658
transform 1 0 4128 0 -1 65772
box -48 -56 144 834
use sg13g2_fill_1  FILLER_85_59
timestamp 1677579658
transform 1 0 6816 0 -1 65772
box -48 -56 144 834
use sg13g2_decap_8  FILLER_85_130
timestamp 1679581782
transform 1 0 13632 0 -1 65772
box -48 -56 720 834
use sg13g2_fill_1  FILLER_85_137
timestamp 1677579658
transform 1 0 14304 0 -1 65772
box -48 -56 144 834
use sg13g2_decap_8  FILLER_85_176
timestamp 1679581782
transform 1 0 18048 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_183
timestamp 1679581782
transform 1 0 18720 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_190
timestamp 1679581782
transform 1 0 19392 0 -1 65772
box -48 -56 720 834
use sg13g2_fill_2  FILLER_85_197
timestamp 1677580104
transform 1 0 20064 0 -1 65772
box -48 -56 240 834
use sg13g2_fill_1  FILLER_85_199
timestamp 1677579658
transform 1 0 20256 0 -1 65772
box -48 -56 144 834
use sg13g2_decap_4  FILLER_86_17
timestamp 1679577901
transform 1 0 2784 0 1 65772
box -48 -56 432 834
use sg13g2_fill_2  FILLER_86_21
timestamp 1677580104
transform 1 0 3168 0 1 65772
box -48 -56 240 834
use sg13g2_fill_2  FILLER_86_64
timestamp 1677580104
transform 1 0 7296 0 1 65772
box -48 -56 240 834
use sg13g2_fill_1  FILLER_86_66
timestamp 1677579658
transform 1 0 7488 0 1 65772
box -48 -56 144 834
use sg13g2_fill_1  FILLER_86_84
timestamp 1677579658
transform 1 0 9216 0 1 65772
box -48 -56 144 834
use sg13g2_decap_8  FILLER_86_95
timestamp 1679581782
transform 1 0 10272 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_102
timestamp 1679581782
transform 1 0 10944 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_109
timestamp 1679581782
transform 1 0 11616 0 1 65772
box -48 -56 720 834
use sg13g2_fill_2  FILLER_86_133
timestamp 1677580104
transform 1 0 13920 0 1 65772
box -48 -56 240 834
use sg13g2_decap_8  FILLER_86_140
timestamp 1679581782
transform 1 0 14592 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_147
timestamp 1679581782
transform 1 0 15264 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_166
timestamp 1679581782
transform 1 0 17088 0 1 65772
box -48 -56 720 834
use sg13g2_decap_4  FILLER_86_173
timestamp 1679577901
transform 1 0 17760 0 1 65772
box -48 -56 432 834
use sg13g2_fill_2  FILLER_86_177
timestamp 1677580104
transform 1 0 18144 0 1 65772
box -48 -56 240 834
use sg13g2_decap_4  FILLER_86_196
timestamp 1679577901
transform 1 0 19968 0 1 65772
box -48 -56 432 834
use sg13g2_decap_4  FILLER_87_0
timestamp 1679577901
transform 1 0 1152 0 -1 67284
box -48 -56 432 834
use sg13g2_fill_1  FILLER_87_4
timestamp 1677579658
transform 1 0 1536 0 -1 67284
box -48 -56 144 834
use sg13g2_fill_2  FILLER_87_22
timestamp 1677580104
transform 1 0 3264 0 -1 67284
box -48 -56 240 834
use sg13g2_fill_2  FILLER_87_75
timestamp 1677580104
transform 1 0 8352 0 -1 67284
box -48 -56 240 834
use sg13g2_fill_2  FILLER_87_91
timestamp 1677580104
transform 1 0 9888 0 -1 67284
box -48 -56 240 834
use sg13g2_fill_1  FILLER_87_93
timestamp 1677579658
transform 1 0 10080 0 -1 67284
box -48 -56 144 834
use sg13g2_fill_1  FILLER_87_111
timestamp 1677579658
transform 1 0 11808 0 -1 67284
box -48 -56 144 834
use sg13g2_fill_2  FILLER_87_172
timestamp 1677580104
transform 1 0 17664 0 -1 67284
box -48 -56 240 834
use sg13g2_fill_1  FILLER_87_174
timestamp 1677579658
transform 1 0 17856 0 -1 67284
box -48 -56 144 834
use sg13g2_fill_2  FILLER_87_197
timestamp 1677580104
transform 1 0 20064 0 -1 67284
box -48 -56 240 834
use sg13g2_fill_1  FILLER_87_199
timestamp 1677579658
transform 1 0 20256 0 -1 67284
box -48 -56 144 834
use sg13g2_decap_8  FILLER_88_0
timestamp 1679581782
transform 1 0 1152 0 1 67284
box -48 -56 720 834
use sg13g2_decap_4  FILLER_88_7
timestamp 1679577901
transform 1 0 1824 0 1 67284
box -48 -56 432 834
use sg13g2_fill_2  FILLER_88_66
timestamp 1677580104
transform 1 0 7488 0 1 67284
box -48 -56 240 834
use sg13g2_fill_1  FILLER_88_68
timestamp 1677579658
transform 1 0 7680 0 1 67284
box -48 -56 144 834
use sg13g2_decap_4  FILLER_88_107
timestamp 1679577901
transform 1 0 11424 0 1 67284
box -48 -56 432 834
use sg13g2_fill_2  FILLER_88_111
timestamp 1677580104
transform 1 0 11808 0 1 67284
box -48 -56 240 834
use sg13g2_decap_4  FILLER_88_130
timestamp 1679577901
transform 1 0 13632 0 1 67284
box -48 -56 432 834
use sg13g2_fill_2  FILLER_88_138
timestamp 1677580104
transform 1 0 14400 0 1 67284
box -48 -56 240 834
use sg13g2_fill_1  FILLER_88_140
timestamp 1677579658
transform 1 0 14592 0 1 67284
box -48 -56 144 834
use sg13g2_fill_2  FILLER_88_167
timestamp 1677580104
transform 1 0 17184 0 1 67284
box -48 -56 240 834
use sg13g2_decap_8  FILLER_89_0
timestamp 1679581782
transform 1 0 1152 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_4  FILLER_89_7
timestamp 1679577901
transform 1 0 1824 0 -1 68796
box -48 -56 432 834
use sg13g2_fill_1  FILLER_89_11
timestamp 1677579658
transform 1 0 2208 0 -1 68796
box -48 -56 144 834
use sg13g2_fill_1  FILLER_89_29
timestamp 1677579658
transform 1 0 3936 0 -1 68796
box -48 -56 144 834
use sg13g2_decap_8  FILLER_89_97
timestamp 1679581782
transform 1 0 10464 0 -1 68796
box -48 -56 720 834
use sg13g2_fill_2  FILLER_89_104
timestamp 1677580104
transform 1 0 11136 0 -1 68796
box -48 -56 240 834
use sg13g2_fill_1  FILLER_89_106
timestamp 1677579658
transform 1 0 11328 0 -1 68796
box -48 -56 144 834
use sg13g2_decap_4  FILLER_89_124
timestamp 1679577901
transform 1 0 13056 0 -1 68796
box -48 -56 432 834
use sg13g2_fill_2  FILLER_89_128
timestamp 1677580104
transform 1 0 13440 0 -1 68796
box -48 -56 240 834
use sg13g2_decap_8  FILLER_89_191
timestamp 1679581782
transform 1 0 19488 0 -1 68796
box -48 -56 720 834
use sg13g2_fill_2  FILLER_89_198
timestamp 1677580104
transform 1 0 20160 0 -1 68796
box -48 -56 240 834
use sg13g2_decap_4  FILLER_90_0
timestamp 1679577901
transform 1 0 1152 0 1 68796
box -48 -56 432 834
use sg13g2_fill_2  FILLER_90_4
timestamp 1677580104
transform 1 0 1536 0 1 68796
box -48 -56 240 834
use sg13g2_decap_8  FILLER_90_66
timestamp 1679581782
transform 1 0 7488 0 1 68796
box -48 -56 720 834
use sg13g2_fill_1  FILLER_90_111
timestamp 1677579658
transform 1 0 11808 0 1 68796
box -48 -56 144 834
use sg13g2_fill_1  FILLER_90_129
timestamp 1677579658
transform 1 0 13536 0 1 68796
box -48 -56 144 834
use sg13g2_fill_1  FILLER_90_157
timestamp 1677579658
transform 1 0 16224 0 1 68796
box -48 -56 144 834
use sg13g2_fill_2  FILLER_90_175
timestamp 1677580104
transform 1 0 17952 0 1 68796
box -48 -56 240 834
use sg13g2_fill_2  FILLER_90_197
timestamp 1677580104
transform 1 0 20064 0 1 68796
box -48 -56 240 834
use sg13g2_fill_1  FILLER_90_199
timestamp 1677579658
transform 1 0 20256 0 1 68796
box -48 -56 144 834
use sg13g2_fill_2  FILLER_91_56
timestamp 1677580104
transform 1 0 6528 0 -1 70308
box -48 -56 240 834
use sg13g2_decap_8  FILLER_91_62
timestamp 1679581782
transform 1 0 7104 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_4  FILLER_91_69
timestamp 1679577901
transform 1 0 7776 0 -1 70308
box -48 -56 432 834
use sg13g2_decap_8  FILLER_91_128
timestamp 1679581782
transform 1 0 13440 0 -1 70308
box -48 -56 720 834
use sg13g2_fill_2  FILLER_91_135
timestamp 1677580104
transform 1 0 14112 0 -1 70308
box -48 -56 240 834
use sg13g2_fill_2  FILLER_91_168
timestamp 1677580104
transform 1 0 17280 0 -1 70308
box -48 -56 240 834
use sg13g2_decap_8  FILLER_92_0
timestamp 1679581782
transform 1 0 1152 0 1 70308
box -48 -56 720 834
use sg13g2_decap_4  FILLER_92_7
timestamp 1679577901
transform 1 0 1824 0 1 70308
box -48 -56 432 834
use sg13g2_fill_1  FILLER_92_11
timestamp 1677579658
transform 1 0 2208 0 1 70308
box -48 -56 144 834
use sg13g2_decap_4  FILLER_92_33
timestamp 1679577901
transform 1 0 4320 0 1 70308
box -48 -56 432 834
use sg13g2_fill_2  FILLER_92_37
timestamp 1677580104
transform 1 0 4704 0 1 70308
box -48 -56 240 834
use sg13g2_fill_1  FILLER_92_69
timestamp 1677579658
transform 1 0 7776 0 1 70308
box -48 -56 144 834
use sg13g2_fill_2  FILLER_92_91
timestamp 1677580104
transform 1 0 9888 0 1 70308
box -48 -56 240 834
use sg13g2_fill_1  FILLER_92_93
timestamp 1677579658
transform 1 0 10080 0 1 70308
box -48 -56 144 834
use sg13g2_decap_8  FILLER_92_116
timestamp 1679581782
transform 1 0 12288 0 1 70308
box -48 -56 720 834
use sg13g2_fill_1  FILLER_92_140
timestamp 1677579658
transform 1 0 14592 0 1 70308
box -48 -56 144 834
use sg13g2_fill_2  FILLER_92_168
timestamp 1677580104
transform 1 0 17280 0 1 70308
box -48 -56 240 834
use sg13g2_fill_1  FILLER_92_170
timestamp 1677579658
transform 1 0 17472 0 1 70308
box -48 -56 144 834
use sg13g2_fill_2  FILLER_92_198
timestamp 1677580104
transform 1 0 20160 0 1 70308
box -48 -56 240 834
use sg13g2_decap_8  FILLER_93_34
timestamp 1679581782
transform 1 0 4416 0 -1 71820
box -48 -56 720 834
use sg13g2_fill_2  FILLER_93_41
timestamp 1677580104
transform 1 0 5088 0 -1 71820
box -48 -56 240 834
use sg13g2_fill_1  FILLER_93_43
timestamp 1677579658
transform 1 0 5280 0 -1 71820
box -48 -56 144 834
use sg13g2_fill_2  FILLER_93_66
timestamp 1677580104
transform 1 0 7488 0 -1 71820
box -48 -56 240 834
use sg13g2_decap_8  FILLER_93_102
timestamp 1679581782
transform 1 0 10944 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_4  FILLER_93_109
timestamp 1679577901
transform 1 0 11616 0 -1 71820
box -48 -56 432 834
use sg13g2_fill_1  FILLER_93_113
timestamp 1677579658
transform 1 0 12000 0 -1 71820
box -48 -56 144 834
use sg13g2_fill_1  FILLER_93_148
timestamp 1677579658
transform 1 0 15360 0 -1 71820
box -48 -56 144 834
use sg13g2_fill_2  FILLER_93_187
timestamp 1677580104
transform 1 0 19104 0 -1 71820
box -48 -56 240 834
use sg13g2_decap_8  FILLER_93_192
timestamp 1679581782
transform 1 0 19584 0 -1 71820
box -48 -56 720 834
use sg13g2_fill_1  FILLER_93_199
timestamp 1677579658
transform 1 0 20256 0 -1 71820
box -48 -56 144 834
use sg13g2_decap_8  FILLER_94_0
timestamp 1679581782
transform 1 0 1152 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_28
timestamp 1679581782
transform 1 0 3840 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_97
timestamp 1679581782
transform 1 0 10464 0 1 71820
box -48 -56 720 834
use sg13g2_decap_4  FILLER_94_104
timestamp 1679577901
transform 1 0 11136 0 1 71820
box -48 -56 432 834
use sg13g2_fill_2  FILLER_94_108
timestamp 1677580104
transform 1 0 11520 0 1 71820
box -48 -56 240 834
use sg13g2_fill_2  FILLER_94_131
timestamp 1677580104
transform 1 0 13728 0 1 71820
box -48 -56 240 834
use sg13g2_decap_8  FILLER_94_171
timestamp 1679581782
transform 1 0 17568 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_178
timestamp 1679581782
transform 1 0 18240 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_185
timestamp 1679581782
transform 1 0 18912 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_192
timestamp 1679581782
transform 1 0 19584 0 1 71820
box -48 -56 720 834
use sg13g2_fill_1  FILLER_94_199
timestamp 1677579658
transform 1 0 20256 0 1 71820
box -48 -56 144 834
use sg13g2_fill_2  FILLER_95_51
timestamp 1677580104
transform 1 0 6048 0 -1 73332
box -48 -56 240 834
use sg13g2_decap_8  FILLER_95_118
timestamp 1679581782
transform 1 0 12480 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_125
timestamp 1679581782
transform 1 0 13152 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_132
timestamp 1679581782
transform 1 0 13824 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_139
timestamp 1679581782
transform 1 0 14496 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_146
timestamp 1679581782
transform 1 0 15168 0 -1 73332
box -48 -56 720 834
use sg13g2_fill_1  FILLER_95_153
timestamp 1677579658
transform 1 0 15840 0 -1 73332
box -48 -56 144 834
use sg13g2_decap_8  FILLER_95_158
timestamp 1679581782
transform 1 0 16320 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_165
timestamp 1679581782
transform 1 0 16992 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_172
timestamp 1679581782
transform 1 0 17664 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_179
timestamp 1679581782
transform 1 0 18336 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_186
timestamp 1679581782
transform 1 0 19008 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_193
timestamp 1679581782
transform 1 0 19680 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_4  FILLER_96_0
timestamp 1679577901
transform 1 0 1152 0 1 73332
box -48 -56 432 834
use sg13g2_fill_1  FILLER_96_4
timestamp 1677579658
transform 1 0 1536 0 1 73332
box -48 -56 144 834
use sg13g2_decap_8  FILLER_96_26
timestamp 1679581782
transform 1 0 3648 0 1 73332
box -48 -56 720 834
use sg13g2_fill_2  FILLER_96_33
timestamp 1677580104
transform 1 0 4320 0 1 73332
box -48 -56 240 834
use sg13g2_fill_1  FILLER_96_35
timestamp 1677579658
transform 1 0 4512 0 1 73332
box -48 -56 144 834
use sg13g2_fill_1  FILLER_96_57
timestamp 1677579658
transform 1 0 6624 0 1 73332
box -48 -56 144 834
use sg13g2_fill_2  FILLER_96_66
timestamp 1677580104
transform 1 0 7488 0 1 73332
box -48 -56 240 834
use sg13g2_fill_2  FILLER_96_90
timestamp 1677580104
transform 1 0 9792 0 1 73332
box -48 -56 240 834
use sg13g2_decap_8  FILLER_96_117
timestamp 1679581782
transform 1 0 12384 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_124
timestamp 1679581782
transform 1 0 13056 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_131
timestamp 1679581782
transform 1 0 13728 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_138
timestamp 1679581782
transform 1 0 14400 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_145
timestamp 1679581782
transform 1 0 15072 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_152
timestamp 1679581782
transform 1 0 15744 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_159
timestamp 1679581782
transform 1 0 16416 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_166
timestamp 1679581782
transform 1 0 17088 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_173
timestamp 1679581782
transform 1 0 17760 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_180
timestamp 1679581782
transform 1 0 18432 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_187
timestamp 1679581782
transform 1 0 19104 0 1 73332
box -48 -56 720 834
use sg13g2_decap_4  FILLER_96_194
timestamp 1679577901
transform 1 0 19776 0 1 73332
box -48 -56 432 834
use sg13g2_fill_2  FILLER_96_198
timestamp 1677580104
transform 1 0 20160 0 1 73332
box -48 -56 240 834
use sg13g2_decap_8  FILLER_97_34
timestamp 1679581782
transform 1 0 4416 0 -1 74844
box -48 -56 720 834
use sg13g2_fill_2  FILLER_97_41
timestamp 1677580104
transform 1 0 5088 0 -1 74844
box -48 -56 240 834
use sg13g2_fill_1  FILLER_97_43
timestamp 1677579658
transform 1 0 5280 0 -1 74844
box -48 -56 144 834
use sg13g2_decap_8  FILLER_97_69
timestamp 1679581782
transform 1 0 7776 0 -1 74844
box -48 -56 720 834
use sg13g2_fill_1  FILLER_97_76
timestamp 1677579658
transform 1 0 8448 0 -1 74844
box -48 -56 144 834
use sg13g2_fill_2  FILLER_97_97
timestamp 1677580104
transform 1 0 10464 0 -1 74844
box -48 -56 240 834
use sg13g2_fill_2  FILLER_97_102
timestamp 1677580104
transform 1 0 10944 0 -1 74844
box -48 -56 240 834
use sg13g2_fill_1  FILLER_97_104
timestamp 1677579658
transform 1 0 11136 0 -1 74844
box -48 -56 144 834
use sg13g2_decap_8  FILLER_97_122
timestamp 1679581782
transform 1 0 12864 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_129
timestamp 1679581782
transform 1 0 13536 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_136
timestamp 1679581782
transform 1 0 14208 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_143
timestamp 1679581782
transform 1 0 14880 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_150
timestamp 1679581782
transform 1 0 15552 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_157
timestamp 1679581782
transform 1 0 16224 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_164
timestamp 1679581782
transform 1 0 16896 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_171
timestamp 1679581782
transform 1 0 17568 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_178
timestamp 1679581782
transform 1 0 18240 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_185
timestamp 1679581782
transform 1 0 18912 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_192
timestamp 1679581782
transform 1 0 19584 0 -1 74844
box -48 -56 720 834
use sg13g2_fill_1  FILLER_97_199
timestamp 1677579658
transform 1 0 20256 0 -1 74844
box -48 -56 144 834
use sg13g2_decap_8  FILLER_98_17
timestamp 1679581782
transform 1 0 2784 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_24
timestamp 1679581782
transform 1 0 3456 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_69
timestamp 1679581782
transform 1 0 7776 0 1 74844
box -48 -56 720 834
use sg13g2_decap_4  FILLER_98_76
timestamp 1679577901
transform 1 0 8448 0 1 74844
box -48 -56 432 834
use sg13g2_fill_2  FILLER_98_80
timestamp 1677580104
transform 1 0 8832 0 1 74844
box -48 -56 240 834
use sg13g2_decap_8  FILLER_98_120
timestamp 1679581782
transform 1 0 12672 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_127
timestamp 1679581782
transform 1 0 13344 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_134
timestamp 1679581782
transform 1 0 14016 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_141
timestamp 1679581782
transform 1 0 14688 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_148
timestamp 1679581782
transform 1 0 15360 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_155
timestamp 1679581782
transform 1 0 16032 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_162
timestamp 1679581782
transform 1 0 16704 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_169
timestamp 1679581782
transform 1 0 17376 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_176
timestamp 1679581782
transform 1 0 18048 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_183
timestamp 1679581782
transform 1 0 18720 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_190
timestamp 1679581782
transform 1 0 19392 0 1 74844
box -48 -56 720 834
use sg13g2_fill_2  FILLER_98_197
timestamp 1677580104
transform 1 0 20064 0 1 74844
box -48 -56 240 834
use sg13g2_fill_1  FILLER_98_199
timestamp 1677579658
transform 1 0 20256 0 1 74844
box -48 -56 144 834
use sg13g2_fill_2  FILLER_99_0
timestamp 1677580104
transform 1 0 1152 0 -1 76356
box -48 -56 240 834
use sg13g2_decap_8  FILLER_99_23
timestamp 1679581782
transform 1 0 3360 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_30
timestamp 1679581782
transform 1 0 4032 0 -1 76356
box -48 -56 720 834
use sg13g2_fill_1  FILLER_99_37
timestamp 1677579658
transform 1 0 4704 0 -1 76356
box -48 -56 144 834
use sg13g2_fill_2  FILLER_99_69
timestamp 1677580104
transform 1 0 7776 0 -1 76356
box -48 -56 240 834
use sg13g2_fill_2  FILLER_99_92
timestamp 1677580104
transform 1 0 9984 0 -1 76356
box -48 -56 240 834
use sg13g2_fill_1  FILLER_99_94
timestamp 1677579658
transform 1 0 10176 0 -1 76356
box -48 -56 144 834
use sg13g2_decap_8  FILLER_99_119
timestamp 1679581782
transform 1 0 12576 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_126
timestamp 1679581782
transform 1 0 13248 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_133
timestamp 1679581782
transform 1 0 13920 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_140
timestamp 1679581782
transform 1 0 14592 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_147
timestamp 1679581782
transform 1 0 15264 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_154
timestamp 1679581782
transform 1 0 15936 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_161
timestamp 1679581782
transform 1 0 16608 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_168
timestamp 1679581782
transform 1 0 17280 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_175
timestamp 1679581782
transform 1 0 17952 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_182
timestamp 1679581782
transform 1 0 18624 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_189
timestamp 1679581782
transform 1 0 19296 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_4  FILLER_99_196
timestamp 1679577901
transform 1 0 19968 0 -1 76356
box -48 -56 432 834
use sg13g2_decap_8  FILLER_100_0
timestamp 1679581782
transform 1 0 1152 0 1 76356
box -48 -56 720 834
use sg13g2_fill_2  FILLER_100_7
timestamp 1677580104
transform 1 0 1824 0 1 76356
box -48 -56 240 834
use sg13g2_decap_8  FILLER_100_26
timestamp 1679581782
transform 1 0 3648 0 1 76356
box -48 -56 720 834
use sg13g2_fill_2  FILLER_100_55
timestamp 1677580104
transform 1 0 6432 0 1 76356
box -48 -56 240 834
use sg13g2_decap_8  FILLER_100_112
timestamp 1679581782
transform 1 0 11904 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_119
timestamp 1679581782
transform 1 0 12576 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_126
timestamp 1679581782
transform 1 0 13248 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_133
timestamp 1679581782
transform 1 0 13920 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_140
timestamp 1679581782
transform 1 0 14592 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_147
timestamp 1679581782
transform 1 0 15264 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_154
timestamp 1679581782
transform 1 0 15936 0 1 76356
box -48 -56 720 834
use sg13g2_fill_2  FILLER_100_161
timestamp 1677580104
transform 1 0 16608 0 1 76356
box -48 -56 240 834
use sg13g2_fill_1  FILLER_100_163
timestamp 1677579658
transform 1 0 16800 0 1 76356
box -48 -56 144 834
use sg13g2_decap_8  FILLER_100_168
timestamp 1679581782
transform 1 0 17280 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_175
timestamp 1679581782
transform 1 0 17952 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_182
timestamp 1679581782
transform 1 0 18624 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_189
timestamp 1679581782
transform 1 0 19296 0 1 76356
box -48 -56 720 834
use sg13g2_decap_4  FILLER_100_196
timestamp 1679577901
transform 1 0 19968 0 1 76356
box -48 -56 432 834
use sg13g2_decap_8  FILLER_101_0
timestamp 1679581782
transform 1 0 1152 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_7
timestamp 1679581782
transform 1 0 1824 0 -1 77868
box -48 -56 720 834
use sg13g2_fill_2  FILLER_101_14
timestamp 1677580104
transform 1 0 2496 0 -1 77868
box -48 -56 240 834
use sg13g2_fill_2  FILLER_101_37
timestamp 1677580104
transform 1 0 4704 0 -1 77868
box -48 -56 240 834
use sg13g2_fill_1  FILLER_101_39
timestamp 1677579658
transform 1 0 4896 0 -1 77868
box -48 -56 144 834
use sg13g2_decap_8  FILLER_101_88
timestamp 1679581782
transform 1 0 9600 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_95
timestamp 1679581782
transform 1 0 10272 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_102
timestamp 1679581782
transform 1 0 10944 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_109
timestamp 1679581782
transform 1 0 11616 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_116
timestamp 1679581782
transform 1 0 12288 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_123
timestamp 1679581782
transform 1 0 12960 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_130
timestamp 1679581782
transform 1 0 13632 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_137
timestamp 1679581782
transform 1 0 14304 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_144
timestamp 1679581782
transform 1 0 14976 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_151
timestamp 1679581782
transform 1 0 15648 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_158
timestamp 1679581782
transform 1 0 16320 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_165
timestamp 1679581782
transform 1 0 16992 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_172
timestamp 1679581782
transform 1 0 17664 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_179
timestamp 1679581782
transform 1 0 18336 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_186
timestamp 1679581782
transform 1 0 19008 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_193
timestamp 1679581782
transform 1 0 19680 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_4  FILLER_102_17
timestamp 1679577901
transform 1 0 2784 0 1 77868
box -48 -56 432 834
use sg13g2_fill_1  FILLER_102_21
timestamp 1677579658
transform 1 0 3168 0 1 77868
box -48 -56 144 834
use sg13g2_fill_1  FILLER_102_56
timestamp 1677579658
transform 1 0 6528 0 1 77868
box -48 -56 144 834
use sg13g2_decap_8  FILLER_102_95
timestamp 1679581782
transform 1 0 10272 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_102
timestamp 1679581782
transform 1 0 10944 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_109
timestamp 1679581782
transform 1 0 11616 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_116
timestamp 1679581782
transform 1 0 12288 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_123
timestamp 1679581782
transform 1 0 12960 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_130
timestamp 1679581782
transform 1 0 13632 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_137
timestamp 1679581782
transform 1 0 14304 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_144
timestamp 1679581782
transform 1 0 14976 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_151
timestamp 1679581782
transform 1 0 15648 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_158
timestamp 1679581782
transform 1 0 16320 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_165
timestamp 1679581782
transform 1 0 16992 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_172
timestamp 1679581782
transform 1 0 17664 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_179
timestamp 1679581782
transform 1 0 18336 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_186
timestamp 1679581782
transform 1 0 19008 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_193
timestamp 1679581782
transform 1 0 19680 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_0
timestamp 1679581782
transform 1 0 1152 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_24
timestamp 1679581782
transform 1 0 3456 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_4  FILLER_103_74
timestamp 1679577901
transform 1 0 8256 0 -1 79380
box -48 -56 432 834
use sg13g2_fill_2  FILLER_103_78
timestamp 1677580104
transform 1 0 8640 0 -1 79380
box -48 -56 240 834
use sg13g2_decap_8  FILLER_103_97
timestamp 1679581782
transform 1 0 10464 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_104
timestamp 1679581782
transform 1 0 11136 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_111
timestamp 1679581782
transform 1 0 11808 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_118
timestamp 1679581782
transform 1 0 12480 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_125
timestamp 1679581782
transform 1 0 13152 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_132
timestamp 1679581782
transform 1 0 13824 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_139
timestamp 1679581782
transform 1 0 14496 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_146
timestamp 1679581782
transform 1 0 15168 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_153
timestamp 1679581782
transform 1 0 15840 0 -1 79380
box -48 -56 720 834
use sg13g2_fill_2  FILLER_103_160
timestamp 1677580104
transform 1 0 16512 0 -1 79380
box -48 -56 240 834
use sg13g2_decap_8  FILLER_103_166
timestamp 1679581782
transform 1 0 17088 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_173
timestamp 1679581782
transform 1 0 17760 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_180
timestamp 1679581782
transform 1 0 18432 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_187
timestamp 1679581782
transform 1 0 19104 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_4  FILLER_103_194
timestamp 1679577901
transform 1 0 19776 0 -1 79380
box -48 -56 432 834
use sg13g2_fill_2  FILLER_103_198
timestamp 1677580104
transform 1 0 20160 0 -1 79380
box -48 -56 240 834
use sg13g2_decap_8  FILLER_104_17
timestamp 1679581782
transform 1 0 2784 0 1 79380
box -48 -56 720 834
use sg13g2_decap_4  FILLER_104_66
timestamp 1679577901
transform 1 0 7488 0 1 79380
box -48 -56 432 834
use sg13g2_decap_8  FILLER_104_87
timestamp 1679581782
transform 1 0 9504 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_94
timestamp 1679581782
transform 1 0 10176 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_101
timestamp 1679581782
transform 1 0 10848 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_108
timestamp 1679581782
transform 1 0 11520 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_115
timestamp 1679581782
transform 1 0 12192 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_122
timestamp 1679581782
transform 1 0 12864 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_129
timestamp 1679581782
transform 1 0 13536 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_136
timestamp 1679581782
transform 1 0 14208 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_143
timestamp 1679581782
transform 1 0 14880 0 1 79380
box -48 -56 720 834
use sg13g2_fill_2  FILLER_104_150
timestamp 1677580104
transform 1 0 15552 0 1 79380
box -48 -56 240 834
use sg13g2_decap_8  FILLER_104_156
timestamp 1679581782
transform 1 0 16128 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_163
timestamp 1679581782
transform 1 0 16800 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_170
timestamp 1679581782
transform 1 0 17472 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_177
timestamp 1679581782
transform 1 0 18144 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_184
timestamp 1679581782
transform 1 0 18816 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_191
timestamp 1679581782
transform 1 0 19488 0 1 79380
box -48 -56 720 834
use sg13g2_fill_2  FILLER_104_198
timestamp 1677580104
transform 1 0 20160 0 1 79380
box -48 -56 240 834
use sg13g2_decap_4  FILLER_105_0
timestamp 1679577901
transform 1 0 1152 0 -1 80892
box -48 -56 432 834
use sg13g2_decap_4  FILLER_105_21
timestamp 1679577901
transform 1 0 3168 0 -1 80892
box -48 -56 432 834
use sg13g2_fill_1  FILLER_105_25
timestamp 1677579658
transform 1 0 3552 0 -1 80892
box -48 -56 144 834
use sg13g2_decap_8  FILLER_105_64
timestamp 1679581782
transform 1 0 7296 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_71
timestamp 1679581782
transform 1 0 7968 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_78
timestamp 1679581782
transform 1 0 8640 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_85
timestamp 1679581782
transform 1 0 9312 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_92
timestamp 1679581782
transform 1 0 9984 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_99
timestamp 1679581782
transform 1 0 10656 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_106
timestamp 1679581782
transform 1 0 11328 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_113
timestamp 1679581782
transform 1 0 12000 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_120
timestamp 1679581782
transform 1 0 12672 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_127
timestamp 1679581782
transform 1 0 13344 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_134
timestamp 1679581782
transform 1 0 14016 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_141
timestamp 1679581782
transform 1 0 14688 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_148
timestamp 1679581782
transform 1 0 15360 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_155
timestamp 1679581782
transform 1 0 16032 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_162
timestamp 1679581782
transform 1 0 16704 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_169
timestamp 1679581782
transform 1 0 17376 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_176
timestamp 1679581782
transform 1 0 18048 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_183
timestamp 1679581782
transform 1 0 18720 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_190
timestamp 1679581782
transform 1 0 19392 0 -1 80892
box -48 -56 720 834
use sg13g2_fill_2  FILLER_105_197
timestamp 1677580104
transform 1 0 20064 0 -1 80892
box -48 -56 240 834
use sg13g2_fill_1  FILLER_105_199
timestamp 1677579658
transform 1 0 20256 0 -1 80892
box -48 -56 144 834
use sg13g2_decap_8  FILLER_106_68
timestamp 1679581782
transform 1 0 7680 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_75
timestamp 1679581782
transform 1 0 8352 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_82
timestamp 1679581782
transform 1 0 9024 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_89
timestamp 1679581782
transform 1 0 9696 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_96
timestamp 1679581782
transform 1 0 10368 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_103
timestamp 1679581782
transform 1 0 11040 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_110
timestamp 1679581782
transform 1 0 11712 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_117
timestamp 1679581782
transform 1 0 12384 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_124
timestamp 1679581782
transform 1 0 13056 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_131
timestamp 1679581782
transform 1 0 13728 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_138
timestamp 1679581782
transform 1 0 14400 0 1 80892
box -48 -56 720 834
use sg13g2_decap_4  FILLER_106_145
timestamp 1679577901
transform 1 0 15072 0 1 80892
box -48 -56 432 834
use sg13g2_fill_1  FILLER_106_149
timestamp 1677579658
transform 1 0 15456 0 1 80892
box -48 -56 144 834
use sg13g2_decap_8  FILLER_106_154
timestamp 1679581782
transform 1 0 15936 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_161
timestamp 1679581782
transform 1 0 16608 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_168
timestamp 1679581782
transform 1 0 17280 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_175
timestamp 1679581782
transform 1 0 17952 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_182
timestamp 1679581782
transform 1 0 18624 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_189
timestamp 1679581782
transform 1 0 19296 0 1 80892
box -48 -56 720 834
use sg13g2_decap_4  FILLER_106_196
timestamp 1679577901
transform 1 0 19968 0 1 80892
box -48 -56 432 834
use sg13g2_decap_8  FILLER_107_17
timestamp 1679581782
transform 1 0 2784 0 -1 82404
box -48 -56 720 834
use sg13g2_fill_2  FILLER_107_24
timestamp 1677580104
transform 1 0 3456 0 -1 82404
box -48 -56 240 834
use sg13g2_decap_8  FILLER_107_43
timestamp 1679581782
transform 1 0 5280 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_50
timestamp 1679581782
transform 1 0 5952 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_57
timestamp 1679581782
transform 1 0 6624 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_64
timestamp 1679581782
transform 1 0 7296 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_71
timestamp 1679581782
transform 1 0 7968 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_78
timestamp 1679581782
transform 1 0 8640 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_85
timestamp 1679581782
transform 1 0 9312 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_92
timestamp 1679581782
transform 1 0 9984 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_99
timestamp 1679581782
transform 1 0 10656 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_106
timestamp 1679581782
transform 1 0 11328 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_113
timestamp 1679581782
transform 1 0 12000 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_120
timestamp 1679581782
transform 1 0 12672 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_127
timestamp 1679581782
transform 1 0 13344 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_134
timestamp 1679581782
transform 1 0 14016 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_141
timestamp 1679581782
transform 1 0 14688 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_148
timestamp 1679581782
transform 1 0 15360 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_155
timestamp 1679581782
transform 1 0 16032 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_107_162
timestamp 1679581782
transform 1 0 16704 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_4  FILLER_107_169
timestamp 1679577901
transform 1 0 17376 0 -1 82404
box -48 -56 432 834
use sg13g2_fill_2  FILLER_107_173
timestamp 1677580104
transform 1 0 17760 0 -1 82404
box -48 -56 240 834
use sg13g2_fill_1  FILLER_107_178
timestamp 1677579658
transform 1 0 18240 0 -1 82404
box -48 -56 144 834
use sg13g2_fill_1  FILLER_107_182
timestamp 1677579658
transform 1 0 18624 0 -1 82404
box -48 -56 144 834
use sg13g2_fill_1  FILLER_107_186
timestamp 1677579658
transform 1 0 19008 0 -1 82404
box -48 -56 144 834
use sg13g2_decap_8  FILLER_107_190
timestamp 1679581782
transform 1 0 19392 0 -1 82404
box -48 -56 720 834
use sg13g2_fill_2  FILLER_107_197
timestamp 1677580104
transform 1 0 20064 0 -1 82404
box -48 -56 240 834
use sg13g2_fill_1  FILLER_107_199
timestamp 1677579658
transform 1 0 20256 0 -1 82404
box -48 -56 144 834
use sg13g2_decap_8  FILLER_108_0
timestamp 1679581782
transform 1 0 1152 0 1 82404
box -48 -56 720 834
use sg13g2_fill_1  FILLER_108_24
timestamp 1677579658
transform 1 0 3456 0 1 82404
box -48 -56 144 834
use sg13g2_fill_1  FILLER_108_29
timestamp 1677579658
transform 1 0 3936 0 1 82404
box -48 -56 144 834
use sg13g2_decap_8  FILLER_108_47
timestamp 1679581782
transform 1 0 5664 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_108_54
timestamp 1679581782
transform 1 0 6336 0 1 82404
box -48 -56 720 834
use sg13g2_fill_2  FILLER_108_61
timestamp 1677580104
transform 1 0 7008 0 1 82404
box -48 -56 240 834
use sg13g2_decap_8  FILLER_108_67
timestamp 1679581782
transform 1 0 7584 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_108_74
timestamp 1679581782
transform 1 0 8256 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_108_81
timestamp 1679581782
transform 1 0 8928 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_108_88
timestamp 1679581782
transform 1 0 9600 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_108_95
timestamp 1679581782
transform 1 0 10272 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_108_102
timestamp 1679581782
transform 1 0 10944 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_108_109
timestamp 1679581782
transform 1 0 11616 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_108_116
timestamp 1679581782
transform 1 0 12288 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_108_123
timestamp 1679581782
transform 1 0 12960 0 1 82404
box -48 -56 720 834
use sg13g2_decap_4  FILLER_108_130
timestamp 1679577901
transform 1 0 13632 0 1 82404
box -48 -56 432 834
use sg13g2_fill_1  FILLER_108_134
timestamp 1677579658
transform 1 0 14016 0 1 82404
box -48 -56 144 834
use sg13g2_decap_8  FILLER_108_143
timestamp 1679581782
transform 1 0 14880 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_108_150
timestamp 1679581782
transform 1 0 15552 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_108_157
timestamp 1679581782
transform 1 0 16224 0 1 82404
box -48 -56 720 834
use sg13g2_decap_4  FILLER_108_164
timestamp 1679577901
transform 1 0 16896 0 1 82404
box -48 -56 432 834
use sg13g2_fill_1  FILLER_108_171
timestamp 1677579658
transform 1 0 17568 0 1 82404
box -48 -56 144 834
use sg13g2_fill_1  FILLER_108_191
timestamp 1677579658
transform 1 0 19488 0 1 82404
box -48 -56 144 834
use sg13g2_fill_1  FILLER_108_195
timestamp 1677579658
transform 1 0 19872 0 1 82404
box -48 -56 144 834
use sg13g2_fill_1  FILLER_108_199
timestamp 1677579658
transform 1 0 20256 0 1 82404
box -48 -56 144 834
use sg13g2_decap_4  FILLER_109_0
timestamp 1679577901
transform 1 0 1152 0 -1 83916
box -48 -56 432 834
use sg13g2_fill_1  FILLER_109_4
timestamp 1677579658
transform 1 0 1536 0 -1 83916
box -48 -56 144 834
use sg13g2_fill_1  FILLER_109_49
timestamp 1677579658
transform 1 0 5856 0 -1 83916
box -48 -56 144 834
use sg13g2_fill_1  FILLER_109_74
timestamp 1677579658
transform 1 0 8256 0 -1 83916
box -48 -56 144 834
use sg13g2_decap_4  FILLER_109_83
timestamp 1679577901
transform 1 0 9120 0 -1 83916
box -48 -56 432 834
use sg13g2_fill_1  FILLER_109_91
timestamp 1677579658
transform 1 0 9888 0 -1 83916
box -48 -56 144 834
use sg13g2_decap_4  FILLER_109_100
timestamp 1679577901
transform 1 0 10752 0 -1 83916
box -48 -56 432 834
use sg13g2_fill_1  FILLER_109_104
timestamp 1677579658
transform 1 0 11136 0 -1 83916
box -48 -56 144 834
use sg13g2_decap_8  FILLER_109_109
timestamp 1679581782
transform 1 0 11616 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_109_116
timestamp 1679581782
transform 1 0 12288 0 -1 83916
box -48 -56 720 834
use sg13g2_fill_1  FILLER_109_123
timestamp 1677579658
transform 1 0 12960 0 -1 83916
box -48 -56 144 834
use sg13g2_fill_2  FILLER_109_148
timestamp 1677580104
transform 1 0 15360 0 -1 83916
box -48 -56 240 834
use sg13g2_fill_1  FILLER_109_150
timestamp 1677579658
transform 1 0 15552 0 -1 83916
box -48 -56 144 834
use sg13g2_decap_4  FILLER_109_155
timestamp 1679577901
transform 1 0 16032 0 -1 83916
box -48 -56 432 834
use sg13g2_fill_1  FILLER_109_159
timestamp 1677579658
transform 1 0 16416 0 -1 83916
box -48 -56 144 834
use sg13g2_decap_8  FILLER_110_0
timestamp 1679581782
transform 1 0 1152 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_7
timestamp 1679581782
transform 1 0 1824 0 1 83916
box -48 -56 720 834
use sg13g2_decap_4  FILLER_110_14
timestamp 1679577901
transform 1 0 2496 0 1 83916
box -48 -56 432 834
use sg13g2_fill_1  FILLER_110_18
timestamp 1677579658
transform 1 0 2880 0 1 83916
box -48 -56 144 834
use sg13g2_decap_8  FILLER_110_27
timestamp 1679581782
transform 1 0 3744 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_34
timestamp 1679581782
transform 1 0 4416 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_41
timestamp 1679581782
transform 1 0 5088 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_48
timestamp 1679581782
transform 1 0 5760 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_55
timestamp 1679581782
transform 1 0 6432 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_62
timestamp 1679581782
transform 1 0 7104 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_69
timestamp 1679581782
transform 1 0 7776 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_76
timestamp 1679581782
transform 1 0 8448 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_83
timestamp 1679581782
transform 1 0 9120 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_90
timestamp 1679581782
transform 1 0 9792 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_97
timestamp 1679581782
transform 1 0 10464 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_104
timestamp 1679581782
transform 1 0 11136 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_111
timestamp 1679581782
transform 1 0 11808 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_118
timestamp 1679581782
transform 1 0 12480 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_125
timestamp 1679581782
transform 1 0 13152 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_132
timestamp 1679581782
transform 1 0 13824 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_139
timestamp 1679581782
transform 1 0 14496 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_146
timestamp 1679581782
transform 1 0 15168 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_153
timestamp 1679581782
transform 1 0 15840 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_160
timestamp 1679581782
transform 1 0 16512 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_110_167
timestamp 1679581782
transform 1 0 17184 0 1 83916
box -48 -56 720 834
use sg13g2_fill_2  FILLER_110_174
timestamp 1677580104
transform 1 0 17856 0 1 83916
box -48 -56 240 834
use sg13g2_fill_1  FILLER_110_179
timestamp 1677579658
transform 1 0 18336 0 1 83916
box -48 -56 144 834
use sg13g2_fill_1  FILLER_110_183
timestamp 1677579658
transform 1 0 18720 0 1 83916
box -48 -56 144 834
use sg13g2_fill_1  FILLER_110_187
timestamp 1677579658
transform 1 0 19104 0 1 83916
box -48 -56 144 834
use sg13g2_decap_8  FILLER_110_191
timestamp 1679581782
transform 1 0 19488 0 1 83916
box -48 -56 720 834
use sg13g2_fill_2  FILLER_110_198
timestamp 1677580104
transform 1 0 20160 0 1 83916
box -48 -56 240 834
<< labels >>
flabel metal3 s 21424 34820 21504 34900 0 FreeSans 320 0 0 0 CLK_TT_PROJECT
port 0 nsew signal output
flabel metal3 s 21424 34148 21504 34228 0 FreeSans 320 0 0 0 ENA_TT_PROJECT
port 1 nsew signal output
flabel metal3 s 21424 35492 21504 35572 0 FreeSans 320 0 0 0 RST_N_TT_PROJECT
port 2 nsew signal output
flabel metal3 s 0 59180 80 59260 0 FreeSans 320 0 0 0 Tile_X0Y0_E1END[0]
port 3 nsew signal input
flabel metal3 s 0 59516 80 59596 0 FreeSans 320 0 0 0 Tile_X0Y0_E1END[1]
port 4 nsew signal input
flabel metal3 s 0 59852 80 59932 0 FreeSans 320 0 0 0 Tile_X0Y0_E1END[2]
port 5 nsew signal input
flabel metal3 s 0 60188 80 60268 0 FreeSans 320 0 0 0 Tile_X0Y0_E1END[3]
port 6 nsew signal input
flabel metal3 s 0 63212 80 63292 0 FreeSans 320 0 0 0 Tile_X0Y0_E2END[0]
port 7 nsew signal input
flabel metal3 s 0 63548 80 63628 0 FreeSans 320 0 0 0 Tile_X0Y0_E2END[1]
port 8 nsew signal input
flabel metal3 s 0 63884 80 63964 0 FreeSans 320 0 0 0 Tile_X0Y0_E2END[2]
port 9 nsew signal input
flabel metal3 s 0 64220 80 64300 0 FreeSans 320 0 0 0 Tile_X0Y0_E2END[3]
port 10 nsew signal input
flabel metal3 s 0 64556 80 64636 0 FreeSans 320 0 0 0 Tile_X0Y0_E2END[4]
port 11 nsew signal input
flabel metal3 s 0 64892 80 64972 0 FreeSans 320 0 0 0 Tile_X0Y0_E2END[5]
port 12 nsew signal input
flabel metal3 s 0 65228 80 65308 0 FreeSans 320 0 0 0 Tile_X0Y0_E2END[6]
port 13 nsew signal input
flabel metal3 s 0 65564 80 65644 0 FreeSans 320 0 0 0 Tile_X0Y0_E2END[7]
port 14 nsew signal input
flabel metal3 s 0 60524 80 60604 0 FreeSans 320 0 0 0 Tile_X0Y0_E2MID[0]
port 15 nsew signal input
flabel metal3 s 0 60860 80 60940 0 FreeSans 320 0 0 0 Tile_X0Y0_E2MID[1]
port 16 nsew signal input
flabel metal3 s 0 61196 80 61276 0 FreeSans 320 0 0 0 Tile_X0Y0_E2MID[2]
port 17 nsew signal input
flabel metal3 s 0 61532 80 61612 0 FreeSans 320 0 0 0 Tile_X0Y0_E2MID[3]
port 18 nsew signal input
flabel metal3 s 0 61868 80 61948 0 FreeSans 320 0 0 0 Tile_X0Y0_E2MID[4]
port 19 nsew signal input
flabel metal3 s 0 62204 80 62284 0 FreeSans 320 0 0 0 Tile_X0Y0_E2MID[5]
port 20 nsew signal input
flabel metal3 s 0 62540 80 62620 0 FreeSans 320 0 0 0 Tile_X0Y0_E2MID[6]
port 21 nsew signal input
flabel metal3 s 0 62876 80 62956 0 FreeSans 320 0 0 0 Tile_X0Y0_E2MID[7]
port 22 nsew signal input
flabel metal3 s 0 71276 80 71356 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[0]
port 23 nsew signal input
flabel metal3 s 0 74636 80 74716 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[10]
port 24 nsew signal input
flabel metal3 s 0 74972 80 75052 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[11]
port 25 nsew signal input
flabel metal3 s 0 71612 80 71692 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[1]
port 26 nsew signal input
flabel metal3 s 0 71948 80 72028 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[2]
port 27 nsew signal input
flabel metal3 s 0 72284 80 72364 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[3]
port 28 nsew signal input
flabel metal3 s 0 72620 80 72700 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[4]
port 29 nsew signal input
flabel metal3 s 0 72956 80 73036 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[5]
port 30 nsew signal input
flabel metal3 s 0 73292 80 73372 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[6]
port 31 nsew signal input
flabel metal3 s 0 73628 80 73708 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[7]
port 32 nsew signal input
flabel metal3 s 0 73964 80 74044 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[8]
port 33 nsew signal input
flabel metal3 s 0 74300 80 74380 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[9]
port 34 nsew signal input
flabel metal3 s 0 65900 80 65980 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[0]
port 35 nsew signal input
flabel metal3 s 0 69260 80 69340 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[10]
port 36 nsew signal input
flabel metal3 s 0 69596 80 69676 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[11]
port 37 nsew signal input
flabel metal3 s 0 69932 80 70012 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[12]
port 38 nsew signal input
flabel metal3 s 0 70268 80 70348 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[13]
port 39 nsew signal input
flabel metal3 s 0 70604 80 70684 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[14]
port 40 nsew signal input
flabel metal3 s 0 70940 80 71020 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[15]
port 41 nsew signal input
flabel metal3 s 0 66236 80 66316 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[1]
port 42 nsew signal input
flabel metal3 s 0 66572 80 66652 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[2]
port 43 nsew signal input
flabel metal3 s 0 66908 80 66988 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[3]
port 44 nsew signal input
flabel metal3 s 0 67244 80 67324 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[4]
port 45 nsew signal input
flabel metal3 s 0 67580 80 67660 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[5]
port 46 nsew signal input
flabel metal3 s 0 67916 80 67996 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[6]
port 47 nsew signal input
flabel metal3 s 0 68252 80 68332 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[7]
port 48 nsew signal input
flabel metal3 s 0 68588 80 68668 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[8]
port 49 nsew signal input
flabel metal3 s 0 68924 80 69004 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[9]
port 50 nsew signal input
flabel metal3 s 0 75308 80 75388 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[0]
port 51 nsew signal input
flabel metal3 s 0 78668 80 78748 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[10]
port 52 nsew signal input
flabel metal3 s 0 79004 80 79084 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[11]
port 53 nsew signal input
flabel metal3 s 0 79340 80 79420 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[12]
port 54 nsew signal input
flabel metal3 s 0 79676 80 79756 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[13]
port 55 nsew signal input
flabel metal3 s 0 80012 80 80092 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[14]
port 56 nsew signal input
flabel metal3 s 0 80348 80 80428 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[15]
port 57 nsew signal input
flabel metal3 s 0 80684 80 80764 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[16]
port 58 nsew signal input
flabel metal3 s 0 81020 80 81100 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[17]
port 59 nsew signal input
flabel metal3 s 0 81356 80 81436 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[18]
port 60 nsew signal input
flabel metal3 s 0 81692 80 81772 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[19]
port 61 nsew signal input
flabel metal3 s 0 75644 80 75724 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[1]
port 62 nsew signal input
flabel metal3 s 0 82028 80 82108 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[20]
port 63 nsew signal input
flabel metal3 s 0 82364 80 82444 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[21]
port 64 nsew signal input
flabel metal3 s 0 82700 80 82780 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[22]
port 65 nsew signal input
flabel metal3 s 0 83036 80 83116 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[23]
port 66 nsew signal input
flabel metal3 s 0 83372 80 83452 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[24]
port 67 nsew signal input
flabel metal3 s 0 83708 80 83788 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[25]
port 68 nsew signal input
flabel metal3 s 0 84044 80 84124 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[26]
port 69 nsew signal input
flabel metal3 s 0 84380 80 84460 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[27]
port 70 nsew signal input
flabel metal3 s 0 84716 80 84796 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[28]
port 71 nsew signal input
flabel metal3 s 0 85052 80 85132 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[29]
port 72 nsew signal input
flabel metal3 s 0 75980 80 76060 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[2]
port 73 nsew signal input
flabel metal3 s 0 85388 80 85468 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[30]
port 74 nsew signal input
flabel metal3 s 0 85724 80 85804 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[31]
port 75 nsew signal input
flabel metal3 s 0 76316 80 76396 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[3]
port 76 nsew signal input
flabel metal3 s 0 76652 80 76732 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[4]
port 77 nsew signal input
flabel metal3 s 0 76988 80 77068 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[5]
port 78 nsew signal input
flabel metal3 s 0 77324 80 77404 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[6]
port 79 nsew signal input
flabel metal3 s 0 77660 80 77740 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[7]
port 80 nsew signal input
flabel metal3 s 0 77996 80 78076 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[8]
port 81 nsew signal input
flabel metal3 s 0 78332 80 78412 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[9]
port 82 nsew signal input
flabel metal3 s 21424 36164 21504 36244 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[0]
port 83 nsew signal output
flabel metal3 s 21424 42884 21504 42964 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[10]
port 84 nsew signal output
flabel metal3 s 21424 43556 21504 43636 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[11]
port 85 nsew signal output
flabel metal3 s 21424 44228 21504 44308 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[12]
port 86 nsew signal output
flabel metal3 s 21424 44900 21504 44980 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[13]
port 87 nsew signal output
flabel metal3 s 21424 45572 21504 45652 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[14]
port 88 nsew signal output
flabel metal3 s 21424 46244 21504 46324 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[15]
port 89 nsew signal output
flabel metal3 s 21424 46916 21504 46996 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[16]
port 90 nsew signal output
flabel metal3 s 21424 47588 21504 47668 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[17]
port 91 nsew signal output
flabel metal3 s 21424 48260 21504 48340 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[18]
port 92 nsew signal output
flabel metal3 s 21424 48932 21504 49012 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[19]
port 93 nsew signal output
flabel metal3 s 21424 36836 21504 36916 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[1]
port 94 nsew signal output
flabel metal3 s 21424 49604 21504 49684 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[20]
port 95 nsew signal output
flabel metal3 s 21424 50276 21504 50356 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[21]
port 96 nsew signal output
flabel metal3 s 21424 50948 21504 51028 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[22]
port 97 nsew signal output
flabel metal3 s 21424 51620 21504 51700 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[23]
port 98 nsew signal output
flabel metal3 s 21424 52292 21504 52372 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[24]
port 99 nsew signal output
flabel metal3 s 21424 52964 21504 53044 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[25]
port 100 nsew signal output
flabel metal3 s 21424 53636 21504 53716 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[26]
port 101 nsew signal output
flabel metal3 s 21424 54308 21504 54388 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[27]
port 102 nsew signal output
flabel metal3 s 21424 54980 21504 55060 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[28]
port 103 nsew signal output
flabel metal3 s 21424 55652 21504 55732 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[29]
port 104 nsew signal output
flabel metal3 s 21424 37508 21504 37588 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[2]
port 105 nsew signal output
flabel metal3 s 21424 56324 21504 56404 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[30]
port 106 nsew signal output
flabel metal3 s 21424 56996 21504 57076 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[31]
port 107 nsew signal output
flabel metal3 s 21424 38180 21504 38260 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[3]
port 108 nsew signal output
flabel metal3 s 21424 38852 21504 38932 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[4]
port 109 nsew signal output
flabel metal3 s 21424 39524 21504 39604 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[5]
port 110 nsew signal output
flabel metal3 s 21424 40196 21504 40276 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[6]
port 111 nsew signal output
flabel metal3 s 21424 40868 21504 40948 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[7]
port 112 nsew signal output
flabel metal3 s 21424 41540 21504 41620 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[8]
port 113 nsew signal output
flabel metal3 s 21424 42212 21504 42292 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[9]
port 114 nsew signal output
flabel metal2 s 15800 85936 15880 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[0]
port 115 nsew signal output
flabel metal2 s 17720 85936 17800 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[10]
port 116 nsew signal output
flabel metal2 s 17912 85936 17992 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[11]
port 117 nsew signal output
flabel metal2 s 18104 85936 18184 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[12]
port 118 nsew signal output
flabel metal2 s 18296 85936 18376 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[13]
port 119 nsew signal output
flabel metal2 s 18488 85936 18568 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[14]
port 120 nsew signal output
flabel metal2 s 18680 85936 18760 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[15]
port 121 nsew signal output
flabel metal2 s 18872 85936 18952 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[16]
port 122 nsew signal output
flabel metal2 s 19064 85936 19144 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[17]
port 123 nsew signal output
flabel metal2 s 19256 85936 19336 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[18]
port 124 nsew signal output
flabel metal2 s 19448 85936 19528 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[19]
port 125 nsew signal output
flabel metal2 s 15992 85936 16072 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[1]
port 126 nsew signal output
flabel metal2 s 16184 85936 16264 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[2]
port 127 nsew signal output
flabel metal2 s 16376 85936 16456 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[3]
port 128 nsew signal output
flabel metal2 s 16568 85936 16648 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[4]
port 129 nsew signal output
flabel metal2 s 16760 85936 16840 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[5]
port 130 nsew signal output
flabel metal2 s 16952 85936 17032 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[6]
port 131 nsew signal output
flabel metal2 s 17144 85936 17224 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[7]
port 132 nsew signal output
flabel metal2 s 17336 85936 17416 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[8]
port 133 nsew signal output
flabel metal2 s 17528 85936 17608 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[9]
port 134 nsew signal output
flabel metal2 s 1784 85936 1864 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N1BEG[0]
port 135 nsew signal output
flabel metal2 s 1976 85936 2056 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N1BEG[1]
port 136 nsew signal output
flabel metal2 s 2168 85936 2248 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N1BEG[2]
port 137 nsew signal output
flabel metal2 s 2360 85936 2440 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N1BEG[3]
port 138 nsew signal output
flabel metal2 s 2552 85936 2632 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEG[0]
port 139 nsew signal output
flabel metal2 s 2744 85936 2824 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEG[1]
port 140 nsew signal output
flabel metal2 s 2936 85936 3016 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEG[2]
port 141 nsew signal output
flabel metal2 s 3128 85936 3208 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEG[3]
port 142 nsew signal output
flabel metal2 s 3320 85936 3400 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEG[4]
port 143 nsew signal output
flabel metal2 s 3512 85936 3592 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEG[5]
port 144 nsew signal output
flabel metal2 s 3704 85936 3784 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEG[6]
port 145 nsew signal output
flabel metal2 s 3896 85936 3976 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEG[7]
port 146 nsew signal output
flabel metal2 s 4088 85936 4168 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEGb[0]
port 147 nsew signal output
flabel metal2 s 4280 85936 4360 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEGb[1]
port 148 nsew signal output
flabel metal2 s 4472 85936 4552 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEGb[2]
port 149 nsew signal output
flabel metal2 s 4664 85936 4744 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEGb[3]
port 150 nsew signal output
flabel metal2 s 4856 85936 4936 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEGb[4]
port 151 nsew signal output
flabel metal2 s 5048 85936 5128 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEGb[5]
port 152 nsew signal output
flabel metal2 s 5240 85936 5320 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEGb[6]
port 153 nsew signal output
flabel metal2 s 5432 85936 5512 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEGb[7]
port 154 nsew signal output
flabel metal2 s 5624 85936 5704 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[0]
port 155 nsew signal output
flabel metal2 s 7544 85936 7624 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[10]
port 156 nsew signal output
flabel metal2 s 7736 85936 7816 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[11]
port 157 nsew signal output
flabel metal2 s 7928 85936 8008 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[12]
port 158 nsew signal output
flabel metal2 s 8120 85936 8200 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[13]
port 159 nsew signal output
flabel metal2 s 8312 85936 8392 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[14]
port 160 nsew signal output
flabel metal2 s 8504 85936 8584 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[15]
port 161 nsew signal output
flabel metal2 s 5816 85936 5896 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[1]
port 162 nsew signal output
flabel metal2 s 6008 85936 6088 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[2]
port 163 nsew signal output
flabel metal2 s 6200 85936 6280 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[3]
port 164 nsew signal output
flabel metal2 s 6392 85936 6472 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[4]
port 165 nsew signal output
flabel metal2 s 6584 85936 6664 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[5]
port 166 nsew signal output
flabel metal2 s 6776 85936 6856 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[6]
port 167 nsew signal output
flabel metal2 s 6968 85936 7048 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[7]
port 168 nsew signal output
flabel metal2 s 7160 85936 7240 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[8]
port 169 nsew signal output
flabel metal2 s 7352 85936 7432 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[9]
port 170 nsew signal output
flabel metal2 s 8696 85936 8776 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S1END[0]
port 171 nsew signal input
flabel metal2 s 8888 85936 8968 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S1END[1]
port 172 nsew signal input
flabel metal2 s 9080 85936 9160 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S1END[2]
port 173 nsew signal input
flabel metal2 s 9272 85936 9352 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S1END[3]
port 174 nsew signal input
flabel metal2 s 11000 85936 11080 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2END[0]
port 175 nsew signal input
flabel metal2 s 11192 85936 11272 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2END[1]
port 176 nsew signal input
flabel metal2 s 11384 85936 11464 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2END[2]
port 177 nsew signal input
flabel metal2 s 11576 85936 11656 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2END[3]
port 178 nsew signal input
flabel metal2 s 11768 85936 11848 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2END[4]
port 179 nsew signal input
flabel metal2 s 11960 85936 12040 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2END[5]
port 180 nsew signal input
flabel metal2 s 12152 85936 12232 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2END[6]
port 181 nsew signal input
flabel metal2 s 12344 85936 12424 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2END[7]
port 182 nsew signal input
flabel metal2 s 9464 85936 9544 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2MID[0]
port 183 nsew signal input
flabel metal2 s 9656 85936 9736 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2MID[1]
port 184 nsew signal input
flabel metal2 s 9848 85936 9928 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2MID[2]
port 185 nsew signal input
flabel metal2 s 10040 85936 10120 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2MID[3]
port 186 nsew signal input
flabel metal2 s 10232 85936 10312 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2MID[4]
port 187 nsew signal input
flabel metal2 s 10424 85936 10504 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2MID[5]
port 188 nsew signal input
flabel metal2 s 10616 85936 10696 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2MID[6]
port 189 nsew signal input
flabel metal2 s 10808 85936 10888 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2MID[7]
port 190 nsew signal input
flabel metal2 s 12536 85936 12616 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[0]
port 191 nsew signal input
flabel metal2 s 14456 85936 14536 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[10]
port 192 nsew signal input
flabel metal2 s 14648 85936 14728 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[11]
port 193 nsew signal input
flabel metal2 s 14840 85936 14920 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[12]
port 194 nsew signal input
flabel metal2 s 15032 85936 15112 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[13]
port 195 nsew signal input
flabel metal2 s 15224 85936 15304 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[14]
port 196 nsew signal input
flabel metal2 s 15416 85936 15496 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[15]
port 197 nsew signal input
flabel metal2 s 12728 85936 12808 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[1]
port 198 nsew signal input
flabel metal2 s 12920 85936 13000 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[2]
port 199 nsew signal input
flabel metal2 s 13112 85936 13192 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[3]
port 200 nsew signal input
flabel metal2 s 13304 85936 13384 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[4]
port 201 nsew signal input
flabel metal2 s 13496 85936 13576 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[5]
port 202 nsew signal input
flabel metal2 s 13688 85936 13768 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[6]
port 203 nsew signal input
flabel metal2 s 13880 85936 13960 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[7]
port 204 nsew signal input
flabel metal2 s 14072 85936 14152 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[8]
port 205 nsew signal input
flabel metal2 s 14264 85936 14344 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[9]
port 206 nsew signal input
flabel metal2 s 15608 85936 15688 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_UserCLKo
port 207 nsew signal output
flabel metal3 s 0 43052 80 43132 0 FreeSans 320 0 0 0 Tile_X0Y0_W1BEG[0]
port 208 nsew signal output
flabel metal3 s 0 43388 80 43468 0 FreeSans 320 0 0 0 Tile_X0Y0_W1BEG[1]
port 209 nsew signal output
flabel metal3 s 0 43724 80 43804 0 FreeSans 320 0 0 0 Tile_X0Y0_W1BEG[2]
port 210 nsew signal output
flabel metal3 s 0 44060 80 44140 0 FreeSans 320 0 0 0 Tile_X0Y0_W1BEG[3]
port 211 nsew signal output
flabel metal3 s 0 44396 80 44476 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEG[0]
port 212 nsew signal output
flabel metal3 s 0 44732 80 44812 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEG[1]
port 213 nsew signal output
flabel metal3 s 0 45068 80 45148 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEG[2]
port 214 nsew signal output
flabel metal3 s 0 45404 80 45484 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEG[3]
port 215 nsew signal output
flabel metal3 s 0 45740 80 45820 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEG[4]
port 216 nsew signal output
flabel metal3 s 0 46076 80 46156 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEG[5]
port 217 nsew signal output
flabel metal3 s 0 46412 80 46492 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEG[6]
port 218 nsew signal output
flabel metal3 s 0 46748 80 46828 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEG[7]
port 219 nsew signal output
flabel metal3 s 0 47084 80 47164 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEGb[0]
port 220 nsew signal output
flabel metal3 s 0 47420 80 47500 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEGb[1]
port 221 nsew signal output
flabel metal3 s 0 47756 80 47836 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEGb[2]
port 222 nsew signal output
flabel metal3 s 0 48092 80 48172 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEGb[3]
port 223 nsew signal output
flabel metal3 s 0 48428 80 48508 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEGb[4]
port 224 nsew signal output
flabel metal3 s 0 48764 80 48844 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEGb[5]
port 225 nsew signal output
flabel metal3 s 0 49100 80 49180 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEGb[6]
port 226 nsew signal output
flabel metal3 s 0 49436 80 49516 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEGb[7]
port 227 nsew signal output
flabel metal3 s 0 55148 80 55228 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[0]
port 228 nsew signal output
flabel metal3 s 0 58508 80 58588 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[10]
port 229 nsew signal output
flabel metal3 s 0 58844 80 58924 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[11]
port 230 nsew signal output
flabel metal3 s 0 55484 80 55564 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[1]
port 231 nsew signal output
flabel metal3 s 0 55820 80 55900 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[2]
port 232 nsew signal output
flabel metal3 s 0 56156 80 56236 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[3]
port 233 nsew signal output
flabel metal3 s 0 56492 80 56572 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[4]
port 234 nsew signal output
flabel metal3 s 0 56828 80 56908 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[5]
port 235 nsew signal output
flabel metal3 s 0 57164 80 57244 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[6]
port 236 nsew signal output
flabel metal3 s 0 57500 80 57580 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[7]
port 237 nsew signal output
flabel metal3 s 0 57836 80 57916 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[8]
port 238 nsew signal output
flabel metal3 s 0 58172 80 58252 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[9]
port 239 nsew signal output
flabel metal3 s 0 49772 80 49852 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[0]
port 240 nsew signal output
flabel metal3 s 0 53132 80 53212 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[10]
port 241 nsew signal output
flabel metal3 s 0 53468 80 53548 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[11]
port 242 nsew signal output
flabel metal3 s 0 53804 80 53884 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[12]
port 243 nsew signal output
flabel metal3 s 0 54140 80 54220 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[13]
port 244 nsew signal output
flabel metal3 s 0 54476 80 54556 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[14]
port 245 nsew signal output
flabel metal3 s 0 54812 80 54892 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[15]
port 246 nsew signal output
flabel metal3 s 0 50108 80 50188 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[1]
port 247 nsew signal output
flabel metal3 s 0 50444 80 50524 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[2]
port 248 nsew signal output
flabel metal3 s 0 50780 80 50860 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[3]
port 249 nsew signal output
flabel metal3 s 0 51116 80 51196 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[4]
port 250 nsew signal output
flabel metal3 s 0 51452 80 51532 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[5]
port 251 nsew signal output
flabel metal3 s 0 51788 80 51868 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[6]
port 252 nsew signal output
flabel metal3 s 0 52124 80 52204 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[7]
port 253 nsew signal output
flabel metal3 s 0 52460 80 52540 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[8]
port 254 nsew signal output
flabel metal3 s 0 52796 80 52876 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[9]
port 255 nsew signal output
flabel metal3 s 0 16172 80 16252 0 FreeSans 320 0 0 0 Tile_X0Y1_E1END[0]
port 256 nsew signal input
flabel metal3 s 0 16508 80 16588 0 FreeSans 320 0 0 0 Tile_X0Y1_E1END[1]
port 257 nsew signal input
flabel metal3 s 0 16844 80 16924 0 FreeSans 320 0 0 0 Tile_X0Y1_E1END[2]
port 258 nsew signal input
flabel metal3 s 0 17180 80 17260 0 FreeSans 320 0 0 0 Tile_X0Y1_E1END[3]
port 259 nsew signal input
flabel metal3 s 0 20204 80 20284 0 FreeSans 320 0 0 0 Tile_X0Y1_E2END[0]
port 260 nsew signal input
flabel metal3 s 0 20540 80 20620 0 FreeSans 320 0 0 0 Tile_X0Y1_E2END[1]
port 261 nsew signal input
flabel metal3 s 0 20876 80 20956 0 FreeSans 320 0 0 0 Tile_X0Y1_E2END[2]
port 262 nsew signal input
flabel metal3 s 0 21212 80 21292 0 FreeSans 320 0 0 0 Tile_X0Y1_E2END[3]
port 263 nsew signal input
flabel metal3 s 0 21548 80 21628 0 FreeSans 320 0 0 0 Tile_X0Y1_E2END[4]
port 264 nsew signal input
flabel metal3 s 0 21884 80 21964 0 FreeSans 320 0 0 0 Tile_X0Y1_E2END[5]
port 265 nsew signal input
flabel metal3 s 0 22220 80 22300 0 FreeSans 320 0 0 0 Tile_X0Y1_E2END[6]
port 266 nsew signal input
flabel metal3 s 0 22556 80 22636 0 FreeSans 320 0 0 0 Tile_X0Y1_E2END[7]
port 267 nsew signal input
flabel metal3 s 0 17516 80 17596 0 FreeSans 320 0 0 0 Tile_X0Y1_E2MID[0]
port 268 nsew signal input
flabel metal3 s 0 17852 80 17932 0 FreeSans 320 0 0 0 Tile_X0Y1_E2MID[1]
port 269 nsew signal input
flabel metal3 s 0 18188 80 18268 0 FreeSans 320 0 0 0 Tile_X0Y1_E2MID[2]
port 270 nsew signal input
flabel metal3 s 0 18524 80 18604 0 FreeSans 320 0 0 0 Tile_X0Y1_E2MID[3]
port 271 nsew signal input
flabel metal3 s 0 18860 80 18940 0 FreeSans 320 0 0 0 Tile_X0Y1_E2MID[4]
port 272 nsew signal input
flabel metal3 s 0 19196 80 19276 0 FreeSans 320 0 0 0 Tile_X0Y1_E2MID[5]
port 273 nsew signal input
flabel metal3 s 0 19532 80 19612 0 FreeSans 320 0 0 0 Tile_X0Y1_E2MID[6]
port 274 nsew signal input
flabel metal3 s 0 19868 80 19948 0 FreeSans 320 0 0 0 Tile_X0Y1_E2MID[7]
port 275 nsew signal input
flabel metal3 s 0 28268 80 28348 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[0]
port 276 nsew signal input
flabel metal3 s 0 31628 80 31708 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[10]
port 277 nsew signal input
flabel metal3 s 0 31964 80 32044 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[11]
port 278 nsew signal input
flabel metal3 s 0 28604 80 28684 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[1]
port 279 nsew signal input
flabel metal3 s 0 28940 80 29020 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[2]
port 280 nsew signal input
flabel metal3 s 0 29276 80 29356 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[3]
port 281 nsew signal input
flabel metal3 s 0 29612 80 29692 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[4]
port 282 nsew signal input
flabel metal3 s 0 29948 80 30028 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[5]
port 283 nsew signal input
flabel metal3 s 0 30284 80 30364 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[6]
port 284 nsew signal input
flabel metal3 s 0 30620 80 30700 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[7]
port 285 nsew signal input
flabel metal3 s 0 30956 80 31036 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[8]
port 286 nsew signal input
flabel metal3 s 0 31292 80 31372 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[9]
port 287 nsew signal input
flabel metal3 s 0 22892 80 22972 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[0]
port 288 nsew signal input
flabel metal3 s 0 26252 80 26332 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[10]
port 289 nsew signal input
flabel metal3 s 0 26588 80 26668 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[11]
port 290 nsew signal input
flabel metal3 s 0 26924 80 27004 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[12]
port 291 nsew signal input
flabel metal3 s 0 27260 80 27340 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[13]
port 292 nsew signal input
flabel metal3 s 0 27596 80 27676 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[14]
port 293 nsew signal input
flabel metal3 s 0 27932 80 28012 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[15]
port 294 nsew signal input
flabel metal3 s 0 23228 80 23308 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[1]
port 295 nsew signal input
flabel metal3 s 0 23564 80 23644 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[2]
port 296 nsew signal input
flabel metal3 s 0 23900 80 23980 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[3]
port 297 nsew signal input
flabel metal3 s 0 24236 80 24316 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[4]
port 298 nsew signal input
flabel metal3 s 0 24572 80 24652 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[5]
port 299 nsew signal input
flabel metal3 s 0 24908 80 24988 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[6]
port 300 nsew signal input
flabel metal3 s 0 25244 80 25324 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[7]
port 301 nsew signal input
flabel metal3 s 0 25580 80 25660 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[8]
port 302 nsew signal input
flabel metal3 s 0 25916 80 25996 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[9]
port 303 nsew signal input
flabel metal3 s 0 32300 80 32380 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[0]
port 304 nsew signal input
flabel metal3 s 0 35660 80 35740 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[10]
port 305 nsew signal input
flabel metal3 s 0 35996 80 36076 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[11]
port 306 nsew signal input
flabel metal3 s 0 36332 80 36412 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[12]
port 307 nsew signal input
flabel metal3 s 0 36668 80 36748 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[13]
port 308 nsew signal input
flabel metal3 s 0 37004 80 37084 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[14]
port 309 nsew signal input
flabel metal3 s 0 37340 80 37420 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[15]
port 310 nsew signal input
flabel metal3 s 0 37676 80 37756 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[16]
port 311 nsew signal input
flabel metal3 s 0 38012 80 38092 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[17]
port 312 nsew signal input
flabel metal3 s 0 38348 80 38428 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[18]
port 313 nsew signal input
flabel metal3 s 0 38684 80 38764 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[19]
port 314 nsew signal input
flabel metal3 s 0 32636 80 32716 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[1]
port 315 nsew signal input
flabel metal3 s 0 39020 80 39100 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[20]
port 316 nsew signal input
flabel metal3 s 0 39356 80 39436 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[21]
port 317 nsew signal input
flabel metal3 s 0 39692 80 39772 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[22]
port 318 nsew signal input
flabel metal3 s 0 40028 80 40108 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[23]
port 319 nsew signal input
flabel metal3 s 0 40364 80 40444 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[24]
port 320 nsew signal input
flabel metal3 s 0 40700 80 40780 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[25]
port 321 nsew signal input
flabel metal3 s 0 41036 80 41116 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[26]
port 322 nsew signal input
flabel metal3 s 0 41372 80 41452 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[27]
port 323 nsew signal input
flabel metal3 s 0 41708 80 41788 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[28]
port 324 nsew signal input
flabel metal3 s 0 42044 80 42124 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[29]
port 325 nsew signal input
flabel metal3 s 0 32972 80 33052 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[2]
port 326 nsew signal input
flabel metal3 s 0 42380 80 42460 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[30]
port 327 nsew signal input
flabel metal3 s 0 42716 80 42796 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[31]
port 328 nsew signal input
flabel metal3 s 0 33308 80 33388 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[3]
port 329 nsew signal input
flabel metal3 s 0 33644 80 33724 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[4]
port 330 nsew signal input
flabel metal3 s 0 33980 80 34060 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[5]
port 331 nsew signal input
flabel metal3 s 0 34316 80 34396 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[6]
port 332 nsew signal input
flabel metal3 s 0 34652 80 34732 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[7]
port 333 nsew signal input
flabel metal3 s 0 34988 80 35068 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[8]
port 334 nsew signal input
flabel metal3 s 0 35324 80 35404 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[9]
port 335 nsew signal input
flabel metal3 s 21424 57668 21504 57748 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[0]
port 336 nsew signal output
flabel metal3 s 21424 64388 21504 64468 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[10]
port 337 nsew signal output
flabel metal3 s 21424 65060 21504 65140 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[11]
port 338 nsew signal output
flabel metal3 s 21424 65732 21504 65812 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[12]
port 339 nsew signal output
flabel metal3 s 21424 66404 21504 66484 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[13]
port 340 nsew signal output
flabel metal3 s 21424 67076 21504 67156 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[14]
port 341 nsew signal output
flabel metal3 s 21424 67748 21504 67828 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[15]
port 342 nsew signal output
flabel metal3 s 21424 68420 21504 68500 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[16]
port 343 nsew signal output
flabel metal3 s 21424 69092 21504 69172 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[17]
port 344 nsew signal output
flabel metal3 s 21424 69764 21504 69844 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[18]
port 345 nsew signal output
flabel metal3 s 21424 70436 21504 70516 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[19]
port 346 nsew signal output
flabel metal3 s 21424 58340 21504 58420 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[1]
port 347 nsew signal output
flabel metal3 s 21424 71108 21504 71188 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[20]
port 348 nsew signal output
flabel metal3 s 21424 71780 21504 71860 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[21]
port 349 nsew signal output
flabel metal3 s 21424 72452 21504 72532 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[22]
port 350 nsew signal output
flabel metal3 s 21424 73124 21504 73204 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[23]
port 351 nsew signal output
flabel metal3 s 21424 73796 21504 73876 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[24]
port 352 nsew signal output
flabel metal3 s 21424 74468 21504 74548 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[25]
port 353 nsew signal output
flabel metal3 s 21424 75140 21504 75220 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[26]
port 354 nsew signal output
flabel metal3 s 21424 75812 21504 75892 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[27]
port 355 nsew signal output
flabel metal3 s 21424 76484 21504 76564 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[28]
port 356 nsew signal output
flabel metal3 s 21424 77156 21504 77236 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[29]
port 357 nsew signal output
flabel metal3 s 21424 59012 21504 59092 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[2]
port 358 nsew signal output
flabel metal3 s 21424 77828 21504 77908 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[30]
port 359 nsew signal output
flabel metal3 s 21424 78500 21504 78580 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[31]
port 360 nsew signal output
flabel metal3 s 21424 59684 21504 59764 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[3]
port 361 nsew signal output
flabel metal3 s 21424 60356 21504 60436 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[4]
port 362 nsew signal output
flabel metal3 s 21424 61028 21504 61108 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[5]
port 363 nsew signal output
flabel metal3 s 21424 61700 21504 61780 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[6]
port 364 nsew signal output
flabel metal3 s 21424 62372 21504 62452 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[7]
port 365 nsew signal output
flabel metal3 s 21424 63044 21504 63124 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[8]
port 366 nsew signal output
flabel metal3 s 21424 63716 21504 63796 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[9]
port 367 nsew signal output
flabel metal2 s 15800 0 15880 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[0]
port 368 nsew signal input
flabel metal2 s 17720 0 17800 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[10]
port 369 nsew signal input
flabel metal2 s 17912 0 17992 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[11]
port 370 nsew signal input
flabel metal2 s 18104 0 18184 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[12]
port 371 nsew signal input
flabel metal2 s 18296 0 18376 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[13]
port 372 nsew signal input
flabel metal2 s 18488 0 18568 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[14]
port 373 nsew signal input
flabel metal2 s 18680 0 18760 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[15]
port 374 nsew signal input
flabel metal2 s 18872 0 18952 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[16]
port 375 nsew signal input
flabel metal2 s 19064 0 19144 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[17]
port 376 nsew signal input
flabel metal2 s 19256 0 19336 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[18]
port 377 nsew signal input
flabel metal2 s 19448 0 19528 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[19]
port 378 nsew signal input
flabel metal2 s 15992 0 16072 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[1]
port 379 nsew signal input
flabel metal2 s 16184 0 16264 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[2]
port 380 nsew signal input
flabel metal2 s 16376 0 16456 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[3]
port 381 nsew signal input
flabel metal2 s 16568 0 16648 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[4]
port 382 nsew signal input
flabel metal2 s 16760 0 16840 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[5]
port 383 nsew signal input
flabel metal2 s 16952 0 17032 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[6]
port 384 nsew signal input
flabel metal2 s 17144 0 17224 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[7]
port 385 nsew signal input
flabel metal2 s 17336 0 17416 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[8]
port 386 nsew signal input
flabel metal2 s 17528 0 17608 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[9]
port 387 nsew signal input
flabel metal2 s 1784 0 1864 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N1END[0]
port 388 nsew signal input
flabel metal2 s 1976 0 2056 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N1END[1]
port 389 nsew signal input
flabel metal2 s 2168 0 2248 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N1END[2]
port 390 nsew signal input
flabel metal2 s 2360 0 2440 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N1END[3]
port 391 nsew signal input
flabel metal2 s 4088 0 4168 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2END[0]
port 392 nsew signal input
flabel metal2 s 4280 0 4360 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2END[1]
port 393 nsew signal input
flabel metal2 s 4472 0 4552 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2END[2]
port 394 nsew signal input
flabel metal2 s 4664 0 4744 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2END[3]
port 395 nsew signal input
flabel metal2 s 4856 0 4936 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2END[4]
port 396 nsew signal input
flabel metal2 s 5048 0 5128 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2END[5]
port 397 nsew signal input
flabel metal2 s 5240 0 5320 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2END[6]
port 398 nsew signal input
flabel metal2 s 5432 0 5512 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2END[7]
port 399 nsew signal input
flabel metal2 s 2552 0 2632 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2MID[0]
port 400 nsew signal input
flabel metal2 s 2744 0 2824 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2MID[1]
port 401 nsew signal input
flabel metal2 s 2936 0 3016 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2MID[2]
port 402 nsew signal input
flabel metal2 s 3128 0 3208 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2MID[3]
port 403 nsew signal input
flabel metal2 s 3320 0 3400 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2MID[4]
port 404 nsew signal input
flabel metal2 s 3512 0 3592 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2MID[5]
port 405 nsew signal input
flabel metal2 s 3704 0 3784 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2MID[6]
port 406 nsew signal input
flabel metal2 s 3896 0 3976 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2MID[7]
port 407 nsew signal input
flabel metal2 s 5624 0 5704 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[0]
port 408 nsew signal input
flabel metal2 s 7544 0 7624 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[10]
port 409 nsew signal input
flabel metal2 s 7736 0 7816 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[11]
port 410 nsew signal input
flabel metal2 s 7928 0 8008 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[12]
port 411 nsew signal input
flabel metal2 s 8120 0 8200 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[13]
port 412 nsew signal input
flabel metal2 s 8312 0 8392 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[14]
port 413 nsew signal input
flabel metal2 s 8504 0 8584 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[15]
port 414 nsew signal input
flabel metal2 s 5816 0 5896 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[1]
port 415 nsew signal input
flabel metal2 s 6008 0 6088 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[2]
port 416 nsew signal input
flabel metal2 s 6200 0 6280 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[3]
port 417 nsew signal input
flabel metal2 s 6392 0 6472 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[4]
port 418 nsew signal input
flabel metal2 s 6584 0 6664 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[5]
port 419 nsew signal input
flabel metal2 s 6776 0 6856 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[6]
port 420 nsew signal input
flabel metal2 s 6968 0 7048 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[7]
port 421 nsew signal input
flabel metal2 s 7160 0 7240 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[8]
port 422 nsew signal input
flabel metal2 s 7352 0 7432 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[9]
port 423 nsew signal input
flabel metal2 s 8696 0 8776 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S1BEG[0]
port 424 nsew signal output
flabel metal2 s 8888 0 8968 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S1BEG[1]
port 425 nsew signal output
flabel metal2 s 9080 0 9160 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S1BEG[2]
port 426 nsew signal output
flabel metal2 s 9272 0 9352 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S1BEG[3]
port 427 nsew signal output
flabel metal2 s 9464 0 9544 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEG[0]
port 428 nsew signal output
flabel metal2 s 9656 0 9736 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEG[1]
port 429 nsew signal output
flabel metal2 s 9848 0 9928 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEG[2]
port 430 nsew signal output
flabel metal2 s 10040 0 10120 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEG[3]
port 431 nsew signal output
flabel metal2 s 10232 0 10312 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEG[4]
port 432 nsew signal output
flabel metal2 s 10424 0 10504 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEG[5]
port 433 nsew signal output
flabel metal2 s 10616 0 10696 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEG[6]
port 434 nsew signal output
flabel metal2 s 10808 0 10888 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEG[7]
port 435 nsew signal output
flabel metal2 s 11000 0 11080 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEGb[0]
port 436 nsew signal output
flabel metal2 s 11192 0 11272 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEGb[1]
port 437 nsew signal output
flabel metal2 s 11384 0 11464 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEGb[2]
port 438 nsew signal output
flabel metal2 s 11576 0 11656 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEGb[3]
port 439 nsew signal output
flabel metal2 s 11768 0 11848 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEGb[4]
port 440 nsew signal output
flabel metal2 s 11960 0 12040 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEGb[5]
port 441 nsew signal output
flabel metal2 s 12152 0 12232 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEGb[6]
port 442 nsew signal output
flabel metal2 s 12344 0 12424 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEGb[7]
port 443 nsew signal output
flabel metal2 s 12536 0 12616 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[0]
port 444 nsew signal output
flabel metal2 s 14456 0 14536 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[10]
port 445 nsew signal output
flabel metal2 s 14648 0 14728 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[11]
port 446 nsew signal output
flabel metal2 s 14840 0 14920 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[12]
port 447 nsew signal output
flabel metal2 s 15032 0 15112 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[13]
port 448 nsew signal output
flabel metal2 s 15224 0 15304 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[14]
port 449 nsew signal output
flabel metal2 s 15416 0 15496 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[15]
port 450 nsew signal output
flabel metal2 s 12728 0 12808 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[1]
port 451 nsew signal output
flabel metal2 s 12920 0 13000 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[2]
port 452 nsew signal output
flabel metal2 s 13112 0 13192 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[3]
port 453 nsew signal output
flabel metal2 s 13304 0 13384 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[4]
port 454 nsew signal output
flabel metal2 s 13496 0 13576 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[5]
port 455 nsew signal output
flabel metal2 s 13688 0 13768 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[6]
port 456 nsew signal output
flabel metal2 s 13880 0 13960 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[7]
port 457 nsew signal output
flabel metal2 s 14072 0 14152 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[8]
port 458 nsew signal output
flabel metal2 s 14264 0 14344 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[9]
port 459 nsew signal output
flabel metal2 s 15608 0 15688 80 0 FreeSans 320 0 0 0 Tile_X0Y1_UserCLK
port 460 nsew signal input
flabel metal3 s 0 44 80 124 0 FreeSans 320 0 0 0 Tile_X0Y1_W1BEG[0]
port 461 nsew signal output
flabel metal3 s 0 380 80 460 0 FreeSans 320 0 0 0 Tile_X0Y1_W1BEG[1]
port 462 nsew signal output
flabel metal3 s 0 716 80 796 0 FreeSans 320 0 0 0 Tile_X0Y1_W1BEG[2]
port 463 nsew signal output
flabel metal3 s 0 1052 80 1132 0 FreeSans 320 0 0 0 Tile_X0Y1_W1BEG[3]
port 464 nsew signal output
flabel metal3 s 0 1388 80 1468 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEG[0]
port 465 nsew signal output
flabel metal3 s 0 1724 80 1804 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEG[1]
port 466 nsew signal output
flabel metal3 s 0 2060 80 2140 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEG[2]
port 467 nsew signal output
flabel metal3 s 0 2396 80 2476 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEG[3]
port 468 nsew signal output
flabel metal3 s 0 2732 80 2812 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEG[4]
port 469 nsew signal output
flabel metal3 s 0 3068 80 3148 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEG[5]
port 470 nsew signal output
flabel metal3 s 0 3404 80 3484 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEG[6]
port 471 nsew signal output
flabel metal3 s 0 3740 80 3820 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEG[7]
port 472 nsew signal output
flabel metal3 s 0 4076 80 4156 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEGb[0]
port 473 nsew signal output
flabel metal3 s 0 4412 80 4492 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEGb[1]
port 474 nsew signal output
flabel metal3 s 0 4748 80 4828 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEGb[2]
port 475 nsew signal output
flabel metal3 s 0 5084 80 5164 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEGb[3]
port 476 nsew signal output
flabel metal3 s 0 5420 80 5500 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEGb[4]
port 477 nsew signal output
flabel metal3 s 0 5756 80 5836 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEGb[5]
port 478 nsew signal output
flabel metal3 s 0 6092 80 6172 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEGb[6]
port 479 nsew signal output
flabel metal3 s 0 6428 80 6508 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEGb[7]
port 480 nsew signal output
flabel metal3 s 0 12140 80 12220 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[0]
port 481 nsew signal output
flabel metal3 s 0 15500 80 15580 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[10]
port 482 nsew signal output
flabel metal3 s 0 15836 80 15916 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[11]
port 483 nsew signal output
flabel metal3 s 0 12476 80 12556 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[1]
port 484 nsew signal output
flabel metal3 s 0 12812 80 12892 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[2]
port 485 nsew signal output
flabel metal3 s 0 13148 80 13228 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[3]
port 486 nsew signal output
flabel metal3 s 0 13484 80 13564 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[4]
port 487 nsew signal output
flabel metal3 s 0 13820 80 13900 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[5]
port 488 nsew signal output
flabel metal3 s 0 14156 80 14236 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[6]
port 489 nsew signal output
flabel metal3 s 0 14492 80 14572 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[7]
port 490 nsew signal output
flabel metal3 s 0 14828 80 14908 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[8]
port 491 nsew signal output
flabel metal3 s 0 15164 80 15244 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[9]
port 492 nsew signal output
flabel metal3 s 0 6764 80 6844 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[0]
port 493 nsew signal output
flabel metal3 s 0 10124 80 10204 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[10]
port 494 nsew signal output
flabel metal3 s 0 10460 80 10540 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[11]
port 495 nsew signal output
flabel metal3 s 0 10796 80 10876 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[12]
port 496 nsew signal output
flabel metal3 s 0 11132 80 11212 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[13]
port 497 nsew signal output
flabel metal3 s 0 11468 80 11548 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[14]
port 498 nsew signal output
flabel metal3 s 0 11804 80 11884 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[15]
port 499 nsew signal output
flabel metal3 s 0 7100 80 7180 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[1]
port 500 nsew signal output
flabel metal3 s 0 7436 80 7516 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[2]
port 501 nsew signal output
flabel metal3 s 0 7772 80 7852 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[3]
port 502 nsew signal output
flabel metal3 s 0 8108 80 8188 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[4]
port 503 nsew signal output
flabel metal3 s 0 8444 80 8524 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[5]
port 504 nsew signal output
flabel metal3 s 0 8780 80 8860 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[6]
port 505 nsew signal output
flabel metal3 s 0 9116 80 9196 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[7]
port 506 nsew signal output
flabel metal3 s 0 9452 80 9532 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[8]
port 507 nsew signal output
flabel metal3 s 0 9788 80 9868 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[9]
port 508 nsew signal output
flabel metal3 s 21424 28772 21504 28852 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT0
port 509 nsew signal output
flabel metal3 s 21424 29444 21504 29524 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT1
port 510 nsew signal output
flabel metal3 s 21424 30116 21504 30196 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT2
port 511 nsew signal output
flabel metal3 s 21424 30788 21504 30868 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT3
port 512 nsew signal output
flabel metal3 s 21424 31460 21504 31540 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT4
port 513 nsew signal output
flabel metal3 s 21424 32132 21504 32212 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT5
port 514 nsew signal output
flabel metal3 s 21424 32804 21504 32884 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT6
port 515 nsew signal output
flabel metal3 s 21424 33476 21504 33556 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT7
port 516 nsew signal output
flabel metal3 s 21424 18020 21504 18100 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT0
port 517 nsew signal input
flabel metal3 s 21424 18692 21504 18772 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT1
port 518 nsew signal input
flabel metal3 s 21424 19364 21504 19444 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT2
port 519 nsew signal input
flabel metal3 s 21424 20036 21504 20116 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT3
port 520 nsew signal input
flabel metal3 s 21424 20708 21504 20788 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT4
port 521 nsew signal input
flabel metal3 s 21424 21380 21504 21460 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT5
port 522 nsew signal input
flabel metal3 s 21424 22052 21504 22132 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT6
port 523 nsew signal input
flabel metal3 s 21424 22724 21504 22804 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT7
port 524 nsew signal input
flabel metal3 s 21424 12644 21504 12724 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT0
port 525 nsew signal input
flabel metal3 s 21424 13316 21504 13396 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT1
port 526 nsew signal input
flabel metal3 s 21424 13988 21504 14068 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT2
port 527 nsew signal input
flabel metal3 s 21424 14660 21504 14740 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT3
port 528 nsew signal input
flabel metal3 s 21424 15332 21504 15412 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT4
port 529 nsew signal input
flabel metal3 s 21424 16004 21504 16084 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT5
port 530 nsew signal input
flabel metal3 s 21424 16676 21504 16756 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT6
port 531 nsew signal input
flabel metal3 s 21424 17348 21504 17428 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT7
port 532 nsew signal input
flabel metal3 s 21424 23396 21504 23476 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT0
port 533 nsew signal output
flabel metal3 s 21424 24068 21504 24148 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT1
port 534 nsew signal output
flabel metal3 s 21424 24740 21504 24820 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT2
port 535 nsew signal output
flabel metal3 s 21424 25412 21504 25492 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT3
port 536 nsew signal output
flabel metal3 s 21424 26084 21504 26164 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT4
port 537 nsew signal output
flabel metal3 s 21424 26756 21504 26836 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT5
port 538 nsew signal output
flabel metal3 s 21424 27428 21504 27508 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT6
port 539 nsew signal output
flabel metal3 s 21424 28100 21504 28180 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT7
port 540 nsew signal output
flabel metal3 s 21424 7268 21504 7348 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT0
port 541 nsew signal input
flabel metal3 s 21424 7940 21504 8020 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT1
port 542 nsew signal input
flabel metal3 s 21424 8612 21504 8692 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT2
port 543 nsew signal input
flabel metal3 s 21424 9284 21504 9364 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT3
port 544 nsew signal input
flabel metal3 s 21424 9956 21504 10036 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT4
port 545 nsew signal input
flabel metal3 s 21424 10628 21504 10708 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT5
port 546 nsew signal input
flabel metal3 s 21424 11300 21504 11380 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT6
port 547 nsew signal input
flabel metal3 s 21424 11972 21504 12052 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT7
port 548 nsew signal input
flabel metal6 s 4892 0 5332 86016 0 FreeSans 2624 90 0 0 VGND
port 549 nsew ground bidirectional
flabel metal6 s 4892 0 5332 328 0 FreeSans 2624 0 0 0 VGND
port 549 nsew ground bidirectional
flabel metal6 s 4892 85688 5332 86016 0 FreeSans 2624 0 0 0 VGND
port 549 nsew ground bidirectional
flabel metal6 s 20012 0 20452 86016 0 FreeSans 2624 90 0 0 VGND
port 549 nsew ground bidirectional
flabel metal6 s 20012 0 20452 328 0 FreeSans 2624 0 0 0 VGND
port 549 nsew ground bidirectional
flabel metal6 s 20012 85688 20452 86016 0 FreeSans 2624 0 0 0 VGND
port 549 nsew ground bidirectional
flabel metal6 s 3652 0 4092 86016 0 FreeSans 2624 90 0 0 VPWR
port 550 nsew power bidirectional
flabel metal6 s 3652 0 4092 328 0 FreeSans 2624 0 0 0 VPWR
port 550 nsew power bidirectional
flabel metal6 s 3652 85688 4092 86016 0 FreeSans 2624 0 0 0 VPWR
port 550 nsew power bidirectional
flabel metal6 s 18772 0 19212 86016 0 FreeSans 2624 90 0 0 VPWR
port 550 nsew power bidirectional
flabel metal6 s 18772 0 19212 328 0 FreeSans 2624 0 0 0 VPWR
port 550 nsew power bidirectional
flabel metal6 s 18772 85688 19212 86016 0 FreeSans 2624 0 0 0 VPWR
port 550 nsew power bidirectional
rlabel metal1 10802 83916 10802 83916 0 VGND
rlabel metal1 10752 84672 10752 84672 0 VPWR
rlabel metal3 18384 34944 18384 34944 0 CLK_TT_PROJECT
rlabel metal3 20658 34188 20658 34188 0 ENA_TT_PROJECT
rlabel metal3 13440 35826 13440 35826 0 RST_N_TT_PROJECT
rlabel metal3 480 59178 480 59178 0 Tile_X0Y0_E1END[0]
rlabel metal2 12384 59766 12384 59766 0 Tile_X0Y0_E1END[1]
rlabel metal3 126 59892 126 59892 0 Tile_X0Y0_E1END[2]
rlabel metal2 4848 68628 4848 68628 0 Tile_X0Y0_E1END[3]
rlabel metal3 2112 63126 2112 63126 0 Tile_X0Y0_E2END[0]
rlabel metal2 9696 61152 9696 61152 0 Tile_X0Y0_E2END[1]
rlabel metal4 1440 67326 1440 67326 0 Tile_X0Y0_E2END[2]
rlabel metal3 2112 64302 2112 64302 0 Tile_X0Y0_E2END[3]
rlabel metal2 2496 72114 2496 72114 0 Tile_X0Y0_E2END[4]
rlabel metal2 10080 66318 10080 66318 0 Tile_X0Y0_E2END[5]
rlabel metal2 2448 68712 2448 68712 0 Tile_X0Y0_E2END[6]
rlabel metal2 2256 71904 2256 71904 0 Tile_X0Y0_E2END[7]
rlabel metal2 2304 61068 2304 61068 0 Tile_X0Y0_E2MID[0]
rlabel metal3 78 60900 78 60900 0 Tile_X0Y0_E2MID[1]
rlabel metal3 1134 61236 1134 61236 0 Tile_X0Y0_E2MID[2]
rlabel metal2 2400 62790 2400 62790 0 Tile_X0Y0_E2MID[3]
rlabel metal3 1776 72156 1776 72156 0 Tile_X0Y0_E2MID[4]
rlabel metal2 9696 67830 9696 67830 0 Tile_X0Y0_E2MID[5]
rlabel metal3 1038 62580 1038 62580 0 Tile_X0Y0_E2MID[6]
rlabel metal2 1728 65394 1728 65394 0 Tile_X0Y0_E2MID[7]
rlabel metal2 6144 69930 6144 69930 0 Tile_X0Y0_E6END[0]
rlabel metal3 6336 74718 6336 74718 0 Tile_X0Y0_E6END[10]
rlabel metal2 6480 72660 6480 72660 0 Tile_X0Y0_E6END[11]
rlabel metal2 13056 66066 13056 66066 0 Tile_X0Y0_E6END[1]
rlabel metal3 2304 71904 2304 71904 0 Tile_X0Y0_E6END[2]
rlabel metal3 558 72324 558 72324 0 Tile_X0Y0_E6END[3]
rlabel metal3 846 72660 846 72660 0 Tile_X0Y0_E6END[4]
rlabel metal3 126 72996 126 72996 0 Tile_X0Y0_E6END[5]
rlabel metal3 1824 69216 1824 69216 0 Tile_X0Y0_E6END[6]
rlabel metal2 1920 74634 1920 74634 0 Tile_X0Y0_E6END[7]
rlabel metal2 1968 71568 1968 71568 0 Tile_X0Y0_E6END[8]
rlabel metal3 318 74340 318 74340 0 Tile_X0Y0_E6END[9]
rlabel metal3 1290 65940 1290 65940 0 Tile_X0Y0_EE4END[0]
rlabel metal2 15360 67746 15360 67746 0 Tile_X0Y0_EE4END[10]
rlabel metal2 5568 70140 5568 70140 0 Tile_X0Y0_EE4END[11]
rlabel metal3 606 69972 606 69972 0 Tile_X0Y0_EE4END[12]
rlabel metal2 14400 69888 14400 69888 0 Tile_X0Y0_EE4END[13]
rlabel metal3 702 70644 702 70644 0 Tile_X0Y0_EE4END[14]
rlabel metal2 9120 71568 9120 71568 0 Tile_X0Y0_EE4END[15]
rlabel metal2 12192 66864 12192 66864 0 Tile_X0Y0_EE4END[1]
rlabel metal3 606 66612 606 66612 0 Tile_X0Y0_EE4END[2]
rlabel metal3 462 66948 462 66948 0 Tile_X0Y0_EE4END[3]
rlabel metal2 8064 65520 8064 65520 0 Tile_X0Y0_EE4END[4]
rlabel metal3 606 67620 606 67620 0 Tile_X0Y0_EE4END[5]
rlabel metal2 18048 67830 18048 67830 0 Tile_X0Y0_EE4END[6]
rlabel metal4 4800 68922 4800 68922 0 Tile_X0Y0_EE4END[7]
rlabel metal2 5184 68544 5184 68544 0 Tile_X0Y0_EE4END[8]
rlabel metal3 11958 66864 11958 66864 0 Tile_X0Y0_EE4END[9]
rlabel metal2 7488 56574 7488 56574 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit0.Q
rlabel metal2 9024 56403 9024 56403 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit1.Q
rlabel via2 11520 69134 11520 69134 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit10.Q
rlabel metal2 9984 69426 9984 69426 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit11.Q
rlabel metal2 13584 71652 13584 71652 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit12.Q
rlabel metal2 11904 72450 11904 72450 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit13.Q
rlabel via1 5232 79720 5232 79720 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit14.Q
rlabel metal2 3456 82572 3456 82572 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit15.Q
rlabel metal2 6720 42420 6720 42420 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit16.Q
rlabel metal2 4992 42798 4992 42798 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit17.Q
rlabel metal2 12768 74928 12768 74928 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit18.Q
rlabel metal2 10848 75138 10848 75138 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit19.Q
rlabel metal2 13248 48846 13248 48846 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit2.Q
rlabel metal2 13440 69804 13440 69804 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit20.Q
rlabel metal2 11616 70224 11616 70224 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit21.Q
rlabel metal2 7008 80805 7008 80805 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit22.Q
rlabel metal2 5520 82572 5520 82572 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit23.Q
rlabel metal2 7008 59724 7008 59724 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit24.Q
rlabel metal3 7920 60900 7920 60900 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit25.Q
rlabel metal2 13536 59724 13536 59724 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit26.Q
rlabel metal2 12720 59556 12720 59556 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit27.Q
rlabel metal3 17853 63924 17853 63924 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit28.Q
rlabel metal3 17760 63336 17760 63336 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit29.Q
rlabel via1 14832 48799 14832 48799 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit3.Q
rlabel metal2 7301 73542 7301 73542 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit30.Q
rlabel metal2 7104 73752 7104 73752 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit31.Q
rlabel metal2 16752 56532 16752 56532 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit4.Q
rlabel metal2 18336 57715 18336 57715 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit5.Q
rlabel metal2 8160 76272 8160 76272 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit6.Q
rlabel metal2 9696 76059 9696 76059 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit7.Q
rlabel metal2 4416 79293 4416 79293 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit8.Q
rlabel metal2 2832 77532 2832 77532 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit9.Q
rlabel metal2 14832 63336 14832 63336 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit0.Q
rlabel metal2 16224 64176 16224 64176 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit1.Q
rlabel metal2 13056 54894 13056 54894 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit10.Q
rlabel metal2 14592 55101 14592 55101 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit11.Q
rlabel metal3 17424 59388 17424 59388 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit12.Q
rlabel metal2 19872 58968 19872 58968 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit13.Q
rlabel metal2 8448 78162 8448 78162 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit14.Q
rlabel metal2 9984 78505 9984 78505 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit15.Q
rlabel metal2 6912 53550 6912 53550 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit16.Q
rlabel metal2 8448 53179 8448 53179 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit17.Q
rlabel metal2 12624 52500 12624 52500 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit18.Q
rlabel metal2 14208 52843 14208 52843 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit19.Q
rlabel metal3 18000 68208 18000 68208 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit2.Q
rlabel metal2 17568 60312 17568 60312 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit20.Q
rlabel metal2 19104 60109 19104 60109 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit21.Q
rlabel metal2 7728 77532 7728 77532 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit22.Q
rlabel via1 9360 77527 9360 77527 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit23.Q
rlabel metal2 7584 53382 7584 53382 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit24.Q
rlabel via2 9120 53337 9120 53337 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit25.Q
rlabel metal2 13248 51282 13248 51282 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit26.Q
rlabel metal2 14832 51051 14832 51051 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit27.Q
rlabel metal2 17472 56994 17472 56994 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit28.Q
rlabel metal2 19008 56487 19008 56487 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit29.Q
rlabel metal2 19920 67620 19920 67620 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit3.Q
rlabel metal2 8448 76986 8448 76986 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit30.Q
rlabel via1 10032 76696 10032 76696 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit31.Q
rlabel metal2 19104 67370 19104 67370 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit4.Q
rlabel metal3 8256 71988 8256 71988 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit5.Q
rlabel metal2 9312 72114 9312 72114 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit6.Q
rlabel metal2 9216 71736 9216 71736 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit7.Q
rlabel metal2 7200 57918 7200 57918 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit8.Q
rlabel metal2 8736 57715 8736 57715 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit9.Q
rlabel via1 6576 47287 6576 47287 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit0.Q
rlabel metal2 4896 47292 4896 47292 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit1.Q
rlabel metal2 16704 53589 16704 53589 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit10.Q
rlabel metal2 15168 53592 15168 53592 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit11.Q
rlabel metal2 13152 57337 13152 57337 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit12.Q
rlabel metal3 11616 56994 11616 56994 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit13.Q
rlabel metal2 5400 57866 5400 57866 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit14.Q
rlabel metal3 3408 57876 3408 57876 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit15.Q
rlabel metal3 5856 69300 5856 69300 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit16.Q
rlabel metal2 7200 68502 7200 68502 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit17.Q
rlabel metal2 4464 68460 4464 68460 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit18.Q
rlabel metal3 12528 66948 12528 66948 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit19.Q
rlabel via1 19152 50311 19152 50311 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit2.Q
rlabel metal2 14160 66780 14160 66780 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit20.Q
rlabel metal2 13632 67197 13632 67197 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit21.Q
rlabel metal2 14880 67662 14880 67662 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit22.Q
rlabel metal2 17040 66696 17040 66696 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit23.Q
rlabel metal2 16800 67914 16800 67914 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit24.Q
rlabel via2 5469 71484 5469 71484 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit25.Q
rlabel metal2 7680 70980 7680 70980 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit26.Q
rlabel metal2 5760 71442 5760 71442 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit27.Q
rlabel metal2 8256 66696 8256 66696 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit28.Q
rlabel metal2 9504 65772 9504 65772 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit29.Q
rlabel metal2 17280 50106 17280 50106 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit3.Q
rlabel metal2 9120 66654 9120 66654 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit30.Q
rlabel metal2 14688 63630 14688 63630 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit31.Q
rlabel metal3 10896 55524 10896 55524 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit4.Q
rlabel metal2 12288 55825 12288 55825 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit5.Q
rlabel metal2 3264 54012 3264 54012 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit6.Q
rlabel metal2 4896 54355 4896 54355 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit7.Q
rlabel metal2 9072 50484 9072 50484 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit8.Q
rlabel metal2 7296 50148 7296 50148 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit9.Q
rlabel metal2 7008 47922 7008 47922 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit0.Q
rlabel metal3 5712 47964 5712 47964 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit1.Q
rlabel metal2 18048 48510 18048 48510 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit10.Q
rlabel metal2 19680 48468 19680 48468 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit11.Q
rlabel metal2 10368 52794 10368 52794 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit12.Q
rlabel metal2 11904 53179 11904 53179 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit13.Q
rlabel metal3 3888 54348 3888 54348 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit14.Q
rlabel via1 3312 53335 3312 53335 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit15.Q
rlabel metal2 5376 51660 5376 51660 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit16.Q
rlabel metal2 6912 51289 6912 51289 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit17.Q
rlabel metal2 15744 52080 15744 52080 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit18.Q
rlabel metal3 17472 51240 17472 51240 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit19.Q
rlabel metal2 15360 49518 15360 49518 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit2.Q
rlabel metal3 17040 54852 17040 54852 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit20.Q
rlabel metal2 19344 54264 19344 54264 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit21.Q
rlabel metal2 4800 58128 4800 58128 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit22.Q
rlabel metal2 3264 56613 3264 56613 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit23.Q
rlabel metal2 7920 55524 7920 55524 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit24.Q
rlabel metal2 9456 55020 9456 55020 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit25.Q
rlabel metal2 14976 54852 14976 54852 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit26.Q
rlabel metal2 16560 54847 16560 54847 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit27.Q
rlabel metal2 13824 57372 13824 57372 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit28.Q
rlabel metal2 15360 57211 15360 57211 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit29.Q
rlabel metal2 17040 48972 17040 48972 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit3.Q
rlabel metal2 8400 57876 8400 57876 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit30.Q
rlabel metal2 9984 58125 9984 58125 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit31.Q
rlabel metal3 10272 50988 10272 50988 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit4.Q
rlabel metal2 12000 51289 12000 51289 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit5.Q
rlabel metal2 4128 51954 4128 51954 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit6.Q
rlabel metal2 2160 52164 2160 52164 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit7.Q
rlabel metal3 8880 47964 8880 47964 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit8.Q
rlabel metal2 8016 47460 8016 47460 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit9.Q
rlabel metal2 2688 41286 2688 41286 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit0.Q
rlabel metal2 2496 41708 2496 41708 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit1.Q
rlabel metal2 17952 45066 17952 45066 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit10.Q
rlabel metal2 19584 44688 19584 44688 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit11.Q
rlabel metal2 9456 45192 9456 45192 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit12.Q
rlabel metal2 11040 45479 11040 45479 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit13.Q
rlabel metal2 2304 47922 2304 47922 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit14.Q
rlabel metal2 3840 47541 3840 47541 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit15.Q
rlabel metal3 3456 42840 3456 42840 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit16.Q
rlabel metal2 2688 43729 2688 43729 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit17.Q
rlabel metal2 15072 47544 15072 47544 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit18.Q
rlabel metal2 16704 46956 16704 46956 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit19.Q
rlabel metal2 15168 45822 15168 45822 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit2.Q
rlabel metal2 11712 43722 11712 43722 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit20.Q
rlabel via1 13296 43432 13296 43432 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit21.Q
rlabel metal2 4080 49476 4080 49476 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit22.Q
rlabel metal2 2496 49777 2496 49777 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit23.Q
rlabel metal2 6432 50568 6432 50568 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit24.Q
rlabel metal2 4896 50183 4896 50183 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit25.Q
rlabel metal2 18336 51870 18336 51870 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit26.Q
rlabel metal2 19872 52455 19872 52455 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit27.Q
rlabel metal2 11616 49560 11616 49560 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit28.Q
rlabel metal2 13152 49777 13152 49777 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit29.Q
rlabel metal2 16704 45479 16704 45479 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit3.Q
rlabel metal2 5184 55860 5184 55860 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit30.Q
rlabel metal2 6720 56161 6720 56161 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit31.Q
rlabel metal2 11424 43974 11424 43974 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit4.Q
rlabel metal2 13824 43218 13824 43218 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit5.Q
rlabel metal2 4128 45276 4128 45276 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit6.Q
rlabel metal2 2496 45276 2496 45276 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit7.Q
rlabel metal2 5616 44940 5616 44940 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit8.Q
rlabel metal2 7200 45241 7200 45241 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit9.Q
rlabel metal2 9120 60060 9120 60060 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit0.Q
rlabel metal2 10896 59556 10896 59556 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit1.Q
rlabel metal2 18720 69426 18720 69426 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit10.Q
rlabel metal2 18912 69258 18912 69258 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit11.Q
rlabel metal2 19296 70938 19296 70938 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit12.Q
rlabel metal2 8544 73038 8544 73038 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit13.Q
rlabel metal2 10848 74214 10848 74214 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit14.Q
rlabel metal3 9888 73500 9888 73500 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit15.Q
rlabel metal2 9600 43176 9600 43176 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit16.Q
rlabel metal2 7968 43386 7968 43386 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit17.Q
rlabel metal2 14184 46536 14184 46536 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit18.Q
rlabel metal2 12576 46746 12576 46746 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit19.Q
rlabel metal3 2784 65940 2784 65940 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit2.Q
rlabel metal2 17280 43967 17280 43967 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit20.Q
rlabel metal2 15744 44352 15744 44352 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit21.Q
rlabel via1 10416 48799 10416 48799 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit22.Q
rlabel metal2 8832 49056 8832 49056 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit23.Q
rlabel metal2 5568 44184 5568 44184 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit24.Q
rlabel metal2 7104 45273 7104 45273 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit25.Q
rlabel metal3 18192 47040 18192 47040 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit26.Q
rlabel metal2 19824 46788 19824 46788 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit27.Q
rlabel metal2 9888 46368 9888 46368 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit28.Q
rlabel metal2 11592 46452 11592 46452 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit29.Q
rlabel metal2 4896 64428 4896 64428 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit3.Q
rlabel metal3 3360 55356 3360 55356 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit30.Q
rlabel via1 2352 54847 2352 54847 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit31.Q
rlabel metal2 10272 63231 10272 63231 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit4.Q
rlabel metal2 10464 63378 10464 63378 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit5.Q
rlabel metal3 7968 64302 7968 64302 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit6.Q
rlabel metal2 13920 61278 13920 61278 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit7.Q
rlabel metal2 14400 61320 14400 61320 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit8.Q
rlabel metal2 16032 58590 16032 58590 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit9.Q
rlabel metal2 3744 66234 3744 66234 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit0.Q
rlabel metal2 5184 64932 5184 64932 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit1.Q
rlabel metal2 7008 79170 7008 79170 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit10.Q
rlabel metal2 5184 77616 5184 77616 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit11.Q
rlabel metal2 7296 61950 7296 61950 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit12.Q
rlabel metal2 5664 61866 5664 61866 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit13.Q
rlabel metal2 12288 60270 12288 60270 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit14.Q
rlabel metal3 14112 59556 14112 59556 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit15.Q
rlabel metal2 16224 65478 16224 65478 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit16.Q
rlabel metal2 17712 64848 17712 64848 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit17.Q
rlabel metal2 4752 73668 4752 73668 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit18.Q
rlabel metal2 6336 74641 6336 74641 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit19.Q
rlabel metal2 4128 66192 4128 66192 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit2.Q
rlabel metal3 1872 65436 1872 65436 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit20.Q
rlabel metal2 3168 65517 3168 65517 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit21.Q
rlabel metal3 2304 68208 2304 68208 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit22.Q
rlabel via1 3984 67624 3984 67624 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit23.Q
rlabel metal2 9600 67578 9600 67578 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit24.Q
rlabel metal2 11712 67158 11712 67158 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit25.Q
rlabel metal2 2016 72618 2016 72618 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit26.Q
rlabel metal2 3552 72625 3552 72625 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit27.Q
rlabel metal2 4320 64015 4320 64015 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit28.Q
rlabel metal4 2688 66990 2688 66990 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit29.Q
rlabel metal2 12768 65352 12768 65352 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit3.Q
rlabel metal2 2640 64428 2640 64428 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit30.Q
rlabel via1 4176 59383 4176 59383 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit31.Q
rlabel metal2 12576 65310 12576 65310 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit4.Q
rlabel metal2 12864 64514 12864 64514 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit5.Q
rlabel metal2 14496 70224 14496 70224 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit6.Q
rlabel metal2 15552 71526 15552 71526 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit7.Q
rlabel metal2 16032 69258 16032 69258 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit8.Q
rlabel metal2 8064 79170 8064 79170 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit9.Q
rlabel metal2 12000 62328 12000 62328 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit10.Q
rlabel metal2 13584 61824 13584 61824 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit11.Q
rlabel metal2 15744 72114 15744 72114 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit12.Q
rlabel metal2 17376 71904 17376 71904 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit13.Q
rlabel metal2 4320 76608 4320 76608 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit14.Q
rlabel metal2 5856 75775 5856 75775 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit15.Q
rlabel metal2 1536 78582 1536 78582 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit16.Q
rlabel metal2 3072 78159 3072 78159 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit17.Q
rlabel metal2 1824 69132 1824 69132 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit18.Q
rlabel metal2 3456 70945 3456 70945 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit19.Q
rlabel metal2 8496 68460 8496 68460 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit20.Q
rlabel metal2 10176 68709 10176 68709 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit21.Q
rlabel metal2 1824 74256 1824 74256 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit22.Q
rlabel metal2 3360 75061 3360 75061 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit23.Q
rlabel metal2 2304 64218 2304 64218 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit24.Q
rlabel metal3 3984 68208 3984 68208 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit25.Q
rlabel via1 2496 70651 2496 70651 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit26.Q
rlabel metal2 4032 70693 4032 70693 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit27.Q
rlabel metal2 9216 60942 9216 60942 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit28.Q
rlabel via1 10800 60895 10800 60895 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit29.Q
rlabel metal3 2364 61572 2364 61572 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit30.Q
rlabel metal3 3600 61824 3600 61824 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit31.Q
rlabel metal2 7008 64173 7008 64173 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit8.Q
rlabel metal2 5472 64008 5472 64008 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit9.Q
rlabel metal2 3072 52500 3072 52500 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG0
rlabel metal3 11664 50988 11664 50988 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG1
rlabel metal2 16800 51954 16800 51954 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG2
rlabel metal2 3360 54894 3360 54894 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG3
rlabel metal2 3840 53214 3840 53214 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG4
rlabel metal2 11424 52542 11424 52542 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG5
rlabel metal2 13056 52416 13056 52416 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG6
rlabel metal2 5376 50568 5376 50568 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG7
rlabel metal3 16992 49560 16992 49560 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG10
rlabel metal2 6432 49098 6432 49098 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG11
rlabel metal2 6240 65184 6240 65184 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG12
rlabel metal3 12960 49560 12960 49560 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG13
rlabel metal3 18768 54264 18768 54264 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG14
rlabel metal3 7296 50232 7296 50232 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG15
rlabel metal2 4320 53172 4320 53172 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG4
rlabel metal2 14352 52416 14352 52416 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG5
rlabel metal3 16944 53256 16944 53256 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG6
rlabel metal2 8064 51408 8064 51408 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG7
rlabel metal2 3936 53970 3936 53970 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG8
rlabel metal2 14592 53676 14592 53676 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG9
rlabel metal3 7392 64092 7392 64092 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1BEG0
rlabel metal3 1728 83538 1728 83538 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1BEG1
rlabel metal2 17472 72576 17472 72576 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1BEG2
rlabel metal3 5904 83496 5904 83496 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1BEG3
rlabel metal2 8112 35952 8112 35952 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END0
rlabel metal2 15504 30660 15504 30660 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END1
rlabel metal3 18144 31248 18144 31248 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END2
rlabel metal3 9024 48804 9024 48804 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END3
rlabel metal2 2160 83496 2160 83496 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG0
rlabel metal3 3456 69384 3456 69384 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG1
rlabel metal2 3648 84252 3648 84252 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG2
rlabel metal3 2112 82236 2112 82236 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG3
rlabel metal2 3840 82362 3840 82362 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG4
rlabel metal2 4224 74088 4224 74088 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG5
rlabel metal3 10560 83160 10560 83160 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG6
rlabel metal3 3120 83328 3120 83328 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG7
rlabel metal3 2928 83496 2928 83496 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb0
rlabel metal4 15168 46326 15168 46326 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb1
rlabel metal2 4992 83412 4992 83412 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb2
rlabel metal2 4128 83496 4128 83496 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb3
rlabel metal3 4752 42756 4752 42756 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb4
rlabel metal3 10848 83496 10848 83496 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb5
rlabel metal3 11616 83496 11616 83496 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb6
rlabel metal2 5424 83496 5424 83496 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb7
rlabel metal3 7104 82824 7104 82824 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N4BEG0
rlabel metal2 12384 66528 12384 66528 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N4BEG1
rlabel metal2 9072 83496 9072 83496 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N4BEG2
rlabel metal2 7200 82698 7200 82698 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N4BEG3
rlabel metal2 13248 35784 13248 35784 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG0
rlabel metal4 1104 63336 1104 63336 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG1
rlabel metal3 11856 31332 11856 31332 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG2
rlabel metal4 11520 18606 11520 18606 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG3
rlabel metal3 528 39312 528 39312 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG4
rlabel metal4 16608 21000 16608 21000 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG5
rlabel metal4 16896 21168 16896 21168 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG6
rlabel metal4 2496 51114 2496 51114 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG7
rlabel metal2 13248 2184 13248 2184 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S4BEG0
rlabel metal3 15600 1848 15600 1848 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S4BEG1
rlabel metal3 15984 1176 15984 1176 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S4BEG2
rlabel metal3 14016 1848 14016 1848 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S4BEG3
rlabel metal2 9216 43974 9216 43974 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W1BEG0
rlabel metal2 14112 44898 14112 44898 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W1BEG1
rlabel metal2 17664 43932 17664 43932 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W1BEG2
rlabel metal2 10560 47754 10560 47754 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W1BEG3
rlabel metal2 7296 44730 7296 44730 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG0
rlabel metal3 19344 45696 19344 45696 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG1
rlabel metal2 11616 45990 11616 45990 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG2
rlabel metal3 1776 52668 1776 52668 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG3
rlabel metal2 2112 41916 2112 41916 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG4
rlabel metal2 17040 45024 17040 45024 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG5
rlabel metal2 13536 44520 13536 44520 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG6
rlabel metal3 2064 45696 2064 45696 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG7
rlabel metal2 2112 45486 2112 45486 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb0
rlabel metal2 19392 45612 19392 45612 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb1
rlabel metal2 10848 46914 10848 46914 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb2
rlabel metal2 4032 47292 4032 47292 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb3
rlabel metal3 2256 44184 2256 44184 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb4
rlabel metal3 16608 47460 16608 47460 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb5
rlabel metal2 13152 44478 13152 44478 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb6
rlabel metal2 1728 49476 1728 49476 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb7
rlabel metal2 10080 55655 10080 55655 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG0
rlabel metal2 16800 55188 16800 55188 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG1
rlabel metal2 11520 57624 11520 57624 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG10
rlabel metal3 2112 59346 2112 59346 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG11
rlabel metal3 15312 56280 15312 56280 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG2
rlabel metal3 9936 57120 9936 57120 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG3
rlabel metal2 6720 47754 6720 47754 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG4
rlabel metal3 19536 50484 19536 50484 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG5
rlabel metal2 12528 55440 12528 55440 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG6
rlabel metal2 2016 56112 2016 56112 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG7
rlabel metal3 6192 51072 6192 51072 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG8
rlabel metal3 17136 53508 17136 53508 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG9
rlabel metal2 2112 51156 2112 51156 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG0
rlabel metal3 19824 51996 19824 51996 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG1
rlabel metal2 12144 54096 12144 54096 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG10
rlabel metal3 2268 54768 2268 54768 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG11
rlabel metal2 6816 51702 6816 51702 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG12
rlabel metal2 17472 52038 17472 52038 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG13
rlabel metal2 19488 54852 19488 54852 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG14
rlabel metal2 3216 55608 3216 55608 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG15
rlabel metal2 13440 50022 13440 50022 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG2
rlabel metal2 2112 54012 2112 54012 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG3
rlabel metal3 4176 48720 4176 48720 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG4
rlabel metal3 16560 50232 16560 50232 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG5
rlabel metal2 12576 51030 12576 51030 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG6
rlabel metal2 2400 51828 2400 51828 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG7
rlabel metal2 2400 49224 2400 49224 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG8
rlabel metal3 19488 48972 19488 48972 0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG9
rlabel metal2 14640 82740 14640 82740 0 Tile_X0Y0_E_TT_IF2_top.N4BEG_outbuf_10.A
rlabel metal3 7248 83244 7248 83244 0 Tile_X0Y0_E_TT_IF2_top.N4BEG_outbuf_11.A
rlabel metal4 480 46998 480 46998 0 Tile_X0Y0_E_TT_IF2_top.N4BEG_outbuf_8.A
rlabel metal5 7928 83496 7928 83496 0 Tile_X0Y0_E_TT_IF2_top.N4BEG_outbuf_9.A
rlabel metal3 19344 37296 19344 37296 0 Tile_X0Y0_FrameData[0]
rlabel metal2 15552 54222 15552 54222 0 Tile_X0Y0_FrameData[10]
rlabel metal2 18288 47964 18288 47964 0 Tile_X0Y0_FrameData[11]
rlabel metal2 14016 71778 14016 71778 0 Tile_X0Y0_FrameData[12]
rlabel metal3 1056 72744 1056 72744 0 Tile_X0Y0_FrameData[13]
rlabel metal2 1440 54054 1440 54054 0 Tile_X0Y0_FrameData[14]
rlabel metal4 1536 51870 1536 51870 0 Tile_X0Y0_FrameData[15]
rlabel metal2 14496 65268 14496 65268 0 Tile_X0Y0_FrameData[16]
rlabel metal2 19968 48594 19968 48594 0 Tile_X0Y0_FrameData[17]
rlabel metal2 14592 52962 14592 52962 0 Tile_X0Y0_FrameData[18]
rlabel metal2 12768 53676 12768 53676 0 Tile_X0Y0_FrameData[19]
rlabel metal2 19152 37464 19152 37464 0 Tile_X0Y0_FrameData[1]
rlabel metal2 1248 71022 1248 71022 0 Tile_X0Y0_FrameData[20]
rlabel metal3 2190 82404 2190 82404 0 Tile_X0Y0_FrameData[21]
rlabel metal2 1248 51912 1248 51912 0 Tile_X0Y0_FrameData[22]
rlabel metal2 2208 57162 2208 57162 0 Tile_X0Y0_FrameData[23]
rlabel metal3 3582 83412 3582 83412 0 Tile_X0Y0_FrameData[24]
rlabel metal3 1728 68460 1728 68460 0 Tile_X0Y0_FrameData[25]
rlabel metal3 702 84084 702 84084 0 Tile_X0Y0_FrameData[26]
rlabel metal3 1086 84420 1086 84420 0 Tile_X0Y0_FrameData[27]
rlabel via3 78 84756 78 84756 0 Tile_X0Y0_FrameData[28]
rlabel metal2 1296 69972 1296 69972 0 Tile_X0Y0_FrameData[29]
rlabel metal2 1248 66486 1248 66486 0 Tile_X0Y0_FrameData[2]
rlabel metal2 1392 58548 1392 58548 0 Tile_X0Y0_FrameData[30]
rlabel metal3 1344 66948 1344 66948 0 Tile_X0Y0_FrameData[31]
rlabel metal3 13248 49476 13248 49476 0 Tile_X0Y0_FrameData[3]
rlabel metal3 16896 64344 16896 64344 0 Tile_X0Y0_FrameData[4]
rlabel metal2 12384 42000 12384 42000 0 Tile_X0Y0_FrameData[5]
rlabel metal2 1248 53970 1248 53970 0 Tile_X0Y0_FrameData[6]
rlabel metal3 13200 71484 13200 71484 0 Tile_X0Y0_FrameData[7]
rlabel metal2 13728 68964 13728 68964 0 Tile_X0Y0_FrameData[8]
rlabel metal2 1248 82026 1248 82026 0 Tile_X0Y0_FrameData[9]
rlabel metal2 19296 36330 19296 36330 0 Tile_X0Y0_FrameData_O[0]
rlabel metal2 18048 43092 18048 43092 0 Tile_X0Y0_FrameData_O[10]
rlabel metal2 19968 43806 19968 43806 0 Tile_X0Y0_FrameData_O[11]
rlabel metal2 19968 44520 19968 44520 0 Tile_X0Y0_FrameData_O[12]
rlabel metal2 19776 45234 19776 45234 0 Tile_X0Y0_FrameData_O[13]
rlabel metal3 21426 45612 21426 45612 0 Tile_X0Y0_FrameData_O[14]
rlabel metal3 20754 46284 20754 46284 0 Tile_X0Y0_FrameData_O[15]
rlabel metal2 19968 47376 19968 47376 0 Tile_X0Y0_FrameData_O[16]
rlabel metal3 21378 47628 21378 47628 0 Tile_X0Y0_FrameData_O[17]
rlabel metal2 19872 48804 19872 48804 0 Tile_X0Y0_FrameData_O[18]
rlabel metal2 19968 49140 19968 49140 0 Tile_X0Y0_FrameData_O[19]
rlabel metal2 19200 37044 19200 37044 0 Tile_X0Y0_FrameData_O[1]
rlabel metal2 19680 49854 19680 49854 0 Tile_X0Y0_FrameData_O[20]
rlabel metal2 20064 50232 20064 50232 0 Tile_X0Y0_FrameData_O[21]
rlabel metal3 20802 50988 20802 50988 0 Tile_X0Y0_FrameData_O[22]
rlabel metal2 19968 51996 19968 51996 0 Tile_X0Y0_FrameData_O[23]
rlabel metal2 19680 53088 19680 53088 0 Tile_X0Y0_FrameData_O[24]
rlabel metal3 21378 53004 21378 53004 0 Tile_X0Y0_FrameData_O[25]
rlabel metal3 21426 53676 21426 53676 0 Tile_X0Y0_FrameData_O[26]
rlabel metal2 19872 54474 19872 54474 0 Tile_X0Y0_FrameData_O[27]
rlabel metal3 20850 55020 20850 55020 0 Tile_X0Y0_FrameData_O[28]
rlabel metal3 20514 55692 20514 55692 0 Tile_X0Y0_FrameData_O[29]
rlabel metal2 18768 37968 18768 37968 0 Tile_X0Y0_FrameData_O[2]
rlabel metal3 21426 56364 21426 56364 0 Tile_X0Y0_FrameData_O[30]
rlabel metal2 19584 56784 19584 56784 0 Tile_X0Y0_FrameData_O[31]
rlabel metal2 19584 38472 19584 38472 0 Tile_X0Y0_FrameData_O[3]
rlabel metal2 19296 39186 19296 39186 0 Tile_X0Y0_FrameData_O[4]
rlabel metal3 20994 39564 20994 39564 0 Tile_X0Y0_FrameData_O[5]
rlabel metal3 20658 40236 20658 40236 0 Tile_X0Y0_FrameData_O[6]
rlabel metal3 20802 40908 20802 40908 0 Tile_X0Y0_FrameData_O[7]
rlabel metal3 21234 41580 21234 41580 0 Tile_X0Y0_FrameData_O[8]
rlabel metal2 19680 42756 19680 42756 0 Tile_X0Y0_FrameData_O[9]
rlabel metal2 15840 83718 15840 83718 0 Tile_X0Y0_FrameStrobe_O[0]
rlabel metal2 18096 83328 18096 83328 0 Tile_X0Y0_FrameStrobe_O[10]
rlabel metal2 18480 83328 18480 83328 0 Tile_X0Y0_FrameStrobe_O[11]
rlabel metal2 18240 83622 18240 83622 0 Tile_X0Y0_FrameStrobe_O[12]
rlabel metal3 18624 83748 18624 83748 0 Tile_X0Y0_FrameStrobe_O[13]
rlabel metal2 18624 83622 18624 83622 0 Tile_X0Y0_FrameStrobe_O[14]
rlabel metal3 19056 83328 19056 83328 0 Tile_X0Y0_FrameStrobe_O[15]
rlabel metal2 19152 82992 19152 82992 0 Tile_X0Y0_FrameStrobe_O[16]
rlabel metal2 19680 84378 19680 84378 0 Tile_X0Y0_FrameStrobe_O[17]
rlabel metal2 19488 82908 19488 82908 0 Tile_X0Y0_FrameStrobe_O[18]
rlabel metal2 20016 83748 20016 83748 0 Tile_X0Y0_FrameStrobe_O[19]
rlabel metal2 16032 82962 16032 82962 0 Tile_X0Y0_FrameStrobe_O[1]
rlabel metal2 16224 79392 16224 79392 0 Tile_X0Y0_FrameStrobe_O[2]
rlabel metal2 16416 85188 16416 85188 0 Tile_X0Y0_FrameStrobe_O[3]
rlabel metal2 16608 85188 16608 85188 0 Tile_X0Y0_FrameStrobe_O[4]
rlabel metal2 16800 84852 16800 84852 0 Tile_X0Y0_FrameStrobe_O[5]
rlabel metal2 17040 83496 17040 83496 0 Tile_X0Y0_FrameStrobe_O[6]
rlabel metal2 17232 83664 17232 83664 0 Tile_X0Y0_FrameStrobe_O[7]
rlabel metal2 17376 84852 17376 84852 0 Tile_X0Y0_FrameStrobe_O[8]
rlabel metal2 17760 84084 17760 84084 0 Tile_X0Y0_FrameStrobe_O[9]
rlabel metal2 1824 84978 1824 84978 0 Tile_X0Y0_N1BEG[0]
rlabel metal2 1968 83748 1968 83748 0 Tile_X0Y0_N1BEG[1]
rlabel via2 2208 85944 2208 85944 0 Tile_X0Y0_N1BEG[2]
rlabel metal2 5568 83790 5568 83790 0 Tile_X0Y0_N1BEG[3]
rlabel metal2 2304 84084 2304 84084 0 Tile_X0Y0_N2BEG[0]
rlabel metal2 2928 84420 2928 84420 0 Tile_X0Y0_N2BEG[1]
rlabel metal2 3456 84504 3456 84504 0 Tile_X0Y0_N2BEG[2]
rlabel metal2 2688 84504 2688 84504 0 Tile_X0Y0_N2BEG[3]
rlabel metal2 3600 82992 3600 82992 0 Tile_X0Y0_N2BEG[4]
rlabel metal2 3504 83748 3504 83748 0 Tile_X0Y0_N2BEG[5]
rlabel metal2 3744 85902 3744 85902 0 Tile_X0Y0_N2BEG[6]
rlabel metal2 3984 83748 3984 83748 0 Tile_X0Y0_N2BEG[7]
rlabel metal3 3696 83748 3696 83748 0 Tile_X0Y0_N2BEGb[0]
rlabel metal2 4320 85860 4320 85860 0 Tile_X0Y0_N2BEGb[1]
rlabel metal2 4800 83286 4800 83286 0 Tile_X0Y0_N2BEGb[2]
rlabel metal2 4224 84294 4224 84294 0 Tile_X0Y0_N2BEGb[3]
rlabel metal2 4608 84042 4608 84042 0 Tile_X0Y0_N2BEGb[4]
rlabel metal2 5088 85020 5088 85020 0 Tile_X0Y0_N2BEGb[5]
rlabel metal2 5280 85188 5280 85188 0 Tile_X0Y0_N2BEGb[6]
rlabel metal2 5424 83748 5424 83748 0 Tile_X0Y0_N2BEGb[7]
rlabel metal2 5664 85272 5664 85272 0 Tile_X0Y0_N4BEG[0]
rlabel metal2 7968 83286 7968 83286 0 Tile_X0Y0_N4BEG[10]
rlabel metal3 7392 83748 7392 83748 0 Tile_X0Y0_N4BEG[11]
rlabel metal2 7488 83076 7488 83076 0 Tile_X0Y0_N4BEG[12]
rlabel metal3 8304 83748 8304 83748 0 Tile_X0Y0_N4BEG[13]
rlabel metal2 8832 84042 8832 84042 0 Tile_X0Y0_N4BEG[14]
rlabel metal3 7968 83412 7968 83412 0 Tile_X0Y0_N4BEG[15]
rlabel metal4 1008 59220 1008 59220 0 Tile_X0Y0_N4BEG[1]
rlabel metal2 6048 85230 6048 85230 0 Tile_X0Y0_N4BEG[2]
rlabel metal4 2352 7812 2352 7812 0 Tile_X0Y0_N4BEG[3]
rlabel metal2 6432 85188 6432 85188 0 Tile_X0Y0_N4BEG[4]
rlabel metal2 6624 85230 6624 85230 0 Tile_X0Y0_N4BEG[5]
rlabel metal2 6816 85188 6816 85188 0 Tile_X0Y0_N4BEG[6]
rlabel metal2 7008 85188 7008 85188 0 Tile_X0Y0_N4BEG[7]
rlabel metal2 6240 83790 6240 83790 0 Tile_X0Y0_N4BEG[8]
rlabel metal2 7584 83790 7584 83790 0 Tile_X0Y0_N4BEG[9]
rlabel metal2 8736 85440 8736 85440 0 Tile_X0Y0_S1END[0]
rlabel metal2 8928 84852 8928 84852 0 Tile_X0Y0_S1END[1]
rlabel metal2 9120 85440 9120 85440 0 Tile_X0Y0_S1END[2]
rlabel metal3 9120 82236 9120 82236 0 Tile_X0Y0_S1END[3]
rlabel metal3 7488 78456 7488 78456 0 Tile_X0Y0_S2END[0]
rlabel metal2 11232 83928 11232 83928 0 Tile_X0Y0_S2END[1]
rlabel metal3 12192 76776 12192 76776 0 Tile_X0Y0_S2END[2]
rlabel metal2 11616 84222 11616 84222 0 Tile_X0Y0_S2END[3]
rlabel metal2 11808 85188 11808 85188 0 Tile_X0Y0_S2END[4]
rlabel metal2 12000 83928 12000 83928 0 Tile_X0Y0_S2END[5]
rlabel metal2 12768 69972 12768 69972 0 Tile_X0Y0_S2END[6]
rlabel metal2 12384 84516 12384 84516 0 Tile_X0Y0_S2END[7]
rlabel metal2 9504 84012 9504 84012 0 Tile_X0Y0_S2MID[0]
rlabel metal2 9696 85188 9696 85188 0 Tile_X0Y0_S2MID[1]
rlabel metal2 9888 85230 9888 85230 0 Tile_X0Y0_S2MID[2]
rlabel metal2 10080 85902 10080 85902 0 Tile_X0Y0_S2MID[3]
rlabel metal2 10272 85188 10272 85188 0 Tile_X0Y0_S2MID[4]
rlabel metal2 10464 85188 10464 85188 0 Tile_X0Y0_S2MID[5]
rlabel metal2 10656 85608 10656 85608 0 Tile_X0Y0_S2MID[6]
rlabel metal3 6624 41244 6624 41244 0 Tile_X0Y0_S2MID[7]
rlabel metal2 12336 64428 12336 64428 0 Tile_X0Y0_S4END[0]
rlabel metal2 14496 85356 14496 85356 0 Tile_X0Y0_S4END[10]
rlabel metal2 14688 84726 14688 84726 0 Tile_X0Y0_S4END[11]
rlabel metal2 14880 84726 14880 84726 0 Tile_X0Y0_S4END[12]
rlabel metal2 15072 85146 15072 85146 0 Tile_X0Y0_S4END[13]
rlabel metal2 15264 84726 15264 84726 0 Tile_X0Y0_S4END[14]
rlabel metal2 15456 85188 15456 85188 0 Tile_X0Y0_S4END[15]
rlabel metal2 14304 49896 14304 49896 0 Tile_X0Y0_S4END[1]
rlabel metal2 12960 85188 12960 85188 0 Tile_X0Y0_S4END[2]
rlabel metal2 13104 83496 13104 83496 0 Tile_X0Y0_S4END[3]
rlabel metal2 13344 85188 13344 85188 0 Tile_X0Y0_S4END[4]
rlabel metal2 13536 85776 13536 85776 0 Tile_X0Y0_S4END[5]
rlabel metal2 13728 85230 13728 85230 0 Tile_X0Y0_S4END[6]
rlabel metal2 13920 85188 13920 85188 0 Tile_X0Y0_S4END[7]
rlabel metal2 14112 85944 14112 85944 0 Tile_X0Y0_S4END[8]
rlabel metal2 14304 84726 14304 84726 0 Tile_X0Y0_S4END[9]
rlabel metal2 15696 83748 15696 83748 0 Tile_X0Y0_UserCLKo
rlabel metal3 1290 43092 1290 43092 0 Tile_X0Y0_W1BEG[0]
rlabel metal2 13920 43344 13920 43344 0 Tile_X0Y0_W1BEG[1]
rlabel metal2 17472 43722 17472 43722 0 Tile_X0Y0_W1BEG[2]
rlabel metal3 3552 44268 3552 44268 0 Tile_X0Y0_W1BEG[3]
rlabel metal3 990 44436 990 44436 0 Tile_X0Y0_W2BEG[0]
rlabel metal4 16416 45024 16416 45024 0 Tile_X0Y0_W2BEG[1]
rlabel metal2 11424 45318 11424 45318 0 Tile_X0Y0_W2BEG[2]
rlabel metal2 1536 45318 1536 45318 0 Tile_X0Y0_W2BEG[3]
rlabel metal2 1776 42168 1776 42168 0 Tile_X0Y0_W2BEG[4]
rlabel metal3 1290 46116 1290 46116 0 Tile_X0Y0_W2BEG[5]
rlabel metal2 13728 45780 13728 45780 0 Tile_X0Y0_W2BEG[6]
rlabel metal3 798 46788 798 46788 0 Tile_X0Y0_W2BEG[7]
rlabel metal3 990 47124 990 47124 0 Tile_X0Y0_W2BEGb[0]
rlabel metal3 15264 47418 15264 47418 0 Tile_X0Y0_W2BEGb[1]
rlabel metal3 1290 47796 1290 47796 0 Tile_X0Y0_W2BEGb[2]
rlabel metal2 1776 47460 1776 47460 0 Tile_X0Y0_W2BEGb[3]
rlabel metal2 1488 46956 1488 46956 0 Tile_X0Y0_W2BEGb[4]
rlabel metal2 16224 48552 16224 48552 0 Tile_X0Y0_W2BEGb[5]
rlabel metal3 318 49140 318 49140 0 Tile_X0Y0_W2BEGb[6]
rlabel metal3 798 49476 798 49476 0 Tile_X0Y0_W2BEGb[7]
rlabel metal3 1290 55188 1290 55188 0 Tile_X0Y0_W6BEG[0]
rlabel metal2 11328 58128 11328 58128 0 Tile_X0Y0_W6BEG[10]
rlabel metal3 990 58884 990 58884 0 Tile_X0Y0_W6BEG[11]
rlabel metal2 15840 56196 15840 56196 0 Tile_X0Y0_W6BEG[1]
rlabel metal2 14880 55986 14880 55986 0 Tile_X0Y0_W6BEG[2]
rlabel metal2 9504 56532 9504 56532 0 Tile_X0Y0_W6BEG[3]
rlabel metal3 846 56532 846 56532 0 Tile_X0Y0_W6BEG[4]
rlabel metal3 414 56868 414 56868 0 Tile_X0Y0_W6BEG[5]
rlabel metal2 12384 56868 12384 56868 0 Tile_X0Y0_W6BEG[6]
rlabel metal2 1824 57414 1824 57414 0 Tile_X0Y0_W6BEG[7]
rlabel metal2 2880 51786 2880 51786 0 Tile_X0Y0_W6BEG[8]
rlabel metal2 17184 54138 17184 54138 0 Tile_X0Y0_W6BEG[9]
rlabel metal3 990 49812 990 49812 0 Tile_X0Y0_WW4BEG[0]
rlabel metal2 12000 53508 12000 53508 0 Tile_X0Y0_WW4BEG[10]
rlabel metal3 942 53508 942 53508 0 Tile_X0Y0_WW4BEG[11]
rlabel metal2 1776 52752 1776 52752 0 Tile_X0Y0_WW4BEG[12]
rlabel metal3 16848 53088 16848 53088 0 Tile_X0Y0_WW4BEG[13]
rlabel metal3 1290 54516 1290 54516 0 Tile_X0Y0_WW4BEG[14]
rlabel metal2 3072 55104 3072 55104 0 Tile_X0Y0_WW4BEG[15]
rlabel metal3 15360 50232 15360 50232 0 Tile_X0Y0_WW4BEG[1]
rlabel metal2 13248 50316 13248 50316 0 Tile_X0Y0_WW4BEG[2]
rlabel metal3 798 50820 798 50820 0 Tile_X0Y0_WW4BEG[3]
rlabel metal2 2832 48972 2832 48972 0 Tile_X0Y0_WW4BEG[4]
rlabel metal4 6624 50778 6624 50778 0 Tile_X0Y0_WW4BEG[5]
rlabel metal2 12384 51576 12384 51576 0 Tile_X0Y0_WW4BEG[6]
rlabel metal3 750 52164 750 52164 0 Tile_X0Y0_WW4BEG[7]
rlabel metal3 942 52500 942 52500 0 Tile_X0Y0_WW4BEG[8]
rlabel metal3 18288 49728 18288 49728 0 Tile_X0Y0_WW4BEG[9]
rlabel metal2 2784 17472 2784 17472 0 Tile_X0Y1_E1END[0]
rlabel metal2 13632 18396 13632 18396 0 Tile_X0Y1_E1END[1]
rlabel metal2 17664 30030 17664 30030 0 Tile_X0Y1_E1END[2]
rlabel metal2 8736 18690 8736 18690 0 Tile_X0Y1_E1END[3]
rlabel metal2 9120 19362 9120 19362 0 Tile_X0Y1_E2END[0]
rlabel metal3 414 20580 414 20580 0 Tile_X0Y1_E2END[1]
rlabel metal2 10704 35196 10704 35196 0 Tile_X0Y1_E2END[2]
rlabel metal4 2112 28686 2112 28686 0 Tile_X0Y1_E2END[3]
rlabel metal3 174 21588 174 21588 0 Tile_X0Y1_E2END[4]
rlabel metal2 13152 34188 13152 34188 0 Tile_X0Y1_E2END[5]
rlabel metal3 1230 22260 1230 22260 0 Tile_X0Y1_E2END[6]
rlabel metal2 1968 20832 1968 20832 0 Tile_X0Y1_E2END[7]
rlabel metal2 2496 37170 2496 37170 0 Tile_X0Y1_E2MID[0]
rlabel metal2 10080 18186 10080 18186 0 Tile_X0Y1_E2MID[1]
rlabel metal2 9984 17640 9984 17640 0 Tile_X0Y1_E2MID[2]
rlabel metal3 270 18564 270 18564 0 Tile_X0Y1_E2MID[3]
rlabel metal3 126 18900 126 18900 0 Tile_X0Y1_E2MID[4]
rlabel metal2 11952 29064 11952 29064 0 Tile_X0Y1_E2MID[5]
rlabel metal2 11808 33768 11808 33768 0 Tile_X0Y1_E2MID[6]
rlabel metal2 1584 26796 1584 26796 0 Tile_X0Y1_E2MID[7]
rlabel metal3 894 28308 894 28308 0 Tile_X0Y1_E6END[0]
rlabel metal2 14208 31206 14208 31206 0 Tile_X0Y1_E6END[10]
rlabel metal2 6048 34860 6048 34860 0 Tile_X0Y1_E6END[11]
rlabel metal3 990 28644 990 28644 0 Tile_X0Y1_E6END[1]
rlabel metal3 270 28980 270 28980 0 Tile_X0Y1_E6END[2]
rlabel metal2 6768 37716 6768 37716 0 Tile_X0Y1_E6END[3]
rlabel metal2 5088 31458 5088 31458 0 Tile_X0Y1_E6END[4]
rlabel metal2 14112 21966 14112 21966 0 Tile_X0Y1_E6END[5]
rlabel metal3 17424 29904 17424 29904 0 Tile_X0Y1_E6END[6]
rlabel metal2 1776 28476 1776 28476 0 Tile_X0Y1_E6END[7]
rlabel metal2 2112 21126 2112 21126 0 Tile_X0Y1_E6END[8]
rlabel metal3 654 31332 654 31332 0 Tile_X0Y1_E6END[9]
rlabel metal2 2112 22344 2112 22344 0 Tile_X0Y1_EE4END[0]
rlabel metal4 4704 26166 4704 26166 0 Tile_X0Y1_EE4END[10]
rlabel metal3 414 26628 414 26628 0 Tile_X0Y1_EE4END[11]
rlabel metal3 1278 26964 1278 26964 0 Tile_X0Y1_EE4END[12]
rlabel metal2 16416 23562 16416 23562 0 Tile_X0Y1_EE4END[13]
rlabel metal2 18144 29400 18144 29400 0 Tile_X0Y1_EE4END[14]
rlabel metal3 78 27972 78 27972 0 Tile_X0Y1_EE4END[15]
rlabel metal2 12864 23184 12864 23184 0 Tile_X0Y1_EE4END[1]
rlabel metal2 14304 29778 14304 29778 0 Tile_X0Y1_EE4END[2]
rlabel metal3 480 24066 480 24066 0 Tile_X0Y1_EE4END[3]
rlabel metal2 3360 24780 3360 24780 0 Tile_X0Y1_EE4END[4]
rlabel metal2 16512 24150 16512 24150 0 Tile_X0Y1_EE4END[5]
rlabel metal4 12480 25956 12480 25956 0 Tile_X0Y1_EE4END[6]
rlabel metal2 9120 25914 9120 25914 0 Tile_X0Y1_EE4END[7]
rlabel metal2 2496 23226 2496 23226 0 Tile_X0Y1_EE4END[8]
rlabel metal3 14064 23772 14064 23772 0 Tile_X0Y1_EE4END[9]
rlabel metal2 6240 26754 6240 26754 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit0.Q
rlabel metal2 7776 26756 7776 26756 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit1.Q
rlabel metal3 9504 2352 9504 2352 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit10.Q
rlabel metal2 10320 1932 10320 1932 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit11.Q
rlabel metal2 12480 32592 12480 32592 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit12.Q
rlabel metal2 13296 31332 13296 31332 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit13.Q
rlabel metal2 4128 35238 4128 35238 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit14.Q
rlabel metal2 4320 35448 4320 35448 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit15.Q
rlabel metal2 3456 39438 3456 39438 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit16.Q
rlabel metal2 5568 39981 5568 39981 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit17.Q
rlabel metal2 9408 41076 9408 41076 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit18.Q
rlabel metal2 10944 40663 10944 40663 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit19.Q
rlabel metal2 15216 5124 15216 5124 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit2.Q
rlabel metal2 10464 41286 10464 41286 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit20.Q
rlabel via1 12048 41239 12048 41239 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit21.Q
rlabel metal2 5376 41286 5376 41286 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit22.Q
rlabel metal2 7392 41076 7392 41076 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit23.Q
rlabel metal2 2112 30576 2112 30576 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit24.Q
rlabel metal3 2364 30660 2364 30660 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit25.Q
rlabel metal2 15168 17640 15168 17640 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit26.Q
rlabel metal3 15360 17976 15360 17976 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit27.Q
rlabel metal2 17472 28476 17472 28476 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit28.Q
rlabel metal2 16992 29190 16992 29190 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit29.Q
rlabel metal2 16896 4410 16896 4410 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit3.Q
rlabel metal2 7584 39900 7584 39900 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit30.Q
rlabel metal2 6720 39438 6720 39438 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit31.Q
rlabel metal2 16704 16254 16704 16254 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit4.Q
rlabel metal2 18144 15708 18144 15708 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit5.Q
rlabel metal3 8736 38220 8736 38220 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit6.Q
rlabel metal2 10464 37506 10464 37506 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit7.Q
rlabel metal2 3168 28602 3168 28602 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit8.Q
rlabel metal2 5664 27678 5664 27678 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit9.Q
rlabel metal2 11424 34440 11424 34440 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit0.Q
rlabel via2 13536 35028 13536 35028 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit1.Q
rlabel metal2 14688 4074 14688 4074 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit10.Q
rlabel metal2 16320 3486 16320 3486 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit11.Q
rlabel metal2 16992 17094 16992 17094 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit12.Q
rlabel metal2 18528 17343 18528 17343 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit13.Q
rlabel metal2 8400 34356 8400 34356 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit14.Q
rlabel metal3 9888 33852 9888 33852 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit15.Q
rlabel metal2 6288 24780 6288 24780 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit16.Q
rlabel metal2 7776 25585 7776 25585 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit17.Q
rlabel metal2 15648 8862 15648 8862 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit18.Q
rlabel metal2 17280 9702 17280 9702 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit19.Q
rlabel metal2 13536 35280 13536 35280 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit2.Q
rlabel metal2 17040 17976 17040 17976 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit20.Q
rlabel via1 18576 18559 18576 18559 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit21.Q
rlabel metal2 8640 38850 8640 38850 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit22.Q
rlabel metal2 10176 38983 10176 38983 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit23.Q
rlabel metal2 5856 28392 5856 28392 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit24.Q
rlabel metal2 7392 28058 7392 28058 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit25.Q
rlabel metal2 14784 7686 14784 7686 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit26.Q
rlabel metal2 16896 7266 16896 7266 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit27.Q
rlabel metal3 17232 13440 17232 13440 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit28.Q
rlabel metal3 18912 14196 18912 14196 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit29.Q
rlabel metal2 14784 33852 14784 33852 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit3.Q
rlabel metal2 8352 35826 8352 35826 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit30.Q
rlabel metal2 9984 35616 9984 35616 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit31.Q
rlabel metal2 10272 36750 10272 36750 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit4.Q
rlabel metal2 13008 38388 13008 38388 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit5.Q
rlabel metal2 12960 39438 12960 39438 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit6.Q
rlabel metal3 14640 37968 14640 37968 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit7.Q
rlabel metal2 5952 19152 5952 19152 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit8.Q
rlabel metal2 7488 19537 7488 19537 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit9.Q
rlabel metal2 8640 14826 8640 14826 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit0.Q
rlabel metal2 7008 15456 7008 15456 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit1.Q
rlabel metal2 2880 23142 2880 23142 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit10.Q
rlabel metal2 14592 24150 14592 24150 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit11.Q
rlabel via2 15072 23774 15072 23774 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit12.Q
rlabel metal3 16464 24780 16464 24780 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit13.Q
rlabel metal3 14352 25536 14352 25536 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit14.Q
rlabel metal2 15840 26754 15840 26754 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit15.Q
rlabel metal2 16704 25578 16704 25578 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit16.Q
rlabel metal2 5856 32298 5856 32298 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit17.Q
rlabel metal3 7632 32676 7632 32676 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit18.Q
rlabel metal2 8208 31584 8208 31584 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit19.Q
rlabel metal2 17472 13307 17472 13307 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit2.Q
rlabel metal2 5856 25326 5856 25326 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit20.Q
rlabel metal2 2496 25158 2496 25158 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit21.Q
rlabel metal2 3072 24780 3072 24780 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit22.Q
rlabel metal3 17856 23268 17856 23268 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit23.Q
rlabel metal2 18048 24108 18048 24108 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit24.Q
rlabel metal3 19440 23604 19440 23604 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit25.Q
rlabel metal2 19296 27006 19296 27006 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit26.Q
rlabel metal2 17376 26754 17376 26754 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit27.Q
rlabel metal2 19632 26124 19632 26124 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit28.Q
rlabel via1 10224 27631 10224 27631 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit29.Q
rlabel metal2 15648 14070 15648 14070 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit3.Q
rlabel metal2 9504 27888 9504 27888 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit30.Q
rlabel metal2 11136 29064 11136 29064 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit31.Q
rlabel metal2 15072 9912 15072 9912 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit4.Q
rlabel metal2 13344 9660 13344 9660 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit5.Q
rlabel metal3 7344 12600 7344 12600 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit6.Q
rlabel metal2 7296 12558 7296 12558 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit7.Q
rlabel metal2 2016 22974 2016 22974 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit8.Q
rlabel metal2 3552 22421 3552 22421 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit9.Q
rlabel metal2 8352 11508 8352 11508 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit0.Q
rlabel metal3 10032 11172 10032 11172 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit1.Q
rlabel metal2 15168 12894 15168 12894 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit10.Q
rlabel metal2 13344 13482 13344 13482 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit11.Q
rlabel metal2 12912 7392 12912 7392 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit12.Q
rlabel metal2 14592 7644 14592 7644 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit13.Q
rlabel metal2 5616 11424 5616 11424 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit14.Q
rlabel metal2 3936 11634 3936 11634 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit15.Q
rlabel metal2 6048 18522 6048 18522 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit16.Q
rlabel metal3 7344 17976 7344 17976 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit17.Q
rlabel metal3 16224 11172 16224 11172 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit18.Q
rlabel metal2 17472 11636 17472 11636 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit19.Q
rlabel metal2 18048 12264 18048 12264 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit2.Q
rlabel metal2 12384 15582 12384 15582 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit20.Q
rlabel metal2 13920 15789 13920 15789 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit21.Q
rlabel metal2 6912 29190 6912 29190 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit22.Q
rlabel via1 8496 29143 8496 29143 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit23.Q
rlabel metal2 7440 16275 7440 16275 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit24.Q
rlabel metal2 5856 16263 5856 16263 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit25.Q
rlabel metal2 15072 15001 15072 15001 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit26.Q
rlabel metal2 13536 14574 13536 14574 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit27.Q
rlabel metal2 12720 11928 12720 11928 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit28.Q
rlabel metal2 11232 12306 11232 12306 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit29.Q
rlabel metal3 19104 10416 19104 10416 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit3.Q
rlabel metal2 5664 14450 5664 14450 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit30.Q
rlabel metal2 4080 14196 4080 14196 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit31.Q
rlabel metal2 12480 10248 12480 10248 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit4.Q
rlabel metal3 10608 9660 10608 9660 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit5.Q
rlabel metal2 7776 10290 7776 10290 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit6.Q
rlabel metal2 6096 10416 6096 10416 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit7.Q
rlabel metal2 9312 13314 9312 13314 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit8.Q
rlabel metal2 11232 13692 11232 13692 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit9.Q
rlabel metal2 2976 6384 2976 6384 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit0.Q
rlabel metal2 2688 6174 2688 6174 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit1.Q
rlabel metal2 12576 4998 12576 4998 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit10.Q
rlabel metal2 12096 5628 12096 5628 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit11.Q
rlabel metal2 6240 6132 6240 6132 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit12.Q
rlabel metal2 7488 5040 7488 5040 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit13.Q
rlabel metal3 4176 6468 4176 6468 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit14.Q
rlabel metal2 4224 6174 4224 6174 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit15.Q
rlabel metal2 3552 17934 3552 17934 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit16.Q
rlabel metal3 4992 17136 4992 17136 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit17.Q
rlabel via1 19056 8656 19056 8656 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit18.Q
rlabel metal3 17232 8148 17232 8148 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit19.Q
rlabel metal3 5328 2100 5328 2100 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit2.Q
rlabel metal2 12768 6090 12768 6090 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit20.Q
rlabel metal2 14400 6174 14400 6174 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit21.Q
rlabel metal3 6336 8148 6336 8148 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit22.Q
rlabel metal2 7488 8610 7488 8610 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit23.Q
rlabel metal2 9408 14952 9408 14952 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit24.Q
rlabel metal2 11232 15582 11232 15582 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit25.Q
rlabel metal2 14760 11676 14760 11676 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit26.Q
rlabel metal2 13152 11424 13152 11424 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit27.Q
rlabel metal2 10752 8148 10752 8148 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit28.Q
rlabel metal2 12480 8400 12480 8400 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit29.Q
rlabel metal2 4896 2100 4896 2100 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit3.Q
rlabel metal2 6096 12684 6096 12684 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit30.Q
rlabel metal2 4608 13146 4608 13146 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit31.Q
rlabel metal2 10368 9030 10368 9030 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit4.Q
rlabel metal3 9216 8820 9216 8820 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit5.Q
rlabel metal2 3840 10290 3840 10290 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit6.Q
rlabel metal2 3552 10248 3552 10248 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit7.Q
rlabel metal3 4656 9492 4656 9492 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit8.Q
rlabel metal2 4704 8232 4704 8232 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit9.Q
rlabel metal2 18048 20706 18048 20706 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit0.Q
rlabel metal2 17040 19908 17040 19908 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit1.Q
rlabel metal2 14400 3143 14400 3143 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit10.Q
rlabel metal2 12864 3486 12864 3486 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit11.Q
rlabel metal2 18720 5929 18720 5929 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit12.Q
rlabel metal2 16992 5166 16992 5166 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit13.Q
rlabel metal2 8064 5929 8064 5929 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit14.Q
rlabel metal2 6528 5670 6528 5670 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit15.Q
rlabel metal3 2028 17724 2028 17724 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit16.Q
rlabel metal2 1632 17430 1632 17430 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit17.Q
rlabel metal2 5664 1428 5664 1428 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit18.Q
rlabel metal2 4992 1848 4992 1848 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit19.Q
rlabel via2 18432 30240 18432 30240 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit2.Q
rlabel metal2 10080 4536 10080 4536 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit20.Q
rlabel metal2 9888 5334 9888 5334 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit21.Q
rlabel metal2 2832 8652 2832 8652 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit22.Q
rlabel metal2 3072 8526 3072 8526 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit23.Q
rlabel metal2 3216 15288 3216 15288 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit24.Q
rlabel metal2 3552 15498 3552 15498 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit25.Q
rlabel metal2 11232 6762 11232 6762 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit26.Q
rlabel metal2 10855 7226 10855 7226 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit27.Q
rlabel metal2 7680 1764 7680 1764 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit28.Q
rlabel metal2 7776 3192 7776 3192 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit29.Q
rlabel metal2 20064 30156 20064 30156 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit3.Q
rlabel metal2 2688 13734 2688 13734 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit30.Q
rlabel metal3 2544 12684 2544 12684 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit31.Q
rlabel metal3 19824 30240 19824 30240 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit4.Q
rlabel metal3 9840 30660 9840 30660 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit5.Q
rlabel metal2 10848 31080 10848 31080 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit6.Q
rlabel metal2 9120 31626 9120 31626 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit7.Q
rlabel metal2 8784 7392 8784 7392 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit8.Q
rlabel metal2 7104 7392 7104 7392 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit9.Q
rlabel metal3 15504 32172 15504 32172 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit0.Q
rlabel metal2 5280 34524 5280 34524 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit1.Q
rlabel via1 6048 37379 6048 37379 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit10.Q
rlabel metal2 7296 36582 7296 36582 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit11.Q
rlabel metal3 2112 20748 2112 20748 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit12.Q
rlabel metal3 2928 19488 2928 19488 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit13.Q
rlabel metal2 9312 21630 9312 21630 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit14.Q
rlabel metal2 11040 21287 11040 21287 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit15.Q
rlabel metal2 11808 27090 11808 27090 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit16.Q
rlabel metal2 13440 26544 13440 26544 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit17.Q
rlabel metal2 2640 30072 2640 30072 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit18.Q
rlabel metal2 4080 32340 4080 32340 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit19.Q
rlabel metal3 6576 33768 6576 33768 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit2.Q
rlabel metal2 8928 20496 8928 20496 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit20.Q
rlabel metal2 7296 20664 7296 20664 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit21.Q
rlabel metal2 10944 17091 10944 17091 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit22.Q
rlabel metal2 9408 17094 9408 17094 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit23.Q
rlabel metal3 12768 17976 12768 17976 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit24.Q
rlabel metal2 10992 18564 10992 18564 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit25.Q
rlabel metal2 10320 17976 10320 17976 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit26.Q
rlabel metal2 8688 17976 8688 17976 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit27.Q
rlabel metal2 6720 24192 6720 24192 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit28.Q
rlabel metal2 7296 23821 7296 23821 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit29.Q
rlabel metal3 7056 34356 7056 34356 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit3.Q
rlabel metal2 8736 23142 8736 23142 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit30.Q
rlabel metal2 15744 21000 15744 21000 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit31.Q
rlabel metal2 3840 29568 3840 29568 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit4.Q
rlabel metal3 5040 30072 5040 30072 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit5.Q
rlabel metal3 13872 19236 13872 19236 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit6.Q
rlabel metal2 15216 18732 15216 18732 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit7.Q
rlabel metal2 14496 28056 14496 28056 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit8.Q
rlabel metal2 16032 28609 16032 28609 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit9.Q
rlabel metal2 6048 30704 6048 30704 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit0.Q
rlabel metal3 4176 30828 4176 30828 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit1.Q
rlabel via1 9312 24602 9312 24602 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit10.Q
rlabel metal2 10896 24024 10896 24024 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit11.Q
rlabel metal2 11904 29410 11904 29410 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit12.Q
rlabel metal2 13536 28770 13536 28770 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit13.Q
rlabel metal4 2208 32928 2208 32928 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit14.Q
rlabel metal2 3168 33894 3168 33894 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit15.Q
rlabel metal2 2016 39396 2016 39396 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit16.Q
rlabel metal2 3120 38388 3120 38388 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit17.Q
rlabel metal2 9504 25914 9504 25914 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit18.Q
rlabel metal2 11232 25825 11232 25825 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit19.Q
rlabel via1 15120 21583 15120 21583 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit2.Q
rlabel metal2 10848 20118 10848 20118 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit20.Q
rlabel metal2 12672 19824 12672 19824 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit21.Q
rlabel metal2 2400 36792 2400 36792 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit22.Q
rlabel metal2 4272 36876 4272 36876 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit23.Q
rlabel metal3 5040 20076 5040 20076 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit24.Q
rlabel metal2 5088 20790 5088 20790 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit25.Q
rlabel metal2 6528 21714 6528 21714 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit26.Q
rlabel metal2 11904 22673 11904 22673 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit27.Q
rlabel metal2 13440 23436 13440 23436 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit28.Q
rlabel metal3 11376 23772 11376 23772 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit29.Q
rlabel metal2 13632 21000 13632 21000 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit3.Q
rlabel metal3 14736 31500 14736 31500 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit30.Q
rlabel metal3 14208 30072 14208 30072 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit31.Q
rlabel metal2 17664 32011 17664 32011 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit4.Q
rlabel metal2 16128 31626 16128 31626 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit5.Q
rlabel metal2 7008 38259 7008 38259 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit6.Q
rlabel metal2 5472 38472 5472 38472 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit7.Q
rlabel metal2 1296 24024 1296 24024 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit8.Q
rlabel metal2 2784 24948 2784 24948 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit9.Q
rlabel metal2 7104 8736 7104 8736 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG12
rlabel metal2 13440 15246 13440 15246 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG13
rlabel metal3 18000 11508 18000 11508 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG14
rlabel metal3 8352 18564 8352 18564 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG15
rlabel metal3 6864 1848 6864 1848 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S1BEG0
rlabel metal2 15264 13482 15264 13482 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S1BEG1
rlabel metal3 16128 27720 16128 27720 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S1BEG2
rlabel metal3 8544 1848 8544 1848 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S1BEG3
rlabel metal3 3216 17808 3216 17808 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG0
rlabel metal2 9360 1176 9360 1176 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG1
rlabel metal3 13248 26628 13248 26628 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG2
rlabel metal3 8928 1176 8928 1176 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG3
rlabel metal2 8640 2184 8640 2184 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG4
rlabel metal3 10512 1176 10512 1176 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG5
rlabel metal2 11856 1848 11856 1848 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG6
rlabel metal2 9552 2184 9552 2184 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG7
rlabel metal5 13344 6972 13344 6972 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S4BEG0
rlabel metal2 15984 1176 15984 1176 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S4BEG1
rlabel metal3 18480 1848 18480 1848 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S4BEG2
rlabel metal2 14688 2142 14688 2142 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S4BEG3
rlabel metal2 2112 1008 2112 1008 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W1BEG0
rlabel metal2 2928 1848 2928 1848 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W1BEG1
rlabel metal3 2496 3990 2496 3990 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W1BEG2
rlabel metal3 1632 2604 1632 2604 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W1BEG3
rlabel metal4 2496 9114 2496 9114 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG0
rlabel metal2 1776 1848 1776 1848 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG1
rlabel metal2 2112 2016 2112 2016 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG2
rlabel metal2 2592 2856 2592 2856 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG3
rlabel metal3 3360 4620 3360 4620 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG4
rlabel metal2 2016 3528 2016 3528 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG5
rlabel metal2 1632 2982 1632 2982 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG6
rlabel metal4 2880 7812 2880 7812 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG7
rlabel metal2 2400 4788 2400 4788 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb0
rlabel metal2 1728 3276 1728 3276 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb1
rlabel metal2 2208 4956 2208 4956 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb2
rlabel metal2 3264 5544 3264 5544 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb3
rlabel metal2 2112 5250 2112 5250 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb4
rlabel metal2 11520 5418 11520 5418 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb5
rlabel metal2 1728 4410 1728 4410 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb6
rlabel metal3 3840 7224 3840 7224 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb7
rlabel metal2 7728 11760 7728 11760 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG0
rlabel metal2 17856 12222 17856 12222 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG1
rlabel metal2 14688 10164 14688 10164 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG10
rlabel metal2 1632 14994 1632 14994 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG11
rlabel metal2 1920 14616 1920 14616 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG2
rlabel metal2 2112 29148 2112 29148 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG3
rlabel metal2 1632 15540 1632 15540 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG4
rlabel metal2 15264 14994 15264 14994 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG5
rlabel metal2 12960 12180 12960 12180 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG6
rlabel metal2 3072 16079 3072 16079 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG7
rlabel metal3 8304 14784 8304 14784 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG8
rlabel metal2 1536 14112 1536 14112 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG9
rlabel metal2 1968 8232 1968 8232 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG0
rlabel metal3 19008 7896 19008 7896 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG1
rlabel metal2 2496 9912 2496 9912 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG10
rlabel metal2 8160 11004 8160 11004 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG11
rlabel metal2 10800 11760 10800 11760 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG12
rlabel metal2 1632 12390 1632 12390 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG13
rlabel metal2 14592 8274 14592 8274 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG14
rlabel metal2 1920 11214 1920 11214 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG15
rlabel metal2 1632 6888 1632 6888 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG2
rlabel metal3 4608 7896 4608 7896 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG3
rlabel metal3 4032 8778 4032 8778 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG4
rlabel metal2 2112 8232 2112 8232 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG5
rlabel metal2 1440 8400 1440 8400 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG6
rlabel metal2 1872 9408 1872 9408 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG7
rlabel metal2 1589 10920 1589 10920 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG8
rlabel metal2 17664 10248 17664 10248 0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG9
rlabel metal2 1392 7728 1392 7728 0 Tile_X0Y1_FrameData[0]
rlabel metal3 702 35700 702 35700 0 Tile_X0Y1_FrameData[10]
rlabel metal2 11904 14616 11904 14616 0 Tile_X0Y1_FrameData[11]
rlabel metal2 1488 21252 1488 21252 0 Tile_X0Y1_FrameData[12]
rlabel metal3 1584 19740 1584 19740 0 Tile_X0Y1_FrameData[13]
rlabel metal3 750 37044 750 37044 0 Tile_X0Y1_FrameData[14]
rlabel metal2 1728 7812 1728 7812 0 Tile_X0Y1_FrameData[15]
rlabel metal2 1296 17052 1296 17052 0 Tile_X0Y1_FrameData[16]
rlabel metal2 1632 38136 1632 38136 0 Tile_X0Y1_FrameData[17]
rlabel metal2 1296 29820 1296 29820 0 Tile_X0Y1_FrameData[18]
rlabel metal2 2496 32004 2496 32004 0 Tile_X0Y1_FrameData[19]
rlabel metal2 1632 4956 1632 4956 0 Tile_X0Y1_FrameData[1]
rlabel metal3 78 39060 78 39060 0 Tile_X0Y1_FrameData[20]
rlabel metal2 1296 22260 1296 22260 0 Tile_X0Y1_FrameData[21]
rlabel metal2 1632 7938 1632 7938 0 Tile_X0Y1_FrameData[22]
rlabel metal3 1536 8022 1536 8022 0 Tile_X0Y1_FrameData[23]
rlabel metal2 1248 28266 1248 28266 0 Tile_X0Y1_FrameData[24]
rlabel metal2 1248 27678 1248 27678 0 Tile_X0Y1_FrameData[25]
rlabel metal2 14304 15414 14304 15414 0 Tile_X0Y1_FrameData[26]
rlabel metal3 12576 17724 12576 17724 0 Tile_X0Y1_FrameData[27]
rlabel metal3 18384 30492 18384 30492 0 Tile_X0Y1_FrameData[28]
rlabel metal2 17712 13944 17712 13944 0 Tile_X0Y1_FrameData[29]
rlabel metal2 16176 12516 16176 12516 0 Tile_X0Y1_FrameData[2]
rlabel metal3 13536 31374 13536 31374 0 Tile_X0Y1_FrameData[30]
rlabel metal2 1296 12516 1296 12516 0 Tile_X0Y1_FrameData[31]
rlabel metal2 13920 14616 13920 14616 0 Tile_X0Y1_FrameData[3]
rlabel metal2 2208 31962 2208 31962 0 Tile_X0Y1_FrameData[4]
rlabel metal2 15360 32256 15360 32256 0 Tile_X0Y1_FrameData[5]
rlabel metal2 2112 10458 2112 10458 0 Tile_X0Y1_FrameData[6]
rlabel metal2 1872 10080 1872 10080 0 Tile_X0Y1_FrameData[7]
rlabel metal3 1872 26124 1872 26124 0 Tile_X0Y1_FrameData[8]
rlabel metal3 702 35364 702 35364 0 Tile_X0Y1_FrameData[9]
rlabel metal3 18432 34608 18432 34608 0 Tile_X0Y1_FrameData_O[0]
rlabel metal3 21330 64428 21330 64428 0 Tile_X0Y1_FrameData_O[10]
rlabel metal2 15312 49308 15312 49308 0 Tile_X0Y1_FrameData_O[11]
rlabel metal3 20994 65772 20994 65772 0 Tile_X0Y1_FrameData_O[12]
rlabel metal3 18048 37632 18048 37632 0 Tile_X0Y1_FrameData_O[13]
rlabel metal2 19584 37506 19584 37506 0 Tile_X0Y1_FrameData_O[14]
rlabel metal3 20802 67788 20802 67788 0 Tile_X0Y1_FrameData_O[15]
rlabel metal3 21042 68460 21042 68460 0 Tile_X0Y1_FrameData_O[16]
rlabel metal3 20802 69132 20802 69132 0 Tile_X0Y1_FrameData_O[17]
rlabel metal2 19440 49056 19440 49056 0 Tile_X0Y1_FrameData_O[18]
rlabel metal3 20802 70476 20802 70476 0 Tile_X0Y1_FrameData_O[19]
rlabel metal2 19968 35658 19968 35658 0 Tile_X0Y1_FrameData_O[1]
rlabel metal2 20064 42420 20064 42420 0 Tile_X0Y1_FrameData_O[20]
rlabel metal3 21378 71820 21378 71820 0 Tile_X0Y1_FrameData_O[21]
rlabel metal3 16392 72492 16392 72492 0 Tile_X0Y1_FrameData_O[22]
rlabel metal3 21234 73164 21234 73164 0 Tile_X0Y1_FrameData_O[23]
rlabel metal5 17904 40656 17904 40656 0 Tile_X0Y1_FrameData_O[24]
rlabel metal3 21090 74508 21090 74508 0 Tile_X0Y1_FrameData_O[25]
rlabel via2 21426 75180 21426 75180 0 Tile_X0Y1_FrameData_O[26]
rlabel metal3 21186 75852 21186 75852 0 Tile_X0Y1_FrameData_O[27]
rlabel metal3 20994 76524 20994 76524 0 Tile_X0Y1_FrameData_O[28]
rlabel via3 21426 77196 21426 77196 0 Tile_X0Y1_FrameData_O[29]
rlabel metal3 21234 59052 21234 59052 0 Tile_X0Y1_FrameData_O[2]
rlabel metal3 21330 77868 21330 77868 0 Tile_X0Y1_FrameData_O[30]
rlabel metal3 21138 78540 21138 78540 0 Tile_X0Y1_FrameData_O[31]
rlabel metal3 21042 59724 21042 59724 0 Tile_X0Y1_FrameData_O[3]
rlabel metal3 21234 60396 21234 60396 0 Tile_X0Y1_FrameData_O[4]
rlabel metal3 21330 61068 21330 61068 0 Tile_X0Y1_FrameData_O[5]
rlabel metal3 21090 61740 21090 61740 0 Tile_X0Y1_FrameData_O[6]
rlabel metal3 21378 62412 21378 62412 0 Tile_X0Y1_FrameData_O[7]
rlabel metal3 21378 63084 21378 63084 0 Tile_X0Y1_FrameData_O[8]
rlabel metal3 21282 63756 21282 63756 0 Tile_X0Y1_FrameData_O[9]
rlabel metal3 15696 336 15696 336 0 Tile_X0Y1_FrameStrobe[0]
rlabel metal2 17760 450 17760 450 0 Tile_X0Y1_FrameStrobe[10]
rlabel metal2 17952 534 17952 534 0 Tile_X0Y1_FrameStrobe[11]
rlabel metal2 18144 660 18144 660 0 Tile_X0Y1_FrameStrobe[12]
rlabel metal2 18336 492 18336 492 0 Tile_X0Y1_FrameStrobe[13]
rlabel metal2 18528 660 18528 660 0 Tile_X0Y1_FrameStrobe[14]
rlabel metal2 18720 324 18720 324 0 Tile_X0Y1_FrameStrobe[15]
rlabel metal2 18912 576 18912 576 0 Tile_X0Y1_FrameStrobe[16]
rlabel metal2 19104 618 19104 618 0 Tile_X0Y1_FrameStrobe[17]
rlabel metal2 19296 660 19296 660 0 Tile_X0Y1_FrameStrobe[18]
rlabel metal2 19488 660 19488 660 0 Tile_X0Y1_FrameStrobe[19]
rlabel metal3 16176 1008 16176 1008 0 Tile_X0Y1_FrameStrobe[1]
rlabel metal2 16224 366 16224 366 0 Tile_X0Y1_FrameStrobe[2]
rlabel metal2 2448 52500 2448 52500 0 Tile_X0Y1_FrameStrobe[3]
rlabel metal2 16608 828 16608 828 0 Tile_X0Y1_FrameStrobe[4]
rlabel metal2 2496 58590 2496 58590 0 Tile_X0Y1_FrameStrobe[5]
rlabel metal2 2496 71694 2496 71694 0 Tile_X0Y1_FrameStrobe[6]
rlabel metal3 1968 23772 1968 23772 0 Tile_X0Y1_FrameStrobe[7]
rlabel metal2 17376 660 17376 660 0 Tile_X0Y1_FrameStrobe[8]
rlabel metal2 17568 660 17568 660 0 Tile_X0Y1_FrameStrobe[9]
rlabel metal2 1968 29820 1968 29820 0 Tile_X0Y1_N1END[0]
rlabel metal2 2016 912 2016 912 0 Tile_X0Y1_N1END[1]
rlabel metal2 2208 366 2208 366 0 Tile_X0Y1_N1END[2]
rlabel metal2 2400 576 2400 576 0 Tile_X0Y1_N1END[3]
rlabel metal2 1152 13902 1152 13902 0 Tile_X0Y1_N2END[0]
rlabel metal2 10176 2436 10176 2436 0 Tile_X0Y1_N2END[1]
rlabel metal2 12960 34440 12960 34440 0 Tile_X0Y1_N2END[2]
rlabel metal4 960 18270 960 18270 0 Tile_X0Y1_N2END[3]
rlabel metal4 192 20664 192 20664 0 Tile_X0Y1_N2END[4]
rlabel metal2 5088 324 5088 324 0 Tile_X0Y1_N2END[5]
rlabel metal2 5280 114 5280 114 0 Tile_X0Y1_N2END[6]
rlabel metal5 2208 10668 2208 10668 0 Tile_X0Y1_N2END[7]
rlabel metal4 2208 15372 2208 15372 0 Tile_X0Y1_N2MID[0]
rlabel metal2 2784 1038 2784 1038 0 Tile_X0Y1_N2MID[1]
rlabel metal5 12284 30660 12284 30660 0 Tile_X0Y1_N2MID[2]
rlabel metal2 1056 12348 1056 12348 0 Tile_X0Y1_N2MID[3]
rlabel metal2 960 21168 960 21168 0 Tile_X0Y1_N2MID[4]
rlabel metal2 11424 75432 11424 75432 0 Tile_X0Y1_N2MID[5]
rlabel metal2 12864 34272 12864 34272 0 Tile_X0Y1_N2MID[6]
rlabel metal2 3936 660 3936 660 0 Tile_X0Y1_N2MID[7]
rlabel metal3 6480 18564 6480 18564 0 Tile_X0Y1_N4END[0]
rlabel metal2 7584 240 7584 240 0 Tile_X0Y1_N4END[10]
rlabel metal2 7776 534 7776 534 0 Tile_X0Y1_N4END[11]
rlabel metal2 7968 492 7968 492 0 Tile_X0Y1_N4END[12]
rlabel metal2 8160 324 8160 324 0 Tile_X0Y1_N4END[13]
rlabel metal2 8352 534 8352 534 0 Tile_X0Y1_N4END[14]
rlabel metal2 8544 618 8544 618 0 Tile_X0Y1_N4END[15]
rlabel metal2 15792 10248 15792 10248 0 Tile_X0Y1_N4END[1]
rlabel metal2 12096 840 12096 840 0 Tile_X0Y1_N4END[2]
rlabel metal2 6240 576 6240 576 0 Tile_X0Y1_N4END[3]
rlabel metal2 6432 408 6432 408 0 Tile_X0Y1_N4END[4]
rlabel metal2 13728 48678 13728 48678 0 Tile_X0Y1_N4END[5]
rlabel metal2 14304 36876 14304 36876 0 Tile_X0Y1_N4END[6]
rlabel metal2 7008 408 7008 408 0 Tile_X0Y1_N4END[7]
rlabel metal2 7200 618 7200 618 0 Tile_X0Y1_N4END[8]
rlabel metal2 7392 324 7392 324 0 Tile_X0Y1_N4END[9]
rlabel metal2 8736 660 8736 660 0 Tile_X0Y1_S1BEG[0]
rlabel metal2 14976 504 14976 504 0 Tile_X0Y1_S1BEG[1]
rlabel metal2 15744 1218 15744 1218 0 Tile_X0Y1_S1BEG[2]
rlabel metal2 9312 576 9312 576 0 Tile_X0Y1_S1BEG[3]
rlabel metal2 9504 786 9504 786 0 Tile_X0Y1_S2BEG[0]
rlabel metal2 9696 492 9696 492 0 Tile_X0Y1_S2BEG[1]
rlabel metal2 12768 1596 12768 1596 0 Tile_X0Y1_S2BEG[2]
rlabel metal2 10080 492 10080 492 0 Tile_X0Y1_S2BEG[3]
rlabel metal2 10272 450 10272 450 0 Tile_X0Y1_S2BEG[4]
rlabel metal2 10464 492 10464 492 0 Tile_X0Y1_S2BEG[5]
rlabel metal2 11712 1512 11712 1512 0 Tile_X0Y1_S2BEG[6]
rlabel metal2 10848 240 10848 240 0 Tile_X0Y1_S2BEG[7]
rlabel metal2 11088 2436 11088 2436 0 Tile_X0Y1_S2BEGb[0]
rlabel metal2 11232 408 11232 408 0 Tile_X0Y1_S2BEGb[1]
rlabel metal2 11424 576 11424 576 0 Tile_X0Y1_S2BEGb[2]
rlabel metal2 11616 282 11616 282 0 Tile_X0Y1_S2BEGb[3]
rlabel metal2 11808 492 11808 492 0 Tile_X0Y1_S2BEGb[4]
rlabel metal2 12000 744 12000 744 0 Tile_X0Y1_S2BEGb[5]
rlabel metal2 12192 660 12192 660 0 Tile_X0Y1_S2BEGb[6]
rlabel metal2 12384 870 12384 870 0 Tile_X0Y1_S2BEGb[7]
rlabel metal2 12576 576 12576 576 0 Tile_X0Y1_S4BEG[0]
rlabel metal2 14496 492 14496 492 0 Tile_X0Y1_S4BEG[10]
rlabel metal2 14688 576 14688 576 0 Tile_X0Y1_S4BEG[11]
rlabel metal2 14880 450 14880 450 0 Tile_X0Y1_S4BEG[12]
rlabel metal2 15840 714 15840 714 0 Tile_X0Y1_S4BEG[13]
rlabel metal2 15264 450 15264 450 0 Tile_X0Y1_S4BEG[14]
rlabel metal2 15456 534 15456 534 0 Tile_X0Y1_S4BEG[15]
rlabel metal2 12768 660 12768 660 0 Tile_X0Y1_S4BEG[1]
rlabel metal2 12960 828 12960 828 0 Tile_X0Y1_S4BEG[2]
rlabel metal3 14400 83328 14400 83328 0 Tile_X0Y1_S4BEG[3]
rlabel metal2 13344 828 13344 828 0 Tile_X0Y1_S4BEG[4]
rlabel metal2 13536 366 13536 366 0 Tile_X0Y1_S4BEG[5]
rlabel metal2 13728 450 13728 450 0 Tile_X0Y1_S4BEG[6]
rlabel metal2 13920 660 13920 660 0 Tile_X0Y1_S4BEG[7]
rlabel metal2 14112 408 14112 408 0 Tile_X0Y1_S4BEG[8]
rlabel metal2 15456 1554 15456 1554 0 Tile_X0Y1_S4BEG[9]
rlabel metal2 15648 660 15648 660 0 Tile_X0Y1_UserCLK
rlabel metal3 990 84 990 84 0 Tile_X0Y1_W1BEG[0]
rlabel metal2 2688 1050 2688 1050 0 Tile_X0Y1_W1BEG[1]
rlabel metal3 1182 756 1182 756 0 Tile_X0Y1_W1BEG[2]
rlabel metal3 798 1092 798 1092 0 Tile_X0Y1_W1BEG[3]
rlabel metal3 1182 1428 1182 1428 0 Tile_X0Y1_W2BEG[0]
rlabel metal3 798 1764 798 1764 0 Tile_X0Y1_W2BEG[1]
rlabel metal3 990 2100 990 2100 0 Tile_X0Y1_W2BEG[2]
rlabel metal3 1230 2436 1230 2436 0 Tile_X0Y1_W2BEG[3]
rlabel metal2 3072 2982 3072 2982 0 Tile_X0Y1_W2BEG[4]
rlabel metal2 1920 2940 1920 2940 0 Tile_X0Y1_W2BEG[5]
rlabel metal2 1488 2856 1488 2856 0 Tile_X0Y1_W2BEG[6]
rlabel metal2 2688 3696 2688 3696 0 Tile_X0Y1_W2BEG[7]
rlabel metal2 2304 3864 2304 3864 0 Tile_X0Y1_W2BEGb[0]
rlabel metal2 1488 3612 1488 3612 0 Tile_X0Y1_W2BEGb[1]
rlabel metal2 1872 3612 1872 3612 0 Tile_X0Y1_W2BEGb[2]
rlabel metal2 3072 4956 3072 4956 0 Tile_X0Y1_W2BEGb[3]
rlabel metal2 1920 4914 1920 4914 0 Tile_X0Y1_W2BEGb[4]
rlabel metal2 2304 5082 2304 5082 0 Tile_X0Y1_W2BEGb[5]
rlabel metal2 1536 4578 1536 4578 0 Tile_X0Y1_W2BEGb[6]
rlabel metal3 846 6468 846 6468 0 Tile_X0Y1_W2BEGb[7]
rlabel metal2 7488 12054 7488 12054 0 Tile_X0Y1_W6BEG[0]
rlabel metal2 1440 10710 1440 10710 0 Tile_X0Y1_W6BEG[10]
rlabel metal2 1488 14952 1488 14952 0 Tile_X0Y1_W6BEG[11]
rlabel metal3 126 12516 126 12516 0 Tile_X0Y1_W6BEG[1]
rlabel metal3 894 12852 894 12852 0 Tile_X0Y1_W6BEG[2]
rlabel via2 78 13188 78 13188 0 Tile_X0Y1_W6BEG[3]
rlabel metal3 654 13524 654 13524 0 Tile_X0Y1_W6BEG[4]
rlabel metal3 1134 13860 1134 13860 0 Tile_X0Y1_W6BEG[5]
rlabel metal2 1824 13062 1824 13062 0 Tile_X0Y1_W6BEG[6]
rlabel metal2 2880 15288 2880 15288 0 Tile_X0Y1_W6BEG[7]
rlabel metal3 3870 14868 3870 14868 0 Tile_X0Y1_W6BEG[8]
rlabel metal2 1344 14700 1344 14700 0 Tile_X0Y1_W6BEG[9]
rlabel metal2 1728 6720 1728 6720 0 Tile_X0Y1_WW4BEG[0]
rlabel metal2 2304 9912 2304 9912 0 Tile_X0Y1_WW4BEG[10]
rlabel metal2 7968 10626 7968 10626 0 Tile_X0Y1_WW4BEG[11]
rlabel metal2 10560 11424 10560 11424 0 Tile_X0Y1_WW4BEG[12]
rlabel metal3 750 11172 750 11172 0 Tile_X0Y1_WW4BEG[13]
rlabel metal3 654 11508 654 11508 0 Tile_X0Y1_WW4BEG[14]
rlabel metal3 894 11844 894 11844 0 Tile_X0Y1_WW4BEG[15]
rlabel metal3 1230 7140 1230 7140 0 Tile_X0Y1_WW4BEG[1]
rlabel metal2 1344 7056 1344 7056 0 Tile_X0Y1_WW4BEG[2]
rlabel metal3 1662 7812 1662 7812 0 Tile_X0Y1_WW4BEG[3]
rlabel metal3 798 8148 798 8148 0 Tile_X0Y1_WW4BEG[4]
rlabel metal3 990 8484 990 8484 0 Tile_X0Y1_WW4BEG[5]
rlabel metal2 1248 8484 1248 8484 0 Tile_X0Y1_WW4BEG[6]
rlabel metal3 798 9156 798 9156 0 Tile_X0Y1_WW4BEG[7]
rlabel metal3 702 9492 702 9492 0 Tile_X0Y1_WW4BEG[8]
rlabel metal2 1920 9744 1920 9744 0 Tile_X0Y1_WW4BEG[9]
rlabel metal3 14370 28812 14370 28812 0 UIO_IN_TT_PROJECT0
rlabel metal3 15552 31416 15552 31416 0 UIO_IN_TT_PROJECT1
rlabel metal4 17568 64428 17568 64428 0 UIO_IN_TT_PROJECT2
rlabel metal3 7104 70728 7104 70728 0 UIO_IN_TT_PROJECT3
rlabel metal3 10272 65940 10272 65940 0 UIO_IN_TT_PROJECT4
rlabel metal4 16992 47922 16992 47922 0 UIO_IN_TT_PROJECT5
rlabel metal4 19968 49812 19968 49812 0 UIO_IN_TT_PROJECT6
rlabel metal3 15360 33600 15360 33600 0 UIO_IN_TT_PROJECT7
rlabel via2 21426 18060 21426 18060 0 UIO_OE_TT_PROJECT0
rlabel metal3 19986 18732 19986 18732 0 UIO_OE_TT_PROJECT1
rlabel metal3 15762 19404 15762 19404 0 UIO_OE_TT_PROJECT2
rlabel metal3 19746 20076 19746 20076 0 UIO_OE_TT_PROJECT3
rlabel metal3 20802 20748 20802 20748 0 UIO_OE_TT_PROJECT4
rlabel metal3 21378 21420 21378 21420 0 UIO_OE_TT_PROJECT5
rlabel metal2 12096 49686 12096 49686 0 UIO_OE_TT_PROJECT6
rlabel metal3 20802 22764 20802 22764 0 UIO_OE_TT_PROJECT7
rlabel metal3 18834 12684 18834 12684 0 UIO_OUT_TT_PROJECT0
rlabel metal3 19890 13356 19890 13356 0 UIO_OUT_TT_PROJECT1
rlabel metal3 14592 55272 14592 55272 0 UIO_OUT_TT_PROJECT2
rlabel metal3 2400 47334 2400 47334 0 UIO_OUT_TT_PROJECT3
rlabel metal3 21378 15372 21378 15372 0 UIO_OUT_TT_PROJECT4
rlabel metal3 21042 16044 21042 16044 0 UIO_OUT_TT_PROJECT5
rlabel metal3 13296 16800 13296 16800 0 UIO_OUT_TT_PROJECT6
rlabel metal3 20994 17388 20994 17388 0 UIO_OUT_TT_PROJECT7
rlabel metal3 21042 23436 21042 23436 0 UI_IN_TT_PROJECT0
rlabel metal2 17280 24360 17280 24360 0 UI_IN_TT_PROJECT1
rlabel metal2 17376 25116 17376 25116 0 UI_IN_TT_PROJECT2
rlabel metal3 21186 25452 21186 25452 0 UI_IN_TT_PROJECT3
rlabel metal4 17664 25662 17664 25662 0 UI_IN_TT_PROJECT4
rlabel metal3 21090 26796 21090 26796 0 UI_IN_TT_PROJECT5
rlabel metal2 19968 27804 19968 27804 0 UI_IN_TT_PROJECT6
rlabel metal3 16626 28140 16626 28140 0 UI_IN_TT_PROJECT7
rlabel metal2 2112 6636 2112 6636 0 UO_OUT_TT_PROJECT0
rlabel metal3 14592 13188 14592 13188 0 UO_OUT_TT_PROJECT1
rlabel via2 21426 8652 21426 8652 0 UO_OUT_TT_PROJECT2
rlabel metal3 20802 9324 20802 9324 0 UO_OUT_TT_PROJECT3
rlabel metal3 3936 16212 3936 16212 0 UO_OUT_TT_PROJECT4
rlabel metal3 13776 13272 13776 13272 0 UO_OUT_TT_PROJECT5
rlabel metal3 20994 11340 20994 11340 0 UO_OUT_TT_PROJECT6
rlabel metal2 2112 14322 2112 14322 0 UO_OUT_TT_PROJECT7
rlabel metal2 8064 15708 8064 15708 0 _0000_
rlabel metal2 13632 6678 13632 6678 0 _0001_
rlabel metal3 12192 29064 12192 29064 0 _0002_
rlabel metal2 9744 19236 9744 19236 0 _0003_
rlabel metal3 7920 59892 7920 59892 0 _0004_
rlabel metal2 8448 59724 8448 59724 0 _0005_
rlabel metal3 7536 61572 7536 61572 0 _0006_
rlabel metal4 6528 17220 6528 17220 0 _0007_
rlabel metal2 2976 31248 2976 31248 0 _0008_
rlabel metal2 2016 31080 2016 31080 0 _0009_
rlabel metal3 4320 31332 4320 31332 0 _0010_
rlabel metal2 5952 51366 5952 51366 0 _0011_
rlabel metal2 15744 69720 15744 69720 0 _0012_
rlabel metal2 17952 54894 17952 54894 0 _0013_
rlabel metal2 4224 57078 4224 57078 0 _0014_
rlabel metal2 5952 65688 5952 65688 0 _0015_
rlabel metal3 3792 66108 3792 66108 0 _0016_
rlabel metal3 4944 65436 4944 65436 0 _0017_
rlabel metal2 6720 65604 6720 65604 0 _0018_
rlabel metal2 6528 65562 6528 65562 0 _0019_
rlabel metal2 5376 65226 5376 65226 0 _0020_
rlabel metal2 5280 64806 5280 64806 0 _0021_
rlabel metal2 13152 63588 13152 63588 0 _0022_
rlabel metal3 13248 64596 13248 64596 0 _0023_
rlabel metal3 13200 65436 13200 65436 0 _0024_
rlabel metal2 13104 64848 13104 64848 0 _0025_
rlabel metal3 12960 65520 12960 65520 0 _0026_
rlabel metal2 13728 64554 13728 64554 0 _0027_
rlabel metal2 13728 65226 13728 65226 0 _0028_
rlabel metal2 16704 70140 16704 70140 0 _0029_
rlabel metal3 15888 70140 15888 70140 0 _0030_
rlabel metal3 15312 70644 15312 70644 0 _0031_
rlabel metal2 14784 69972 14784 69972 0 _0032_
rlabel metal3 15936 70686 15936 70686 0 _0033_
rlabel metal2 16224 70602 16224 70602 0 _0034_
rlabel metal2 15744 70938 15744 70938 0 _0035_
rlabel metal2 6336 76692 6336 76692 0 _0036_
rlabel metal3 7344 76020 7344 76020 0 _0037_
rlabel metal2 7632 76188 7632 76188 0 _0038_
rlabel metal2 8160 78960 8160 78960 0 _0039_
rlabel metal3 7680 79212 7680 79212 0 _0040_
rlabel metal3 6672 76188 6672 76188 0 _0041_
rlabel metal3 6576 79212 6576 79212 0 _0042_
rlabel metal2 9168 64428 9168 64428 0 _0043_
rlabel metal3 10128 62580 10128 62580 0 _0044_
rlabel metal2 10560 63336 10560 63336 0 _0045_
rlabel metal2 9888 63126 9888 63126 0 _0046_
rlabel via1 8444 63924 8444 63924 0 _0047_
rlabel metal2 9312 63042 9312 63042 0 _0048_
rlabel metal3 9552 62580 9552 62580 0 _0049_
rlabel metal2 10752 63252 10752 63252 0 _0050_
rlabel metal3 10080 63042 10080 63042 0 _0051_
rlabel metal2 15360 62328 15360 62328 0 _0052_
rlabel metal2 15360 61351 15360 61351 0 _0053_
rlabel metal2 17520 57876 17520 57876 0 _0054_
rlabel metal3 16848 57876 16848 57876 0 _0055_
rlabel metal2 15840 62076 15840 62076 0 _0056_
rlabel metal2 16512 60354 16512 60354 0 _0057_
rlabel metal2 16608 58674 16608 58674 0 _0058_
rlabel metal3 15120 61068 15120 61068 0 _0059_
rlabel metal3 15840 60942 15840 60942 0 _0060_
rlabel metal2 19968 69132 19968 69132 0 _0061_
rlabel metal2 18672 68964 18672 68964 0 _0062_
rlabel metal2 19008 69174 19008 69174 0 _0063_
rlabel metal2 19680 70434 19680 70434 0 _0064_
rlabel metal2 19872 70392 19872 70392 0 _0065_
rlabel metal3 19488 70602 19488 70602 0 _0066_
rlabel metal2 19584 70224 19584 70224 0 _0067_
rlabel metal2 20064 70014 20064 70014 0 _0068_
rlabel metal2 19920 69972 19920 69972 0 _0069_
rlabel metal2 8928 74697 8928 74697 0 _0070_
rlabel metal3 9792 73668 9792 73668 0 _0071_
rlabel metal3 10464 73668 10464 73668 0 _0072_
rlabel metal2 10560 73038 10560 73038 0 _0073_
rlabel metal2 8064 74004 8064 74004 0 _0074_
rlabel metal2 10272 74550 10272 74550 0 _0075_
rlabel metal2 10416 74508 10416 74508 0 _0076_
rlabel metal2 10272 73122 10272 73122 0 _0077_
rlabel metal2 10800 72996 10800 72996 0 _0078_
rlabel metal2 4512 68208 4512 68208 0 _0079_
rlabel metal3 6768 69132 6768 69132 0 _0080_
rlabel metal2 6480 68628 6480 68628 0 _0081_
rlabel metal2 7344 69132 7344 69132 0 _0082_
rlabel metal2 13248 66066 13248 66066 0 _0083_
rlabel metal3 13776 65940 13776 65940 0 _0084_
rlabel metal2 13824 67242 13824 67242 0 _0085_
rlabel metal2 14496 66948 14496 66948 0 _0086_
rlabel metal2 16512 66780 16512 66780 0 _0087_
rlabel metal3 16944 66108 16944 66108 0 _0088_
rlabel metal2 16800 66234 16800 66234 0 _0089_
rlabel metal3 17184 66192 17184 66192 0 _0090_
rlabel metal2 5664 71904 5664 71904 0 _0091_
rlabel metal2 7008 70980 7008 70980 0 _0092_
rlabel metal2 7488 70602 7488 70602 0 _0093_
rlabel metal2 7296 70728 7296 70728 0 _0094_
rlabel metal3 8112 65268 8112 65268 0 _0095_
rlabel metal2 9408 66990 9408 66990 0 _0096_
rlabel metal2 9360 65604 9360 65604 0 _0097_
rlabel metal2 9936 66108 9936 66108 0 _0098_
rlabel metal3 9696 66276 9696 66276 0 _0099_
rlabel metal3 16176 63924 16176 63924 0 _0100_
rlabel metal3 15840 62580 15840 62580 0 _0101_
rlabel metal2 15696 64596 15696 64596 0 _0102_
rlabel metal3 16368 64092 16368 64092 0 _0103_
rlabel metal3 16656 63756 16656 63756 0 _0104_
rlabel metal3 19008 68460 19008 68460 0 _0105_
rlabel metal2 19776 67578 19776 67578 0 _0106_
rlabel metal2 20256 67578 20256 67578 0 _0107_
rlabel metal2 19776 67158 19776 67158 0 _0108_
rlabel metal2 19680 66780 19680 66780 0 _0109_
rlabel metal3 9312 72156 9312 72156 0 _0110_
rlabel metal2 9408 72240 9408 72240 0 _0111_
rlabel metal2 10080 71358 10080 71358 0 _0112_
rlabel metal2 10320 70644 10320 70644 0 _0113_
rlabel metal2 10368 71400 10368 71400 0 _0114_
rlabel metal2 3168 17892 3168 17892 0 _0115_
rlabel metal2 1440 17304 1440 17304 0 _0116_
rlabel metal3 5712 2604 5712 2604 0 _0117_
rlabel metal2 5376 1344 5376 1344 0 _0118_
rlabel metal2 10464 5376 10464 5376 0 _0119_
rlabel metal2 9792 4704 9792 4704 0 _0120_
rlabel metal2 3264 8568 3264 8568 0 _0121_
rlabel metal2 2976 8988 2976 8988 0 _0122_
rlabel metal2 3744 14742 3744 14742 0 _0123_
rlabel metal2 3456 15790 3456 15790 0 _0124_
rlabel metal2 11136 6552 11136 6552 0 _0125_
rlabel metal2 10848 6594 10848 6594 0 _0126_
rlabel metal2 8352 3696 8352 3696 0 _0127_
rlabel metal2 7440 3276 7440 3276 0 _0128_
rlabel metal2 3936 12600 3936 12600 0 _0129_
rlabel metal2 2208 13230 2208 13230 0 _0130_
rlabel metal2 2832 3948 2832 3948 0 _0131_
rlabel metal3 2364 6552 2364 6552 0 _0132_
rlabel metal2 5568 3696 5568 3696 0 _0133_
rlabel metal2 5280 3138 5280 3138 0 _0134_
rlabel metal2 10656 11130 10656 11130 0 _0135_
rlabel metal3 9120 8652 9120 8652 0 _0136_
rlabel metal3 4128 9996 4128 9996 0 _0137_
rlabel metal2 3456 9912 3456 9912 0 _0138_
rlabel metal2 5472 7266 5472 7266 0 _0139_
rlabel metal2 4560 9492 4560 9492 0 _0140_
rlabel metal2 11904 5796 11904 5796 0 _0141_
rlabel metal2 12960 5250 12960 5250 0 _0142_
rlabel metal2 7680 4998 7680 4998 0 _0143_
rlabel metal2 7152 3948 7152 3948 0 _0144_
rlabel metal2 5376 5586 5376 5586 0 _0145_
rlabel metal2 4080 6468 4080 6468 0 _0146_
rlabel metal3 10848 30744 10848 30744 0 _0147_
rlabel metal2 14016 14826 14016 14826 0 _0148_
rlabel metal2 11424 8400 11424 8400 0 _0149_
rlabel metal2 7536 28140 7536 28140 0 _0150_
rlabel metal2 7488 15750 7488 15750 0 _0151_
rlabel metal2 16128 14070 16128 14070 0 _0152_
rlabel metal2 16464 16464 16464 16464 0 _0153_
rlabel metal3 5472 14784 5472 14784 0 _0154_
rlabel metal2 7632 15456 7632 15456 0 _0155_
rlabel metal2 16224 13818 16224 13818 0 _0156_
rlabel metal3 13296 15876 13296 15876 0 _0157_
rlabel metal2 7968 13104 7968 13104 0 _0158_
rlabel metal3 4992 20748 4992 20748 0 _0159_
rlabel metal2 5376 20685 5376 20685 0 _0160_
rlabel metal2 4704 20118 4704 20118 0 _0161_
rlabel metal3 5472 19908 5472 19908 0 _0162_
rlabel metal3 6048 21588 6048 21588 0 _0163_
rlabel metal2 7200 21630 7200 21630 0 _0164_
rlabel metal2 6048 21504 6048 21504 0 _0165_
rlabel metal2 13056 23142 13056 23142 0 _0166_
rlabel metal2 12576 23688 12576 23688 0 _0167_
rlabel metal3 12336 22260 12336 22260 0 _0168_
rlabel metal2 13152 22302 13152 22302 0 _0169_
rlabel metal3 12384 23772 12384 23772 0 _0170_
rlabel metal2 11712 23520 11712 23520 0 _0171_
rlabel metal2 12384 23814 12384 23814 0 _0172_
rlabel metal3 15792 29820 15792 29820 0 _0173_
rlabel metal2 15264 31248 15264 31248 0 _0174_
rlabel metal2 15936 31458 15936 31458 0 _0175_
rlabel metal2 14880 32088 14880 32088 0 _0176_
rlabel metal2 15168 31458 15168 31458 0 _0177_
rlabel metal2 15504 30828 15504 30828 0 _0178_
rlabel metal2 15456 31416 15456 31416 0 _0179_
rlabel metal2 7584 33558 7584 33558 0 _0180_
rlabel metal2 7776 33936 7776 33936 0 _0181_
rlabel metal2 6336 33936 6336 33936 0 _0182_
rlabel metal3 6864 33852 6864 33852 0 _0183_
rlabel metal3 6960 34608 6960 34608 0 _0184_
rlabel metal2 7968 34314 7968 34314 0 _0185_
rlabel metal2 7968 34650 7968 34650 0 _0186_
rlabel metal2 8256 24864 8256 24864 0 _0187_
rlabel metal2 8448 25074 8448 25074 0 _0188_
rlabel metal2 8064 22680 8064 22680 0 _0189_
rlabel metal2 8352 23142 8352 23142 0 _0190_
rlabel metal2 9120 23730 9120 23730 0 _0191_
rlabel metal2 8928 23856 8928 23856 0 _0192_
rlabel metal3 17520 20748 17520 20748 0 _0193_
rlabel metal2 18336 20454 18336 20454 0 _0194_
rlabel metal2 18048 20097 18048 20097 0 _0195_
rlabel metal2 17664 19950 17664 19950 0 _0196_
rlabel metal2 18528 20790 18528 20790 0 _0197_
rlabel metal3 18000 19824 18000 19824 0 _0198_
rlabel metal2 20256 30366 20256 30366 0 _0199_
rlabel metal2 19488 30744 19488 30744 0 _0200_
rlabel metal2 20544 29778 20544 29778 0 _0201_
rlabel metal2 19920 29316 19920 29316 0 _0202_
rlabel metal2 19728 31332 19728 31332 0 _0203_
rlabel metal2 19296 30828 19296 30828 0 _0204_
rlabel metal2 10944 31332 10944 31332 0 _0205_
rlabel metal2 10752 31710 10752 31710 0 _0206_
rlabel metal3 10560 29148 10560 29148 0 _0207_
rlabel metal2 10752 29568 10752 29568 0 _0208_
rlabel metal3 9888 29820 9888 29820 0 _0209_
rlabel metal2 10464 29904 10464 29904 0 _0210_
rlabel metal2 6240 22218 6240 22218 0 _0211_
rlabel metal2 1728 22512 1728 22512 0 _0212_
rlabel metal2 3744 23352 3744 23352 0 _0213_
rlabel metal2 6144 23058 6144 23058 0 _0214_
rlabel metal2 16368 22932 16368 22932 0 _0215_
rlabel metal2 17184 25032 17184 25032 0 _0216_
rlabel metal2 15552 23724 15552 23724 0 _0217_
rlabel metal3 15648 23982 15648 23982 0 _0218_
rlabel metal2 15792 25536 15792 25536 0 _0219_
rlabel metal3 15648 25536 15648 25536 0 _0220_
rlabel metal2 16992 25746 16992 25746 0 _0221_
rlabel metal2 17088 25956 17088 25956 0 _0222_
rlabel metal2 6720 32172 6720 32172 0 _0223_
rlabel metal2 8064 32886 8064 32886 0 _0224_
rlabel metal2 8352 32214 8352 32214 0 _0225_
rlabel metal2 8448 32340 8448 32340 0 _0226_
rlabel metal3 4896 26124 4896 26124 0 _0227_
rlabel metal2 4992 25284 4992 25284 0 _0228_
rlabel metal2 2208 25284 2208 25284 0 _0229_
rlabel metal2 5664 25284 5664 25284 0 _0230_
rlabel metal2 5184 25326 5184 25326 0 _0231_
rlabel metal2 19872 23730 19872 23730 0 _0232_
rlabel metal3 20064 23562 20064 23562 0 _0233_
rlabel metal2 19584 23268 19584 23268 0 _0234_
rlabel metal2 18624 22596 18624 22596 0 _0235_
rlabel metal3 19248 23100 19248 23100 0 _0236_
rlabel metal2 20064 26922 20064 26922 0 _0237_
rlabel metal2 19488 27048 19488 27048 0 _0238_
rlabel metal3 19776 26628 19776 26628 0 _0239_
rlabel metal2 19488 26376 19488 26376 0 _0240_
rlabel metal2 19296 26376 19296 26376 0 _0241_
rlabel metal2 10368 28140 10368 28140 0 _0242_
rlabel metal2 11424 29148 11424 29148 0 _0243_
rlabel metal4 11616 26838 11616 26838 0 _0244_
rlabel metal2 11328 26922 11328 26922 0 _0245_
rlabel metal2 11616 27552 11616 27552 0 _0246_
rlabel metal2 11520 34314 11520 34314 0 _0247_
rlabel metal2 13824 34440 13824 34440 0 _0248_
rlabel metal2 11712 33894 11712 33894 0 _0249_
rlabel metal2 13008 33684 13008 33684 0 _0250_
rlabel metal3 13104 33852 13104 33852 0 _0251_
rlabel metal2 12384 33936 12384 33936 0 _0252_
rlabel metal2 12480 34104 12480 34104 0 _0253_
rlabel metal2 14304 35616 14304 35616 0 _0254_
rlabel metal2 13728 36078 13728 36078 0 _0255_
rlabel metal3 12576 35196 12576 35196 0 _0256_
rlabel metal2 13248 35406 13248 35406 0 _0257_
rlabel metal2 13248 33978 13248 33978 0 _0258_
rlabel metal2 13392 32844 13392 32844 0 _0259_
rlabel metal2 13536 33054 13536 33054 0 _0260_
rlabel metal3 13824 33012 13824 33012 0 _0261_
rlabel metal2 14304 34314 14304 34314 0 _0262_
rlabel metal2 14016 35994 14016 35994 0 _0263_
rlabel metal2 19776 34440 19776 34440 0 _0264_
rlabel metal2 12288 36414 12288 36414 0 _0265_
rlabel metal2 12384 37464 12384 37464 0 _0266_
rlabel metal2 12288 35280 12288 35280 0 _0267_
rlabel metal2 10560 35322 10560 35322 0 _0268_
rlabel metal2 12384 35322 12384 35322 0 _0269_
rlabel metal2 11904 36960 11904 36960 0 _0270_
rlabel metal2 12096 36708 12096 36708 0 _0271_
rlabel metal2 11088 36120 11088 36120 0 _0272_
rlabel via1 12674 36708 12674 36708 0 _0273_
rlabel metal2 10464 36330 10464 36330 0 _0274_
rlabel metal2 12480 36624 12480 36624 0 _0275_
rlabel metal2 12480 35532 12480 35532 0 _0276_
rlabel metal2 12624 35280 12624 35280 0 _0277_
rlabel metal2 13104 35700 13104 35700 0 _0278_
rlabel metal3 10848 36918 10848 36918 0 _0279_
rlabel metal2 13056 37338 13056 37338 0 _0280_
rlabel metal2 13536 36750 13536 36750 0 _0281_
rlabel metal2 13296 38220 13296 38220 0 _0282_
rlabel metal2 13776 36876 13776 36876 0 _0283_
rlabel metal2 13440 38472 13440 38472 0 _0284_
rlabel metal2 13632 38136 13632 38136 0 _0285_
rlabel metal3 13584 37044 13584 37044 0 _0286_
rlabel metal3 12480 58548 12480 58548 0 _0287_
rlabel metal3 17712 64428 17712 64428 0 _0288_
rlabel metal3 7104 73668 7104 73668 0 _0289_
rlabel metal2 8832 60018 8832 60018 0 _0290_
rlabel metal3 4224 68418 4224 68418 0 _0291_
rlabel metal3 13248 66108 13248 66108 0 _0292_
rlabel metal2 16128 66990 16128 66990 0 _0293_
rlabel metal3 6144 71484 6144 71484 0 _0294_
rlabel metal2 14112 36624 14112 36624 0 _0295_
rlabel metal3 12672 36876 12672 36876 0 _0296_
rlabel metal2 8064 38724 8064 38724 0 _0297_
rlabel metal3 16416 27636 16416 27636 0 _0298_
rlabel metal2 15840 19194 15840 19194 0 _0299_
rlabel metal2 1728 30870 1728 30870 0 _0300_
rlabel metal3 8640 22260 8640 22260 0 _0301_
rlabel metal3 17424 20076 17424 20076 0 _0302_
rlabel metal3 19008 29148 19008 29148 0 _0303_
rlabel metal2 10656 29232 10656 29232 0 _0304_
rlabel metal2 13440 33642 13440 33642 0 _0305_
rlabel metal2 13536 33558 13536 33558 0 _0306_
rlabel metal2 13584 37212 13584 37212 0 _0307_
rlabel metal3 13536 58380 13536 58380 0 _0308_
rlabel metal2 13344 59010 13344 59010 0 _0309_
rlabel metal2 13248 60060 13248 60060 0 _0310_
rlabel metal2 15264 17808 15264 17808 0 _0311_
rlabel metal2 15456 17598 15456 17598 0 _0312_
rlabel metal2 14688 17010 14688 17010 0 _0313_
rlabel metal2 14592 19068 14592 19068 0 _0314_
rlabel metal2 17904 64092 17904 64092 0 _0315_
rlabel metal2 18144 63588 18144 63588 0 _0316_
rlabel metal2 17280 65688 17280 65688 0 _0317_
rlabel metal3 17952 14700 17952 14700 0 _0318_
rlabel metal3 17280 29148 17280 29148 0 _0319_
rlabel metal2 16704 29232 16704 29232 0 _0320_
rlabel metal3 17136 29316 17136 29316 0 _0321_
rlabel metal2 6912 73878 6912 73878 0 _0322_
rlabel metal2 6528 72786 6528 72786 0 _0323_
rlabel metal2 5856 73794 5856 73794 0 _0324_
rlabel metal3 9072 34356 9072 34356 0 _0325_
rlabel metal2 6528 39648 6528 39648 0 _0326_
rlabel metal2 6432 39690 6432 39690 0 _0327_
rlabel metal2 6624 37632 6624 37632 0 _0328_
rlabel metal3 5472 27594 5472 27594 0 _0329_
rlabel metal2 5328 27636 5328 27636 0 _0330_
rlabel metal3 3600 28140 3600 28140 0 _0331_
rlabel metal2 3648 28392 3648 28392 0 _0332_
rlabel metal2 4704 27846 4704 27846 0 _0333_
rlabel via1 3362 12516 3362 12516 0 _0334_
rlabel metal2 3024 17892 3024 17892 0 _0335_
rlabel metal2 10752 2688 10752 2688 0 _0336_
rlabel metal2 10608 3444 10608 3444 0 _0337_
rlabel metal2 9840 2100 9840 2100 0 _0338_
rlabel metal3 10560 1932 10560 1932 0 _0339_
rlabel metal2 10272 2100 10272 2100 0 _0340_
rlabel metal4 13344 13104 13344 13104 0 _0341_
rlabel metal2 14592 14742 14592 14742 0 _0342_
rlabel metal2 13152 30912 13152 30912 0 _0343_
rlabel metal2 12960 30912 12960 30912 0 _0344_
rlabel metal3 13056 32088 13056 32088 0 _0345_
rlabel metal3 12624 32172 12624 32172 0 _0346_
rlabel metal2 13056 31290 13056 31290 0 _0347_
rlabel metal3 13440 18732 13440 18732 0 _0348_
rlabel metal2 12960 29400 12960 29400 0 _0349_
rlabel metal2 3312 35196 3312 35196 0 _0350_
rlabel metal2 4128 34650 4128 34650 0 _0351_
rlabel metal2 4704 36456 4704 36456 0 _0352_
rlabel metal2 4800 36624 4800 36624 0 _0353_
rlabel metal3 4320 34356 4320 34356 0 _0354_
rlabel metal3 3760 8652 3760 8652 0 _0355_
rlabel metal2 5184 14826 5184 14826 0 _0356_
rlabel metal2 17136 53256 17136 53256 0 clknet_0_Tile_X0Y1_UserCLK
rlabel metal2 16512 48342 16512 48342 0 clknet_1_0__leaf_Tile_X0Y1_UserCLK
rlabel metal3 16272 71568 16272 71568 0 clknet_1_1__leaf_Tile_X0Y1_UserCLK
<< properties >>
string FIXED_BBOX 0 0 21504 86016
<< end >>
