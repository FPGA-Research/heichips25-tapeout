magic
tech ihp-sg13g2
magscale 1 2
timestamp 1753456648
<< metal1 >>
rect 576 81668 99360 81692
rect 576 81628 3112 81668
rect 3152 81628 3194 81668
rect 3234 81628 3276 81668
rect 3316 81628 3358 81668
rect 3398 81628 3440 81668
rect 3480 81628 18232 81668
rect 18272 81628 18314 81668
rect 18354 81628 18396 81668
rect 18436 81628 18478 81668
rect 18518 81628 18560 81668
rect 18600 81628 33352 81668
rect 33392 81628 33434 81668
rect 33474 81628 33516 81668
rect 33556 81628 33598 81668
rect 33638 81628 33680 81668
rect 33720 81628 48472 81668
rect 48512 81628 48554 81668
rect 48594 81628 48636 81668
rect 48676 81628 48718 81668
rect 48758 81628 48800 81668
rect 48840 81628 63592 81668
rect 63632 81628 63674 81668
rect 63714 81628 63756 81668
rect 63796 81628 63838 81668
rect 63878 81628 63920 81668
rect 63960 81628 78712 81668
rect 78752 81628 78794 81668
rect 78834 81628 78876 81668
rect 78916 81628 78958 81668
rect 78998 81628 79040 81668
rect 79080 81628 93832 81668
rect 93872 81628 93914 81668
rect 93954 81628 93996 81668
rect 94036 81628 94078 81668
rect 94118 81628 94160 81668
rect 94200 81628 99360 81668
rect 576 81604 99360 81628
rect 576 80912 99360 80936
rect 576 80872 4352 80912
rect 4392 80872 4434 80912
rect 4474 80872 4516 80912
rect 4556 80872 4598 80912
rect 4638 80872 4680 80912
rect 4720 80872 19472 80912
rect 19512 80872 19554 80912
rect 19594 80872 19636 80912
rect 19676 80872 19718 80912
rect 19758 80872 19800 80912
rect 19840 80872 34592 80912
rect 34632 80872 34674 80912
rect 34714 80872 34756 80912
rect 34796 80872 34838 80912
rect 34878 80872 34920 80912
rect 34960 80872 49712 80912
rect 49752 80872 49794 80912
rect 49834 80872 49876 80912
rect 49916 80872 49958 80912
rect 49998 80872 50040 80912
rect 50080 80872 64832 80912
rect 64872 80872 64914 80912
rect 64954 80872 64996 80912
rect 65036 80872 65078 80912
rect 65118 80872 65160 80912
rect 65200 80872 79952 80912
rect 79992 80872 80034 80912
rect 80074 80872 80116 80912
rect 80156 80872 80198 80912
rect 80238 80872 80280 80912
rect 80320 80872 95072 80912
rect 95112 80872 95154 80912
rect 95194 80872 95236 80912
rect 95276 80872 95318 80912
rect 95358 80872 95400 80912
rect 95440 80872 99360 80912
rect 576 80848 99360 80872
rect 576 80156 99360 80180
rect 576 80116 3112 80156
rect 3152 80116 3194 80156
rect 3234 80116 3276 80156
rect 3316 80116 3358 80156
rect 3398 80116 3440 80156
rect 3480 80116 18232 80156
rect 18272 80116 18314 80156
rect 18354 80116 18396 80156
rect 18436 80116 18478 80156
rect 18518 80116 18560 80156
rect 18600 80116 33352 80156
rect 33392 80116 33434 80156
rect 33474 80116 33516 80156
rect 33556 80116 33598 80156
rect 33638 80116 33680 80156
rect 33720 80116 48472 80156
rect 48512 80116 48554 80156
rect 48594 80116 48636 80156
rect 48676 80116 48718 80156
rect 48758 80116 48800 80156
rect 48840 80116 63592 80156
rect 63632 80116 63674 80156
rect 63714 80116 63756 80156
rect 63796 80116 63838 80156
rect 63878 80116 63920 80156
rect 63960 80116 78712 80156
rect 78752 80116 78794 80156
rect 78834 80116 78876 80156
rect 78916 80116 78958 80156
rect 78998 80116 79040 80156
rect 79080 80116 93832 80156
rect 93872 80116 93914 80156
rect 93954 80116 93996 80156
rect 94036 80116 94078 80156
rect 94118 80116 94160 80156
rect 94200 80116 99360 80156
rect 576 80092 99360 80116
rect 576 79400 99360 79424
rect 576 79360 4352 79400
rect 4392 79360 4434 79400
rect 4474 79360 4516 79400
rect 4556 79360 4598 79400
rect 4638 79360 4680 79400
rect 4720 79360 19472 79400
rect 19512 79360 19554 79400
rect 19594 79360 19636 79400
rect 19676 79360 19718 79400
rect 19758 79360 19800 79400
rect 19840 79360 34592 79400
rect 34632 79360 34674 79400
rect 34714 79360 34756 79400
rect 34796 79360 34838 79400
rect 34878 79360 34920 79400
rect 34960 79360 49712 79400
rect 49752 79360 49794 79400
rect 49834 79360 49876 79400
rect 49916 79360 49958 79400
rect 49998 79360 50040 79400
rect 50080 79360 64832 79400
rect 64872 79360 64914 79400
rect 64954 79360 64996 79400
rect 65036 79360 65078 79400
rect 65118 79360 65160 79400
rect 65200 79360 79952 79400
rect 79992 79360 80034 79400
rect 80074 79360 80116 79400
rect 80156 79360 80198 79400
rect 80238 79360 80280 79400
rect 80320 79360 95072 79400
rect 95112 79360 95154 79400
rect 95194 79360 95236 79400
rect 95276 79360 95318 79400
rect 95358 79360 95400 79400
rect 95440 79360 99360 79400
rect 576 79336 99360 79360
rect 576 78644 99360 78668
rect 576 78604 3112 78644
rect 3152 78604 3194 78644
rect 3234 78604 3276 78644
rect 3316 78604 3358 78644
rect 3398 78604 3440 78644
rect 3480 78604 18232 78644
rect 18272 78604 18314 78644
rect 18354 78604 18396 78644
rect 18436 78604 18478 78644
rect 18518 78604 18560 78644
rect 18600 78604 33352 78644
rect 33392 78604 33434 78644
rect 33474 78604 33516 78644
rect 33556 78604 33598 78644
rect 33638 78604 33680 78644
rect 33720 78604 48472 78644
rect 48512 78604 48554 78644
rect 48594 78604 48636 78644
rect 48676 78604 48718 78644
rect 48758 78604 48800 78644
rect 48840 78604 63592 78644
rect 63632 78604 63674 78644
rect 63714 78604 63756 78644
rect 63796 78604 63838 78644
rect 63878 78604 63920 78644
rect 63960 78604 78712 78644
rect 78752 78604 78794 78644
rect 78834 78604 78876 78644
rect 78916 78604 78958 78644
rect 78998 78604 79040 78644
rect 79080 78604 93832 78644
rect 93872 78604 93914 78644
rect 93954 78604 93996 78644
rect 94036 78604 94078 78644
rect 94118 78604 94160 78644
rect 94200 78604 99360 78644
rect 576 78580 99360 78604
rect 576 77888 99360 77912
rect 576 77848 4352 77888
rect 4392 77848 4434 77888
rect 4474 77848 4516 77888
rect 4556 77848 4598 77888
rect 4638 77848 4680 77888
rect 4720 77848 19472 77888
rect 19512 77848 19554 77888
rect 19594 77848 19636 77888
rect 19676 77848 19718 77888
rect 19758 77848 19800 77888
rect 19840 77848 34592 77888
rect 34632 77848 34674 77888
rect 34714 77848 34756 77888
rect 34796 77848 34838 77888
rect 34878 77848 34920 77888
rect 34960 77848 49712 77888
rect 49752 77848 49794 77888
rect 49834 77848 49876 77888
rect 49916 77848 49958 77888
rect 49998 77848 50040 77888
rect 50080 77848 64832 77888
rect 64872 77848 64914 77888
rect 64954 77848 64996 77888
rect 65036 77848 65078 77888
rect 65118 77848 65160 77888
rect 65200 77848 79952 77888
rect 79992 77848 80034 77888
rect 80074 77848 80116 77888
rect 80156 77848 80198 77888
rect 80238 77848 80280 77888
rect 80320 77848 95072 77888
rect 95112 77848 95154 77888
rect 95194 77848 95236 77888
rect 95276 77848 95318 77888
rect 95358 77848 95400 77888
rect 95440 77848 99360 77888
rect 576 77824 99360 77848
rect 576 77132 99360 77156
rect 576 77092 3112 77132
rect 3152 77092 3194 77132
rect 3234 77092 3276 77132
rect 3316 77092 3358 77132
rect 3398 77092 3440 77132
rect 3480 77092 18232 77132
rect 18272 77092 18314 77132
rect 18354 77092 18396 77132
rect 18436 77092 18478 77132
rect 18518 77092 18560 77132
rect 18600 77092 33352 77132
rect 33392 77092 33434 77132
rect 33474 77092 33516 77132
rect 33556 77092 33598 77132
rect 33638 77092 33680 77132
rect 33720 77092 48472 77132
rect 48512 77092 48554 77132
rect 48594 77092 48636 77132
rect 48676 77092 48718 77132
rect 48758 77092 48800 77132
rect 48840 77092 63592 77132
rect 63632 77092 63674 77132
rect 63714 77092 63756 77132
rect 63796 77092 63838 77132
rect 63878 77092 63920 77132
rect 63960 77092 78712 77132
rect 78752 77092 78794 77132
rect 78834 77092 78876 77132
rect 78916 77092 78958 77132
rect 78998 77092 79040 77132
rect 79080 77092 93832 77132
rect 93872 77092 93914 77132
rect 93954 77092 93996 77132
rect 94036 77092 94078 77132
rect 94118 77092 94160 77132
rect 94200 77092 99360 77132
rect 576 77068 99360 77092
rect 576 76376 99360 76400
rect 576 76336 4352 76376
rect 4392 76336 4434 76376
rect 4474 76336 4516 76376
rect 4556 76336 4598 76376
rect 4638 76336 4680 76376
rect 4720 76336 19472 76376
rect 19512 76336 19554 76376
rect 19594 76336 19636 76376
rect 19676 76336 19718 76376
rect 19758 76336 19800 76376
rect 19840 76336 34592 76376
rect 34632 76336 34674 76376
rect 34714 76336 34756 76376
rect 34796 76336 34838 76376
rect 34878 76336 34920 76376
rect 34960 76336 49712 76376
rect 49752 76336 49794 76376
rect 49834 76336 49876 76376
rect 49916 76336 49958 76376
rect 49998 76336 50040 76376
rect 50080 76336 64832 76376
rect 64872 76336 64914 76376
rect 64954 76336 64996 76376
rect 65036 76336 65078 76376
rect 65118 76336 65160 76376
rect 65200 76336 79952 76376
rect 79992 76336 80034 76376
rect 80074 76336 80116 76376
rect 80156 76336 80198 76376
rect 80238 76336 80280 76376
rect 80320 76336 95072 76376
rect 95112 76336 95154 76376
rect 95194 76336 95236 76376
rect 95276 76336 95318 76376
rect 95358 76336 95400 76376
rect 95440 76336 99360 76376
rect 576 76312 99360 76336
rect 576 75620 99360 75644
rect 576 75580 3112 75620
rect 3152 75580 3194 75620
rect 3234 75580 3276 75620
rect 3316 75580 3358 75620
rect 3398 75580 3440 75620
rect 3480 75580 18232 75620
rect 18272 75580 18314 75620
rect 18354 75580 18396 75620
rect 18436 75580 18478 75620
rect 18518 75580 18560 75620
rect 18600 75580 33352 75620
rect 33392 75580 33434 75620
rect 33474 75580 33516 75620
rect 33556 75580 33598 75620
rect 33638 75580 33680 75620
rect 33720 75580 48472 75620
rect 48512 75580 48554 75620
rect 48594 75580 48636 75620
rect 48676 75580 48718 75620
rect 48758 75580 48800 75620
rect 48840 75580 63592 75620
rect 63632 75580 63674 75620
rect 63714 75580 63756 75620
rect 63796 75580 63838 75620
rect 63878 75580 63920 75620
rect 63960 75580 78712 75620
rect 78752 75580 78794 75620
rect 78834 75580 78876 75620
rect 78916 75580 78958 75620
rect 78998 75580 79040 75620
rect 79080 75580 93832 75620
rect 93872 75580 93914 75620
rect 93954 75580 93996 75620
rect 94036 75580 94078 75620
rect 94118 75580 94160 75620
rect 94200 75580 99360 75620
rect 576 75556 99360 75580
rect 643 75284 701 75285
rect 643 75244 652 75284
rect 692 75244 701 75284
rect 643 75243 701 75244
rect 843 75032 885 75041
rect 843 74992 844 75032
rect 884 74992 885 75032
rect 843 74983 885 74992
rect 576 74864 99360 74888
rect 576 74824 4352 74864
rect 4392 74824 4434 74864
rect 4474 74824 4516 74864
rect 4556 74824 4598 74864
rect 4638 74824 4680 74864
rect 4720 74824 19472 74864
rect 19512 74824 19554 74864
rect 19594 74824 19636 74864
rect 19676 74824 19718 74864
rect 19758 74824 19800 74864
rect 19840 74824 34592 74864
rect 34632 74824 34674 74864
rect 34714 74824 34756 74864
rect 34796 74824 34838 74864
rect 34878 74824 34920 74864
rect 34960 74824 49712 74864
rect 49752 74824 49794 74864
rect 49834 74824 49876 74864
rect 49916 74824 49958 74864
rect 49998 74824 50040 74864
rect 50080 74824 64832 74864
rect 64872 74824 64914 74864
rect 64954 74824 64996 74864
rect 65036 74824 65078 74864
rect 65118 74824 65160 74864
rect 65200 74824 79952 74864
rect 79992 74824 80034 74864
rect 80074 74824 80116 74864
rect 80156 74824 80198 74864
rect 80238 74824 80280 74864
rect 80320 74824 95072 74864
rect 95112 74824 95154 74864
rect 95194 74824 95236 74864
rect 95276 74824 95318 74864
rect 95358 74824 95400 74864
rect 95440 74824 99360 74864
rect 576 74800 99360 74824
rect 576 74108 99360 74132
rect 576 74068 3112 74108
rect 3152 74068 3194 74108
rect 3234 74068 3276 74108
rect 3316 74068 3358 74108
rect 3398 74068 3440 74108
rect 3480 74068 18232 74108
rect 18272 74068 18314 74108
rect 18354 74068 18396 74108
rect 18436 74068 18478 74108
rect 18518 74068 18560 74108
rect 18600 74068 33352 74108
rect 33392 74068 33434 74108
rect 33474 74068 33516 74108
rect 33556 74068 33598 74108
rect 33638 74068 33680 74108
rect 33720 74068 48472 74108
rect 48512 74068 48554 74108
rect 48594 74068 48636 74108
rect 48676 74068 48718 74108
rect 48758 74068 48800 74108
rect 48840 74068 63592 74108
rect 63632 74068 63674 74108
rect 63714 74068 63756 74108
rect 63796 74068 63838 74108
rect 63878 74068 63920 74108
rect 63960 74068 78712 74108
rect 78752 74068 78794 74108
rect 78834 74068 78876 74108
rect 78916 74068 78958 74108
rect 78998 74068 79040 74108
rect 79080 74068 93832 74108
rect 93872 74068 93914 74108
rect 93954 74068 93996 74108
rect 94036 74068 94078 74108
rect 94118 74068 94160 74108
rect 94200 74068 99360 74108
rect 576 74044 99360 74068
rect 576 73352 99360 73376
rect 576 73312 4352 73352
rect 4392 73312 4434 73352
rect 4474 73312 4516 73352
rect 4556 73312 4598 73352
rect 4638 73312 4680 73352
rect 4720 73312 19472 73352
rect 19512 73312 19554 73352
rect 19594 73312 19636 73352
rect 19676 73312 19718 73352
rect 19758 73312 19800 73352
rect 19840 73312 34592 73352
rect 34632 73312 34674 73352
rect 34714 73312 34756 73352
rect 34796 73312 34838 73352
rect 34878 73312 34920 73352
rect 34960 73312 49712 73352
rect 49752 73312 49794 73352
rect 49834 73312 49876 73352
rect 49916 73312 49958 73352
rect 49998 73312 50040 73352
rect 50080 73312 64832 73352
rect 64872 73312 64914 73352
rect 64954 73312 64996 73352
rect 65036 73312 65078 73352
rect 65118 73312 65160 73352
rect 65200 73312 79952 73352
rect 79992 73312 80034 73352
rect 80074 73312 80116 73352
rect 80156 73312 80198 73352
rect 80238 73312 80280 73352
rect 80320 73312 95072 73352
rect 95112 73312 95154 73352
rect 95194 73312 95236 73352
rect 95276 73312 95318 73352
rect 95358 73312 95400 73352
rect 95440 73312 99360 73352
rect 576 73288 99360 73312
rect 643 72932 701 72933
rect 643 72892 652 72932
rect 692 72892 701 72932
rect 643 72891 701 72892
rect 843 72764 885 72773
rect 843 72724 844 72764
rect 884 72724 885 72764
rect 843 72715 885 72724
rect 576 72596 99360 72620
rect 576 72556 3112 72596
rect 3152 72556 3194 72596
rect 3234 72556 3276 72596
rect 3316 72556 3358 72596
rect 3398 72556 3440 72596
rect 3480 72556 18232 72596
rect 18272 72556 18314 72596
rect 18354 72556 18396 72596
rect 18436 72556 18478 72596
rect 18518 72556 18560 72596
rect 18600 72556 33352 72596
rect 33392 72556 33434 72596
rect 33474 72556 33516 72596
rect 33556 72556 33598 72596
rect 33638 72556 33680 72596
rect 33720 72556 48472 72596
rect 48512 72556 48554 72596
rect 48594 72556 48636 72596
rect 48676 72556 48718 72596
rect 48758 72556 48800 72596
rect 48840 72556 63592 72596
rect 63632 72556 63674 72596
rect 63714 72556 63756 72596
rect 63796 72556 63838 72596
rect 63878 72556 63920 72596
rect 63960 72556 78712 72596
rect 78752 72556 78794 72596
rect 78834 72556 78876 72596
rect 78916 72556 78958 72596
rect 78998 72556 79040 72596
rect 79080 72556 93832 72596
rect 93872 72556 93914 72596
rect 93954 72556 93996 72596
rect 94036 72556 94078 72596
rect 94118 72556 94160 72596
rect 94200 72556 99360 72596
rect 576 72532 99360 72556
rect 576 71840 99360 71864
rect 576 71800 4352 71840
rect 4392 71800 4434 71840
rect 4474 71800 4516 71840
rect 4556 71800 4598 71840
rect 4638 71800 4680 71840
rect 4720 71800 19472 71840
rect 19512 71800 19554 71840
rect 19594 71800 19636 71840
rect 19676 71800 19718 71840
rect 19758 71800 19800 71840
rect 19840 71800 34592 71840
rect 34632 71800 34674 71840
rect 34714 71800 34756 71840
rect 34796 71800 34838 71840
rect 34878 71800 34920 71840
rect 34960 71800 49712 71840
rect 49752 71800 49794 71840
rect 49834 71800 49876 71840
rect 49916 71800 49958 71840
rect 49998 71800 50040 71840
rect 50080 71800 64832 71840
rect 64872 71800 64914 71840
rect 64954 71800 64996 71840
rect 65036 71800 65078 71840
rect 65118 71800 65160 71840
rect 65200 71800 79952 71840
rect 79992 71800 80034 71840
rect 80074 71800 80116 71840
rect 80156 71800 80198 71840
rect 80238 71800 80280 71840
rect 80320 71800 95072 71840
rect 95112 71800 95154 71840
rect 95194 71800 95236 71840
rect 95276 71800 95318 71840
rect 95358 71800 95400 71840
rect 95440 71800 99360 71840
rect 576 71776 99360 71800
rect 643 71504 701 71505
rect 643 71464 652 71504
rect 692 71464 701 71504
rect 643 71463 701 71464
rect 835 71504 893 71505
rect 835 71464 844 71504
rect 884 71464 893 71504
rect 835 71463 893 71464
rect 576 71084 99360 71108
rect 576 71044 3112 71084
rect 3152 71044 3194 71084
rect 3234 71044 3276 71084
rect 3316 71044 3358 71084
rect 3398 71044 3440 71084
rect 3480 71044 18232 71084
rect 18272 71044 18314 71084
rect 18354 71044 18396 71084
rect 18436 71044 18478 71084
rect 18518 71044 18560 71084
rect 18600 71044 33352 71084
rect 33392 71044 33434 71084
rect 33474 71044 33516 71084
rect 33556 71044 33598 71084
rect 33638 71044 33680 71084
rect 33720 71044 48472 71084
rect 48512 71044 48554 71084
rect 48594 71044 48636 71084
rect 48676 71044 48718 71084
rect 48758 71044 48800 71084
rect 48840 71044 63592 71084
rect 63632 71044 63674 71084
rect 63714 71044 63756 71084
rect 63796 71044 63838 71084
rect 63878 71044 63920 71084
rect 63960 71044 78712 71084
rect 78752 71044 78794 71084
rect 78834 71044 78876 71084
rect 78916 71044 78958 71084
rect 78998 71044 79040 71084
rect 79080 71044 93832 71084
rect 93872 71044 93914 71084
rect 93954 71044 93996 71084
rect 94036 71044 94078 71084
rect 94118 71044 94160 71084
rect 94200 71044 99360 71084
rect 576 71020 99360 71044
rect 576 70328 99360 70352
rect 576 70288 4352 70328
rect 4392 70288 4434 70328
rect 4474 70288 4516 70328
rect 4556 70288 4598 70328
rect 4638 70288 4680 70328
rect 4720 70288 19472 70328
rect 19512 70288 19554 70328
rect 19594 70288 19636 70328
rect 19676 70288 19718 70328
rect 19758 70288 19800 70328
rect 19840 70288 34592 70328
rect 34632 70288 34674 70328
rect 34714 70288 34756 70328
rect 34796 70288 34838 70328
rect 34878 70288 34920 70328
rect 34960 70288 49712 70328
rect 49752 70288 49794 70328
rect 49834 70288 49876 70328
rect 49916 70288 49958 70328
rect 49998 70288 50040 70328
rect 50080 70288 64832 70328
rect 64872 70288 64914 70328
rect 64954 70288 64996 70328
rect 65036 70288 65078 70328
rect 65118 70288 65160 70328
rect 65200 70288 79952 70328
rect 79992 70288 80034 70328
rect 80074 70288 80116 70328
rect 80156 70288 80198 70328
rect 80238 70288 80280 70328
rect 80320 70288 95072 70328
rect 95112 70288 95154 70328
rect 95194 70288 95236 70328
rect 95276 70288 95318 70328
rect 95358 70288 95400 70328
rect 95440 70288 99360 70328
rect 576 70264 99360 70288
rect 576 69572 99360 69596
rect 576 69532 3112 69572
rect 3152 69532 3194 69572
rect 3234 69532 3276 69572
rect 3316 69532 3358 69572
rect 3398 69532 3440 69572
rect 3480 69532 18232 69572
rect 18272 69532 18314 69572
rect 18354 69532 18396 69572
rect 18436 69532 18478 69572
rect 18518 69532 18560 69572
rect 18600 69532 33352 69572
rect 33392 69532 33434 69572
rect 33474 69532 33516 69572
rect 33556 69532 33598 69572
rect 33638 69532 33680 69572
rect 33720 69532 48472 69572
rect 48512 69532 48554 69572
rect 48594 69532 48636 69572
rect 48676 69532 48718 69572
rect 48758 69532 48800 69572
rect 48840 69532 63592 69572
rect 63632 69532 63674 69572
rect 63714 69532 63756 69572
rect 63796 69532 63838 69572
rect 63878 69532 63920 69572
rect 63960 69532 78712 69572
rect 78752 69532 78794 69572
rect 78834 69532 78876 69572
rect 78916 69532 78958 69572
rect 78998 69532 79040 69572
rect 79080 69532 93832 69572
rect 93872 69532 93914 69572
rect 93954 69532 93996 69572
rect 94036 69532 94078 69572
rect 94118 69532 94160 69572
rect 94200 69532 99360 69572
rect 576 69508 99360 69532
rect 643 69236 701 69237
rect 643 69196 652 69236
rect 692 69196 701 69236
rect 643 69195 701 69196
rect 843 68984 885 68993
rect 843 68944 844 68984
rect 884 68944 885 68984
rect 843 68935 885 68944
rect 576 68816 99360 68840
rect 576 68776 4352 68816
rect 4392 68776 4434 68816
rect 4474 68776 4516 68816
rect 4556 68776 4598 68816
rect 4638 68776 4680 68816
rect 4720 68776 19472 68816
rect 19512 68776 19554 68816
rect 19594 68776 19636 68816
rect 19676 68776 19718 68816
rect 19758 68776 19800 68816
rect 19840 68776 34592 68816
rect 34632 68776 34674 68816
rect 34714 68776 34756 68816
rect 34796 68776 34838 68816
rect 34878 68776 34920 68816
rect 34960 68776 49712 68816
rect 49752 68776 49794 68816
rect 49834 68776 49876 68816
rect 49916 68776 49958 68816
rect 49998 68776 50040 68816
rect 50080 68776 64832 68816
rect 64872 68776 64914 68816
rect 64954 68776 64996 68816
rect 65036 68776 65078 68816
rect 65118 68776 65160 68816
rect 65200 68776 79952 68816
rect 79992 68776 80034 68816
rect 80074 68776 80116 68816
rect 80156 68776 80198 68816
rect 80238 68776 80280 68816
rect 80320 68776 95072 68816
rect 95112 68776 95154 68816
rect 95194 68776 95236 68816
rect 95276 68776 95318 68816
rect 95358 68776 95400 68816
rect 95440 68776 99360 68816
rect 576 68752 99360 68776
rect 576 68060 99360 68084
rect 576 68020 3112 68060
rect 3152 68020 3194 68060
rect 3234 68020 3276 68060
rect 3316 68020 3358 68060
rect 3398 68020 3440 68060
rect 3480 68020 18232 68060
rect 18272 68020 18314 68060
rect 18354 68020 18396 68060
rect 18436 68020 18478 68060
rect 18518 68020 18560 68060
rect 18600 68020 33352 68060
rect 33392 68020 33434 68060
rect 33474 68020 33516 68060
rect 33556 68020 33598 68060
rect 33638 68020 33680 68060
rect 33720 68020 48472 68060
rect 48512 68020 48554 68060
rect 48594 68020 48636 68060
rect 48676 68020 48718 68060
rect 48758 68020 48800 68060
rect 48840 68020 63592 68060
rect 63632 68020 63674 68060
rect 63714 68020 63756 68060
rect 63796 68020 63838 68060
rect 63878 68020 63920 68060
rect 63960 68020 78712 68060
rect 78752 68020 78794 68060
rect 78834 68020 78876 68060
rect 78916 68020 78958 68060
rect 78998 68020 79040 68060
rect 79080 68020 93832 68060
rect 93872 68020 93914 68060
rect 93954 68020 93996 68060
rect 94036 68020 94078 68060
rect 94118 68020 94160 68060
rect 94200 68020 99360 68060
rect 576 67996 99360 68020
rect 643 67724 701 67725
rect 643 67684 652 67724
rect 692 67684 701 67724
rect 643 67683 701 67684
rect 843 67472 885 67481
rect 843 67432 844 67472
rect 884 67432 885 67472
rect 843 67423 885 67432
rect 576 67304 99360 67328
rect 576 67264 4352 67304
rect 4392 67264 4434 67304
rect 4474 67264 4516 67304
rect 4556 67264 4598 67304
rect 4638 67264 4680 67304
rect 4720 67264 19472 67304
rect 19512 67264 19554 67304
rect 19594 67264 19636 67304
rect 19676 67264 19718 67304
rect 19758 67264 19800 67304
rect 19840 67264 34592 67304
rect 34632 67264 34674 67304
rect 34714 67264 34756 67304
rect 34796 67264 34838 67304
rect 34878 67264 34920 67304
rect 34960 67264 49712 67304
rect 49752 67264 49794 67304
rect 49834 67264 49876 67304
rect 49916 67264 49958 67304
rect 49998 67264 50040 67304
rect 50080 67264 64832 67304
rect 64872 67264 64914 67304
rect 64954 67264 64996 67304
rect 65036 67264 65078 67304
rect 65118 67264 65160 67304
rect 65200 67264 79952 67304
rect 79992 67264 80034 67304
rect 80074 67264 80116 67304
rect 80156 67264 80198 67304
rect 80238 67264 80280 67304
rect 80320 67264 95072 67304
rect 95112 67264 95154 67304
rect 95194 67264 95236 67304
rect 95276 67264 95318 67304
rect 95358 67264 95400 67304
rect 95440 67264 99360 67304
rect 576 67240 99360 67264
rect 576 66548 99360 66572
rect 576 66508 3112 66548
rect 3152 66508 3194 66548
rect 3234 66508 3276 66548
rect 3316 66508 3358 66548
rect 3398 66508 3440 66548
rect 3480 66508 18232 66548
rect 18272 66508 18314 66548
rect 18354 66508 18396 66548
rect 18436 66508 18478 66548
rect 18518 66508 18560 66548
rect 18600 66508 33352 66548
rect 33392 66508 33434 66548
rect 33474 66508 33516 66548
rect 33556 66508 33598 66548
rect 33638 66508 33680 66548
rect 33720 66508 48472 66548
rect 48512 66508 48554 66548
rect 48594 66508 48636 66548
rect 48676 66508 48718 66548
rect 48758 66508 48800 66548
rect 48840 66508 63592 66548
rect 63632 66508 63674 66548
rect 63714 66508 63756 66548
rect 63796 66508 63838 66548
rect 63878 66508 63920 66548
rect 63960 66508 78712 66548
rect 78752 66508 78794 66548
rect 78834 66508 78876 66548
rect 78916 66508 78958 66548
rect 78998 66508 79040 66548
rect 79080 66508 93832 66548
rect 93872 66508 93914 66548
rect 93954 66508 93996 66548
rect 94036 66508 94078 66548
rect 94118 66508 94160 66548
rect 94200 66508 99360 66548
rect 576 66484 99360 66508
rect 643 66212 701 66213
rect 643 66172 652 66212
rect 692 66172 701 66212
rect 643 66171 701 66172
rect 843 65960 885 65969
rect 843 65920 844 65960
rect 884 65920 885 65960
rect 843 65911 885 65920
rect 576 65792 99360 65816
rect 576 65752 4352 65792
rect 4392 65752 4434 65792
rect 4474 65752 4516 65792
rect 4556 65752 4598 65792
rect 4638 65752 4680 65792
rect 4720 65752 19472 65792
rect 19512 65752 19554 65792
rect 19594 65752 19636 65792
rect 19676 65752 19718 65792
rect 19758 65752 19800 65792
rect 19840 65752 34592 65792
rect 34632 65752 34674 65792
rect 34714 65752 34756 65792
rect 34796 65752 34838 65792
rect 34878 65752 34920 65792
rect 34960 65752 49712 65792
rect 49752 65752 49794 65792
rect 49834 65752 49876 65792
rect 49916 65752 49958 65792
rect 49998 65752 50040 65792
rect 50080 65752 64832 65792
rect 64872 65752 64914 65792
rect 64954 65752 64996 65792
rect 65036 65752 65078 65792
rect 65118 65752 65160 65792
rect 65200 65752 79952 65792
rect 79992 65752 80034 65792
rect 80074 65752 80116 65792
rect 80156 65752 80198 65792
rect 80238 65752 80280 65792
rect 80320 65752 95072 65792
rect 95112 65752 95154 65792
rect 95194 65752 95236 65792
rect 95276 65752 95318 65792
rect 95358 65752 95400 65792
rect 95440 65752 99360 65792
rect 576 65728 99360 65752
rect 576 65036 99360 65060
rect 576 64996 3112 65036
rect 3152 64996 3194 65036
rect 3234 64996 3276 65036
rect 3316 64996 3358 65036
rect 3398 64996 3440 65036
rect 3480 64996 18232 65036
rect 18272 64996 18314 65036
rect 18354 64996 18396 65036
rect 18436 64996 18478 65036
rect 18518 64996 18560 65036
rect 18600 64996 33352 65036
rect 33392 64996 33434 65036
rect 33474 64996 33516 65036
rect 33556 64996 33598 65036
rect 33638 64996 33680 65036
rect 33720 64996 48472 65036
rect 48512 64996 48554 65036
rect 48594 64996 48636 65036
rect 48676 64996 48718 65036
rect 48758 64996 48800 65036
rect 48840 64996 63592 65036
rect 63632 64996 63674 65036
rect 63714 64996 63756 65036
rect 63796 64996 63838 65036
rect 63878 64996 63920 65036
rect 63960 64996 78712 65036
rect 78752 64996 78794 65036
rect 78834 64996 78876 65036
rect 78916 64996 78958 65036
rect 78998 64996 79040 65036
rect 79080 64996 93832 65036
rect 93872 64996 93914 65036
rect 93954 64996 93996 65036
rect 94036 64996 94078 65036
rect 94118 64996 94160 65036
rect 94200 64996 99360 65036
rect 576 64972 99360 64996
rect 576 64280 99360 64304
rect 576 64240 4352 64280
rect 4392 64240 4434 64280
rect 4474 64240 4516 64280
rect 4556 64240 4598 64280
rect 4638 64240 4680 64280
rect 4720 64240 19472 64280
rect 19512 64240 19554 64280
rect 19594 64240 19636 64280
rect 19676 64240 19718 64280
rect 19758 64240 19800 64280
rect 19840 64240 34592 64280
rect 34632 64240 34674 64280
rect 34714 64240 34756 64280
rect 34796 64240 34838 64280
rect 34878 64240 34920 64280
rect 34960 64240 49712 64280
rect 49752 64240 49794 64280
rect 49834 64240 49876 64280
rect 49916 64240 49958 64280
rect 49998 64240 50040 64280
rect 50080 64240 64832 64280
rect 64872 64240 64914 64280
rect 64954 64240 64996 64280
rect 65036 64240 65078 64280
rect 65118 64240 65160 64280
rect 65200 64240 79952 64280
rect 79992 64240 80034 64280
rect 80074 64240 80116 64280
rect 80156 64240 80198 64280
rect 80238 64240 80280 64280
rect 80320 64240 95072 64280
rect 95112 64240 95154 64280
rect 95194 64240 95236 64280
rect 95276 64240 95318 64280
rect 95358 64240 95400 64280
rect 95440 64240 99360 64280
rect 576 64216 99360 64240
rect 643 63860 701 63861
rect 643 63820 652 63860
rect 692 63820 701 63860
rect 643 63819 701 63820
rect 843 63692 885 63701
rect 843 63652 844 63692
rect 884 63652 885 63692
rect 843 63643 885 63652
rect 576 63524 99360 63548
rect 576 63484 3112 63524
rect 3152 63484 3194 63524
rect 3234 63484 3276 63524
rect 3316 63484 3358 63524
rect 3398 63484 3440 63524
rect 3480 63484 18232 63524
rect 18272 63484 18314 63524
rect 18354 63484 18396 63524
rect 18436 63484 18478 63524
rect 18518 63484 18560 63524
rect 18600 63484 33352 63524
rect 33392 63484 33434 63524
rect 33474 63484 33516 63524
rect 33556 63484 33598 63524
rect 33638 63484 33680 63524
rect 33720 63484 48472 63524
rect 48512 63484 48554 63524
rect 48594 63484 48636 63524
rect 48676 63484 48718 63524
rect 48758 63484 48800 63524
rect 48840 63484 63592 63524
rect 63632 63484 63674 63524
rect 63714 63484 63756 63524
rect 63796 63484 63838 63524
rect 63878 63484 63920 63524
rect 63960 63484 78712 63524
rect 78752 63484 78794 63524
rect 78834 63484 78876 63524
rect 78916 63484 78958 63524
rect 78998 63484 79040 63524
rect 79080 63484 93832 63524
rect 93872 63484 93914 63524
rect 93954 63484 93996 63524
rect 94036 63484 94078 63524
rect 94118 63484 94160 63524
rect 94200 63484 99360 63524
rect 576 63460 99360 63484
rect 576 62768 99360 62792
rect 576 62728 4352 62768
rect 4392 62728 4434 62768
rect 4474 62728 4516 62768
rect 4556 62728 4598 62768
rect 4638 62728 4680 62768
rect 4720 62728 19472 62768
rect 19512 62728 19554 62768
rect 19594 62728 19636 62768
rect 19676 62728 19718 62768
rect 19758 62728 19800 62768
rect 19840 62728 34592 62768
rect 34632 62728 34674 62768
rect 34714 62728 34756 62768
rect 34796 62728 34838 62768
rect 34878 62728 34920 62768
rect 34960 62728 49712 62768
rect 49752 62728 49794 62768
rect 49834 62728 49876 62768
rect 49916 62728 49958 62768
rect 49998 62728 50040 62768
rect 50080 62728 64832 62768
rect 64872 62728 64914 62768
rect 64954 62728 64996 62768
rect 65036 62728 65078 62768
rect 65118 62728 65160 62768
rect 65200 62728 79952 62768
rect 79992 62728 80034 62768
rect 80074 62728 80116 62768
rect 80156 62728 80198 62768
rect 80238 62728 80280 62768
rect 80320 62728 95072 62768
rect 95112 62728 95154 62768
rect 95194 62728 95236 62768
rect 95276 62728 95318 62768
rect 95358 62728 95400 62768
rect 95440 62728 99360 62768
rect 576 62704 99360 62728
rect 643 62348 701 62349
rect 643 62308 652 62348
rect 692 62308 701 62348
rect 643 62307 701 62308
rect 843 62180 885 62189
rect 843 62140 844 62180
rect 884 62140 885 62180
rect 843 62131 885 62140
rect 576 62012 99360 62036
rect 576 61972 3112 62012
rect 3152 61972 3194 62012
rect 3234 61972 3276 62012
rect 3316 61972 3358 62012
rect 3398 61972 3440 62012
rect 3480 61972 18232 62012
rect 18272 61972 18314 62012
rect 18354 61972 18396 62012
rect 18436 61972 18478 62012
rect 18518 61972 18560 62012
rect 18600 61972 33352 62012
rect 33392 61972 33434 62012
rect 33474 61972 33516 62012
rect 33556 61972 33598 62012
rect 33638 61972 33680 62012
rect 33720 61972 48472 62012
rect 48512 61972 48554 62012
rect 48594 61972 48636 62012
rect 48676 61972 48718 62012
rect 48758 61972 48800 62012
rect 48840 61972 63592 62012
rect 63632 61972 63674 62012
rect 63714 61972 63756 62012
rect 63796 61972 63838 62012
rect 63878 61972 63920 62012
rect 63960 61972 78712 62012
rect 78752 61972 78794 62012
rect 78834 61972 78876 62012
rect 78916 61972 78958 62012
rect 78998 61972 79040 62012
rect 79080 61972 93832 62012
rect 93872 61972 93914 62012
rect 93954 61972 93996 62012
rect 94036 61972 94078 62012
rect 94118 61972 94160 62012
rect 94200 61972 99360 62012
rect 576 61948 99360 61972
rect 576 61256 99360 61280
rect 576 61216 4352 61256
rect 4392 61216 4434 61256
rect 4474 61216 4516 61256
rect 4556 61216 4598 61256
rect 4638 61216 4680 61256
rect 4720 61216 19472 61256
rect 19512 61216 19554 61256
rect 19594 61216 19636 61256
rect 19676 61216 19718 61256
rect 19758 61216 19800 61256
rect 19840 61216 34592 61256
rect 34632 61216 34674 61256
rect 34714 61216 34756 61256
rect 34796 61216 34838 61256
rect 34878 61216 34920 61256
rect 34960 61216 49712 61256
rect 49752 61216 49794 61256
rect 49834 61216 49876 61256
rect 49916 61216 49958 61256
rect 49998 61216 50040 61256
rect 50080 61216 64832 61256
rect 64872 61216 64914 61256
rect 64954 61216 64996 61256
rect 65036 61216 65078 61256
rect 65118 61216 65160 61256
rect 65200 61216 79952 61256
rect 79992 61216 80034 61256
rect 80074 61216 80116 61256
rect 80156 61216 80198 61256
rect 80238 61216 80280 61256
rect 80320 61216 95072 61256
rect 95112 61216 95154 61256
rect 95194 61216 95236 61256
rect 95276 61216 95318 61256
rect 95358 61216 95400 61256
rect 95440 61216 99360 61256
rect 576 61192 99360 61216
rect 6507 60920 6549 60929
rect 6507 60880 6508 60920
rect 6548 60880 6549 60920
rect 6507 60871 6549 60880
rect 6595 60920 6653 60921
rect 6595 60880 6604 60920
rect 6644 60880 6653 60920
rect 6595 60879 6653 60880
rect 6883 60836 6941 60837
rect 6883 60796 6892 60836
rect 6932 60796 6941 60836
rect 6883 60795 6941 60796
rect 576 60500 99360 60524
rect 576 60460 3112 60500
rect 3152 60460 3194 60500
rect 3234 60460 3276 60500
rect 3316 60460 3358 60500
rect 3398 60460 3440 60500
rect 3480 60460 18232 60500
rect 18272 60460 18314 60500
rect 18354 60460 18396 60500
rect 18436 60460 18478 60500
rect 18518 60460 18560 60500
rect 18600 60460 33352 60500
rect 33392 60460 33434 60500
rect 33474 60460 33516 60500
rect 33556 60460 33598 60500
rect 33638 60460 33680 60500
rect 33720 60460 48472 60500
rect 48512 60460 48554 60500
rect 48594 60460 48636 60500
rect 48676 60460 48718 60500
rect 48758 60460 48800 60500
rect 48840 60460 63592 60500
rect 63632 60460 63674 60500
rect 63714 60460 63756 60500
rect 63796 60460 63838 60500
rect 63878 60460 63920 60500
rect 63960 60460 78712 60500
rect 78752 60460 78794 60500
rect 78834 60460 78876 60500
rect 78916 60460 78958 60500
rect 78998 60460 79040 60500
rect 79080 60460 93832 60500
rect 93872 60460 93914 60500
rect 93954 60460 93996 60500
rect 94036 60460 94078 60500
rect 94118 60460 94160 60500
rect 94200 60460 99360 60500
rect 576 60436 99360 60460
rect 843 60332 885 60341
rect 843 60292 844 60332
rect 884 60292 885 60332
rect 843 60283 885 60292
rect 643 60164 701 60165
rect 643 60124 652 60164
rect 692 60124 701 60164
rect 643 60123 701 60124
rect 6787 60080 6845 60081
rect 6787 60040 6796 60080
rect 6836 60040 6845 60080
rect 6787 60039 6845 60040
rect 6891 60080 6933 60089
rect 6891 60040 6892 60080
rect 6932 60040 6933 60080
rect 6891 60031 6933 60040
rect 6507 59912 6549 59921
rect 6507 59872 6508 59912
rect 6548 59872 6549 59912
rect 6507 59863 6549 59872
rect 576 59744 99360 59768
rect 576 59704 4352 59744
rect 4392 59704 4434 59744
rect 4474 59704 4516 59744
rect 4556 59704 4598 59744
rect 4638 59704 4680 59744
rect 4720 59704 19472 59744
rect 19512 59704 19554 59744
rect 19594 59704 19636 59744
rect 19676 59704 19718 59744
rect 19758 59704 19800 59744
rect 19840 59704 34592 59744
rect 34632 59704 34674 59744
rect 34714 59704 34756 59744
rect 34796 59704 34838 59744
rect 34878 59704 34920 59744
rect 34960 59704 49712 59744
rect 49752 59704 49794 59744
rect 49834 59704 49876 59744
rect 49916 59704 49958 59744
rect 49998 59704 50040 59744
rect 50080 59704 64832 59744
rect 64872 59704 64914 59744
rect 64954 59704 64996 59744
rect 65036 59704 65078 59744
rect 65118 59704 65160 59744
rect 65200 59704 79952 59744
rect 79992 59704 80034 59744
rect 80074 59704 80116 59744
rect 80156 59704 80198 59744
rect 80238 59704 80280 59744
rect 80320 59704 95072 59744
rect 95112 59704 95154 59744
rect 95194 59704 95236 59744
rect 95276 59704 95318 59744
rect 95358 59704 95400 59744
rect 95440 59704 99360 59744
rect 576 59680 99360 59704
rect 576 58988 99360 59012
rect 576 58948 3112 58988
rect 3152 58948 3194 58988
rect 3234 58948 3276 58988
rect 3316 58948 3358 58988
rect 3398 58948 3440 58988
rect 3480 58948 18232 58988
rect 18272 58948 18314 58988
rect 18354 58948 18396 58988
rect 18436 58948 18478 58988
rect 18518 58948 18560 58988
rect 18600 58948 33352 58988
rect 33392 58948 33434 58988
rect 33474 58948 33516 58988
rect 33556 58948 33598 58988
rect 33638 58948 33680 58988
rect 33720 58948 48472 58988
rect 48512 58948 48554 58988
rect 48594 58948 48636 58988
rect 48676 58948 48718 58988
rect 48758 58948 48800 58988
rect 48840 58948 63592 58988
rect 63632 58948 63674 58988
rect 63714 58948 63756 58988
rect 63796 58948 63838 58988
rect 63878 58948 63920 58988
rect 63960 58948 78712 58988
rect 78752 58948 78794 58988
rect 78834 58948 78876 58988
rect 78916 58948 78958 58988
rect 78998 58948 79040 58988
rect 79080 58948 93832 58988
rect 93872 58948 93914 58988
rect 93954 58948 93996 58988
rect 94036 58948 94078 58988
rect 94118 58948 94160 58988
rect 94200 58948 99360 58988
rect 576 58924 99360 58948
rect 643 58652 701 58653
rect 643 58612 652 58652
rect 692 58612 701 58652
rect 643 58611 701 58612
rect 843 58400 885 58409
rect 843 58360 844 58400
rect 884 58360 885 58400
rect 843 58351 885 58360
rect 576 58232 99360 58256
rect 576 58192 4352 58232
rect 4392 58192 4434 58232
rect 4474 58192 4516 58232
rect 4556 58192 4598 58232
rect 4638 58192 4680 58232
rect 4720 58192 19472 58232
rect 19512 58192 19554 58232
rect 19594 58192 19636 58232
rect 19676 58192 19718 58232
rect 19758 58192 19800 58232
rect 19840 58192 34592 58232
rect 34632 58192 34674 58232
rect 34714 58192 34756 58232
rect 34796 58192 34838 58232
rect 34878 58192 34920 58232
rect 34960 58192 49712 58232
rect 49752 58192 49794 58232
rect 49834 58192 49876 58232
rect 49916 58192 49958 58232
rect 49998 58192 50040 58232
rect 50080 58192 64832 58232
rect 64872 58192 64914 58232
rect 64954 58192 64996 58232
rect 65036 58192 65078 58232
rect 65118 58192 65160 58232
rect 65200 58192 79952 58232
rect 79992 58192 80034 58232
rect 80074 58192 80116 58232
rect 80156 58192 80198 58232
rect 80238 58192 80280 58232
rect 80320 58192 95072 58232
rect 95112 58192 95154 58232
rect 95194 58192 95236 58232
rect 95276 58192 95318 58232
rect 95358 58192 95400 58232
rect 95440 58192 99360 58232
rect 576 58168 99360 58192
rect 6315 57896 6357 57905
rect 6315 57856 6316 57896
rect 6356 57856 6357 57896
rect 6315 57847 6357 57856
rect 6507 57896 6549 57905
rect 6507 57856 6508 57896
rect 6548 57856 6549 57896
rect 6507 57847 6549 57856
rect 6507 57644 6549 57653
rect 6507 57604 6508 57644
rect 6548 57604 6549 57644
rect 6507 57595 6549 57604
rect 576 57476 99360 57500
rect 576 57436 3112 57476
rect 3152 57436 3194 57476
rect 3234 57436 3276 57476
rect 3316 57436 3358 57476
rect 3398 57436 3440 57476
rect 3480 57436 18232 57476
rect 18272 57436 18314 57476
rect 18354 57436 18396 57476
rect 18436 57436 18478 57476
rect 18518 57436 18560 57476
rect 18600 57436 33352 57476
rect 33392 57436 33434 57476
rect 33474 57436 33516 57476
rect 33556 57436 33598 57476
rect 33638 57436 33680 57476
rect 33720 57436 48472 57476
rect 48512 57436 48554 57476
rect 48594 57436 48636 57476
rect 48676 57436 48718 57476
rect 48758 57436 48800 57476
rect 48840 57436 63592 57476
rect 63632 57436 63674 57476
rect 63714 57436 63756 57476
rect 63796 57436 63838 57476
rect 63878 57436 63920 57476
rect 63960 57436 78712 57476
rect 78752 57436 78794 57476
rect 78834 57436 78876 57476
rect 78916 57436 78958 57476
rect 78998 57436 79040 57476
rect 79080 57436 93832 57476
rect 93872 57436 93914 57476
rect 93954 57436 93996 57476
rect 94036 57436 94078 57476
rect 94118 57436 94160 57476
rect 94200 57436 99360 57476
rect 576 57412 99360 57436
rect 6022 57079 6080 57080
rect 5835 57056 5877 57065
rect 5835 57016 5836 57056
rect 5876 57016 5877 57056
rect 5835 57007 5877 57016
rect 5931 57056 5973 57065
rect 5931 57016 5932 57056
rect 5972 57016 5973 57056
rect 6022 57039 6031 57079
rect 6071 57039 6080 57079
rect 6022 57038 6080 57039
rect 6211 57056 6269 57057
rect 5931 57007 5973 57016
rect 6211 57016 6220 57056
rect 6260 57016 6269 57056
rect 6211 57015 6269 57016
rect 6499 57056 6557 57057
rect 6499 57016 6508 57056
rect 6548 57016 6557 57056
rect 6499 57015 6557 57016
rect 6987 57056 7029 57065
rect 6987 57016 6988 57056
rect 7028 57016 7029 57056
rect 6987 57007 7029 57016
rect 7083 57056 7125 57065
rect 7083 57016 7084 57056
rect 7124 57016 7125 57056
rect 7083 57007 7125 57016
rect 7179 57056 7221 57065
rect 7179 57016 7180 57056
rect 7220 57016 7221 57056
rect 7179 57007 7221 57016
rect 7275 57056 7317 57065
rect 7275 57016 7276 57056
rect 7316 57016 7317 57056
rect 7275 57007 7317 57016
rect 6699 56888 6741 56897
rect 6699 56848 6700 56888
rect 6740 56848 6741 56888
rect 6699 56839 6741 56848
rect 576 56720 99360 56744
rect 576 56680 4352 56720
rect 4392 56680 4434 56720
rect 4474 56680 4516 56720
rect 4556 56680 4598 56720
rect 4638 56680 4680 56720
rect 4720 56680 19472 56720
rect 19512 56680 19554 56720
rect 19594 56680 19636 56720
rect 19676 56680 19718 56720
rect 19758 56680 19800 56720
rect 19840 56680 34592 56720
rect 34632 56680 34674 56720
rect 34714 56680 34756 56720
rect 34796 56680 34838 56720
rect 34878 56680 34920 56720
rect 34960 56680 49712 56720
rect 49752 56680 49794 56720
rect 49834 56680 49876 56720
rect 49916 56680 49958 56720
rect 49998 56680 50040 56720
rect 50080 56680 64832 56720
rect 64872 56680 64914 56720
rect 64954 56680 64996 56720
rect 65036 56680 65078 56720
rect 65118 56680 65160 56720
rect 65200 56680 79952 56720
rect 79992 56680 80034 56720
rect 80074 56680 80116 56720
rect 80156 56680 80198 56720
rect 80238 56680 80280 56720
rect 80320 56680 95072 56720
rect 95112 56680 95154 56720
rect 95194 56680 95236 56720
rect 95276 56680 95318 56720
rect 95358 56680 95400 56720
rect 95440 56680 99360 56720
rect 576 56656 99360 56680
rect 6595 56384 6653 56385
rect 6595 56344 6604 56384
rect 6644 56344 6653 56384
rect 6595 56343 6653 56344
rect 6699 56384 6741 56393
rect 6699 56344 6700 56384
rect 6740 56344 6741 56384
rect 6699 56335 6741 56344
rect 643 56300 701 56301
rect 643 56260 652 56300
rect 692 56260 701 56300
rect 643 56259 701 56260
rect 843 56132 885 56141
rect 843 56092 844 56132
rect 884 56092 885 56132
rect 843 56083 885 56092
rect 6411 56132 6453 56141
rect 6411 56092 6412 56132
rect 6452 56092 6453 56132
rect 6411 56083 6453 56092
rect 576 55964 99360 55988
rect 576 55924 3112 55964
rect 3152 55924 3194 55964
rect 3234 55924 3276 55964
rect 3316 55924 3358 55964
rect 3398 55924 3440 55964
rect 3480 55924 18232 55964
rect 18272 55924 18314 55964
rect 18354 55924 18396 55964
rect 18436 55924 18478 55964
rect 18518 55924 18560 55964
rect 18600 55924 33352 55964
rect 33392 55924 33434 55964
rect 33474 55924 33516 55964
rect 33556 55924 33598 55964
rect 33638 55924 33680 55964
rect 33720 55924 48472 55964
rect 48512 55924 48554 55964
rect 48594 55924 48636 55964
rect 48676 55924 48718 55964
rect 48758 55924 48800 55964
rect 48840 55924 63592 55964
rect 63632 55924 63674 55964
rect 63714 55924 63756 55964
rect 63796 55924 63838 55964
rect 63878 55924 63920 55964
rect 63960 55924 78712 55964
rect 78752 55924 78794 55964
rect 78834 55924 78876 55964
rect 78916 55924 78958 55964
rect 78998 55924 79040 55964
rect 79080 55924 93832 55964
rect 93872 55924 93914 55964
rect 93954 55924 93996 55964
rect 94036 55924 94078 55964
rect 94118 55924 94160 55964
rect 94200 55924 99360 55964
rect 576 55900 99360 55924
rect 576 55208 99360 55232
rect 576 55168 4352 55208
rect 4392 55168 4434 55208
rect 4474 55168 4516 55208
rect 4556 55168 4598 55208
rect 4638 55168 4680 55208
rect 4720 55168 19472 55208
rect 19512 55168 19554 55208
rect 19594 55168 19636 55208
rect 19676 55168 19718 55208
rect 19758 55168 19800 55208
rect 19840 55168 34592 55208
rect 34632 55168 34674 55208
rect 34714 55168 34756 55208
rect 34796 55168 34838 55208
rect 34878 55168 34920 55208
rect 34960 55168 49712 55208
rect 49752 55168 49794 55208
rect 49834 55168 49876 55208
rect 49916 55168 49958 55208
rect 49998 55168 50040 55208
rect 50080 55168 64832 55208
rect 64872 55168 64914 55208
rect 64954 55168 64996 55208
rect 65036 55168 65078 55208
rect 65118 55168 65160 55208
rect 65200 55168 79952 55208
rect 79992 55168 80034 55208
rect 80074 55168 80116 55208
rect 80156 55168 80198 55208
rect 80238 55168 80280 55208
rect 80320 55168 95072 55208
rect 95112 55168 95154 55208
rect 95194 55168 95236 55208
rect 95276 55168 95318 55208
rect 95358 55168 95400 55208
rect 95440 55168 99360 55208
rect 576 55144 99360 55168
rect 643 54788 701 54789
rect 643 54748 652 54788
rect 692 54748 701 54788
rect 643 54747 701 54748
rect 843 54620 885 54629
rect 843 54580 844 54620
rect 884 54580 885 54620
rect 843 54571 885 54580
rect 576 54452 99360 54476
rect 576 54412 3112 54452
rect 3152 54412 3194 54452
rect 3234 54412 3276 54452
rect 3316 54412 3358 54452
rect 3398 54412 3440 54452
rect 3480 54412 18232 54452
rect 18272 54412 18314 54452
rect 18354 54412 18396 54452
rect 18436 54412 18478 54452
rect 18518 54412 18560 54452
rect 18600 54412 33352 54452
rect 33392 54412 33434 54452
rect 33474 54412 33516 54452
rect 33556 54412 33598 54452
rect 33638 54412 33680 54452
rect 33720 54412 48472 54452
rect 48512 54412 48554 54452
rect 48594 54412 48636 54452
rect 48676 54412 48718 54452
rect 48758 54412 48800 54452
rect 48840 54412 63592 54452
rect 63632 54412 63674 54452
rect 63714 54412 63756 54452
rect 63796 54412 63838 54452
rect 63878 54412 63920 54452
rect 63960 54412 78712 54452
rect 78752 54412 78794 54452
rect 78834 54412 78876 54452
rect 78916 54412 78958 54452
rect 78998 54412 79040 54452
rect 79080 54412 93832 54452
rect 93872 54412 93914 54452
rect 93954 54412 93996 54452
rect 94036 54412 94078 54452
rect 94118 54412 94160 54452
rect 94200 54412 99360 54452
rect 576 54388 99360 54412
rect 576 53696 99360 53720
rect 576 53656 4352 53696
rect 4392 53656 4434 53696
rect 4474 53656 4516 53696
rect 4556 53656 4598 53696
rect 4638 53656 4680 53696
rect 4720 53656 19472 53696
rect 19512 53656 19554 53696
rect 19594 53656 19636 53696
rect 19676 53656 19718 53696
rect 19758 53656 19800 53696
rect 19840 53656 34592 53696
rect 34632 53656 34674 53696
rect 34714 53656 34756 53696
rect 34796 53656 34838 53696
rect 34878 53656 34920 53696
rect 34960 53656 49712 53696
rect 49752 53656 49794 53696
rect 49834 53656 49876 53696
rect 49916 53656 49958 53696
rect 49998 53656 50040 53696
rect 50080 53656 64832 53696
rect 64872 53656 64914 53696
rect 64954 53656 64996 53696
rect 65036 53656 65078 53696
rect 65118 53656 65160 53696
rect 65200 53656 79952 53696
rect 79992 53656 80034 53696
rect 80074 53656 80116 53696
rect 80156 53656 80198 53696
rect 80238 53656 80280 53696
rect 80320 53656 95072 53696
rect 95112 53656 95154 53696
rect 95194 53656 95236 53696
rect 95276 53656 95318 53696
rect 95358 53656 95400 53696
rect 95440 53656 99360 53696
rect 576 53632 99360 53656
rect 6411 53360 6453 53369
rect 6411 53320 6412 53360
rect 6452 53320 6453 53360
rect 6411 53311 6453 53320
rect 6603 53360 6645 53369
rect 6603 53320 6604 53360
rect 6644 53320 6645 53360
rect 6603 53311 6645 53320
rect 6411 53108 6453 53117
rect 6411 53068 6412 53108
rect 6452 53068 6453 53108
rect 6411 53059 6453 53068
rect 576 52940 99360 52964
rect 576 52900 3112 52940
rect 3152 52900 3194 52940
rect 3234 52900 3276 52940
rect 3316 52900 3358 52940
rect 3398 52900 3440 52940
rect 3480 52900 18232 52940
rect 18272 52900 18314 52940
rect 18354 52900 18396 52940
rect 18436 52900 18478 52940
rect 18518 52900 18560 52940
rect 18600 52900 33352 52940
rect 33392 52900 33434 52940
rect 33474 52900 33516 52940
rect 33556 52900 33598 52940
rect 33638 52900 33680 52940
rect 33720 52900 48472 52940
rect 48512 52900 48554 52940
rect 48594 52900 48636 52940
rect 48676 52900 48718 52940
rect 48758 52900 48800 52940
rect 48840 52900 63592 52940
rect 63632 52900 63674 52940
rect 63714 52900 63756 52940
rect 63796 52900 63838 52940
rect 63878 52900 63920 52940
rect 63960 52900 78712 52940
rect 78752 52900 78794 52940
rect 78834 52900 78876 52940
rect 78916 52900 78958 52940
rect 78998 52900 79040 52940
rect 79080 52900 93832 52940
rect 93872 52900 93914 52940
rect 93954 52900 93996 52940
rect 94036 52900 94078 52940
rect 94118 52900 94160 52940
rect 94200 52900 99360 52940
rect 576 52876 99360 52900
rect 5643 52772 5685 52781
rect 5643 52732 5644 52772
rect 5684 52732 5685 52772
rect 5643 52723 5685 52732
rect 643 52604 701 52605
rect 643 52564 652 52604
rect 692 52564 701 52604
rect 643 52563 701 52564
rect 6184 52535 6226 52544
rect 5635 52520 5693 52521
rect 5635 52480 5644 52520
rect 5684 52480 5693 52520
rect 5635 52479 5693 52480
rect 5731 52520 5789 52521
rect 5731 52480 5740 52520
rect 5780 52480 5789 52520
rect 5731 52479 5789 52480
rect 5931 52520 5973 52529
rect 5931 52480 5932 52520
rect 5972 52480 5973 52520
rect 5931 52471 5973 52480
rect 6027 52520 6069 52529
rect 6027 52480 6028 52520
rect 6068 52480 6069 52520
rect 6184 52495 6185 52535
rect 6225 52495 6226 52535
rect 6184 52486 6226 52495
rect 6595 52520 6653 52521
rect 6027 52471 6069 52480
rect 6595 52480 6604 52520
rect 6644 52480 6653 52520
rect 6595 52479 6653 52480
rect 6691 52520 6749 52521
rect 6691 52480 6700 52520
rect 6740 52480 6749 52520
rect 6691 52479 6749 52480
rect 843 52352 885 52361
rect 843 52312 844 52352
rect 884 52312 885 52352
rect 843 52303 885 52312
rect 6411 52352 6453 52361
rect 6411 52312 6412 52352
rect 6452 52312 6453 52352
rect 6411 52303 6453 52312
rect 576 52184 99360 52208
rect 576 52144 4352 52184
rect 4392 52144 4434 52184
rect 4474 52144 4516 52184
rect 4556 52144 4598 52184
rect 4638 52144 4680 52184
rect 4720 52144 19472 52184
rect 19512 52144 19554 52184
rect 19594 52144 19636 52184
rect 19676 52144 19718 52184
rect 19758 52144 19800 52184
rect 19840 52144 34592 52184
rect 34632 52144 34674 52184
rect 34714 52144 34756 52184
rect 34796 52144 34838 52184
rect 34878 52144 34920 52184
rect 34960 52144 49712 52184
rect 49752 52144 49794 52184
rect 49834 52144 49876 52184
rect 49916 52144 49958 52184
rect 49998 52144 50040 52184
rect 50080 52144 64832 52184
rect 64872 52144 64914 52184
rect 64954 52144 64996 52184
rect 65036 52144 65078 52184
rect 65118 52144 65160 52184
rect 65200 52144 79952 52184
rect 79992 52144 80034 52184
rect 80074 52144 80116 52184
rect 80156 52144 80198 52184
rect 80238 52144 80280 52184
rect 80320 52144 95072 52184
rect 95112 52144 95154 52184
rect 95194 52144 95236 52184
rect 95276 52144 95318 52184
rect 95358 52144 95400 52184
rect 95440 52144 99360 52184
rect 576 52120 99360 52144
rect 5643 52016 5685 52025
rect 5643 51976 5644 52016
rect 5684 51976 5685 52016
rect 5643 51967 5685 51976
rect 6315 52016 6357 52025
rect 6315 51976 6316 52016
rect 6356 51976 6357 52016
rect 6315 51967 6357 51976
rect 2187 51932 2229 51941
rect 2187 51892 2188 51932
rect 2228 51892 2229 51932
rect 2187 51883 2229 51892
rect 2947 51932 3005 51933
rect 2947 51892 2956 51932
rect 2996 51892 3005 51932
rect 2947 51891 3005 51892
rect 2091 51848 2133 51857
rect 2091 51808 2092 51848
rect 2132 51808 2133 51848
rect 2091 51799 2133 51808
rect 2275 51848 2333 51849
rect 2275 51808 2284 51848
rect 2324 51808 2333 51848
rect 2275 51807 2333 51808
rect 2467 51848 2525 51849
rect 2467 51808 2476 51848
rect 2516 51808 2525 51848
rect 2467 51807 2525 51808
rect 2755 51848 2813 51849
rect 2755 51808 2764 51848
rect 2804 51808 2813 51848
rect 2755 51807 2813 51808
rect 3235 51848 3293 51849
rect 3235 51808 3244 51848
rect 3284 51808 3293 51848
rect 3235 51807 3293 51808
rect 3435 51848 3477 51857
rect 3435 51808 3436 51848
rect 3476 51808 3477 51848
rect 3435 51799 3477 51808
rect 3915 51848 3957 51857
rect 3915 51808 3916 51848
rect 3956 51808 3957 51848
rect 3915 51799 3957 51808
rect 4011 51848 4053 51857
rect 4011 51808 4012 51848
rect 4052 51808 4053 51848
rect 4011 51799 4053 51808
rect 4099 51848 4157 51849
rect 4099 51808 4108 51848
rect 4148 51808 4157 51848
rect 4099 51807 4157 51808
rect 5251 51848 5309 51849
rect 5251 51808 5260 51848
rect 5300 51808 5309 51848
rect 5251 51807 5309 51808
rect 5355 51848 5397 51857
rect 5355 51808 5356 51848
rect 5396 51808 5397 51848
rect 5355 51799 5397 51808
rect 5547 51848 5589 51857
rect 5547 51808 5548 51848
rect 5588 51808 5589 51848
rect 5547 51799 5589 51808
rect 5739 51848 5781 51857
rect 5739 51808 5740 51848
rect 5780 51808 5781 51848
rect 5739 51799 5781 51808
rect 6219 51848 6261 51857
rect 6219 51808 6220 51848
rect 6260 51808 6261 51848
rect 6219 51799 6261 51808
rect 6411 51848 6453 51857
rect 6411 51808 6412 51848
rect 6452 51808 6453 51848
rect 6411 51799 6453 51808
rect 6787 51848 6845 51849
rect 6787 51808 6796 51848
rect 6836 51808 6845 51848
rect 6787 51807 6845 51808
rect 6883 51848 6941 51849
rect 6883 51808 6892 51848
rect 6932 51808 6941 51848
rect 6883 51807 6941 51808
rect 3339 51596 3381 51605
rect 3339 51556 3340 51596
rect 3380 51556 3381 51596
rect 3339 51547 3381 51556
rect 6699 51596 6741 51605
rect 6699 51556 6700 51596
rect 6740 51556 6741 51596
rect 6699 51547 6741 51556
rect 576 51428 99360 51452
rect 576 51388 3112 51428
rect 3152 51388 3194 51428
rect 3234 51388 3276 51428
rect 3316 51388 3358 51428
rect 3398 51388 3440 51428
rect 3480 51388 18232 51428
rect 18272 51388 18314 51428
rect 18354 51388 18396 51428
rect 18436 51388 18478 51428
rect 18518 51388 18560 51428
rect 18600 51388 33352 51428
rect 33392 51388 33434 51428
rect 33474 51388 33516 51428
rect 33556 51388 33598 51428
rect 33638 51388 33680 51428
rect 33720 51388 48472 51428
rect 48512 51388 48554 51428
rect 48594 51388 48636 51428
rect 48676 51388 48718 51428
rect 48758 51388 48800 51428
rect 48840 51388 63592 51428
rect 63632 51388 63674 51428
rect 63714 51388 63756 51428
rect 63796 51388 63838 51428
rect 63878 51388 63920 51428
rect 63960 51388 78712 51428
rect 78752 51388 78794 51428
rect 78834 51388 78876 51428
rect 78916 51388 78958 51428
rect 78998 51388 79040 51428
rect 79080 51388 93832 51428
rect 93872 51388 93914 51428
rect 93954 51388 93996 51428
rect 94036 51388 94078 51428
rect 94118 51388 94160 51428
rect 94200 51388 99360 51428
rect 576 51364 99360 51388
rect 643 51092 701 51093
rect 643 51052 652 51092
rect 692 51052 701 51092
rect 643 51051 701 51052
rect 2755 51008 2813 51009
rect 2755 50968 2764 51008
rect 2804 50968 2813 51008
rect 2755 50967 2813 50968
rect 2859 51008 2901 51017
rect 2859 50968 2860 51008
rect 2900 50968 2901 51008
rect 2859 50959 2901 50968
rect 843 50840 885 50849
rect 843 50800 844 50840
rect 884 50800 885 50840
rect 843 50791 885 50800
rect 2475 50840 2517 50849
rect 2475 50800 2476 50840
rect 2516 50800 2517 50840
rect 2475 50791 2517 50800
rect 576 50672 99360 50696
rect 576 50632 4352 50672
rect 4392 50632 4434 50672
rect 4474 50632 4516 50672
rect 4556 50632 4598 50672
rect 4638 50632 4680 50672
rect 4720 50632 19472 50672
rect 19512 50632 19554 50672
rect 19594 50632 19636 50672
rect 19676 50632 19718 50672
rect 19758 50632 19800 50672
rect 19840 50632 34592 50672
rect 34632 50632 34674 50672
rect 34714 50632 34756 50672
rect 34796 50632 34838 50672
rect 34878 50632 34920 50672
rect 34960 50632 49712 50672
rect 49752 50632 49794 50672
rect 49834 50632 49876 50672
rect 49916 50632 49958 50672
rect 49998 50632 50040 50672
rect 50080 50632 64832 50672
rect 64872 50632 64914 50672
rect 64954 50632 64996 50672
rect 65036 50632 65078 50672
rect 65118 50632 65160 50672
rect 65200 50632 79952 50672
rect 79992 50632 80034 50672
rect 80074 50632 80116 50672
rect 80156 50632 80198 50672
rect 80238 50632 80280 50672
rect 80320 50632 95072 50672
rect 95112 50632 95154 50672
rect 95194 50632 95236 50672
rect 95276 50632 95318 50672
rect 95358 50632 95400 50672
rect 95440 50632 99360 50672
rect 576 50608 99360 50632
rect 576 49916 99360 49940
rect 576 49876 3112 49916
rect 3152 49876 3194 49916
rect 3234 49876 3276 49916
rect 3316 49876 3358 49916
rect 3398 49876 3440 49916
rect 3480 49876 18232 49916
rect 18272 49876 18314 49916
rect 18354 49876 18396 49916
rect 18436 49876 18478 49916
rect 18518 49876 18560 49916
rect 18600 49876 33352 49916
rect 33392 49876 33434 49916
rect 33474 49876 33516 49916
rect 33556 49876 33598 49916
rect 33638 49876 33680 49916
rect 33720 49876 48472 49916
rect 48512 49876 48554 49916
rect 48594 49876 48636 49916
rect 48676 49876 48718 49916
rect 48758 49876 48800 49916
rect 48840 49876 63592 49916
rect 63632 49876 63674 49916
rect 63714 49876 63756 49916
rect 63796 49876 63838 49916
rect 63878 49876 63920 49916
rect 63960 49876 78712 49916
rect 78752 49876 78794 49916
rect 78834 49876 78876 49916
rect 78916 49876 78958 49916
rect 78998 49876 79040 49916
rect 79080 49876 93832 49916
rect 93872 49876 93914 49916
rect 93954 49876 93996 49916
rect 94036 49876 94078 49916
rect 94118 49876 94160 49916
rect 94200 49876 99360 49916
rect 576 49852 99360 49876
rect 643 49580 701 49581
rect 643 49540 652 49580
rect 692 49540 701 49580
rect 643 49539 701 49540
rect 843 49328 885 49337
rect 843 49288 844 49328
rect 884 49288 885 49328
rect 843 49279 885 49288
rect 576 49160 99360 49184
rect 576 49120 4352 49160
rect 4392 49120 4434 49160
rect 4474 49120 4516 49160
rect 4556 49120 4598 49160
rect 4638 49120 4680 49160
rect 4720 49120 19472 49160
rect 19512 49120 19554 49160
rect 19594 49120 19636 49160
rect 19676 49120 19718 49160
rect 19758 49120 19800 49160
rect 19840 49120 34592 49160
rect 34632 49120 34674 49160
rect 34714 49120 34756 49160
rect 34796 49120 34838 49160
rect 34878 49120 34920 49160
rect 34960 49120 49712 49160
rect 49752 49120 49794 49160
rect 49834 49120 49876 49160
rect 49916 49120 49958 49160
rect 49998 49120 50040 49160
rect 50080 49120 64832 49160
rect 64872 49120 64914 49160
rect 64954 49120 64996 49160
rect 65036 49120 65078 49160
rect 65118 49120 65160 49160
rect 65200 49120 79952 49160
rect 79992 49120 80034 49160
rect 80074 49120 80116 49160
rect 80156 49120 80198 49160
rect 80238 49120 80280 49160
rect 80320 49120 95072 49160
rect 95112 49120 95154 49160
rect 95194 49120 95236 49160
rect 95276 49120 95318 49160
rect 95358 49120 95400 49160
rect 95440 49120 99360 49160
rect 576 49096 99360 49120
rect 576 48404 99360 48428
rect 576 48364 3112 48404
rect 3152 48364 3194 48404
rect 3234 48364 3276 48404
rect 3316 48364 3358 48404
rect 3398 48364 3440 48404
rect 3480 48364 18232 48404
rect 18272 48364 18314 48404
rect 18354 48364 18396 48404
rect 18436 48364 18478 48404
rect 18518 48364 18560 48404
rect 18600 48364 33352 48404
rect 33392 48364 33434 48404
rect 33474 48364 33516 48404
rect 33556 48364 33598 48404
rect 33638 48364 33680 48404
rect 33720 48364 48472 48404
rect 48512 48364 48554 48404
rect 48594 48364 48636 48404
rect 48676 48364 48718 48404
rect 48758 48364 48800 48404
rect 48840 48364 63592 48404
rect 63632 48364 63674 48404
rect 63714 48364 63756 48404
rect 63796 48364 63838 48404
rect 63878 48364 63920 48404
rect 63960 48364 78712 48404
rect 78752 48364 78794 48404
rect 78834 48364 78876 48404
rect 78916 48364 78958 48404
rect 78998 48364 79040 48404
rect 79080 48364 93832 48404
rect 93872 48364 93914 48404
rect 93954 48364 93996 48404
rect 94036 48364 94078 48404
rect 94118 48364 94160 48404
rect 94200 48364 99360 48404
rect 576 48340 99360 48364
rect 6123 47984 6165 47993
rect 6123 47944 6124 47984
rect 6164 47944 6165 47984
rect 6123 47935 6165 47944
rect 6219 47984 6261 47993
rect 6219 47944 6220 47984
rect 6260 47944 6261 47984
rect 6219 47935 6261 47944
rect 6315 47984 6357 47993
rect 6315 47944 6316 47984
rect 6356 47944 6357 47984
rect 6315 47935 6357 47944
rect 6411 47984 6453 47993
rect 6411 47944 6412 47984
rect 6452 47944 6453 47984
rect 6411 47935 6453 47944
rect 9475 47984 9533 47985
rect 9475 47944 9484 47984
rect 9524 47944 9533 47984
rect 9475 47943 9533 47944
rect 9859 47984 9917 47985
rect 9859 47944 9868 47984
rect 9908 47944 9917 47984
rect 9859 47943 9917 47944
rect 9379 47900 9437 47901
rect 9379 47860 9388 47900
rect 9428 47860 9437 47900
rect 9379 47859 9437 47860
rect 576 47648 99360 47672
rect 576 47608 4352 47648
rect 4392 47608 4434 47648
rect 4474 47608 4516 47648
rect 4556 47608 4598 47648
rect 4638 47608 4680 47648
rect 4720 47608 19472 47648
rect 19512 47608 19554 47648
rect 19594 47608 19636 47648
rect 19676 47608 19718 47648
rect 19758 47608 19800 47648
rect 19840 47608 34592 47648
rect 34632 47608 34674 47648
rect 34714 47608 34756 47648
rect 34796 47608 34838 47648
rect 34878 47608 34920 47648
rect 34960 47608 49712 47648
rect 49752 47608 49794 47648
rect 49834 47608 49876 47648
rect 49916 47608 49958 47648
rect 49998 47608 50040 47648
rect 50080 47608 64832 47648
rect 64872 47608 64914 47648
rect 64954 47608 64996 47648
rect 65036 47608 65078 47648
rect 65118 47608 65160 47648
rect 65200 47608 79952 47648
rect 79992 47608 80034 47648
rect 80074 47608 80116 47648
rect 80156 47608 80198 47648
rect 80238 47608 80280 47648
rect 80320 47608 95072 47648
rect 95112 47608 95154 47648
rect 95194 47608 95236 47648
rect 95276 47608 95318 47648
rect 95358 47608 95400 47648
rect 95440 47608 99360 47648
rect 576 47584 99360 47608
rect 1987 47480 2045 47481
rect 1987 47440 1996 47480
rect 2036 47440 2045 47480
rect 1987 47439 2045 47440
rect 2275 47480 2333 47481
rect 2275 47440 2284 47480
rect 2324 47440 2333 47480
rect 2275 47439 2333 47440
rect 3907 47480 3965 47481
rect 3907 47440 3916 47480
rect 3956 47440 3965 47480
rect 3907 47439 3965 47440
rect 6307 47480 6365 47481
rect 6307 47440 6316 47480
rect 6356 47440 6365 47480
rect 6307 47439 6365 47440
rect 13123 47480 13181 47481
rect 13123 47440 13132 47480
rect 13172 47440 13181 47480
rect 13123 47439 13181 47440
rect 2947 47396 3005 47397
rect 2947 47356 2956 47396
rect 2996 47356 3005 47396
rect 2947 47355 3005 47356
rect 14083 47396 14141 47397
rect 14083 47356 14092 47396
rect 14132 47356 14141 47396
rect 14083 47355 14141 47356
rect 14467 47396 14525 47397
rect 14467 47356 14476 47396
rect 14516 47356 14525 47396
rect 14467 47355 14525 47356
rect 2083 47312 2141 47313
rect 2083 47272 2092 47312
rect 2132 47272 2141 47312
rect 2083 47271 2141 47272
rect 2467 47312 2525 47313
rect 2467 47272 2476 47312
rect 2516 47272 2525 47312
rect 2467 47271 2525 47272
rect 2755 47312 2813 47313
rect 2755 47272 2764 47312
rect 2804 47272 2813 47312
rect 2755 47271 2813 47272
rect 3715 47312 3773 47313
rect 3715 47272 3724 47312
rect 3764 47272 3773 47312
rect 3715 47271 3773 47272
rect 3819 47312 3861 47321
rect 3819 47272 3820 47312
rect 3860 47272 3861 47312
rect 3819 47263 3861 47272
rect 4011 47312 4053 47321
rect 4011 47272 4012 47312
rect 4052 47272 4053 47312
rect 4011 47263 4053 47272
rect 5827 47312 5885 47313
rect 5827 47272 5836 47312
rect 5876 47272 5885 47312
rect 5827 47271 5885 47272
rect 5931 47312 5973 47321
rect 5931 47272 5932 47312
rect 5972 47272 5973 47312
rect 5931 47263 5973 47272
rect 6507 47312 6549 47321
rect 6507 47272 6508 47312
rect 6548 47272 6549 47312
rect 6507 47263 6549 47272
rect 6603 47312 6645 47321
rect 6603 47272 6604 47312
rect 6644 47272 6645 47312
rect 6603 47263 6645 47272
rect 6795 47312 6837 47321
rect 6795 47272 6796 47312
rect 6836 47272 6837 47312
rect 6795 47263 6837 47272
rect 6987 47312 7029 47321
rect 6987 47272 6988 47312
rect 7028 47272 7029 47312
rect 6987 47263 7029 47272
rect 7371 47312 7413 47321
rect 7371 47272 7372 47312
rect 7412 47272 7413 47312
rect 7371 47263 7413 47272
rect 7563 47312 7605 47321
rect 7563 47272 7564 47312
rect 7604 47272 7605 47312
rect 7563 47263 7605 47272
rect 13219 47312 13277 47313
rect 13219 47272 13228 47312
rect 13268 47272 13277 47312
rect 13219 47271 13277 47272
rect 13603 47312 13661 47313
rect 13603 47272 13612 47312
rect 13652 47272 13661 47312
rect 13603 47271 13661 47272
rect 13891 47312 13949 47313
rect 13891 47272 13900 47312
rect 13940 47272 13949 47312
rect 13891 47271 13949 47272
rect 14563 47312 14621 47313
rect 14563 47272 14572 47312
rect 14612 47272 14621 47312
rect 14563 47271 14621 47272
rect 14947 47312 15005 47313
rect 14947 47272 14956 47312
rect 14996 47272 15005 47312
rect 14947 47271 15005 47272
rect 643 47228 701 47229
rect 643 47188 652 47228
rect 692 47188 701 47228
rect 643 47187 701 47188
rect 6891 47228 6933 47237
rect 6891 47188 6892 47228
rect 6932 47188 6933 47228
rect 6891 47179 6933 47188
rect 7371 47144 7413 47153
rect 7371 47104 7372 47144
rect 7412 47104 7413 47144
rect 7371 47095 7413 47104
rect 843 47060 885 47069
rect 843 47020 844 47060
rect 884 47020 885 47060
rect 843 47011 885 47020
rect 5643 47060 5685 47069
rect 5643 47020 5644 47060
rect 5684 47020 5685 47060
rect 5643 47011 5685 47020
rect 13411 47060 13469 47061
rect 13411 47020 13420 47060
rect 13460 47020 13469 47060
rect 13411 47019 13469 47020
rect 576 46892 99360 46916
rect 576 46852 3112 46892
rect 3152 46852 3194 46892
rect 3234 46852 3276 46892
rect 3316 46852 3358 46892
rect 3398 46852 3440 46892
rect 3480 46852 18232 46892
rect 18272 46852 18314 46892
rect 18354 46852 18396 46892
rect 18436 46852 18478 46892
rect 18518 46852 18560 46892
rect 18600 46852 33352 46892
rect 33392 46852 33434 46892
rect 33474 46852 33516 46892
rect 33556 46852 33598 46892
rect 33638 46852 33680 46892
rect 33720 46852 48472 46892
rect 48512 46852 48554 46892
rect 48594 46852 48636 46892
rect 48676 46852 48718 46892
rect 48758 46852 48800 46892
rect 48840 46852 63592 46892
rect 63632 46852 63674 46892
rect 63714 46852 63756 46892
rect 63796 46852 63838 46892
rect 63878 46852 63920 46892
rect 63960 46852 78712 46892
rect 78752 46852 78794 46892
rect 78834 46852 78876 46892
rect 78916 46852 78958 46892
rect 78998 46852 79040 46892
rect 79080 46852 93832 46892
rect 93872 46852 93914 46892
rect 93954 46852 93996 46892
rect 94036 46852 94078 46892
rect 94118 46852 94160 46892
rect 94200 46852 99360 46892
rect 576 46828 99360 46852
rect 2859 46724 2901 46733
rect 2859 46684 2860 46724
rect 2900 46684 2901 46724
rect 2859 46675 2901 46684
rect 2667 46640 2709 46649
rect 2667 46600 2668 46640
rect 2708 46600 2709 46640
rect 2667 46591 2709 46600
rect 13803 46640 13845 46649
rect 13803 46600 13804 46640
rect 13844 46600 13845 46640
rect 13803 46591 13845 46600
rect 13707 46556 13749 46565
rect 13707 46516 13708 46556
rect 13748 46516 13749 46556
rect 13707 46507 13749 46516
rect 14275 46556 14333 46557
rect 14275 46516 14284 46556
rect 14324 46516 14333 46556
rect 14275 46515 14333 46516
rect 2667 46472 2709 46481
rect 2667 46432 2668 46472
rect 2708 46432 2709 46472
rect 2667 46423 2709 46432
rect 14083 46472 14141 46473
rect 14083 46432 14092 46472
rect 14132 46432 14141 46472
rect 14083 46431 14141 46432
rect 576 46136 99360 46160
rect 576 46096 4352 46136
rect 4392 46096 4434 46136
rect 4474 46096 4516 46136
rect 4556 46096 4598 46136
rect 4638 46096 4680 46136
rect 4720 46096 19472 46136
rect 19512 46096 19554 46136
rect 19594 46096 19636 46136
rect 19676 46096 19718 46136
rect 19758 46096 19800 46136
rect 19840 46096 34592 46136
rect 34632 46096 34674 46136
rect 34714 46096 34756 46136
rect 34796 46096 34838 46136
rect 34878 46096 34920 46136
rect 34960 46096 49712 46136
rect 49752 46096 49794 46136
rect 49834 46096 49876 46136
rect 49916 46096 49958 46136
rect 49998 46096 50040 46136
rect 50080 46096 64832 46136
rect 64872 46096 64914 46136
rect 64954 46096 64996 46136
rect 65036 46096 65078 46136
rect 65118 46096 65160 46136
rect 65200 46096 79952 46136
rect 79992 46096 80034 46136
rect 80074 46096 80116 46136
rect 80156 46096 80198 46136
rect 80238 46096 80280 46136
rect 80320 46096 95072 46136
rect 95112 46096 95154 46136
rect 95194 46096 95236 46136
rect 95276 46096 95318 46136
rect 95358 46096 95400 46136
rect 95440 46096 99360 46136
rect 576 46072 99360 46096
rect 643 45968 701 45969
rect 643 45928 652 45968
rect 692 45928 701 45968
rect 643 45927 701 45928
rect 7555 45968 7613 45969
rect 7555 45928 7564 45968
rect 7604 45928 7613 45968
rect 7555 45927 7613 45928
rect 7843 45968 7901 45969
rect 7843 45928 7852 45968
rect 7892 45928 7901 45968
rect 7843 45927 7901 45928
rect 8043 45968 8085 45977
rect 8043 45928 8044 45968
rect 8084 45928 8085 45968
rect 8043 45919 8085 45928
rect 14083 45968 14141 45969
rect 14083 45928 14092 45968
rect 14132 45928 14141 45968
rect 14083 45927 14141 45928
rect 14371 45968 14429 45969
rect 14371 45928 14380 45968
rect 14420 45928 14429 45968
rect 14371 45927 14429 45928
rect 7747 45800 7805 45801
rect 7747 45760 7756 45800
rect 7796 45760 7805 45800
rect 7747 45759 7805 45760
rect 8227 45800 8285 45801
rect 8227 45760 8236 45800
rect 8276 45760 8285 45800
rect 8227 45759 8285 45760
rect 8323 45800 8381 45801
rect 8323 45760 8332 45800
rect 8372 45760 8381 45800
rect 8323 45759 8381 45760
rect 14179 45800 14237 45801
rect 14179 45760 14188 45800
rect 14228 45760 14237 45800
rect 14179 45759 14237 45760
rect 576 45380 99360 45404
rect 576 45340 3112 45380
rect 3152 45340 3194 45380
rect 3234 45340 3276 45380
rect 3316 45340 3358 45380
rect 3398 45340 3440 45380
rect 3480 45340 18232 45380
rect 18272 45340 18314 45380
rect 18354 45340 18396 45380
rect 18436 45340 18478 45380
rect 18518 45340 18560 45380
rect 18600 45340 33352 45380
rect 33392 45340 33434 45380
rect 33474 45340 33516 45380
rect 33556 45340 33598 45380
rect 33638 45340 33680 45380
rect 33720 45340 48472 45380
rect 48512 45340 48554 45380
rect 48594 45340 48636 45380
rect 48676 45340 48718 45380
rect 48758 45340 48800 45380
rect 48840 45340 63592 45380
rect 63632 45340 63674 45380
rect 63714 45340 63756 45380
rect 63796 45340 63838 45380
rect 63878 45340 63920 45380
rect 63960 45340 78712 45380
rect 78752 45340 78794 45380
rect 78834 45340 78876 45380
rect 78916 45340 78958 45380
rect 78998 45340 79040 45380
rect 79080 45340 93832 45380
rect 93872 45340 93914 45380
rect 93954 45340 93996 45380
rect 94036 45340 94078 45380
rect 94118 45340 94160 45380
rect 94200 45340 99360 45380
rect 576 45316 99360 45340
rect 14179 44960 14237 44961
rect 14179 44920 14188 44960
rect 14228 44920 14237 44960
rect 14179 44919 14237 44920
rect 14563 44960 14621 44961
rect 14563 44920 14572 44960
rect 14612 44920 14621 44960
rect 14563 44919 14621 44920
rect 14091 44792 14133 44801
rect 14091 44752 14092 44792
rect 14132 44752 14133 44792
rect 14091 44743 14133 44752
rect 576 44624 99360 44648
rect 576 44584 4352 44624
rect 4392 44584 4434 44624
rect 4474 44584 4516 44624
rect 4556 44584 4598 44624
rect 4638 44584 4680 44624
rect 4720 44584 19472 44624
rect 19512 44584 19554 44624
rect 19594 44584 19636 44624
rect 19676 44584 19718 44624
rect 19758 44584 19800 44624
rect 19840 44584 34592 44624
rect 34632 44584 34674 44624
rect 34714 44584 34756 44624
rect 34796 44584 34838 44624
rect 34878 44584 34920 44624
rect 34960 44584 49712 44624
rect 49752 44584 49794 44624
rect 49834 44584 49876 44624
rect 49916 44584 49958 44624
rect 49998 44584 50040 44624
rect 50080 44584 64832 44624
rect 64872 44584 64914 44624
rect 64954 44584 64996 44624
rect 65036 44584 65078 44624
rect 65118 44584 65160 44624
rect 65200 44584 79952 44624
rect 79992 44584 80034 44624
rect 80074 44584 80116 44624
rect 80156 44584 80198 44624
rect 80238 44584 80280 44624
rect 80320 44584 95072 44624
rect 95112 44584 95154 44624
rect 95194 44584 95236 44624
rect 95276 44584 95318 44624
rect 95358 44584 95400 44624
rect 95440 44584 99360 44624
rect 576 44560 99360 44584
rect 576 43868 99360 43892
rect 576 43828 3112 43868
rect 3152 43828 3194 43868
rect 3234 43828 3276 43868
rect 3316 43828 3358 43868
rect 3398 43828 3440 43868
rect 3480 43828 18232 43868
rect 18272 43828 18314 43868
rect 18354 43828 18396 43868
rect 18436 43828 18478 43868
rect 18518 43828 18560 43868
rect 18600 43828 33352 43868
rect 33392 43828 33434 43868
rect 33474 43828 33516 43868
rect 33556 43828 33598 43868
rect 33638 43828 33680 43868
rect 33720 43828 48472 43868
rect 48512 43828 48554 43868
rect 48594 43828 48636 43868
rect 48676 43828 48718 43868
rect 48758 43828 48800 43868
rect 48840 43828 63592 43868
rect 63632 43828 63674 43868
rect 63714 43828 63756 43868
rect 63796 43828 63838 43868
rect 63878 43828 63920 43868
rect 63960 43828 78712 43868
rect 78752 43828 78794 43868
rect 78834 43828 78876 43868
rect 78916 43828 78958 43868
rect 78998 43828 79040 43868
rect 79080 43828 93832 43868
rect 93872 43828 93914 43868
rect 93954 43828 93996 43868
rect 94036 43828 94078 43868
rect 94118 43828 94160 43868
rect 94200 43828 99360 43868
rect 576 43804 99360 43828
rect 643 43280 701 43281
rect 643 43240 652 43280
rect 692 43240 701 43280
rect 643 43239 701 43240
rect 576 43112 99360 43136
rect 576 43072 4352 43112
rect 4392 43072 4434 43112
rect 4474 43072 4516 43112
rect 4556 43072 4598 43112
rect 4638 43072 4680 43112
rect 4720 43072 19472 43112
rect 19512 43072 19554 43112
rect 19594 43072 19636 43112
rect 19676 43072 19718 43112
rect 19758 43072 19800 43112
rect 19840 43072 34592 43112
rect 34632 43072 34674 43112
rect 34714 43072 34756 43112
rect 34796 43072 34838 43112
rect 34878 43072 34920 43112
rect 34960 43072 49712 43112
rect 49752 43072 49794 43112
rect 49834 43072 49876 43112
rect 49916 43072 49958 43112
rect 49998 43072 50040 43112
rect 50080 43072 64832 43112
rect 64872 43072 64914 43112
rect 64954 43072 64996 43112
rect 65036 43072 65078 43112
rect 65118 43072 65160 43112
rect 65200 43072 79952 43112
rect 79992 43072 80034 43112
rect 80074 43072 80116 43112
rect 80156 43072 80198 43112
rect 80238 43072 80280 43112
rect 80320 43072 95072 43112
rect 95112 43072 95154 43112
rect 95194 43072 95236 43112
rect 95276 43072 95318 43112
rect 95358 43072 95400 43112
rect 95440 43072 99360 43112
rect 576 43048 99360 43072
rect 576 42356 99360 42380
rect 576 42316 3112 42356
rect 3152 42316 3194 42356
rect 3234 42316 3276 42356
rect 3316 42316 3358 42356
rect 3398 42316 3440 42356
rect 3480 42316 18232 42356
rect 18272 42316 18314 42356
rect 18354 42316 18396 42356
rect 18436 42316 18478 42356
rect 18518 42316 18560 42356
rect 18600 42316 33352 42356
rect 33392 42316 33434 42356
rect 33474 42316 33516 42356
rect 33556 42316 33598 42356
rect 33638 42316 33680 42356
rect 33720 42316 48472 42356
rect 48512 42316 48554 42356
rect 48594 42316 48636 42356
rect 48676 42316 48718 42356
rect 48758 42316 48800 42356
rect 48840 42316 63592 42356
rect 63632 42316 63674 42356
rect 63714 42316 63756 42356
rect 63796 42316 63838 42356
rect 63878 42316 63920 42356
rect 63960 42316 78712 42356
rect 78752 42316 78794 42356
rect 78834 42316 78876 42356
rect 78916 42316 78958 42356
rect 78998 42316 79040 42356
rect 79080 42316 93832 42356
rect 93872 42316 93914 42356
rect 93954 42316 93996 42356
rect 94036 42316 94078 42356
rect 94118 42316 94160 42356
rect 94200 42316 99360 42356
rect 576 42292 99360 42316
rect 643 41768 701 41769
rect 643 41728 652 41768
rect 692 41728 701 41768
rect 643 41727 701 41728
rect 576 41600 99360 41624
rect 576 41560 4352 41600
rect 4392 41560 4434 41600
rect 4474 41560 4516 41600
rect 4556 41560 4598 41600
rect 4638 41560 4680 41600
rect 4720 41560 19472 41600
rect 19512 41560 19554 41600
rect 19594 41560 19636 41600
rect 19676 41560 19718 41600
rect 19758 41560 19800 41600
rect 19840 41560 34592 41600
rect 34632 41560 34674 41600
rect 34714 41560 34756 41600
rect 34796 41560 34838 41600
rect 34878 41560 34920 41600
rect 34960 41560 49712 41600
rect 49752 41560 49794 41600
rect 49834 41560 49876 41600
rect 49916 41560 49958 41600
rect 49998 41560 50040 41600
rect 50080 41560 64832 41600
rect 64872 41560 64914 41600
rect 64954 41560 64996 41600
rect 65036 41560 65078 41600
rect 65118 41560 65160 41600
rect 65200 41560 79952 41600
rect 79992 41560 80034 41600
rect 80074 41560 80116 41600
rect 80156 41560 80198 41600
rect 80238 41560 80280 41600
rect 80320 41560 95072 41600
rect 95112 41560 95154 41600
rect 95194 41560 95236 41600
rect 95276 41560 95318 41600
rect 95358 41560 95400 41600
rect 95440 41560 99360 41600
rect 576 41536 99360 41560
rect 576 40844 99360 40868
rect 576 40804 3112 40844
rect 3152 40804 3194 40844
rect 3234 40804 3276 40844
rect 3316 40804 3358 40844
rect 3398 40804 3440 40844
rect 3480 40804 18232 40844
rect 18272 40804 18314 40844
rect 18354 40804 18396 40844
rect 18436 40804 18478 40844
rect 18518 40804 18560 40844
rect 18600 40804 33352 40844
rect 33392 40804 33434 40844
rect 33474 40804 33516 40844
rect 33556 40804 33598 40844
rect 33638 40804 33680 40844
rect 33720 40804 48472 40844
rect 48512 40804 48554 40844
rect 48594 40804 48636 40844
rect 48676 40804 48718 40844
rect 48758 40804 48800 40844
rect 48840 40804 63592 40844
rect 63632 40804 63674 40844
rect 63714 40804 63756 40844
rect 63796 40804 63838 40844
rect 63878 40804 63920 40844
rect 63960 40804 78712 40844
rect 78752 40804 78794 40844
rect 78834 40804 78876 40844
rect 78916 40804 78958 40844
rect 78998 40804 79040 40844
rect 79080 40804 93832 40844
rect 93872 40804 93914 40844
rect 93954 40804 93996 40844
rect 94036 40804 94078 40844
rect 94118 40804 94160 40844
rect 94200 40804 99360 40844
rect 576 40780 99360 40804
rect 576 40088 99360 40112
rect 576 40048 4352 40088
rect 4392 40048 4434 40088
rect 4474 40048 4516 40088
rect 4556 40048 4598 40088
rect 4638 40048 4680 40088
rect 4720 40048 19472 40088
rect 19512 40048 19554 40088
rect 19594 40048 19636 40088
rect 19676 40048 19718 40088
rect 19758 40048 19800 40088
rect 19840 40048 34592 40088
rect 34632 40048 34674 40088
rect 34714 40048 34756 40088
rect 34796 40048 34838 40088
rect 34878 40048 34920 40088
rect 34960 40048 49712 40088
rect 49752 40048 49794 40088
rect 49834 40048 49876 40088
rect 49916 40048 49958 40088
rect 49998 40048 50040 40088
rect 50080 40048 64832 40088
rect 64872 40048 64914 40088
rect 64954 40048 64996 40088
rect 65036 40048 65078 40088
rect 65118 40048 65160 40088
rect 65200 40048 79952 40088
rect 79992 40048 80034 40088
rect 80074 40048 80116 40088
rect 80156 40048 80198 40088
rect 80238 40048 80280 40088
rect 80320 40048 95072 40088
rect 95112 40048 95154 40088
rect 95194 40048 95236 40088
rect 95276 40048 95318 40088
rect 95358 40048 95400 40088
rect 95440 40048 99360 40088
rect 576 40024 99360 40048
rect 643 39920 701 39921
rect 643 39880 652 39920
rect 692 39880 701 39920
rect 643 39879 701 39880
rect 576 39332 99360 39356
rect 576 39292 3112 39332
rect 3152 39292 3194 39332
rect 3234 39292 3276 39332
rect 3316 39292 3358 39332
rect 3398 39292 3440 39332
rect 3480 39292 18232 39332
rect 18272 39292 18314 39332
rect 18354 39292 18396 39332
rect 18436 39292 18478 39332
rect 18518 39292 18560 39332
rect 18600 39292 33352 39332
rect 33392 39292 33434 39332
rect 33474 39292 33516 39332
rect 33556 39292 33598 39332
rect 33638 39292 33680 39332
rect 33720 39292 48472 39332
rect 48512 39292 48554 39332
rect 48594 39292 48636 39332
rect 48676 39292 48718 39332
rect 48758 39292 48800 39332
rect 48840 39292 63592 39332
rect 63632 39292 63674 39332
rect 63714 39292 63756 39332
rect 63796 39292 63838 39332
rect 63878 39292 63920 39332
rect 63960 39292 78712 39332
rect 78752 39292 78794 39332
rect 78834 39292 78876 39332
rect 78916 39292 78958 39332
rect 78998 39292 79040 39332
rect 79080 39292 93832 39332
rect 93872 39292 93914 39332
rect 93954 39292 93996 39332
rect 94036 39292 94078 39332
rect 94118 39292 94160 39332
rect 94200 39292 99360 39332
rect 576 39268 99360 39292
rect 576 38576 99360 38600
rect 576 38536 4352 38576
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4720 38536 19472 38576
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19840 38536 34592 38576
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34960 38536 49712 38576
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 50080 38536 64832 38576
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 65200 38536 79952 38576
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 80320 38536 95072 38576
rect 95112 38536 95154 38576
rect 95194 38536 95236 38576
rect 95276 38536 95318 38576
rect 95358 38536 95400 38576
rect 95440 38536 99360 38576
rect 576 38512 99360 38536
rect 643 38408 701 38409
rect 643 38368 652 38408
rect 692 38368 701 38408
rect 643 38367 701 38368
rect 576 37820 99360 37844
rect 576 37780 3112 37820
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3480 37780 18232 37820
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18600 37780 33352 37820
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33720 37780 48472 37820
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48840 37780 63592 37820
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63960 37780 78712 37820
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 79080 37780 93832 37820
rect 93872 37780 93914 37820
rect 93954 37780 93996 37820
rect 94036 37780 94078 37820
rect 94118 37780 94160 37820
rect 94200 37780 99360 37820
rect 576 37756 99360 37780
rect 576 37064 99360 37088
rect 576 37024 4352 37064
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4720 37024 19472 37064
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19840 37024 34592 37064
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34960 37024 49712 37064
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 50080 37024 64832 37064
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 65200 37024 79952 37064
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 80320 37024 95072 37064
rect 95112 37024 95154 37064
rect 95194 37024 95236 37064
rect 95276 37024 95318 37064
rect 95358 37024 95400 37064
rect 95440 37024 99360 37064
rect 576 37000 99360 37024
rect 576 36308 99360 36332
rect 576 36268 3112 36308
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3480 36268 18232 36308
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18600 36268 33352 36308
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33720 36268 48472 36308
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48840 36268 63592 36308
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63960 36268 78712 36308
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 79080 36268 93832 36308
rect 93872 36268 93914 36308
rect 93954 36268 93996 36308
rect 94036 36268 94078 36308
rect 94118 36268 94160 36308
rect 94200 36268 99360 36308
rect 576 36244 99360 36268
rect 643 35720 701 35721
rect 643 35680 652 35720
rect 692 35680 701 35720
rect 643 35679 701 35680
rect 576 35552 99360 35576
rect 576 35512 4352 35552
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4720 35512 19472 35552
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19840 35512 34592 35552
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34960 35512 49712 35552
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 50080 35512 64832 35552
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 65200 35512 79952 35552
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 80320 35512 95072 35552
rect 95112 35512 95154 35552
rect 95194 35512 95236 35552
rect 95276 35512 95318 35552
rect 95358 35512 95400 35552
rect 95440 35512 99360 35552
rect 576 35488 99360 35512
rect 576 34796 99360 34820
rect 576 34756 3112 34796
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3480 34756 18232 34796
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18600 34756 33352 34796
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33720 34756 48472 34796
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48840 34756 63592 34796
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63960 34756 78712 34796
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 79080 34756 93832 34796
rect 93872 34756 93914 34796
rect 93954 34756 93996 34796
rect 94036 34756 94078 34796
rect 94118 34756 94160 34796
rect 94200 34756 99360 34796
rect 576 34732 99360 34756
rect 643 34208 701 34209
rect 643 34168 652 34208
rect 692 34168 701 34208
rect 643 34167 701 34168
rect 576 34040 99360 34064
rect 576 34000 4352 34040
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4720 34000 19472 34040
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19840 34000 34592 34040
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34960 34000 49712 34040
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 50080 34000 64832 34040
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 65200 34000 79952 34040
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 80320 34000 95072 34040
rect 95112 34000 95154 34040
rect 95194 34000 95236 34040
rect 95276 34000 95318 34040
rect 95358 34000 95400 34040
rect 95440 34000 99360 34040
rect 576 33976 99360 34000
rect 576 33284 99360 33308
rect 576 33244 3112 33284
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3480 33244 18232 33284
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18600 33244 33352 33284
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33720 33244 48472 33284
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48840 33244 63592 33284
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63960 33244 78712 33284
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 79080 33244 93832 33284
rect 93872 33244 93914 33284
rect 93954 33244 93996 33284
rect 94036 33244 94078 33284
rect 94118 33244 94160 33284
rect 94200 33244 99360 33284
rect 576 33220 99360 33244
rect 643 32696 701 32697
rect 643 32656 652 32696
rect 692 32656 701 32696
rect 643 32655 701 32656
rect 576 32528 99360 32552
rect 576 32488 4352 32528
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4720 32488 19472 32528
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19840 32488 34592 32528
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34960 32488 49712 32528
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 50080 32488 64832 32528
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 65200 32488 79952 32528
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 80320 32488 95072 32528
rect 95112 32488 95154 32528
rect 95194 32488 95236 32528
rect 95276 32488 95318 32528
rect 95358 32488 95400 32528
rect 95440 32488 99360 32528
rect 576 32464 99360 32488
rect 576 31772 99360 31796
rect 576 31732 3112 31772
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3480 31732 18232 31772
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18600 31732 33352 31772
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33720 31732 48472 31772
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48840 31732 63592 31772
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63960 31732 78712 31772
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 79080 31732 93832 31772
rect 93872 31732 93914 31772
rect 93954 31732 93996 31772
rect 94036 31732 94078 31772
rect 94118 31732 94160 31772
rect 94200 31732 99360 31772
rect 576 31708 99360 31732
rect 576 31016 99360 31040
rect 576 30976 4352 31016
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4720 30976 19472 31016
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19840 30976 34592 31016
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34960 30976 49712 31016
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 50080 30976 64832 31016
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 65200 30976 79952 31016
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 80320 30976 95072 31016
rect 95112 30976 95154 31016
rect 95194 30976 95236 31016
rect 95276 30976 95318 31016
rect 95358 30976 95400 31016
rect 95440 30976 99360 31016
rect 576 30952 99360 30976
rect 643 30848 701 30849
rect 643 30808 652 30848
rect 692 30808 701 30848
rect 643 30807 701 30808
rect 576 30260 99360 30284
rect 576 30220 3112 30260
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3480 30220 18232 30260
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18600 30220 33352 30260
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33720 30220 48472 30260
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48840 30220 63592 30260
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63960 30220 78712 30260
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 79080 30220 93832 30260
rect 93872 30220 93914 30260
rect 93954 30220 93996 30260
rect 94036 30220 94078 30260
rect 94118 30220 94160 30260
rect 94200 30220 99360 30260
rect 576 30196 99360 30220
rect 576 29504 99360 29528
rect 576 29464 4352 29504
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4720 29464 19472 29504
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19840 29464 34592 29504
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34960 29464 49712 29504
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 50080 29464 64832 29504
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 65200 29464 79952 29504
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 80320 29464 95072 29504
rect 95112 29464 95154 29504
rect 95194 29464 95236 29504
rect 95276 29464 95318 29504
rect 95358 29464 95400 29504
rect 95440 29464 99360 29504
rect 576 29440 99360 29464
rect 643 29336 701 29337
rect 643 29296 652 29336
rect 692 29296 701 29336
rect 643 29295 701 29296
rect 576 28748 99360 28772
rect 576 28708 3112 28748
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3480 28708 18232 28748
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18600 28708 33352 28748
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33720 28708 48472 28748
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48840 28708 63592 28748
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63960 28708 78712 28748
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 79080 28708 93832 28748
rect 93872 28708 93914 28748
rect 93954 28708 93996 28748
rect 94036 28708 94078 28748
rect 94118 28708 94160 28748
rect 94200 28708 99360 28748
rect 576 28684 99360 28708
rect 576 27992 99360 28016
rect 576 27952 4352 27992
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4720 27952 19472 27992
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19840 27952 34592 27992
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34960 27952 49712 27992
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 50080 27952 64832 27992
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 65200 27952 79952 27992
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 80320 27952 95072 27992
rect 95112 27952 95154 27992
rect 95194 27952 95236 27992
rect 95276 27952 95318 27992
rect 95358 27952 95400 27992
rect 95440 27952 99360 27992
rect 576 27928 99360 27952
rect 576 27236 99360 27260
rect 576 27196 3112 27236
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3480 27196 18232 27236
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18600 27196 33352 27236
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33720 27196 48472 27236
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48840 27196 63592 27236
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63960 27196 78712 27236
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 79080 27196 93832 27236
rect 93872 27196 93914 27236
rect 93954 27196 93996 27236
rect 94036 27196 94078 27236
rect 94118 27196 94160 27236
rect 94200 27196 99360 27236
rect 576 27172 99360 27196
rect 643 26648 701 26649
rect 643 26608 652 26648
rect 692 26608 701 26648
rect 643 26607 701 26608
rect 576 26480 99360 26504
rect 576 26440 4352 26480
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4720 26440 19472 26480
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19840 26440 34592 26480
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34960 26440 49712 26480
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 50080 26440 64832 26480
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 65200 26440 79952 26480
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 80320 26440 95072 26480
rect 95112 26440 95154 26480
rect 95194 26440 95236 26480
rect 95276 26440 95318 26480
rect 95358 26440 95400 26480
rect 95440 26440 99360 26480
rect 576 26416 99360 26440
rect 576 25724 99360 25748
rect 576 25684 3112 25724
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3480 25684 18232 25724
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18600 25684 33352 25724
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33720 25684 48472 25724
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48840 25684 63592 25724
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63960 25684 78712 25724
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 79080 25684 93832 25724
rect 93872 25684 93914 25724
rect 93954 25684 93996 25724
rect 94036 25684 94078 25724
rect 94118 25684 94160 25724
rect 94200 25684 99360 25724
rect 576 25660 99360 25684
rect 643 25136 701 25137
rect 643 25096 652 25136
rect 692 25096 701 25136
rect 643 25095 701 25096
rect 576 24968 99360 24992
rect 576 24928 4352 24968
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4720 24928 19472 24968
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19840 24928 34592 24968
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34960 24928 49712 24968
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 50080 24928 64832 24968
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 65200 24928 79952 24968
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 80320 24928 95072 24968
rect 95112 24928 95154 24968
rect 95194 24928 95236 24968
rect 95276 24928 95318 24968
rect 95358 24928 95400 24968
rect 95440 24928 99360 24968
rect 576 24904 99360 24928
rect 576 24212 99360 24236
rect 576 24172 3112 24212
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3480 24172 18232 24212
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18600 24172 33352 24212
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33720 24172 48472 24212
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48840 24172 63592 24212
rect 63632 24172 63674 24212
rect 63714 24172 63756 24212
rect 63796 24172 63838 24212
rect 63878 24172 63920 24212
rect 63960 24172 78712 24212
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 79080 24172 93832 24212
rect 93872 24172 93914 24212
rect 93954 24172 93996 24212
rect 94036 24172 94078 24212
rect 94118 24172 94160 24212
rect 94200 24172 99360 24212
rect 576 24148 99360 24172
rect 576 23456 99360 23480
rect 576 23416 4352 23456
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4720 23416 19472 23456
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19840 23416 34592 23456
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34960 23416 49712 23456
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 50080 23416 64832 23456
rect 64872 23416 64914 23456
rect 64954 23416 64996 23456
rect 65036 23416 65078 23456
rect 65118 23416 65160 23456
rect 65200 23416 79952 23456
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 80320 23416 95072 23456
rect 95112 23416 95154 23456
rect 95194 23416 95236 23456
rect 95276 23416 95318 23456
rect 95358 23416 95400 23456
rect 95440 23416 99360 23456
rect 576 23392 99360 23416
rect 643 23288 701 23289
rect 643 23248 652 23288
rect 692 23248 701 23288
rect 643 23247 701 23248
rect 576 22700 99360 22724
rect 576 22660 3112 22700
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3480 22660 18232 22700
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18600 22660 33352 22700
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33720 22660 48472 22700
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48840 22660 63592 22700
rect 63632 22660 63674 22700
rect 63714 22660 63756 22700
rect 63796 22660 63838 22700
rect 63878 22660 63920 22700
rect 63960 22660 78712 22700
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 79080 22660 93832 22700
rect 93872 22660 93914 22700
rect 93954 22660 93996 22700
rect 94036 22660 94078 22700
rect 94118 22660 94160 22700
rect 94200 22660 99360 22700
rect 576 22636 99360 22660
rect 576 21944 99360 21968
rect 576 21904 4352 21944
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4720 21904 19472 21944
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19840 21904 34592 21944
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34960 21904 49712 21944
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 50080 21904 64832 21944
rect 64872 21904 64914 21944
rect 64954 21904 64996 21944
rect 65036 21904 65078 21944
rect 65118 21904 65160 21944
rect 65200 21904 79952 21944
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 80320 21904 95072 21944
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95440 21904 99360 21944
rect 576 21880 99360 21904
rect 643 21776 701 21777
rect 643 21736 652 21776
rect 692 21736 701 21776
rect 643 21735 701 21736
rect 576 21188 99360 21212
rect 576 21148 3112 21188
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3480 21148 18232 21188
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18600 21148 33352 21188
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33720 21148 48472 21188
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48840 21148 63592 21188
rect 63632 21148 63674 21188
rect 63714 21148 63756 21188
rect 63796 21148 63838 21188
rect 63878 21148 63920 21188
rect 63960 21148 78712 21188
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 79080 21148 93832 21188
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 94200 21148 99360 21188
rect 576 21124 99360 21148
rect 576 20432 99360 20456
rect 576 20392 4352 20432
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4720 20392 19472 20432
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19840 20392 34592 20432
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34960 20392 49712 20432
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 50080 20392 64832 20432
rect 64872 20392 64914 20432
rect 64954 20392 64996 20432
rect 65036 20392 65078 20432
rect 65118 20392 65160 20432
rect 65200 20392 79952 20432
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 80320 20392 95072 20432
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95440 20392 99360 20432
rect 576 20368 99360 20392
rect 576 19676 99360 19700
rect 576 19636 3112 19676
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3480 19636 18232 19676
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18600 19636 33352 19676
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33720 19636 48472 19676
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48840 19636 63592 19676
rect 63632 19636 63674 19676
rect 63714 19636 63756 19676
rect 63796 19636 63838 19676
rect 63878 19636 63920 19676
rect 63960 19636 78712 19676
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 79080 19636 93832 19676
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 94200 19636 99360 19676
rect 576 19612 99360 19636
rect 643 19088 701 19089
rect 643 19048 652 19088
rect 692 19048 701 19088
rect 643 19047 701 19048
rect 576 18920 99360 18944
rect 576 18880 4352 18920
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4720 18880 19472 18920
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19840 18880 34592 18920
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34960 18880 49712 18920
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 50080 18880 64832 18920
rect 64872 18880 64914 18920
rect 64954 18880 64996 18920
rect 65036 18880 65078 18920
rect 65118 18880 65160 18920
rect 65200 18880 79952 18920
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 80320 18880 95072 18920
rect 95112 18880 95154 18920
rect 95194 18880 95236 18920
rect 95276 18880 95318 18920
rect 95358 18880 95400 18920
rect 95440 18880 99360 18920
rect 576 18856 99360 18880
rect 576 18164 99360 18188
rect 576 18124 3112 18164
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3480 18124 18232 18164
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18600 18124 33352 18164
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33720 18124 48472 18164
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48840 18124 63592 18164
rect 63632 18124 63674 18164
rect 63714 18124 63756 18164
rect 63796 18124 63838 18164
rect 63878 18124 63920 18164
rect 63960 18124 78712 18164
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 79080 18124 93832 18164
rect 93872 18124 93914 18164
rect 93954 18124 93996 18164
rect 94036 18124 94078 18164
rect 94118 18124 94160 18164
rect 94200 18124 99360 18164
rect 576 18100 99360 18124
rect 643 17576 701 17577
rect 643 17536 652 17576
rect 692 17536 701 17576
rect 643 17535 701 17536
rect 576 17408 99360 17432
rect 576 17368 4352 17408
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4720 17368 19472 17408
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19840 17368 34592 17408
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34960 17368 49712 17408
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 50080 17368 64832 17408
rect 64872 17368 64914 17408
rect 64954 17368 64996 17408
rect 65036 17368 65078 17408
rect 65118 17368 65160 17408
rect 65200 17368 79952 17408
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 80320 17368 95072 17408
rect 95112 17368 95154 17408
rect 95194 17368 95236 17408
rect 95276 17368 95318 17408
rect 95358 17368 95400 17408
rect 95440 17368 99360 17408
rect 576 17344 99360 17368
rect 576 16652 99360 16676
rect 576 16612 3112 16652
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3480 16612 18232 16652
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18600 16612 33352 16652
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33720 16612 48472 16652
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48840 16612 63592 16652
rect 63632 16612 63674 16652
rect 63714 16612 63756 16652
rect 63796 16612 63838 16652
rect 63878 16612 63920 16652
rect 63960 16612 78712 16652
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 79080 16612 93832 16652
rect 93872 16612 93914 16652
rect 93954 16612 93996 16652
rect 94036 16612 94078 16652
rect 94118 16612 94160 16652
rect 94200 16612 99360 16652
rect 576 16588 99360 16612
rect 835 16316 893 16317
rect 835 16276 844 16316
rect 884 16276 893 16316
rect 835 16275 893 16276
rect 651 16064 693 16073
rect 651 16024 652 16064
rect 692 16024 693 16064
rect 651 16015 693 16024
rect 576 15896 99360 15920
rect 576 15856 4352 15896
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4720 15856 19472 15896
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19840 15856 34592 15896
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34960 15856 49712 15896
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 50080 15856 64832 15896
rect 64872 15856 64914 15896
rect 64954 15856 64996 15896
rect 65036 15856 65078 15896
rect 65118 15856 65160 15896
rect 65200 15856 79952 15896
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 80320 15856 95072 15896
rect 95112 15856 95154 15896
rect 95194 15856 95236 15896
rect 95276 15856 95318 15896
rect 95358 15856 95400 15896
rect 95440 15856 99360 15896
rect 576 15832 99360 15856
rect 576 15140 99360 15164
rect 576 15100 3112 15140
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3480 15100 18232 15140
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18600 15100 33352 15140
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 33720 15100 48472 15140
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48840 15100 63592 15140
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63960 15100 78712 15140
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 79080 15100 93832 15140
rect 93872 15100 93914 15140
rect 93954 15100 93996 15140
rect 94036 15100 94078 15140
rect 94118 15100 94160 15140
rect 94200 15100 99360 15140
rect 576 15076 99360 15100
rect 576 14384 99360 14408
rect 576 14344 4352 14384
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4720 14344 19472 14384
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19840 14344 34592 14384
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34960 14344 49712 14384
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 50080 14344 64832 14384
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 65200 14344 79952 14384
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 80320 14344 95072 14384
rect 95112 14344 95154 14384
rect 95194 14344 95236 14384
rect 95276 14344 95318 14384
rect 95358 14344 95400 14384
rect 95440 14344 99360 14384
rect 576 14320 99360 14344
rect 835 13964 893 13965
rect 835 13924 844 13964
rect 884 13924 893 13964
rect 835 13923 893 13924
rect 651 13796 693 13805
rect 651 13756 652 13796
rect 692 13756 693 13796
rect 651 13747 693 13756
rect 576 13628 99360 13652
rect 576 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 18232 13628
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18600 13588 33352 13628
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33720 13588 48472 13628
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48840 13588 63592 13628
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63960 13588 78712 13628
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 79080 13588 93832 13628
rect 93872 13588 93914 13628
rect 93954 13588 93996 13628
rect 94036 13588 94078 13628
rect 94118 13588 94160 13628
rect 94200 13588 99360 13628
rect 576 13564 99360 13588
rect 576 12872 99360 12896
rect 576 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 19472 12872
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19840 12832 34592 12872
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34960 12832 49712 12872
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 50080 12832 64832 12872
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 65200 12832 79952 12872
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 80320 12832 95072 12872
rect 95112 12832 95154 12872
rect 95194 12832 95236 12872
rect 95276 12832 95318 12872
rect 95358 12832 95400 12872
rect 95440 12832 99360 12872
rect 576 12808 99360 12832
rect 835 12452 893 12453
rect 835 12412 844 12452
rect 884 12412 893 12452
rect 835 12411 893 12412
rect 651 12284 693 12293
rect 651 12244 652 12284
rect 692 12244 693 12284
rect 651 12235 693 12244
rect 576 12116 99360 12140
rect 576 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 18232 12116
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18600 12076 33352 12116
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33720 12076 48472 12116
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48840 12076 63592 12116
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63960 12076 78712 12116
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 79080 12076 93832 12116
rect 93872 12076 93914 12116
rect 93954 12076 93996 12116
rect 94036 12076 94078 12116
rect 94118 12076 94160 12116
rect 94200 12076 99360 12116
rect 576 12052 99360 12076
rect 576 11360 99360 11384
rect 576 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 19472 11360
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19840 11320 34592 11360
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34960 11320 49712 11360
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 50080 11320 64832 11360
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 65200 11320 79952 11360
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 80320 11320 95072 11360
rect 95112 11320 95154 11360
rect 95194 11320 95236 11360
rect 95276 11320 95318 11360
rect 95358 11320 95400 11360
rect 95440 11320 99360 11360
rect 576 11296 99360 11320
rect 576 10604 99360 10628
rect 576 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 18232 10604
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18600 10564 33352 10604
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33720 10564 48472 10604
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48840 10564 63592 10604
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63960 10564 78712 10604
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 79080 10564 93832 10604
rect 93872 10564 93914 10604
rect 93954 10564 93996 10604
rect 94036 10564 94078 10604
rect 94118 10564 94160 10604
rect 94200 10564 99360 10604
rect 576 10540 99360 10564
rect 835 10268 893 10269
rect 835 10228 844 10268
rect 884 10228 893 10268
rect 835 10227 893 10228
rect 651 10016 693 10025
rect 651 9976 652 10016
rect 692 9976 693 10016
rect 651 9967 693 9976
rect 576 9848 99360 9872
rect 576 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 19472 9848
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19840 9808 34592 9848
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34960 9808 49712 9848
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 50080 9808 64832 9848
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 65200 9808 79952 9848
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 80320 9808 95072 9848
rect 95112 9808 95154 9848
rect 95194 9808 95236 9848
rect 95276 9808 95318 9848
rect 95358 9808 95400 9848
rect 95440 9808 99360 9848
rect 576 9784 99360 9808
rect 576 9092 99360 9116
rect 576 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 18232 9092
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18600 9052 33352 9092
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33720 9052 48472 9092
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48840 9052 63592 9092
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63960 9052 78712 9092
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 79080 9052 93832 9092
rect 93872 9052 93914 9092
rect 93954 9052 93996 9092
rect 94036 9052 94078 9092
rect 94118 9052 94160 9092
rect 94200 9052 99360 9092
rect 576 9028 99360 9052
rect 835 8756 893 8757
rect 835 8716 844 8756
rect 884 8716 893 8756
rect 835 8715 893 8716
rect 651 8504 693 8513
rect 651 8464 652 8504
rect 692 8464 693 8504
rect 651 8455 693 8464
rect 576 8336 99360 8360
rect 576 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 19472 8336
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19840 8296 34592 8336
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34960 8296 49712 8336
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 50080 8296 64832 8336
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 65200 8296 79952 8336
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 80320 8296 95072 8336
rect 95112 8296 95154 8336
rect 95194 8296 95236 8336
rect 95276 8296 95318 8336
rect 95358 8296 95400 8336
rect 95440 8296 99360 8336
rect 576 8272 99360 8296
rect 576 7580 99360 7604
rect 576 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 18232 7580
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18600 7540 33352 7580
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33720 7540 48472 7580
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48840 7540 63592 7580
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63960 7540 78712 7580
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 79080 7540 93832 7580
rect 93872 7540 93914 7580
rect 93954 7540 93996 7580
rect 94036 7540 94078 7580
rect 94118 7540 94160 7580
rect 94200 7540 99360 7580
rect 576 7516 99360 7540
rect 576 6824 99360 6848
rect 576 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 19472 6824
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19840 6784 34592 6824
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34960 6784 49712 6824
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 50080 6784 64832 6824
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 65200 6784 79952 6824
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 80320 6784 95072 6824
rect 95112 6784 95154 6824
rect 95194 6784 95236 6824
rect 95276 6784 95318 6824
rect 95358 6784 95400 6824
rect 95440 6784 99360 6824
rect 576 6760 99360 6784
rect 835 6404 893 6405
rect 835 6364 844 6404
rect 884 6364 893 6404
rect 835 6363 893 6364
rect 651 6320 693 6329
rect 651 6280 652 6320
rect 692 6280 693 6320
rect 651 6271 693 6280
rect 576 6068 99360 6092
rect 576 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 18232 6068
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18600 6028 33352 6068
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33720 6028 48472 6068
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48840 6028 63592 6068
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63960 6028 78712 6068
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 79080 6028 93832 6068
rect 93872 6028 93914 6068
rect 93954 6028 93996 6068
rect 94036 6028 94078 6068
rect 94118 6028 94160 6068
rect 94200 6028 99360 6068
rect 576 6004 99360 6028
rect 576 5312 99360 5336
rect 576 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 19472 5312
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19840 5272 34592 5312
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34960 5272 49712 5312
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 50080 5272 64832 5312
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 65200 5272 79952 5312
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 80320 5272 95072 5312
rect 95112 5272 95154 5312
rect 95194 5272 95236 5312
rect 95276 5272 95318 5312
rect 95358 5272 95400 5312
rect 95440 5272 99360 5312
rect 576 5248 99360 5272
rect 835 4892 893 4893
rect 835 4852 844 4892
rect 884 4852 893 4892
rect 835 4851 893 4852
rect 651 4724 693 4733
rect 651 4684 652 4724
rect 692 4684 693 4724
rect 651 4675 693 4684
rect 576 4556 99360 4580
rect 576 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 18232 4556
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18600 4516 33352 4556
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33720 4516 48472 4556
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48840 4516 63592 4556
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63960 4516 78712 4556
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 79080 4516 93832 4556
rect 93872 4516 93914 4556
rect 93954 4516 93996 4556
rect 94036 4516 94078 4556
rect 94118 4516 94160 4556
rect 94200 4516 99360 4556
rect 576 4492 99360 4516
rect 576 3800 99360 3824
rect 576 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 19472 3800
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19840 3760 34592 3800
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34960 3760 49712 3800
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 50080 3760 64832 3800
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 65200 3760 79952 3800
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 80320 3760 95072 3800
rect 95112 3760 95154 3800
rect 95194 3760 95236 3800
rect 95276 3760 95318 3800
rect 95358 3760 95400 3800
rect 95440 3760 99360 3800
rect 576 3736 99360 3760
rect 576 3044 99360 3068
rect 576 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 18232 3044
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18600 3004 33352 3044
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33720 3004 48472 3044
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48840 3004 63592 3044
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63960 3004 78712 3044
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 79080 3004 93832 3044
rect 93872 3004 93914 3044
rect 93954 3004 93996 3044
rect 94036 3004 94078 3044
rect 94118 3004 94160 3044
rect 94200 3004 99360 3044
rect 576 2980 99360 3004
rect 651 2792 693 2801
rect 651 2752 652 2792
rect 692 2752 693 2792
rect 651 2743 693 2752
rect 835 2708 893 2709
rect 835 2668 844 2708
rect 884 2668 893 2708
rect 835 2667 893 2668
rect 576 2288 99360 2312
rect 576 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 19472 2288
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19840 2248 34592 2288
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34960 2248 49712 2288
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 50080 2248 64832 2288
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 65200 2248 79952 2288
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 80320 2248 95072 2288
rect 95112 2248 95154 2288
rect 95194 2248 95236 2288
rect 95276 2248 95318 2288
rect 95358 2248 95400 2288
rect 95440 2248 99360 2288
rect 576 2224 99360 2248
rect 576 1532 99360 1556
rect 576 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 18232 1532
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18600 1492 33352 1532
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33720 1492 48472 1532
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48840 1492 63592 1532
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63960 1492 78712 1532
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 79080 1492 93832 1532
rect 93872 1492 93914 1532
rect 93954 1492 93996 1532
rect 94036 1492 94078 1532
rect 94118 1492 94160 1532
rect 94200 1492 99360 1532
rect 576 1468 99360 1492
rect 576 776 99360 800
rect 576 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 19472 776
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19840 736 34592 776
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34960 736 49712 776
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 50080 736 64832 776
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 65200 736 79952 776
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 80320 736 95072 776
rect 95112 736 95154 776
rect 95194 736 95236 776
rect 95276 736 95318 776
rect 95358 736 95400 776
rect 95440 736 99360 776
rect 576 712 99360 736
<< via1 >>
rect 3112 81628 3152 81668
rect 3194 81628 3234 81668
rect 3276 81628 3316 81668
rect 3358 81628 3398 81668
rect 3440 81628 3480 81668
rect 18232 81628 18272 81668
rect 18314 81628 18354 81668
rect 18396 81628 18436 81668
rect 18478 81628 18518 81668
rect 18560 81628 18600 81668
rect 33352 81628 33392 81668
rect 33434 81628 33474 81668
rect 33516 81628 33556 81668
rect 33598 81628 33638 81668
rect 33680 81628 33720 81668
rect 48472 81628 48512 81668
rect 48554 81628 48594 81668
rect 48636 81628 48676 81668
rect 48718 81628 48758 81668
rect 48800 81628 48840 81668
rect 63592 81628 63632 81668
rect 63674 81628 63714 81668
rect 63756 81628 63796 81668
rect 63838 81628 63878 81668
rect 63920 81628 63960 81668
rect 78712 81628 78752 81668
rect 78794 81628 78834 81668
rect 78876 81628 78916 81668
rect 78958 81628 78998 81668
rect 79040 81628 79080 81668
rect 93832 81628 93872 81668
rect 93914 81628 93954 81668
rect 93996 81628 94036 81668
rect 94078 81628 94118 81668
rect 94160 81628 94200 81668
rect 4352 80872 4392 80912
rect 4434 80872 4474 80912
rect 4516 80872 4556 80912
rect 4598 80872 4638 80912
rect 4680 80872 4720 80912
rect 19472 80872 19512 80912
rect 19554 80872 19594 80912
rect 19636 80872 19676 80912
rect 19718 80872 19758 80912
rect 19800 80872 19840 80912
rect 34592 80872 34632 80912
rect 34674 80872 34714 80912
rect 34756 80872 34796 80912
rect 34838 80872 34878 80912
rect 34920 80872 34960 80912
rect 49712 80872 49752 80912
rect 49794 80872 49834 80912
rect 49876 80872 49916 80912
rect 49958 80872 49998 80912
rect 50040 80872 50080 80912
rect 64832 80872 64872 80912
rect 64914 80872 64954 80912
rect 64996 80872 65036 80912
rect 65078 80872 65118 80912
rect 65160 80872 65200 80912
rect 79952 80872 79992 80912
rect 80034 80872 80074 80912
rect 80116 80872 80156 80912
rect 80198 80872 80238 80912
rect 80280 80872 80320 80912
rect 95072 80872 95112 80912
rect 95154 80872 95194 80912
rect 95236 80872 95276 80912
rect 95318 80872 95358 80912
rect 95400 80872 95440 80912
rect 3112 80116 3152 80156
rect 3194 80116 3234 80156
rect 3276 80116 3316 80156
rect 3358 80116 3398 80156
rect 3440 80116 3480 80156
rect 18232 80116 18272 80156
rect 18314 80116 18354 80156
rect 18396 80116 18436 80156
rect 18478 80116 18518 80156
rect 18560 80116 18600 80156
rect 33352 80116 33392 80156
rect 33434 80116 33474 80156
rect 33516 80116 33556 80156
rect 33598 80116 33638 80156
rect 33680 80116 33720 80156
rect 48472 80116 48512 80156
rect 48554 80116 48594 80156
rect 48636 80116 48676 80156
rect 48718 80116 48758 80156
rect 48800 80116 48840 80156
rect 63592 80116 63632 80156
rect 63674 80116 63714 80156
rect 63756 80116 63796 80156
rect 63838 80116 63878 80156
rect 63920 80116 63960 80156
rect 78712 80116 78752 80156
rect 78794 80116 78834 80156
rect 78876 80116 78916 80156
rect 78958 80116 78998 80156
rect 79040 80116 79080 80156
rect 93832 80116 93872 80156
rect 93914 80116 93954 80156
rect 93996 80116 94036 80156
rect 94078 80116 94118 80156
rect 94160 80116 94200 80156
rect 4352 79360 4392 79400
rect 4434 79360 4474 79400
rect 4516 79360 4556 79400
rect 4598 79360 4638 79400
rect 4680 79360 4720 79400
rect 19472 79360 19512 79400
rect 19554 79360 19594 79400
rect 19636 79360 19676 79400
rect 19718 79360 19758 79400
rect 19800 79360 19840 79400
rect 34592 79360 34632 79400
rect 34674 79360 34714 79400
rect 34756 79360 34796 79400
rect 34838 79360 34878 79400
rect 34920 79360 34960 79400
rect 49712 79360 49752 79400
rect 49794 79360 49834 79400
rect 49876 79360 49916 79400
rect 49958 79360 49998 79400
rect 50040 79360 50080 79400
rect 64832 79360 64872 79400
rect 64914 79360 64954 79400
rect 64996 79360 65036 79400
rect 65078 79360 65118 79400
rect 65160 79360 65200 79400
rect 79952 79360 79992 79400
rect 80034 79360 80074 79400
rect 80116 79360 80156 79400
rect 80198 79360 80238 79400
rect 80280 79360 80320 79400
rect 95072 79360 95112 79400
rect 95154 79360 95194 79400
rect 95236 79360 95276 79400
rect 95318 79360 95358 79400
rect 95400 79360 95440 79400
rect 3112 78604 3152 78644
rect 3194 78604 3234 78644
rect 3276 78604 3316 78644
rect 3358 78604 3398 78644
rect 3440 78604 3480 78644
rect 18232 78604 18272 78644
rect 18314 78604 18354 78644
rect 18396 78604 18436 78644
rect 18478 78604 18518 78644
rect 18560 78604 18600 78644
rect 33352 78604 33392 78644
rect 33434 78604 33474 78644
rect 33516 78604 33556 78644
rect 33598 78604 33638 78644
rect 33680 78604 33720 78644
rect 48472 78604 48512 78644
rect 48554 78604 48594 78644
rect 48636 78604 48676 78644
rect 48718 78604 48758 78644
rect 48800 78604 48840 78644
rect 63592 78604 63632 78644
rect 63674 78604 63714 78644
rect 63756 78604 63796 78644
rect 63838 78604 63878 78644
rect 63920 78604 63960 78644
rect 78712 78604 78752 78644
rect 78794 78604 78834 78644
rect 78876 78604 78916 78644
rect 78958 78604 78998 78644
rect 79040 78604 79080 78644
rect 93832 78604 93872 78644
rect 93914 78604 93954 78644
rect 93996 78604 94036 78644
rect 94078 78604 94118 78644
rect 94160 78604 94200 78644
rect 4352 77848 4392 77888
rect 4434 77848 4474 77888
rect 4516 77848 4556 77888
rect 4598 77848 4638 77888
rect 4680 77848 4720 77888
rect 19472 77848 19512 77888
rect 19554 77848 19594 77888
rect 19636 77848 19676 77888
rect 19718 77848 19758 77888
rect 19800 77848 19840 77888
rect 34592 77848 34632 77888
rect 34674 77848 34714 77888
rect 34756 77848 34796 77888
rect 34838 77848 34878 77888
rect 34920 77848 34960 77888
rect 49712 77848 49752 77888
rect 49794 77848 49834 77888
rect 49876 77848 49916 77888
rect 49958 77848 49998 77888
rect 50040 77848 50080 77888
rect 64832 77848 64872 77888
rect 64914 77848 64954 77888
rect 64996 77848 65036 77888
rect 65078 77848 65118 77888
rect 65160 77848 65200 77888
rect 79952 77848 79992 77888
rect 80034 77848 80074 77888
rect 80116 77848 80156 77888
rect 80198 77848 80238 77888
rect 80280 77848 80320 77888
rect 95072 77848 95112 77888
rect 95154 77848 95194 77888
rect 95236 77848 95276 77888
rect 95318 77848 95358 77888
rect 95400 77848 95440 77888
rect 3112 77092 3152 77132
rect 3194 77092 3234 77132
rect 3276 77092 3316 77132
rect 3358 77092 3398 77132
rect 3440 77092 3480 77132
rect 18232 77092 18272 77132
rect 18314 77092 18354 77132
rect 18396 77092 18436 77132
rect 18478 77092 18518 77132
rect 18560 77092 18600 77132
rect 33352 77092 33392 77132
rect 33434 77092 33474 77132
rect 33516 77092 33556 77132
rect 33598 77092 33638 77132
rect 33680 77092 33720 77132
rect 48472 77092 48512 77132
rect 48554 77092 48594 77132
rect 48636 77092 48676 77132
rect 48718 77092 48758 77132
rect 48800 77092 48840 77132
rect 63592 77092 63632 77132
rect 63674 77092 63714 77132
rect 63756 77092 63796 77132
rect 63838 77092 63878 77132
rect 63920 77092 63960 77132
rect 78712 77092 78752 77132
rect 78794 77092 78834 77132
rect 78876 77092 78916 77132
rect 78958 77092 78998 77132
rect 79040 77092 79080 77132
rect 93832 77092 93872 77132
rect 93914 77092 93954 77132
rect 93996 77092 94036 77132
rect 94078 77092 94118 77132
rect 94160 77092 94200 77132
rect 4352 76336 4392 76376
rect 4434 76336 4474 76376
rect 4516 76336 4556 76376
rect 4598 76336 4638 76376
rect 4680 76336 4720 76376
rect 19472 76336 19512 76376
rect 19554 76336 19594 76376
rect 19636 76336 19676 76376
rect 19718 76336 19758 76376
rect 19800 76336 19840 76376
rect 34592 76336 34632 76376
rect 34674 76336 34714 76376
rect 34756 76336 34796 76376
rect 34838 76336 34878 76376
rect 34920 76336 34960 76376
rect 49712 76336 49752 76376
rect 49794 76336 49834 76376
rect 49876 76336 49916 76376
rect 49958 76336 49998 76376
rect 50040 76336 50080 76376
rect 64832 76336 64872 76376
rect 64914 76336 64954 76376
rect 64996 76336 65036 76376
rect 65078 76336 65118 76376
rect 65160 76336 65200 76376
rect 79952 76336 79992 76376
rect 80034 76336 80074 76376
rect 80116 76336 80156 76376
rect 80198 76336 80238 76376
rect 80280 76336 80320 76376
rect 95072 76336 95112 76376
rect 95154 76336 95194 76376
rect 95236 76336 95276 76376
rect 95318 76336 95358 76376
rect 95400 76336 95440 76376
rect 3112 75580 3152 75620
rect 3194 75580 3234 75620
rect 3276 75580 3316 75620
rect 3358 75580 3398 75620
rect 3440 75580 3480 75620
rect 18232 75580 18272 75620
rect 18314 75580 18354 75620
rect 18396 75580 18436 75620
rect 18478 75580 18518 75620
rect 18560 75580 18600 75620
rect 33352 75580 33392 75620
rect 33434 75580 33474 75620
rect 33516 75580 33556 75620
rect 33598 75580 33638 75620
rect 33680 75580 33720 75620
rect 48472 75580 48512 75620
rect 48554 75580 48594 75620
rect 48636 75580 48676 75620
rect 48718 75580 48758 75620
rect 48800 75580 48840 75620
rect 63592 75580 63632 75620
rect 63674 75580 63714 75620
rect 63756 75580 63796 75620
rect 63838 75580 63878 75620
rect 63920 75580 63960 75620
rect 78712 75580 78752 75620
rect 78794 75580 78834 75620
rect 78876 75580 78916 75620
rect 78958 75580 78998 75620
rect 79040 75580 79080 75620
rect 93832 75580 93872 75620
rect 93914 75580 93954 75620
rect 93996 75580 94036 75620
rect 94078 75580 94118 75620
rect 94160 75580 94200 75620
rect 652 75244 692 75284
rect 844 74992 884 75032
rect 4352 74824 4392 74864
rect 4434 74824 4474 74864
rect 4516 74824 4556 74864
rect 4598 74824 4638 74864
rect 4680 74824 4720 74864
rect 19472 74824 19512 74864
rect 19554 74824 19594 74864
rect 19636 74824 19676 74864
rect 19718 74824 19758 74864
rect 19800 74824 19840 74864
rect 34592 74824 34632 74864
rect 34674 74824 34714 74864
rect 34756 74824 34796 74864
rect 34838 74824 34878 74864
rect 34920 74824 34960 74864
rect 49712 74824 49752 74864
rect 49794 74824 49834 74864
rect 49876 74824 49916 74864
rect 49958 74824 49998 74864
rect 50040 74824 50080 74864
rect 64832 74824 64872 74864
rect 64914 74824 64954 74864
rect 64996 74824 65036 74864
rect 65078 74824 65118 74864
rect 65160 74824 65200 74864
rect 79952 74824 79992 74864
rect 80034 74824 80074 74864
rect 80116 74824 80156 74864
rect 80198 74824 80238 74864
rect 80280 74824 80320 74864
rect 95072 74824 95112 74864
rect 95154 74824 95194 74864
rect 95236 74824 95276 74864
rect 95318 74824 95358 74864
rect 95400 74824 95440 74864
rect 3112 74068 3152 74108
rect 3194 74068 3234 74108
rect 3276 74068 3316 74108
rect 3358 74068 3398 74108
rect 3440 74068 3480 74108
rect 18232 74068 18272 74108
rect 18314 74068 18354 74108
rect 18396 74068 18436 74108
rect 18478 74068 18518 74108
rect 18560 74068 18600 74108
rect 33352 74068 33392 74108
rect 33434 74068 33474 74108
rect 33516 74068 33556 74108
rect 33598 74068 33638 74108
rect 33680 74068 33720 74108
rect 48472 74068 48512 74108
rect 48554 74068 48594 74108
rect 48636 74068 48676 74108
rect 48718 74068 48758 74108
rect 48800 74068 48840 74108
rect 63592 74068 63632 74108
rect 63674 74068 63714 74108
rect 63756 74068 63796 74108
rect 63838 74068 63878 74108
rect 63920 74068 63960 74108
rect 78712 74068 78752 74108
rect 78794 74068 78834 74108
rect 78876 74068 78916 74108
rect 78958 74068 78998 74108
rect 79040 74068 79080 74108
rect 93832 74068 93872 74108
rect 93914 74068 93954 74108
rect 93996 74068 94036 74108
rect 94078 74068 94118 74108
rect 94160 74068 94200 74108
rect 4352 73312 4392 73352
rect 4434 73312 4474 73352
rect 4516 73312 4556 73352
rect 4598 73312 4638 73352
rect 4680 73312 4720 73352
rect 19472 73312 19512 73352
rect 19554 73312 19594 73352
rect 19636 73312 19676 73352
rect 19718 73312 19758 73352
rect 19800 73312 19840 73352
rect 34592 73312 34632 73352
rect 34674 73312 34714 73352
rect 34756 73312 34796 73352
rect 34838 73312 34878 73352
rect 34920 73312 34960 73352
rect 49712 73312 49752 73352
rect 49794 73312 49834 73352
rect 49876 73312 49916 73352
rect 49958 73312 49998 73352
rect 50040 73312 50080 73352
rect 64832 73312 64872 73352
rect 64914 73312 64954 73352
rect 64996 73312 65036 73352
rect 65078 73312 65118 73352
rect 65160 73312 65200 73352
rect 79952 73312 79992 73352
rect 80034 73312 80074 73352
rect 80116 73312 80156 73352
rect 80198 73312 80238 73352
rect 80280 73312 80320 73352
rect 95072 73312 95112 73352
rect 95154 73312 95194 73352
rect 95236 73312 95276 73352
rect 95318 73312 95358 73352
rect 95400 73312 95440 73352
rect 652 72892 692 72932
rect 844 72724 884 72764
rect 3112 72556 3152 72596
rect 3194 72556 3234 72596
rect 3276 72556 3316 72596
rect 3358 72556 3398 72596
rect 3440 72556 3480 72596
rect 18232 72556 18272 72596
rect 18314 72556 18354 72596
rect 18396 72556 18436 72596
rect 18478 72556 18518 72596
rect 18560 72556 18600 72596
rect 33352 72556 33392 72596
rect 33434 72556 33474 72596
rect 33516 72556 33556 72596
rect 33598 72556 33638 72596
rect 33680 72556 33720 72596
rect 48472 72556 48512 72596
rect 48554 72556 48594 72596
rect 48636 72556 48676 72596
rect 48718 72556 48758 72596
rect 48800 72556 48840 72596
rect 63592 72556 63632 72596
rect 63674 72556 63714 72596
rect 63756 72556 63796 72596
rect 63838 72556 63878 72596
rect 63920 72556 63960 72596
rect 78712 72556 78752 72596
rect 78794 72556 78834 72596
rect 78876 72556 78916 72596
rect 78958 72556 78998 72596
rect 79040 72556 79080 72596
rect 93832 72556 93872 72596
rect 93914 72556 93954 72596
rect 93996 72556 94036 72596
rect 94078 72556 94118 72596
rect 94160 72556 94200 72596
rect 4352 71800 4392 71840
rect 4434 71800 4474 71840
rect 4516 71800 4556 71840
rect 4598 71800 4638 71840
rect 4680 71800 4720 71840
rect 19472 71800 19512 71840
rect 19554 71800 19594 71840
rect 19636 71800 19676 71840
rect 19718 71800 19758 71840
rect 19800 71800 19840 71840
rect 34592 71800 34632 71840
rect 34674 71800 34714 71840
rect 34756 71800 34796 71840
rect 34838 71800 34878 71840
rect 34920 71800 34960 71840
rect 49712 71800 49752 71840
rect 49794 71800 49834 71840
rect 49876 71800 49916 71840
rect 49958 71800 49998 71840
rect 50040 71800 50080 71840
rect 64832 71800 64872 71840
rect 64914 71800 64954 71840
rect 64996 71800 65036 71840
rect 65078 71800 65118 71840
rect 65160 71800 65200 71840
rect 79952 71800 79992 71840
rect 80034 71800 80074 71840
rect 80116 71800 80156 71840
rect 80198 71800 80238 71840
rect 80280 71800 80320 71840
rect 95072 71800 95112 71840
rect 95154 71800 95194 71840
rect 95236 71800 95276 71840
rect 95318 71800 95358 71840
rect 95400 71800 95440 71840
rect 652 71464 692 71504
rect 844 71464 884 71504
rect 3112 71044 3152 71084
rect 3194 71044 3234 71084
rect 3276 71044 3316 71084
rect 3358 71044 3398 71084
rect 3440 71044 3480 71084
rect 18232 71044 18272 71084
rect 18314 71044 18354 71084
rect 18396 71044 18436 71084
rect 18478 71044 18518 71084
rect 18560 71044 18600 71084
rect 33352 71044 33392 71084
rect 33434 71044 33474 71084
rect 33516 71044 33556 71084
rect 33598 71044 33638 71084
rect 33680 71044 33720 71084
rect 48472 71044 48512 71084
rect 48554 71044 48594 71084
rect 48636 71044 48676 71084
rect 48718 71044 48758 71084
rect 48800 71044 48840 71084
rect 63592 71044 63632 71084
rect 63674 71044 63714 71084
rect 63756 71044 63796 71084
rect 63838 71044 63878 71084
rect 63920 71044 63960 71084
rect 78712 71044 78752 71084
rect 78794 71044 78834 71084
rect 78876 71044 78916 71084
rect 78958 71044 78998 71084
rect 79040 71044 79080 71084
rect 93832 71044 93872 71084
rect 93914 71044 93954 71084
rect 93996 71044 94036 71084
rect 94078 71044 94118 71084
rect 94160 71044 94200 71084
rect 4352 70288 4392 70328
rect 4434 70288 4474 70328
rect 4516 70288 4556 70328
rect 4598 70288 4638 70328
rect 4680 70288 4720 70328
rect 19472 70288 19512 70328
rect 19554 70288 19594 70328
rect 19636 70288 19676 70328
rect 19718 70288 19758 70328
rect 19800 70288 19840 70328
rect 34592 70288 34632 70328
rect 34674 70288 34714 70328
rect 34756 70288 34796 70328
rect 34838 70288 34878 70328
rect 34920 70288 34960 70328
rect 49712 70288 49752 70328
rect 49794 70288 49834 70328
rect 49876 70288 49916 70328
rect 49958 70288 49998 70328
rect 50040 70288 50080 70328
rect 64832 70288 64872 70328
rect 64914 70288 64954 70328
rect 64996 70288 65036 70328
rect 65078 70288 65118 70328
rect 65160 70288 65200 70328
rect 79952 70288 79992 70328
rect 80034 70288 80074 70328
rect 80116 70288 80156 70328
rect 80198 70288 80238 70328
rect 80280 70288 80320 70328
rect 95072 70288 95112 70328
rect 95154 70288 95194 70328
rect 95236 70288 95276 70328
rect 95318 70288 95358 70328
rect 95400 70288 95440 70328
rect 3112 69532 3152 69572
rect 3194 69532 3234 69572
rect 3276 69532 3316 69572
rect 3358 69532 3398 69572
rect 3440 69532 3480 69572
rect 18232 69532 18272 69572
rect 18314 69532 18354 69572
rect 18396 69532 18436 69572
rect 18478 69532 18518 69572
rect 18560 69532 18600 69572
rect 33352 69532 33392 69572
rect 33434 69532 33474 69572
rect 33516 69532 33556 69572
rect 33598 69532 33638 69572
rect 33680 69532 33720 69572
rect 48472 69532 48512 69572
rect 48554 69532 48594 69572
rect 48636 69532 48676 69572
rect 48718 69532 48758 69572
rect 48800 69532 48840 69572
rect 63592 69532 63632 69572
rect 63674 69532 63714 69572
rect 63756 69532 63796 69572
rect 63838 69532 63878 69572
rect 63920 69532 63960 69572
rect 78712 69532 78752 69572
rect 78794 69532 78834 69572
rect 78876 69532 78916 69572
rect 78958 69532 78998 69572
rect 79040 69532 79080 69572
rect 93832 69532 93872 69572
rect 93914 69532 93954 69572
rect 93996 69532 94036 69572
rect 94078 69532 94118 69572
rect 94160 69532 94200 69572
rect 652 69196 692 69236
rect 844 68944 884 68984
rect 4352 68776 4392 68816
rect 4434 68776 4474 68816
rect 4516 68776 4556 68816
rect 4598 68776 4638 68816
rect 4680 68776 4720 68816
rect 19472 68776 19512 68816
rect 19554 68776 19594 68816
rect 19636 68776 19676 68816
rect 19718 68776 19758 68816
rect 19800 68776 19840 68816
rect 34592 68776 34632 68816
rect 34674 68776 34714 68816
rect 34756 68776 34796 68816
rect 34838 68776 34878 68816
rect 34920 68776 34960 68816
rect 49712 68776 49752 68816
rect 49794 68776 49834 68816
rect 49876 68776 49916 68816
rect 49958 68776 49998 68816
rect 50040 68776 50080 68816
rect 64832 68776 64872 68816
rect 64914 68776 64954 68816
rect 64996 68776 65036 68816
rect 65078 68776 65118 68816
rect 65160 68776 65200 68816
rect 79952 68776 79992 68816
rect 80034 68776 80074 68816
rect 80116 68776 80156 68816
rect 80198 68776 80238 68816
rect 80280 68776 80320 68816
rect 95072 68776 95112 68816
rect 95154 68776 95194 68816
rect 95236 68776 95276 68816
rect 95318 68776 95358 68816
rect 95400 68776 95440 68816
rect 3112 68020 3152 68060
rect 3194 68020 3234 68060
rect 3276 68020 3316 68060
rect 3358 68020 3398 68060
rect 3440 68020 3480 68060
rect 18232 68020 18272 68060
rect 18314 68020 18354 68060
rect 18396 68020 18436 68060
rect 18478 68020 18518 68060
rect 18560 68020 18600 68060
rect 33352 68020 33392 68060
rect 33434 68020 33474 68060
rect 33516 68020 33556 68060
rect 33598 68020 33638 68060
rect 33680 68020 33720 68060
rect 48472 68020 48512 68060
rect 48554 68020 48594 68060
rect 48636 68020 48676 68060
rect 48718 68020 48758 68060
rect 48800 68020 48840 68060
rect 63592 68020 63632 68060
rect 63674 68020 63714 68060
rect 63756 68020 63796 68060
rect 63838 68020 63878 68060
rect 63920 68020 63960 68060
rect 78712 68020 78752 68060
rect 78794 68020 78834 68060
rect 78876 68020 78916 68060
rect 78958 68020 78998 68060
rect 79040 68020 79080 68060
rect 93832 68020 93872 68060
rect 93914 68020 93954 68060
rect 93996 68020 94036 68060
rect 94078 68020 94118 68060
rect 94160 68020 94200 68060
rect 652 67684 692 67724
rect 844 67432 884 67472
rect 4352 67264 4392 67304
rect 4434 67264 4474 67304
rect 4516 67264 4556 67304
rect 4598 67264 4638 67304
rect 4680 67264 4720 67304
rect 19472 67264 19512 67304
rect 19554 67264 19594 67304
rect 19636 67264 19676 67304
rect 19718 67264 19758 67304
rect 19800 67264 19840 67304
rect 34592 67264 34632 67304
rect 34674 67264 34714 67304
rect 34756 67264 34796 67304
rect 34838 67264 34878 67304
rect 34920 67264 34960 67304
rect 49712 67264 49752 67304
rect 49794 67264 49834 67304
rect 49876 67264 49916 67304
rect 49958 67264 49998 67304
rect 50040 67264 50080 67304
rect 64832 67264 64872 67304
rect 64914 67264 64954 67304
rect 64996 67264 65036 67304
rect 65078 67264 65118 67304
rect 65160 67264 65200 67304
rect 79952 67264 79992 67304
rect 80034 67264 80074 67304
rect 80116 67264 80156 67304
rect 80198 67264 80238 67304
rect 80280 67264 80320 67304
rect 95072 67264 95112 67304
rect 95154 67264 95194 67304
rect 95236 67264 95276 67304
rect 95318 67264 95358 67304
rect 95400 67264 95440 67304
rect 3112 66508 3152 66548
rect 3194 66508 3234 66548
rect 3276 66508 3316 66548
rect 3358 66508 3398 66548
rect 3440 66508 3480 66548
rect 18232 66508 18272 66548
rect 18314 66508 18354 66548
rect 18396 66508 18436 66548
rect 18478 66508 18518 66548
rect 18560 66508 18600 66548
rect 33352 66508 33392 66548
rect 33434 66508 33474 66548
rect 33516 66508 33556 66548
rect 33598 66508 33638 66548
rect 33680 66508 33720 66548
rect 48472 66508 48512 66548
rect 48554 66508 48594 66548
rect 48636 66508 48676 66548
rect 48718 66508 48758 66548
rect 48800 66508 48840 66548
rect 63592 66508 63632 66548
rect 63674 66508 63714 66548
rect 63756 66508 63796 66548
rect 63838 66508 63878 66548
rect 63920 66508 63960 66548
rect 78712 66508 78752 66548
rect 78794 66508 78834 66548
rect 78876 66508 78916 66548
rect 78958 66508 78998 66548
rect 79040 66508 79080 66548
rect 93832 66508 93872 66548
rect 93914 66508 93954 66548
rect 93996 66508 94036 66548
rect 94078 66508 94118 66548
rect 94160 66508 94200 66548
rect 652 66172 692 66212
rect 844 65920 884 65960
rect 4352 65752 4392 65792
rect 4434 65752 4474 65792
rect 4516 65752 4556 65792
rect 4598 65752 4638 65792
rect 4680 65752 4720 65792
rect 19472 65752 19512 65792
rect 19554 65752 19594 65792
rect 19636 65752 19676 65792
rect 19718 65752 19758 65792
rect 19800 65752 19840 65792
rect 34592 65752 34632 65792
rect 34674 65752 34714 65792
rect 34756 65752 34796 65792
rect 34838 65752 34878 65792
rect 34920 65752 34960 65792
rect 49712 65752 49752 65792
rect 49794 65752 49834 65792
rect 49876 65752 49916 65792
rect 49958 65752 49998 65792
rect 50040 65752 50080 65792
rect 64832 65752 64872 65792
rect 64914 65752 64954 65792
rect 64996 65752 65036 65792
rect 65078 65752 65118 65792
rect 65160 65752 65200 65792
rect 79952 65752 79992 65792
rect 80034 65752 80074 65792
rect 80116 65752 80156 65792
rect 80198 65752 80238 65792
rect 80280 65752 80320 65792
rect 95072 65752 95112 65792
rect 95154 65752 95194 65792
rect 95236 65752 95276 65792
rect 95318 65752 95358 65792
rect 95400 65752 95440 65792
rect 3112 64996 3152 65036
rect 3194 64996 3234 65036
rect 3276 64996 3316 65036
rect 3358 64996 3398 65036
rect 3440 64996 3480 65036
rect 18232 64996 18272 65036
rect 18314 64996 18354 65036
rect 18396 64996 18436 65036
rect 18478 64996 18518 65036
rect 18560 64996 18600 65036
rect 33352 64996 33392 65036
rect 33434 64996 33474 65036
rect 33516 64996 33556 65036
rect 33598 64996 33638 65036
rect 33680 64996 33720 65036
rect 48472 64996 48512 65036
rect 48554 64996 48594 65036
rect 48636 64996 48676 65036
rect 48718 64996 48758 65036
rect 48800 64996 48840 65036
rect 63592 64996 63632 65036
rect 63674 64996 63714 65036
rect 63756 64996 63796 65036
rect 63838 64996 63878 65036
rect 63920 64996 63960 65036
rect 78712 64996 78752 65036
rect 78794 64996 78834 65036
rect 78876 64996 78916 65036
rect 78958 64996 78998 65036
rect 79040 64996 79080 65036
rect 93832 64996 93872 65036
rect 93914 64996 93954 65036
rect 93996 64996 94036 65036
rect 94078 64996 94118 65036
rect 94160 64996 94200 65036
rect 4352 64240 4392 64280
rect 4434 64240 4474 64280
rect 4516 64240 4556 64280
rect 4598 64240 4638 64280
rect 4680 64240 4720 64280
rect 19472 64240 19512 64280
rect 19554 64240 19594 64280
rect 19636 64240 19676 64280
rect 19718 64240 19758 64280
rect 19800 64240 19840 64280
rect 34592 64240 34632 64280
rect 34674 64240 34714 64280
rect 34756 64240 34796 64280
rect 34838 64240 34878 64280
rect 34920 64240 34960 64280
rect 49712 64240 49752 64280
rect 49794 64240 49834 64280
rect 49876 64240 49916 64280
rect 49958 64240 49998 64280
rect 50040 64240 50080 64280
rect 64832 64240 64872 64280
rect 64914 64240 64954 64280
rect 64996 64240 65036 64280
rect 65078 64240 65118 64280
rect 65160 64240 65200 64280
rect 79952 64240 79992 64280
rect 80034 64240 80074 64280
rect 80116 64240 80156 64280
rect 80198 64240 80238 64280
rect 80280 64240 80320 64280
rect 95072 64240 95112 64280
rect 95154 64240 95194 64280
rect 95236 64240 95276 64280
rect 95318 64240 95358 64280
rect 95400 64240 95440 64280
rect 652 63820 692 63860
rect 844 63652 884 63692
rect 3112 63484 3152 63524
rect 3194 63484 3234 63524
rect 3276 63484 3316 63524
rect 3358 63484 3398 63524
rect 3440 63484 3480 63524
rect 18232 63484 18272 63524
rect 18314 63484 18354 63524
rect 18396 63484 18436 63524
rect 18478 63484 18518 63524
rect 18560 63484 18600 63524
rect 33352 63484 33392 63524
rect 33434 63484 33474 63524
rect 33516 63484 33556 63524
rect 33598 63484 33638 63524
rect 33680 63484 33720 63524
rect 48472 63484 48512 63524
rect 48554 63484 48594 63524
rect 48636 63484 48676 63524
rect 48718 63484 48758 63524
rect 48800 63484 48840 63524
rect 63592 63484 63632 63524
rect 63674 63484 63714 63524
rect 63756 63484 63796 63524
rect 63838 63484 63878 63524
rect 63920 63484 63960 63524
rect 78712 63484 78752 63524
rect 78794 63484 78834 63524
rect 78876 63484 78916 63524
rect 78958 63484 78998 63524
rect 79040 63484 79080 63524
rect 93832 63484 93872 63524
rect 93914 63484 93954 63524
rect 93996 63484 94036 63524
rect 94078 63484 94118 63524
rect 94160 63484 94200 63524
rect 4352 62728 4392 62768
rect 4434 62728 4474 62768
rect 4516 62728 4556 62768
rect 4598 62728 4638 62768
rect 4680 62728 4720 62768
rect 19472 62728 19512 62768
rect 19554 62728 19594 62768
rect 19636 62728 19676 62768
rect 19718 62728 19758 62768
rect 19800 62728 19840 62768
rect 34592 62728 34632 62768
rect 34674 62728 34714 62768
rect 34756 62728 34796 62768
rect 34838 62728 34878 62768
rect 34920 62728 34960 62768
rect 49712 62728 49752 62768
rect 49794 62728 49834 62768
rect 49876 62728 49916 62768
rect 49958 62728 49998 62768
rect 50040 62728 50080 62768
rect 64832 62728 64872 62768
rect 64914 62728 64954 62768
rect 64996 62728 65036 62768
rect 65078 62728 65118 62768
rect 65160 62728 65200 62768
rect 79952 62728 79992 62768
rect 80034 62728 80074 62768
rect 80116 62728 80156 62768
rect 80198 62728 80238 62768
rect 80280 62728 80320 62768
rect 95072 62728 95112 62768
rect 95154 62728 95194 62768
rect 95236 62728 95276 62768
rect 95318 62728 95358 62768
rect 95400 62728 95440 62768
rect 652 62308 692 62348
rect 844 62140 884 62180
rect 3112 61972 3152 62012
rect 3194 61972 3234 62012
rect 3276 61972 3316 62012
rect 3358 61972 3398 62012
rect 3440 61972 3480 62012
rect 18232 61972 18272 62012
rect 18314 61972 18354 62012
rect 18396 61972 18436 62012
rect 18478 61972 18518 62012
rect 18560 61972 18600 62012
rect 33352 61972 33392 62012
rect 33434 61972 33474 62012
rect 33516 61972 33556 62012
rect 33598 61972 33638 62012
rect 33680 61972 33720 62012
rect 48472 61972 48512 62012
rect 48554 61972 48594 62012
rect 48636 61972 48676 62012
rect 48718 61972 48758 62012
rect 48800 61972 48840 62012
rect 63592 61972 63632 62012
rect 63674 61972 63714 62012
rect 63756 61972 63796 62012
rect 63838 61972 63878 62012
rect 63920 61972 63960 62012
rect 78712 61972 78752 62012
rect 78794 61972 78834 62012
rect 78876 61972 78916 62012
rect 78958 61972 78998 62012
rect 79040 61972 79080 62012
rect 93832 61972 93872 62012
rect 93914 61972 93954 62012
rect 93996 61972 94036 62012
rect 94078 61972 94118 62012
rect 94160 61972 94200 62012
rect 4352 61216 4392 61256
rect 4434 61216 4474 61256
rect 4516 61216 4556 61256
rect 4598 61216 4638 61256
rect 4680 61216 4720 61256
rect 19472 61216 19512 61256
rect 19554 61216 19594 61256
rect 19636 61216 19676 61256
rect 19718 61216 19758 61256
rect 19800 61216 19840 61256
rect 34592 61216 34632 61256
rect 34674 61216 34714 61256
rect 34756 61216 34796 61256
rect 34838 61216 34878 61256
rect 34920 61216 34960 61256
rect 49712 61216 49752 61256
rect 49794 61216 49834 61256
rect 49876 61216 49916 61256
rect 49958 61216 49998 61256
rect 50040 61216 50080 61256
rect 64832 61216 64872 61256
rect 64914 61216 64954 61256
rect 64996 61216 65036 61256
rect 65078 61216 65118 61256
rect 65160 61216 65200 61256
rect 79952 61216 79992 61256
rect 80034 61216 80074 61256
rect 80116 61216 80156 61256
rect 80198 61216 80238 61256
rect 80280 61216 80320 61256
rect 95072 61216 95112 61256
rect 95154 61216 95194 61256
rect 95236 61216 95276 61256
rect 95318 61216 95358 61256
rect 95400 61216 95440 61256
rect 6508 60880 6548 60920
rect 6604 60880 6644 60920
rect 6892 60796 6932 60836
rect 3112 60460 3152 60500
rect 3194 60460 3234 60500
rect 3276 60460 3316 60500
rect 3358 60460 3398 60500
rect 3440 60460 3480 60500
rect 18232 60460 18272 60500
rect 18314 60460 18354 60500
rect 18396 60460 18436 60500
rect 18478 60460 18518 60500
rect 18560 60460 18600 60500
rect 33352 60460 33392 60500
rect 33434 60460 33474 60500
rect 33516 60460 33556 60500
rect 33598 60460 33638 60500
rect 33680 60460 33720 60500
rect 48472 60460 48512 60500
rect 48554 60460 48594 60500
rect 48636 60460 48676 60500
rect 48718 60460 48758 60500
rect 48800 60460 48840 60500
rect 63592 60460 63632 60500
rect 63674 60460 63714 60500
rect 63756 60460 63796 60500
rect 63838 60460 63878 60500
rect 63920 60460 63960 60500
rect 78712 60460 78752 60500
rect 78794 60460 78834 60500
rect 78876 60460 78916 60500
rect 78958 60460 78998 60500
rect 79040 60460 79080 60500
rect 93832 60460 93872 60500
rect 93914 60460 93954 60500
rect 93996 60460 94036 60500
rect 94078 60460 94118 60500
rect 94160 60460 94200 60500
rect 844 60292 884 60332
rect 652 60124 692 60164
rect 6796 60040 6836 60080
rect 6892 60040 6932 60080
rect 6508 59872 6548 59912
rect 4352 59704 4392 59744
rect 4434 59704 4474 59744
rect 4516 59704 4556 59744
rect 4598 59704 4638 59744
rect 4680 59704 4720 59744
rect 19472 59704 19512 59744
rect 19554 59704 19594 59744
rect 19636 59704 19676 59744
rect 19718 59704 19758 59744
rect 19800 59704 19840 59744
rect 34592 59704 34632 59744
rect 34674 59704 34714 59744
rect 34756 59704 34796 59744
rect 34838 59704 34878 59744
rect 34920 59704 34960 59744
rect 49712 59704 49752 59744
rect 49794 59704 49834 59744
rect 49876 59704 49916 59744
rect 49958 59704 49998 59744
rect 50040 59704 50080 59744
rect 64832 59704 64872 59744
rect 64914 59704 64954 59744
rect 64996 59704 65036 59744
rect 65078 59704 65118 59744
rect 65160 59704 65200 59744
rect 79952 59704 79992 59744
rect 80034 59704 80074 59744
rect 80116 59704 80156 59744
rect 80198 59704 80238 59744
rect 80280 59704 80320 59744
rect 95072 59704 95112 59744
rect 95154 59704 95194 59744
rect 95236 59704 95276 59744
rect 95318 59704 95358 59744
rect 95400 59704 95440 59744
rect 3112 58948 3152 58988
rect 3194 58948 3234 58988
rect 3276 58948 3316 58988
rect 3358 58948 3398 58988
rect 3440 58948 3480 58988
rect 18232 58948 18272 58988
rect 18314 58948 18354 58988
rect 18396 58948 18436 58988
rect 18478 58948 18518 58988
rect 18560 58948 18600 58988
rect 33352 58948 33392 58988
rect 33434 58948 33474 58988
rect 33516 58948 33556 58988
rect 33598 58948 33638 58988
rect 33680 58948 33720 58988
rect 48472 58948 48512 58988
rect 48554 58948 48594 58988
rect 48636 58948 48676 58988
rect 48718 58948 48758 58988
rect 48800 58948 48840 58988
rect 63592 58948 63632 58988
rect 63674 58948 63714 58988
rect 63756 58948 63796 58988
rect 63838 58948 63878 58988
rect 63920 58948 63960 58988
rect 78712 58948 78752 58988
rect 78794 58948 78834 58988
rect 78876 58948 78916 58988
rect 78958 58948 78998 58988
rect 79040 58948 79080 58988
rect 93832 58948 93872 58988
rect 93914 58948 93954 58988
rect 93996 58948 94036 58988
rect 94078 58948 94118 58988
rect 94160 58948 94200 58988
rect 652 58612 692 58652
rect 844 58360 884 58400
rect 4352 58192 4392 58232
rect 4434 58192 4474 58232
rect 4516 58192 4556 58232
rect 4598 58192 4638 58232
rect 4680 58192 4720 58232
rect 19472 58192 19512 58232
rect 19554 58192 19594 58232
rect 19636 58192 19676 58232
rect 19718 58192 19758 58232
rect 19800 58192 19840 58232
rect 34592 58192 34632 58232
rect 34674 58192 34714 58232
rect 34756 58192 34796 58232
rect 34838 58192 34878 58232
rect 34920 58192 34960 58232
rect 49712 58192 49752 58232
rect 49794 58192 49834 58232
rect 49876 58192 49916 58232
rect 49958 58192 49998 58232
rect 50040 58192 50080 58232
rect 64832 58192 64872 58232
rect 64914 58192 64954 58232
rect 64996 58192 65036 58232
rect 65078 58192 65118 58232
rect 65160 58192 65200 58232
rect 79952 58192 79992 58232
rect 80034 58192 80074 58232
rect 80116 58192 80156 58232
rect 80198 58192 80238 58232
rect 80280 58192 80320 58232
rect 95072 58192 95112 58232
rect 95154 58192 95194 58232
rect 95236 58192 95276 58232
rect 95318 58192 95358 58232
rect 95400 58192 95440 58232
rect 6316 57856 6356 57896
rect 6508 57856 6548 57896
rect 6508 57604 6548 57644
rect 3112 57436 3152 57476
rect 3194 57436 3234 57476
rect 3276 57436 3316 57476
rect 3358 57436 3398 57476
rect 3440 57436 3480 57476
rect 18232 57436 18272 57476
rect 18314 57436 18354 57476
rect 18396 57436 18436 57476
rect 18478 57436 18518 57476
rect 18560 57436 18600 57476
rect 33352 57436 33392 57476
rect 33434 57436 33474 57476
rect 33516 57436 33556 57476
rect 33598 57436 33638 57476
rect 33680 57436 33720 57476
rect 48472 57436 48512 57476
rect 48554 57436 48594 57476
rect 48636 57436 48676 57476
rect 48718 57436 48758 57476
rect 48800 57436 48840 57476
rect 63592 57436 63632 57476
rect 63674 57436 63714 57476
rect 63756 57436 63796 57476
rect 63838 57436 63878 57476
rect 63920 57436 63960 57476
rect 78712 57436 78752 57476
rect 78794 57436 78834 57476
rect 78876 57436 78916 57476
rect 78958 57436 78998 57476
rect 79040 57436 79080 57476
rect 93832 57436 93872 57476
rect 93914 57436 93954 57476
rect 93996 57436 94036 57476
rect 94078 57436 94118 57476
rect 94160 57436 94200 57476
rect 5836 57016 5876 57056
rect 5932 57016 5972 57056
rect 6031 57039 6071 57079
rect 6220 57016 6260 57056
rect 6508 57016 6548 57056
rect 6988 57016 7028 57056
rect 7084 57016 7124 57056
rect 7180 57016 7220 57056
rect 7276 57016 7316 57056
rect 6700 56848 6740 56888
rect 4352 56680 4392 56720
rect 4434 56680 4474 56720
rect 4516 56680 4556 56720
rect 4598 56680 4638 56720
rect 4680 56680 4720 56720
rect 19472 56680 19512 56720
rect 19554 56680 19594 56720
rect 19636 56680 19676 56720
rect 19718 56680 19758 56720
rect 19800 56680 19840 56720
rect 34592 56680 34632 56720
rect 34674 56680 34714 56720
rect 34756 56680 34796 56720
rect 34838 56680 34878 56720
rect 34920 56680 34960 56720
rect 49712 56680 49752 56720
rect 49794 56680 49834 56720
rect 49876 56680 49916 56720
rect 49958 56680 49998 56720
rect 50040 56680 50080 56720
rect 64832 56680 64872 56720
rect 64914 56680 64954 56720
rect 64996 56680 65036 56720
rect 65078 56680 65118 56720
rect 65160 56680 65200 56720
rect 79952 56680 79992 56720
rect 80034 56680 80074 56720
rect 80116 56680 80156 56720
rect 80198 56680 80238 56720
rect 80280 56680 80320 56720
rect 95072 56680 95112 56720
rect 95154 56680 95194 56720
rect 95236 56680 95276 56720
rect 95318 56680 95358 56720
rect 95400 56680 95440 56720
rect 6604 56344 6644 56384
rect 6700 56344 6740 56384
rect 652 56260 692 56300
rect 844 56092 884 56132
rect 6412 56092 6452 56132
rect 3112 55924 3152 55964
rect 3194 55924 3234 55964
rect 3276 55924 3316 55964
rect 3358 55924 3398 55964
rect 3440 55924 3480 55964
rect 18232 55924 18272 55964
rect 18314 55924 18354 55964
rect 18396 55924 18436 55964
rect 18478 55924 18518 55964
rect 18560 55924 18600 55964
rect 33352 55924 33392 55964
rect 33434 55924 33474 55964
rect 33516 55924 33556 55964
rect 33598 55924 33638 55964
rect 33680 55924 33720 55964
rect 48472 55924 48512 55964
rect 48554 55924 48594 55964
rect 48636 55924 48676 55964
rect 48718 55924 48758 55964
rect 48800 55924 48840 55964
rect 63592 55924 63632 55964
rect 63674 55924 63714 55964
rect 63756 55924 63796 55964
rect 63838 55924 63878 55964
rect 63920 55924 63960 55964
rect 78712 55924 78752 55964
rect 78794 55924 78834 55964
rect 78876 55924 78916 55964
rect 78958 55924 78998 55964
rect 79040 55924 79080 55964
rect 93832 55924 93872 55964
rect 93914 55924 93954 55964
rect 93996 55924 94036 55964
rect 94078 55924 94118 55964
rect 94160 55924 94200 55964
rect 4352 55168 4392 55208
rect 4434 55168 4474 55208
rect 4516 55168 4556 55208
rect 4598 55168 4638 55208
rect 4680 55168 4720 55208
rect 19472 55168 19512 55208
rect 19554 55168 19594 55208
rect 19636 55168 19676 55208
rect 19718 55168 19758 55208
rect 19800 55168 19840 55208
rect 34592 55168 34632 55208
rect 34674 55168 34714 55208
rect 34756 55168 34796 55208
rect 34838 55168 34878 55208
rect 34920 55168 34960 55208
rect 49712 55168 49752 55208
rect 49794 55168 49834 55208
rect 49876 55168 49916 55208
rect 49958 55168 49998 55208
rect 50040 55168 50080 55208
rect 64832 55168 64872 55208
rect 64914 55168 64954 55208
rect 64996 55168 65036 55208
rect 65078 55168 65118 55208
rect 65160 55168 65200 55208
rect 79952 55168 79992 55208
rect 80034 55168 80074 55208
rect 80116 55168 80156 55208
rect 80198 55168 80238 55208
rect 80280 55168 80320 55208
rect 95072 55168 95112 55208
rect 95154 55168 95194 55208
rect 95236 55168 95276 55208
rect 95318 55168 95358 55208
rect 95400 55168 95440 55208
rect 652 54748 692 54788
rect 844 54580 884 54620
rect 3112 54412 3152 54452
rect 3194 54412 3234 54452
rect 3276 54412 3316 54452
rect 3358 54412 3398 54452
rect 3440 54412 3480 54452
rect 18232 54412 18272 54452
rect 18314 54412 18354 54452
rect 18396 54412 18436 54452
rect 18478 54412 18518 54452
rect 18560 54412 18600 54452
rect 33352 54412 33392 54452
rect 33434 54412 33474 54452
rect 33516 54412 33556 54452
rect 33598 54412 33638 54452
rect 33680 54412 33720 54452
rect 48472 54412 48512 54452
rect 48554 54412 48594 54452
rect 48636 54412 48676 54452
rect 48718 54412 48758 54452
rect 48800 54412 48840 54452
rect 63592 54412 63632 54452
rect 63674 54412 63714 54452
rect 63756 54412 63796 54452
rect 63838 54412 63878 54452
rect 63920 54412 63960 54452
rect 78712 54412 78752 54452
rect 78794 54412 78834 54452
rect 78876 54412 78916 54452
rect 78958 54412 78998 54452
rect 79040 54412 79080 54452
rect 93832 54412 93872 54452
rect 93914 54412 93954 54452
rect 93996 54412 94036 54452
rect 94078 54412 94118 54452
rect 94160 54412 94200 54452
rect 4352 53656 4392 53696
rect 4434 53656 4474 53696
rect 4516 53656 4556 53696
rect 4598 53656 4638 53696
rect 4680 53656 4720 53696
rect 19472 53656 19512 53696
rect 19554 53656 19594 53696
rect 19636 53656 19676 53696
rect 19718 53656 19758 53696
rect 19800 53656 19840 53696
rect 34592 53656 34632 53696
rect 34674 53656 34714 53696
rect 34756 53656 34796 53696
rect 34838 53656 34878 53696
rect 34920 53656 34960 53696
rect 49712 53656 49752 53696
rect 49794 53656 49834 53696
rect 49876 53656 49916 53696
rect 49958 53656 49998 53696
rect 50040 53656 50080 53696
rect 64832 53656 64872 53696
rect 64914 53656 64954 53696
rect 64996 53656 65036 53696
rect 65078 53656 65118 53696
rect 65160 53656 65200 53696
rect 79952 53656 79992 53696
rect 80034 53656 80074 53696
rect 80116 53656 80156 53696
rect 80198 53656 80238 53696
rect 80280 53656 80320 53696
rect 95072 53656 95112 53696
rect 95154 53656 95194 53696
rect 95236 53656 95276 53696
rect 95318 53656 95358 53696
rect 95400 53656 95440 53696
rect 6412 53320 6452 53360
rect 6604 53320 6644 53360
rect 6412 53068 6452 53108
rect 3112 52900 3152 52940
rect 3194 52900 3234 52940
rect 3276 52900 3316 52940
rect 3358 52900 3398 52940
rect 3440 52900 3480 52940
rect 18232 52900 18272 52940
rect 18314 52900 18354 52940
rect 18396 52900 18436 52940
rect 18478 52900 18518 52940
rect 18560 52900 18600 52940
rect 33352 52900 33392 52940
rect 33434 52900 33474 52940
rect 33516 52900 33556 52940
rect 33598 52900 33638 52940
rect 33680 52900 33720 52940
rect 48472 52900 48512 52940
rect 48554 52900 48594 52940
rect 48636 52900 48676 52940
rect 48718 52900 48758 52940
rect 48800 52900 48840 52940
rect 63592 52900 63632 52940
rect 63674 52900 63714 52940
rect 63756 52900 63796 52940
rect 63838 52900 63878 52940
rect 63920 52900 63960 52940
rect 78712 52900 78752 52940
rect 78794 52900 78834 52940
rect 78876 52900 78916 52940
rect 78958 52900 78998 52940
rect 79040 52900 79080 52940
rect 93832 52900 93872 52940
rect 93914 52900 93954 52940
rect 93996 52900 94036 52940
rect 94078 52900 94118 52940
rect 94160 52900 94200 52940
rect 5644 52732 5684 52772
rect 652 52564 692 52604
rect 5644 52480 5684 52520
rect 5740 52480 5780 52520
rect 5932 52480 5972 52520
rect 6028 52480 6068 52520
rect 6185 52495 6225 52535
rect 6604 52480 6644 52520
rect 6700 52480 6740 52520
rect 844 52312 884 52352
rect 6412 52312 6452 52352
rect 4352 52144 4392 52184
rect 4434 52144 4474 52184
rect 4516 52144 4556 52184
rect 4598 52144 4638 52184
rect 4680 52144 4720 52184
rect 19472 52144 19512 52184
rect 19554 52144 19594 52184
rect 19636 52144 19676 52184
rect 19718 52144 19758 52184
rect 19800 52144 19840 52184
rect 34592 52144 34632 52184
rect 34674 52144 34714 52184
rect 34756 52144 34796 52184
rect 34838 52144 34878 52184
rect 34920 52144 34960 52184
rect 49712 52144 49752 52184
rect 49794 52144 49834 52184
rect 49876 52144 49916 52184
rect 49958 52144 49998 52184
rect 50040 52144 50080 52184
rect 64832 52144 64872 52184
rect 64914 52144 64954 52184
rect 64996 52144 65036 52184
rect 65078 52144 65118 52184
rect 65160 52144 65200 52184
rect 79952 52144 79992 52184
rect 80034 52144 80074 52184
rect 80116 52144 80156 52184
rect 80198 52144 80238 52184
rect 80280 52144 80320 52184
rect 95072 52144 95112 52184
rect 95154 52144 95194 52184
rect 95236 52144 95276 52184
rect 95318 52144 95358 52184
rect 95400 52144 95440 52184
rect 5644 51976 5684 52016
rect 6316 51976 6356 52016
rect 2188 51892 2228 51932
rect 2956 51892 2996 51932
rect 2092 51808 2132 51848
rect 2284 51808 2324 51848
rect 2476 51808 2516 51848
rect 2764 51808 2804 51848
rect 3244 51808 3284 51848
rect 3436 51808 3476 51848
rect 3916 51808 3956 51848
rect 4012 51808 4052 51848
rect 4108 51808 4148 51848
rect 5260 51808 5300 51848
rect 5356 51808 5396 51848
rect 5548 51808 5588 51848
rect 5740 51808 5780 51848
rect 6220 51808 6260 51848
rect 6412 51808 6452 51848
rect 6796 51808 6836 51848
rect 6892 51808 6932 51848
rect 3340 51556 3380 51596
rect 6700 51556 6740 51596
rect 3112 51388 3152 51428
rect 3194 51388 3234 51428
rect 3276 51388 3316 51428
rect 3358 51388 3398 51428
rect 3440 51388 3480 51428
rect 18232 51388 18272 51428
rect 18314 51388 18354 51428
rect 18396 51388 18436 51428
rect 18478 51388 18518 51428
rect 18560 51388 18600 51428
rect 33352 51388 33392 51428
rect 33434 51388 33474 51428
rect 33516 51388 33556 51428
rect 33598 51388 33638 51428
rect 33680 51388 33720 51428
rect 48472 51388 48512 51428
rect 48554 51388 48594 51428
rect 48636 51388 48676 51428
rect 48718 51388 48758 51428
rect 48800 51388 48840 51428
rect 63592 51388 63632 51428
rect 63674 51388 63714 51428
rect 63756 51388 63796 51428
rect 63838 51388 63878 51428
rect 63920 51388 63960 51428
rect 78712 51388 78752 51428
rect 78794 51388 78834 51428
rect 78876 51388 78916 51428
rect 78958 51388 78998 51428
rect 79040 51388 79080 51428
rect 93832 51388 93872 51428
rect 93914 51388 93954 51428
rect 93996 51388 94036 51428
rect 94078 51388 94118 51428
rect 94160 51388 94200 51428
rect 652 51052 692 51092
rect 2764 50968 2804 51008
rect 2860 50968 2900 51008
rect 844 50800 884 50840
rect 2476 50800 2516 50840
rect 4352 50632 4392 50672
rect 4434 50632 4474 50672
rect 4516 50632 4556 50672
rect 4598 50632 4638 50672
rect 4680 50632 4720 50672
rect 19472 50632 19512 50672
rect 19554 50632 19594 50672
rect 19636 50632 19676 50672
rect 19718 50632 19758 50672
rect 19800 50632 19840 50672
rect 34592 50632 34632 50672
rect 34674 50632 34714 50672
rect 34756 50632 34796 50672
rect 34838 50632 34878 50672
rect 34920 50632 34960 50672
rect 49712 50632 49752 50672
rect 49794 50632 49834 50672
rect 49876 50632 49916 50672
rect 49958 50632 49998 50672
rect 50040 50632 50080 50672
rect 64832 50632 64872 50672
rect 64914 50632 64954 50672
rect 64996 50632 65036 50672
rect 65078 50632 65118 50672
rect 65160 50632 65200 50672
rect 79952 50632 79992 50672
rect 80034 50632 80074 50672
rect 80116 50632 80156 50672
rect 80198 50632 80238 50672
rect 80280 50632 80320 50672
rect 95072 50632 95112 50672
rect 95154 50632 95194 50672
rect 95236 50632 95276 50672
rect 95318 50632 95358 50672
rect 95400 50632 95440 50672
rect 3112 49876 3152 49916
rect 3194 49876 3234 49916
rect 3276 49876 3316 49916
rect 3358 49876 3398 49916
rect 3440 49876 3480 49916
rect 18232 49876 18272 49916
rect 18314 49876 18354 49916
rect 18396 49876 18436 49916
rect 18478 49876 18518 49916
rect 18560 49876 18600 49916
rect 33352 49876 33392 49916
rect 33434 49876 33474 49916
rect 33516 49876 33556 49916
rect 33598 49876 33638 49916
rect 33680 49876 33720 49916
rect 48472 49876 48512 49916
rect 48554 49876 48594 49916
rect 48636 49876 48676 49916
rect 48718 49876 48758 49916
rect 48800 49876 48840 49916
rect 63592 49876 63632 49916
rect 63674 49876 63714 49916
rect 63756 49876 63796 49916
rect 63838 49876 63878 49916
rect 63920 49876 63960 49916
rect 78712 49876 78752 49916
rect 78794 49876 78834 49916
rect 78876 49876 78916 49916
rect 78958 49876 78998 49916
rect 79040 49876 79080 49916
rect 93832 49876 93872 49916
rect 93914 49876 93954 49916
rect 93996 49876 94036 49916
rect 94078 49876 94118 49916
rect 94160 49876 94200 49916
rect 652 49540 692 49580
rect 844 49288 884 49328
rect 4352 49120 4392 49160
rect 4434 49120 4474 49160
rect 4516 49120 4556 49160
rect 4598 49120 4638 49160
rect 4680 49120 4720 49160
rect 19472 49120 19512 49160
rect 19554 49120 19594 49160
rect 19636 49120 19676 49160
rect 19718 49120 19758 49160
rect 19800 49120 19840 49160
rect 34592 49120 34632 49160
rect 34674 49120 34714 49160
rect 34756 49120 34796 49160
rect 34838 49120 34878 49160
rect 34920 49120 34960 49160
rect 49712 49120 49752 49160
rect 49794 49120 49834 49160
rect 49876 49120 49916 49160
rect 49958 49120 49998 49160
rect 50040 49120 50080 49160
rect 64832 49120 64872 49160
rect 64914 49120 64954 49160
rect 64996 49120 65036 49160
rect 65078 49120 65118 49160
rect 65160 49120 65200 49160
rect 79952 49120 79992 49160
rect 80034 49120 80074 49160
rect 80116 49120 80156 49160
rect 80198 49120 80238 49160
rect 80280 49120 80320 49160
rect 95072 49120 95112 49160
rect 95154 49120 95194 49160
rect 95236 49120 95276 49160
rect 95318 49120 95358 49160
rect 95400 49120 95440 49160
rect 3112 48364 3152 48404
rect 3194 48364 3234 48404
rect 3276 48364 3316 48404
rect 3358 48364 3398 48404
rect 3440 48364 3480 48404
rect 18232 48364 18272 48404
rect 18314 48364 18354 48404
rect 18396 48364 18436 48404
rect 18478 48364 18518 48404
rect 18560 48364 18600 48404
rect 33352 48364 33392 48404
rect 33434 48364 33474 48404
rect 33516 48364 33556 48404
rect 33598 48364 33638 48404
rect 33680 48364 33720 48404
rect 48472 48364 48512 48404
rect 48554 48364 48594 48404
rect 48636 48364 48676 48404
rect 48718 48364 48758 48404
rect 48800 48364 48840 48404
rect 63592 48364 63632 48404
rect 63674 48364 63714 48404
rect 63756 48364 63796 48404
rect 63838 48364 63878 48404
rect 63920 48364 63960 48404
rect 78712 48364 78752 48404
rect 78794 48364 78834 48404
rect 78876 48364 78916 48404
rect 78958 48364 78998 48404
rect 79040 48364 79080 48404
rect 93832 48364 93872 48404
rect 93914 48364 93954 48404
rect 93996 48364 94036 48404
rect 94078 48364 94118 48404
rect 94160 48364 94200 48404
rect 6124 47944 6164 47984
rect 6220 47944 6260 47984
rect 6316 47944 6356 47984
rect 6412 47944 6452 47984
rect 9484 47944 9524 47984
rect 9868 47944 9908 47984
rect 9388 47860 9428 47900
rect 4352 47608 4392 47648
rect 4434 47608 4474 47648
rect 4516 47608 4556 47648
rect 4598 47608 4638 47648
rect 4680 47608 4720 47648
rect 19472 47608 19512 47648
rect 19554 47608 19594 47648
rect 19636 47608 19676 47648
rect 19718 47608 19758 47648
rect 19800 47608 19840 47648
rect 34592 47608 34632 47648
rect 34674 47608 34714 47648
rect 34756 47608 34796 47648
rect 34838 47608 34878 47648
rect 34920 47608 34960 47648
rect 49712 47608 49752 47648
rect 49794 47608 49834 47648
rect 49876 47608 49916 47648
rect 49958 47608 49998 47648
rect 50040 47608 50080 47648
rect 64832 47608 64872 47648
rect 64914 47608 64954 47648
rect 64996 47608 65036 47648
rect 65078 47608 65118 47648
rect 65160 47608 65200 47648
rect 79952 47608 79992 47648
rect 80034 47608 80074 47648
rect 80116 47608 80156 47648
rect 80198 47608 80238 47648
rect 80280 47608 80320 47648
rect 95072 47608 95112 47648
rect 95154 47608 95194 47648
rect 95236 47608 95276 47648
rect 95318 47608 95358 47648
rect 95400 47608 95440 47648
rect 1996 47440 2036 47480
rect 2284 47440 2324 47480
rect 3916 47440 3956 47480
rect 6316 47440 6356 47480
rect 13132 47440 13172 47480
rect 2956 47356 2996 47396
rect 14092 47356 14132 47396
rect 14476 47356 14516 47396
rect 2092 47272 2132 47312
rect 2476 47272 2516 47312
rect 2764 47272 2804 47312
rect 3724 47272 3764 47312
rect 3820 47272 3860 47312
rect 4012 47272 4052 47312
rect 5836 47272 5876 47312
rect 5932 47272 5972 47312
rect 6508 47272 6548 47312
rect 6604 47272 6644 47312
rect 6796 47272 6836 47312
rect 6988 47272 7028 47312
rect 7372 47272 7412 47312
rect 7564 47272 7604 47312
rect 13228 47272 13268 47312
rect 13612 47272 13652 47312
rect 13900 47272 13940 47312
rect 14572 47272 14612 47312
rect 14956 47272 14996 47312
rect 652 47188 692 47228
rect 6892 47188 6932 47228
rect 7372 47104 7412 47144
rect 844 47020 884 47060
rect 5644 47020 5684 47060
rect 13420 47020 13460 47060
rect 3112 46852 3152 46892
rect 3194 46852 3234 46892
rect 3276 46852 3316 46892
rect 3358 46852 3398 46892
rect 3440 46852 3480 46892
rect 18232 46852 18272 46892
rect 18314 46852 18354 46892
rect 18396 46852 18436 46892
rect 18478 46852 18518 46892
rect 18560 46852 18600 46892
rect 33352 46852 33392 46892
rect 33434 46852 33474 46892
rect 33516 46852 33556 46892
rect 33598 46852 33638 46892
rect 33680 46852 33720 46892
rect 48472 46852 48512 46892
rect 48554 46852 48594 46892
rect 48636 46852 48676 46892
rect 48718 46852 48758 46892
rect 48800 46852 48840 46892
rect 63592 46852 63632 46892
rect 63674 46852 63714 46892
rect 63756 46852 63796 46892
rect 63838 46852 63878 46892
rect 63920 46852 63960 46892
rect 78712 46852 78752 46892
rect 78794 46852 78834 46892
rect 78876 46852 78916 46892
rect 78958 46852 78998 46892
rect 79040 46852 79080 46892
rect 93832 46852 93872 46892
rect 93914 46852 93954 46892
rect 93996 46852 94036 46892
rect 94078 46852 94118 46892
rect 94160 46852 94200 46892
rect 2860 46684 2900 46724
rect 2668 46600 2708 46640
rect 13804 46600 13844 46640
rect 13708 46516 13748 46556
rect 14284 46516 14324 46556
rect 2668 46432 2708 46472
rect 14092 46432 14132 46472
rect 4352 46096 4392 46136
rect 4434 46096 4474 46136
rect 4516 46096 4556 46136
rect 4598 46096 4638 46136
rect 4680 46096 4720 46136
rect 19472 46096 19512 46136
rect 19554 46096 19594 46136
rect 19636 46096 19676 46136
rect 19718 46096 19758 46136
rect 19800 46096 19840 46136
rect 34592 46096 34632 46136
rect 34674 46096 34714 46136
rect 34756 46096 34796 46136
rect 34838 46096 34878 46136
rect 34920 46096 34960 46136
rect 49712 46096 49752 46136
rect 49794 46096 49834 46136
rect 49876 46096 49916 46136
rect 49958 46096 49998 46136
rect 50040 46096 50080 46136
rect 64832 46096 64872 46136
rect 64914 46096 64954 46136
rect 64996 46096 65036 46136
rect 65078 46096 65118 46136
rect 65160 46096 65200 46136
rect 79952 46096 79992 46136
rect 80034 46096 80074 46136
rect 80116 46096 80156 46136
rect 80198 46096 80238 46136
rect 80280 46096 80320 46136
rect 95072 46096 95112 46136
rect 95154 46096 95194 46136
rect 95236 46096 95276 46136
rect 95318 46096 95358 46136
rect 95400 46096 95440 46136
rect 652 45928 692 45968
rect 7564 45928 7604 45968
rect 7852 45928 7892 45968
rect 8044 45928 8084 45968
rect 14092 45928 14132 45968
rect 14380 45928 14420 45968
rect 7756 45760 7796 45800
rect 8236 45760 8276 45800
rect 8332 45760 8372 45800
rect 14188 45760 14228 45800
rect 3112 45340 3152 45380
rect 3194 45340 3234 45380
rect 3276 45340 3316 45380
rect 3358 45340 3398 45380
rect 3440 45340 3480 45380
rect 18232 45340 18272 45380
rect 18314 45340 18354 45380
rect 18396 45340 18436 45380
rect 18478 45340 18518 45380
rect 18560 45340 18600 45380
rect 33352 45340 33392 45380
rect 33434 45340 33474 45380
rect 33516 45340 33556 45380
rect 33598 45340 33638 45380
rect 33680 45340 33720 45380
rect 48472 45340 48512 45380
rect 48554 45340 48594 45380
rect 48636 45340 48676 45380
rect 48718 45340 48758 45380
rect 48800 45340 48840 45380
rect 63592 45340 63632 45380
rect 63674 45340 63714 45380
rect 63756 45340 63796 45380
rect 63838 45340 63878 45380
rect 63920 45340 63960 45380
rect 78712 45340 78752 45380
rect 78794 45340 78834 45380
rect 78876 45340 78916 45380
rect 78958 45340 78998 45380
rect 79040 45340 79080 45380
rect 93832 45340 93872 45380
rect 93914 45340 93954 45380
rect 93996 45340 94036 45380
rect 94078 45340 94118 45380
rect 94160 45340 94200 45380
rect 14188 44920 14228 44960
rect 14572 44920 14612 44960
rect 14092 44752 14132 44792
rect 4352 44584 4392 44624
rect 4434 44584 4474 44624
rect 4516 44584 4556 44624
rect 4598 44584 4638 44624
rect 4680 44584 4720 44624
rect 19472 44584 19512 44624
rect 19554 44584 19594 44624
rect 19636 44584 19676 44624
rect 19718 44584 19758 44624
rect 19800 44584 19840 44624
rect 34592 44584 34632 44624
rect 34674 44584 34714 44624
rect 34756 44584 34796 44624
rect 34838 44584 34878 44624
rect 34920 44584 34960 44624
rect 49712 44584 49752 44624
rect 49794 44584 49834 44624
rect 49876 44584 49916 44624
rect 49958 44584 49998 44624
rect 50040 44584 50080 44624
rect 64832 44584 64872 44624
rect 64914 44584 64954 44624
rect 64996 44584 65036 44624
rect 65078 44584 65118 44624
rect 65160 44584 65200 44624
rect 79952 44584 79992 44624
rect 80034 44584 80074 44624
rect 80116 44584 80156 44624
rect 80198 44584 80238 44624
rect 80280 44584 80320 44624
rect 95072 44584 95112 44624
rect 95154 44584 95194 44624
rect 95236 44584 95276 44624
rect 95318 44584 95358 44624
rect 95400 44584 95440 44624
rect 3112 43828 3152 43868
rect 3194 43828 3234 43868
rect 3276 43828 3316 43868
rect 3358 43828 3398 43868
rect 3440 43828 3480 43868
rect 18232 43828 18272 43868
rect 18314 43828 18354 43868
rect 18396 43828 18436 43868
rect 18478 43828 18518 43868
rect 18560 43828 18600 43868
rect 33352 43828 33392 43868
rect 33434 43828 33474 43868
rect 33516 43828 33556 43868
rect 33598 43828 33638 43868
rect 33680 43828 33720 43868
rect 48472 43828 48512 43868
rect 48554 43828 48594 43868
rect 48636 43828 48676 43868
rect 48718 43828 48758 43868
rect 48800 43828 48840 43868
rect 63592 43828 63632 43868
rect 63674 43828 63714 43868
rect 63756 43828 63796 43868
rect 63838 43828 63878 43868
rect 63920 43828 63960 43868
rect 78712 43828 78752 43868
rect 78794 43828 78834 43868
rect 78876 43828 78916 43868
rect 78958 43828 78998 43868
rect 79040 43828 79080 43868
rect 93832 43828 93872 43868
rect 93914 43828 93954 43868
rect 93996 43828 94036 43868
rect 94078 43828 94118 43868
rect 94160 43828 94200 43868
rect 652 43240 692 43280
rect 4352 43072 4392 43112
rect 4434 43072 4474 43112
rect 4516 43072 4556 43112
rect 4598 43072 4638 43112
rect 4680 43072 4720 43112
rect 19472 43072 19512 43112
rect 19554 43072 19594 43112
rect 19636 43072 19676 43112
rect 19718 43072 19758 43112
rect 19800 43072 19840 43112
rect 34592 43072 34632 43112
rect 34674 43072 34714 43112
rect 34756 43072 34796 43112
rect 34838 43072 34878 43112
rect 34920 43072 34960 43112
rect 49712 43072 49752 43112
rect 49794 43072 49834 43112
rect 49876 43072 49916 43112
rect 49958 43072 49998 43112
rect 50040 43072 50080 43112
rect 64832 43072 64872 43112
rect 64914 43072 64954 43112
rect 64996 43072 65036 43112
rect 65078 43072 65118 43112
rect 65160 43072 65200 43112
rect 79952 43072 79992 43112
rect 80034 43072 80074 43112
rect 80116 43072 80156 43112
rect 80198 43072 80238 43112
rect 80280 43072 80320 43112
rect 95072 43072 95112 43112
rect 95154 43072 95194 43112
rect 95236 43072 95276 43112
rect 95318 43072 95358 43112
rect 95400 43072 95440 43112
rect 3112 42316 3152 42356
rect 3194 42316 3234 42356
rect 3276 42316 3316 42356
rect 3358 42316 3398 42356
rect 3440 42316 3480 42356
rect 18232 42316 18272 42356
rect 18314 42316 18354 42356
rect 18396 42316 18436 42356
rect 18478 42316 18518 42356
rect 18560 42316 18600 42356
rect 33352 42316 33392 42356
rect 33434 42316 33474 42356
rect 33516 42316 33556 42356
rect 33598 42316 33638 42356
rect 33680 42316 33720 42356
rect 48472 42316 48512 42356
rect 48554 42316 48594 42356
rect 48636 42316 48676 42356
rect 48718 42316 48758 42356
rect 48800 42316 48840 42356
rect 63592 42316 63632 42356
rect 63674 42316 63714 42356
rect 63756 42316 63796 42356
rect 63838 42316 63878 42356
rect 63920 42316 63960 42356
rect 78712 42316 78752 42356
rect 78794 42316 78834 42356
rect 78876 42316 78916 42356
rect 78958 42316 78998 42356
rect 79040 42316 79080 42356
rect 93832 42316 93872 42356
rect 93914 42316 93954 42356
rect 93996 42316 94036 42356
rect 94078 42316 94118 42356
rect 94160 42316 94200 42356
rect 652 41728 692 41768
rect 4352 41560 4392 41600
rect 4434 41560 4474 41600
rect 4516 41560 4556 41600
rect 4598 41560 4638 41600
rect 4680 41560 4720 41600
rect 19472 41560 19512 41600
rect 19554 41560 19594 41600
rect 19636 41560 19676 41600
rect 19718 41560 19758 41600
rect 19800 41560 19840 41600
rect 34592 41560 34632 41600
rect 34674 41560 34714 41600
rect 34756 41560 34796 41600
rect 34838 41560 34878 41600
rect 34920 41560 34960 41600
rect 49712 41560 49752 41600
rect 49794 41560 49834 41600
rect 49876 41560 49916 41600
rect 49958 41560 49998 41600
rect 50040 41560 50080 41600
rect 64832 41560 64872 41600
rect 64914 41560 64954 41600
rect 64996 41560 65036 41600
rect 65078 41560 65118 41600
rect 65160 41560 65200 41600
rect 79952 41560 79992 41600
rect 80034 41560 80074 41600
rect 80116 41560 80156 41600
rect 80198 41560 80238 41600
rect 80280 41560 80320 41600
rect 95072 41560 95112 41600
rect 95154 41560 95194 41600
rect 95236 41560 95276 41600
rect 95318 41560 95358 41600
rect 95400 41560 95440 41600
rect 3112 40804 3152 40844
rect 3194 40804 3234 40844
rect 3276 40804 3316 40844
rect 3358 40804 3398 40844
rect 3440 40804 3480 40844
rect 18232 40804 18272 40844
rect 18314 40804 18354 40844
rect 18396 40804 18436 40844
rect 18478 40804 18518 40844
rect 18560 40804 18600 40844
rect 33352 40804 33392 40844
rect 33434 40804 33474 40844
rect 33516 40804 33556 40844
rect 33598 40804 33638 40844
rect 33680 40804 33720 40844
rect 48472 40804 48512 40844
rect 48554 40804 48594 40844
rect 48636 40804 48676 40844
rect 48718 40804 48758 40844
rect 48800 40804 48840 40844
rect 63592 40804 63632 40844
rect 63674 40804 63714 40844
rect 63756 40804 63796 40844
rect 63838 40804 63878 40844
rect 63920 40804 63960 40844
rect 78712 40804 78752 40844
rect 78794 40804 78834 40844
rect 78876 40804 78916 40844
rect 78958 40804 78998 40844
rect 79040 40804 79080 40844
rect 93832 40804 93872 40844
rect 93914 40804 93954 40844
rect 93996 40804 94036 40844
rect 94078 40804 94118 40844
rect 94160 40804 94200 40844
rect 4352 40048 4392 40088
rect 4434 40048 4474 40088
rect 4516 40048 4556 40088
rect 4598 40048 4638 40088
rect 4680 40048 4720 40088
rect 19472 40048 19512 40088
rect 19554 40048 19594 40088
rect 19636 40048 19676 40088
rect 19718 40048 19758 40088
rect 19800 40048 19840 40088
rect 34592 40048 34632 40088
rect 34674 40048 34714 40088
rect 34756 40048 34796 40088
rect 34838 40048 34878 40088
rect 34920 40048 34960 40088
rect 49712 40048 49752 40088
rect 49794 40048 49834 40088
rect 49876 40048 49916 40088
rect 49958 40048 49998 40088
rect 50040 40048 50080 40088
rect 64832 40048 64872 40088
rect 64914 40048 64954 40088
rect 64996 40048 65036 40088
rect 65078 40048 65118 40088
rect 65160 40048 65200 40088
rect 79952 40048 79992 40088
rect 80034 40048 80074 40088
rect 80116 40048 80156 40088
rect 80198 40048 80238 40088
rect 80280 40048 80320 40088
rect 95072 40048 95112 40088
rect 95154 40048 95194 40088
rect 95236 40048 95276 40088
rect 95318 40048 95358 40088
rect 95400 40048 95440 40088
rect 652 39880 692 39920
rect 3112 39292 3152 39332
rect 3194 39292 3234 39332
rect 3276 39292 3316 39332
rect 3358 39292 3398 39332
rect 3440 39292 3480 39332
rect 18232 39292 18272 39332
rect 18314 39292 18354 39332
rect 18396 39292 18436 39332
rect 18478 39292 18518 39332
rect 18560 39292 18600 39332
rect 33352 39292 33392 39332
rect 33434 39292 33474 39332
rect 33516 39292 33556 39332
rect 33598 39292 33638 39332
rect 33680 39292 33720 39332
rect 48472 39292 48512 39332
rect 48554 39292 48594 39332
rect 48636 39292 48676 39332
rect 48718 39292 48758 39332
rect 48800 39292 48840 39332
rect 63592 39292 63632 39332
rect 63674 39292 63714 39332
rect 63756 39292 63796 39332
rect 63838 39292 63878 39332
rect 63920 39292 63960 39332
rect 78712 39292 78752 39332
rect 78794 39292 78834 39332
rect 78876 39292 78916 39332
rect 78958 39292 78998 39332
rect 79040 39292 79080 39332
rect 93832 39292 93872 39332
rect 93914 39292 93954 39332
rect 93996 39292 94036 39332
rect 94078 39292 94118 39332
rect 94160 39292 94200 39332
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 95072 38536 95112 38576
rect 95154 38536 95194 38576
rect 95236 38536 95276 38576
rect 95318 38536 95358 38576
rect 95400 38536 95440 38576
rect 652 38368 692 38408
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 93832 37780 93872 37820
rect 93914 37780 93954 37820
rect 93996 37780 94036 37820
rect 94078 37780 94118 37820
rect 94160 37780 94200 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 95072 37024 95112 37064
rect 95154 37024 95194 37064
rect 95236 37024 95276 37064
rect 95318 37024 95358 37064
rect 95400 37024 95440 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 93832 36268 93872 36308
rect 93914 36268 93954 36308
rect 93996 36268 94036 36308
rect 94078 36268 94118 36308
rect 94160 36268 94200 36308
rect 652 35680 692 35720
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 95072 35512 95112 35552
rect 95154 35512 95194 35552
rect 95236 35512 95276 35552
rect 95318 35512 95358 35552
rect 95400 35512 95440 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 93832 34756 93872 34796
rect 93914 34756 93954 34796
rect 93996 34756 94036 34796
rect 94078 34756 94118 34796
rect 94160 34756 94200 34796
rect 652 34168 692 34208
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 95072 34000 95112 34040
rect 95154 34000 95194 34040
rect 95236 34000 95276 34040
rect 95318 34000 95358 34040
rect 95400 34000 95440 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 93832 33244 93872 33284
rect 93914 33244 93954 33284
rect 93996 33244 94036 33284
rect 94078 33244 94118 33284
rect 94160 33244 94200 33284
rect 652 32656 692 32696
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 95072 32488 95112 32528
rect 95154 32488 95194 32528
rect 95236 32488 95276 32528
rect 95318 32488 95358 32528
rect 95400 32488 95440 32528
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 93832 31732 93872 31772
rect 93914 31732 93954 31772
rect 93996 31732 94036 31772
rect 94078 31732 94118 31772
rect 94160 31732 94200 31772
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 95072 30976 95112 31016
rect 95154 30976 95194 31016
rect 95236 30976 95276 31016
rect 95318 30976 95358 31016
rect 95400 30976 95440 31016
rect 652 30808 692 30848
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 93832 30220 93872 30260
rect 93914 30220 93954 30260
rect 93996 30220 94036 30260
rect 94078 30220 94118 30260
rect 94160 30220 94200 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 95072 29464 95112 29504
rect 95154 29464 95194 29504
rect 95236 29464 95276 29504
rect 95318 29464 95358 29504
rect 95400 29464 95440 29504
rect 652 29296 692 29336
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 93832 28708 93872 28748
rect 93914 28708 93954 28748
rect 93996 28708 94036 28748
rect 94078 28708 94118 28748
rect 94160 28708 94200 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 95072 27952 95112 27992
rect 95154 27952 95194 27992
rect 95236 27952 95276 27992
rect 95318 27952 95358 27992
rect 95400 27952 95440 27992
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 93832 27196 93872 27236
rect 93914 27196 93954 27236
rect 93996 27196 94036 27236
rect 94078 27196 94118 27236
rect 94160 27196 94200 27236
rect 652 26608 692 26648
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 95072 26440 95112 26480
rect 95154 26440 95194 26480
rect 95236 26440 95276 26480
rect 95318 26440 95358 26480
rect 95400 26440 95440 26480
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 93832 25684 93872 25724
rect 93914 25684 93954 25724
rect 93996 25684 94036 25724
rect 94078 25684 94118 25724
rect 94160 25684 94200 25724
rect 652 25096 692 25136
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 95072 24928 95112 24968
rect 95154 24928 95194 24968
rect 95236 24928 95276 24968
rect 95318 24928 95358 24968
rect 95400 24928 95440 24968
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 63592 24172 63632 24212
rect 63674 24172 63714 24212
rect 63756 24172 63796 24212
rect 63838 24172 63878 24212
rect 63920 24172 63960 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 93832 24172 93872 24212
rect 93914 24172 93954 24212
rect 93996 24172 94036 24212
rect 94078 24172 94118 24212
rect 94160 24172 94200 24212
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 64832 23416 64872 23456
rect 64914 23416 64954 23456
rect 64996 23416 65036 23456
rect 65078 23416 65118 23456
rect 65160 23416 65200 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 95072 23416 95112 23456
rect 95154 23416 95194 23456
rect 95236 23416 95276 23456
rect 95318 23416 95358 23456
rect 95400 23416 95440 23456
rect 652 23248 692 23288
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 63592 22660 63632 22700
rect 63674 22660 63714 22700
rect 63756 22660 63796 22700
rect 63838 22660 63878 22700
rect 63920 22660 63960 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 93832 22660 93872 22700
rect 93914 22660 93954 22700
rect 93996 22660 94036 22700
rect 94078 22660 94118 22700
rect 94160 22660 94200 22700
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 64832 21904 64872 21944
rect 64914 21904 64954 21944
rect 64996 21904 65036 21944
rect 65078 21904 65118 21944
rect 65160 21904 65200 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 652 21736 692 21776
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 63592 21148 63632 21188
rect 63674 21148 63714 21188
rect 63756 21148 63796 21188
rect 63838 21148 63878 21188
rect 63920 21148 63960 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 64832 20392 64872 20432
rect 64914 20392 64954 20432
rect 64996 20392 65036 20432
rect 65078 20392 65118 20432
rect 65160 20392 65200 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 63592 19636 63632 19676
rect 63674 19636 63714 19676
rect 63756 19636 63796 19676
rect 63838 19636 63878 19676
rect 63920 19636 63960 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 652 19048 692 19088
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 64832 18880 64872 18920
rect 64914 18880 64954 18920
rect 64996 18880 65036 18920
rect 65078 18880 65118 18920
rect 65160 18880 65200 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 95072 18880 95112 18920
rect 95154 18880 95194 18920
rect 95236 18880 95276 18920
rect 95318 18880 95358 18920
rect 95400 18880 95440 18920
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 63592 18124 63632 18164
rect 63674 18124 63714 18164
rect 63756 18124 63796 18164
rect 63838 18124 63878 18164
rect 63920 18124 63960 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 93832 18124 93872 18164
rect 93914 18124 93954 18164
rect 93996 18124 94036 18164
rect 94078 18124 94118 18164
rect 94160 18124 94200 18164
rect 652 17536 692 17576
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 64832 17368 64872 17408
rect 64914 17368 64954 17408
rect 64996 17368 65036 17408
rect 65078 17368 65118 17408
rect 65160 17368 65200 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 95072 17368 95112 17408
rect 95154 17368 95194 17408
rect 95236 17368 95276 17408
rect 95318 17368 95358 17408
rect 95400 17368 95440 17408
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 63592 16612 63632 16652
rect 63674 16612 63714 16652
rect 63756 16612 63796 16652
rect 63838 16612 63878 16652
rect 63920 16612 63960 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 93832 16612 93872 16652
rect 93914 16612 93954 16652
rect 93996 16612 94036 16652
rect 94078 16612 94118 16652
rect 94160 16612 94200 16652
rect 844 16276 884 16316
rect 652 16024 692 16064
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 64832 15856 64872 15896
rect 64914 15856 64954 15896
rect 64996 15856 65036 15896
rect 65078 15856 65118 15896
rect 65160 15856 65200 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 95072 15856 95112 15896
rect 95154 15856 95194 15896
rect 95236 15856 95276 15896
rect 95318 15856 95358 15896
rect 95400 15856 95440 15896
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 93832 15100 93872 15140
rect 93914 15100 93954 15140
rect 93996 15100 94036 15140
rect 94078 15100 94118 15140
rect 94160 15100 94200 15140
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 95072 14344 95112 14384
rect 95154 14344 95194 14384
rect 95236 14344 95276 14384
rect 95318 14344 95358 14384
rect 95400 14344 95440 14384
rect 844 13924 884 13964
rect 652 13756 692 13796
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 93832 13588 93872 13628
rect 93914 13588 93954 13628
rect 93996 13588 94036 13628
rect 94078 13588 94118 13628
rect 94160 13588 94200 13628
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 95072 12832 95112 12872
rect 95154 12832 95194 12872
rect 95236 12832 95276 12872
rect 95318 12832 95358 12872
rect 95400 12832 95440 12872
rect 844 12412 884 12452
rect 652 12244 692 12284
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 93832 12076 93872 12116
rect 93914 12076 93954 12116
rect 93996 12076 94036 12116
rect 94078 12076 94118 12116
rect 94160 12076 94200 12116
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 95072 11320 95112 11360
rect 95154 11320 95194 11360
rect 95236 11320 95276 11360
rect 95318 11320 95358 11360
rect 95400 11320 95440 11360
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 93832 10564 93872 10604
rect 93914 10564 93954 10604
rect 93996 10564 94036 10604
rect 94078 10564 94118 10604
rect 94160 10564 94200 10604
rect 844 10228 884 10268
rect 652 9976 692 10016
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 95072 9808 95112 9848
rect 95154 9808 95194 9848
rect 95236 9808 95276 9848
rect 95318 9808 95358 9848
rect 95400 9808 95440 9848
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 93832 9052 93872 9092
rect 93914 9052 93954 9092
rect 93996 9052 94036 9092
rect 94078 9052 94118 9092
rect 94160 9052 94200 9092
rect 844 8716 884 8756
rect 652 8464 692 8504
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 95072 8296 95112 8336
rect 95154 8296 95194 8336
rect 95236 8296 95276 8336
rect 95318 8296 95358 8336
rect 95400 8296 95440 8336
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 93832 7540 93872 7580
rect 93914 7540 93954 7580
rect 93996 7540 94036 7580
rect 94078 7540 94118 7580
rect 94160 7540 94200 7580
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 95072 6784 95112 6824
rect 95154 6784 95194 6824
rect 95236 6784 95276 6824
rect 95318 6784 95358 6824
rect 95400 6784 95440 6824
rect 844 6364 884 6404
rect 652 6280 692 6320
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 93832 6028 93872 6068
rect 93914 6028 93954 6068
rect 93996 6028 94036 6068
rect 94078 6028 94118 6068
rect 94160 6028 94200 6068
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 95072 5272 95112 5312
rect 95154 5272 95194 5312
rect 95236 5272 95276 5312
rect 95318 5272 95358 5312
rect 95400 5272 95440 5312
rect 844 4852 884 4892
rect 652 4684 692 4724
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 93832 4516 93872 4556
rect 93914 4516 93954 4556
rect 93996 4516 94036 4556
rect 94078 4516 94118 4556
rect 94160 4516 94200 4556
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 95072 3760 95112 3800
rect 95154 3760 95194 3800
rect 95236 3760 95276 3800
rect 95318 3760 95358 3800
rect 95400 3760 95440 3800
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 93832 3004 93872 3044
rect 93914 3004 93954 3044
rect 93996 3004 94036 3044
rect 94078 3004 94118 3044
rect 94160 3004 94200 3044
rect 652 2752 692 2792
rect 844 2668 884 2708
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 95072 2248 95112 2288
rect 95154 2248 95194 2288
rect 95236 2248 95276 2288
rect 95318 2248 95358 2288
rect 95400 2248 95440 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 93832 1492 93872 1532
rect 93914 1492 93954 1532
rect 93996 1492 94036 1532
rect 94078 1492 94118 1532
rect 94160 1492 94200 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
rect 95072 736 95112 776
rect 95154 736 95194 776
rect 95236 736 95276 776
rect 95318 736 95358 776
rect 95400 736 95440 776
<< metal2 >>
rect 3112 81668 3480 81677
rect 3152 81628 3194 81668
rect 3234 81628 3276 81668
rect 3316 81628 3358 81668
rect 3398 81628 3440 81668
rect 3112 81619 3480 81628
rect 18232 81668 18600 81677
rect 18272 81628 18314 81668
rect 18354 81628 18396 81668
rect 18436 81628 18478 81668
rect 18518 81628 18560 81668
rect 18232 81619 18600 81628
rect 33352 81668 33720 81677
rect 33392 81628 33434 81668
rect 33474 81628 33516 81668
rect 33556 81628 33598 81668
rect 33638 81628 33680 81668
rect 33352 81619 33720 81628
rect 48472 81668 48840 81677
rect 48512 81628 48554 81668
rect 48594 81628 48636 81668
rect 48676 81628 48718 81668
rect 48758 81628 48800 81668
rect 48472 81619 48840 81628
rect 63592 81668 63960 81677
rect 63632 81628 63674 81668
rect 63714 81628 63756 81668
rect 63796 81628 63838 81668
rect 63878 81628 63920 81668
rect 63592 81619 63960 81628
rect 78712 81668 79080 81677
rect 78752 81628 78794 81668
rect 78834 81628 78876 81668
rect 78916 81628 78958 81668
rect 78998 81628 79040 81668
rect 78712 81619 79080 81628
rect 93832 81668 94200 81677
rect 93872 81628 93914 81668
rect 93954 81628 93996 81668
rect 94036 81628 94078 81668
rect 94118 81628 94160 81668
rect 93832 81619 94200 81628
rect 4352 80912 4720 80921
rect 4392 80872 4434 80912
rect 4474 80872 4516 80912
rect 4556 80872 4598 80912
rect 4638 80872 4680 80912
rect 4352 80863 4720 80872
rect 19472 80912 19840 80921
rect 19512 80872 19554 80912
rect 19594 80872 19636 80912
rect 19676 80872 19718 80912
rect 19758 80872 19800 80912
rect 19472 80863 19840 80872
rect 34592 80912 34960 80921
rect 34632 80872 34674 80912
rect 34714 80872 34756 80912
rect 34796 80872 34838 80912
rect 34878 80872 34920 80912
rect 34592 80863 34960 80872
rect 49712 80912 50080 80921
rect 49752 80872 49794 80912
rect 49834 80872 49876 80912
rect 49916 80872 49958 80912
rect 49998 80872 50040 80912
rect 49712 80863 50080 80872
rect 64832 80912 65200 80921
rect 64872 80872 64914 80912
rect 64954 80872 64996 80912
rect 65036 80872 65078 80912
rect 65118 80872 65160 80912
rect 64832 80863 65200 80872
rect 79952 80912 80320 80921
rect 79992 80872 80034 80912
rect 80074 80872 80116 80912
rect 80156 80872 80198 80912
rect 80238 80872 80280 80912
rect 79952 80863 80320 80872
rect 95072 80912 95440 80921
rect 95112 80872 95154 80912
rect 95194 80872 95236 80912
rect 95276 80872 95318 80912
rect 95358 80872 95400 80912
rect 95072 80863 95440 80872
rect 3112 80156 3480 80165
rect 3152 80116 3194 80156
rect 3234 80116 3276 80156
rect 3316 80116 3358 80156
rect 3398 80116 3440 80156
rect 3112 80107 3480 80116
rect 18232 80156 18600 80165
rect 18272 80116 18314 80156
rect 18354 80116 18396 80156
rect 18436 80116 18478 80156
rect 18518 80116 18560 80156
rect 18232 80107 18600 80116
rect 33352 80156 33720 80165
rect 33392 80116 33434 80156
rect 33474 80116 33516 80156
rect 33556 80116 33598 80156
rect 33638 80116 33680 80156
rect 33352 80107 33720 80116
rect 48472 80156 48840 80165
rect 48512 80116 48554 80156
rect 48594 80116 48636 80156
rect 48676 80116 48718 80156
rect 48758 80116 48800 80156
rect 48472 80107 48840 80116
rect 63592 80156 63960 80165
rect 63632 80116 63674 80156
rect 63714 80116 63756 80156
rect 63796 80116 63838 80156
rect 63878 80116 63920 80156
rect 63592 80107 63960 80116
rect 78712 80156 79080 80165
rect 78752 80116 78794 80156
rect 78834 80116 78876 80156
rect 78916 80116 78958 80156
rect 78998 80116 79040 80156
rect 78712 80107 79080 80116
rect 93832 80156 94200 80165
rect 93872 80116 93914 80156
rect 93954 80116 93996 80156
rect 94036 80116 94078 80156
rect 94118 80116 94160 80156
rect 93832 80107 94200 80116
rect 4352 79400 4720 79409
rect 4392 79360 4434 79400
rect 4474 79360 4516 79400
rect 4556 79360 4598 79400
rect 4638 79360 4680 79400
rect 4352 79351 4720 79360
rect 19472 79400 19840 79409
rect 19512 79360 19554 79400
rect 19594 79360 19636 79400
rect 19676 79360 19718 79400
rect 19758 79360 19800 79400
rect 19472 79351 19840 79360
rect 34592 79400 34960 79409
rect 34632 79360 34674 79400
rect 34714 79360 34756 79400
rect 34796 79360 34838 79400
rect 34878 79360 34920 79400
rect 34592 79351 34960 79360
rect 49712 79400 50080 79409
rect 49752 79360 49794 79400
rect 49834 79360 49876 79400
rect 49916 79360 49958 79400
rect 49998 79360 50040 79400
rect 49712 79351 50080 79360
rect 64832 79400 65200 79409
rect 64872 79360 64914 79400
rect 64954 79360 64996 79400
rect 65036 79360 65078 79400
rect 65118 79360 65160 79400
rect 64832 79351 65200 79360
rect 79952 79400 80320 79409
rect 79992 79360 80034 79400
rect 80074 79360 80116 79400
rect 80156 79360 80198 79400
rect 80238 79360 80280 79400
rect 79952 79351 80320 79360
rect 95072 79400 95440 79409
rect 95112 79360 95154 79400
rect 95194 79360 95236 79400
rect 95276 79360 95318 79400
rect 95358 79360 95400 79400
rect 95072 79351 95440 79360
rect 3112 78644 3480 78653
rect 3152 78604 3194 78644
rect 3234 78604 3276 78644
rect 3316 78604 3358 78644
rect 3398 78604 3440 78644
rect 3112 78595 3480 78604
rect 18232 78644 18600 78653
rect 18272 78604 18314 78644
rect 18354 78604 18396 78644
rect 18436 78604 18478 78644
rect 18518 78604 18560 78644
rect 18232 78595 18600 78604
rect 33352 78644 33720 78653
rect 33392 78604 33434 78644
rect 33474 78604 33516 78644
rect 33556 78604 33598 78644
rect 33638 78604 33680 78644
rect 33352 78595 33720 78604
rect 48472 78644 48840 78653
rect 48512 78604 48554 78644
rect 48594 78604 48636 78644
rect 48676 78604 48718 78644
rect 48758 78604 48800 78644
rect 48472 78595 48840 78604
rect 63592 78644 63960 78653
rect 63632 78604 63674 78644
rect 63714 78604 63756 78644
rect 63796 78604 63838 78644
rect 63878 78604 63920 78644
rect 63592 78595 63960 78604
rect 78712 78644 79080 78653
rect 78752 78604 78794 78644
rect 78834 78604 78876 78644
rect 78916 78604 78958 78644
rect 78998 78604 79040 78644
rect 78712 78595 79080 78604
rect 93832 78644 94200 78653
rect 93872 78604 93914 78644
rect 93954 78604 93996 78644
rect 94036 78604 94078 78644
rect 94118 78604 94160 78644
rect 93832 78595 94200 78604
rect 4352 77888 4720 77897
rect 4392 77848 4434 77888
rect 4474 77848 4516 77888
rect 4556 77848 4598 77888
rect 4638 77848 4680 77888
rect 4352 77839 4720 77848
rect 19472 77888 19840 77897
rect 19512 77848 19554 77888
rect 19594 77848 19636 77888
rect 19676 77848 19718 77888
rect 19758 77848 19800 77888
rect 19472 77839 19840 77848
rect 34592 77888 34960 77897
rect 34632 77848 34674 77888
rect 34714 77848 34756 77888
rect 34796 77848 34838 77888
rect 34878 77848 34920 77888
rect 34592 77839 34960 77848
rect 49712 77888 50080 77897
rect 49752 77848 49794 77888
rect 49834 77848 49876 77888
rect 49916 77848 49958 77888
rect 49998 77848 50040 77888
rect 49712 77839 50080 77848
rect 64832 77888 65200 77897
rect 64872 77848 64914 77888
rect 64954 77848 64996 77888
rect 65036 77848 65078 77888
rect 65118 77848 65160 77888
rect 64832 77839 65200 77848
rect 79952 77888 80320 77897
rect 79992 77848 80034 77888
rect 80074 77848 80116 77888
rect 80156 77848 80198 77888
rect 80238 77848 80280 77888
rect 79952 77839 80320 77848
rect 95072 77888 95440 77897
rect 95112 77848 95154 77888
rect 95194 77848 95236 77888
rect 95276 77848 95318 77888
rect 95358 77848 95400 77888
rect 95072 77839 95440 77848
rect 3112 77132 3480 77141
rect 3152 77092 3194 77132
rect 3234 77092 3276 77132
rect 3316 77092 3358 77132
rect 3398 77092 3440 77132
rect 3112 77083 3480 77092
rect 18232 77132 18600 77141
rect 18272 77092 18314 77132
rect 18354 77092 18396 77132
rect 18436 77092 18478 77132
rect 18518 77092 18560 77132
rect 18232 77083 18600 77092
rect 33352 77132 33720 77141
rect 33392 77092 33434 77132
rect 33474 77092 33516 77132
rect 33556 77092 33598 77132
rect 33638 77092 33680 77132
rect 33352 77083 33720 77092
rect 48472 77132 48840 77141
rect 48512 77092 48554 77132
rect 48594 77092 48636 77132
rect 48676 77092 48718 77132
rect 48758 77092 48800 77132
rect 48472 77083 48840 77092
rect 63592 77132 63960 77141
rect 63632 77092 63674 77132
rect 63714 77092 63756 77132
rect 63796 77092 63838 77132
rect 63878 77092 63920 77132
rect 63592 77083 63960 77092
rect 78712 77132 79080 77141
rect 78752 77092 78794 77132
rect 78834 77092 78876 77132
rect 78916 77092 78958 77132
rect 78998 77092 79040 77132
rect 78712 77083 79080 77092
rect 93832 77132 94200 77141
rect 93872 77092 93914 77132
rect 93954 77092 93996 77132
rect 94036 77092 94078 77132
rect 94118 77092 94160 77132
rect 93832 77083 94200 77092
rect 4352 76376 4720 76385
rect 4392 76336 4434 76376
rect 4474 76336 4516 76376
rect 4556 76336 4598 76376
rect 4638 76336 4680 76376
rect 4352 76327 4720 76336
rect 19472 76376 19840 76385
rect 19512 76336 19554 76376
rect 19594 76336 19636 76376
rect 19676 76336 19718 76376
rect 19758 76336 19800 76376
rect 19472 76327 19840 76336
rect 34592 76376 34960 76385
rect 34632 76336 34674 76376
rect 34714 76336 34756 76376
rect 34796 76336 34838 76376
rect 34878 76336 34920 76376
rect 34592 76327 34960 76336
rect 49712 76376 50080 76385
rect 49752 76336 49794 76376
rect 49834 76336 49876 76376
rect 49916 76336 49958 76376
rect 49998 76336 50040 76376
rect 49712 76327 50080 76336
rect 64832 76376 65200 76385
rect 64872 76336 64914 76376
rect 64954 76336 64996 76376
rect 65036 76336 65078 76376
rect 65118 76336 65160 76376
rect 64832 76327 65200 76336
rect 79952 76376 80320 76385
rect 79992 76336 80034 76376
rect 80074 76336 80116 76376
rect 80156 76336 80198 76376
rect 80238 76336 80280 76376
rect 79952 76327 80320 76336
rect 95072 76376 95440 76385
rect 95112 76336 95154 76376
rect 95194 76336 95236 76376
rect 95276 76336 95318 76376
rect 95358 76336 95400 76376
rect 95072 76327 95440 76336
rect 3112 75620 3480 75629
rect 3152 75580 3194 75620
rect 3234 75580 3276 75620
rect 3316 75580 3358 75620
rect 3398 75580 3440 75620
rect 3112 75571 3480 75580
rect 18232 75620 18600 75629
rect 18272 75580 18314 75620
rect 18354 75580 18396 75620
rect 18436 75580 18478 75620
rect 18518 75580 18560 75620
rect 18232 75571 18600 75580
rect 33352 75620 33720 75629
rect 33392 75580 33434 75620
rect 33474 75580 33516 75620
rect 33556 75580 33598 75620
rect 33638 75580 33680 75620
rect 33352 75571 33720 75580
rect 48472 75620 48840 75629
rect 48512 75580 48554 75620
rect 48594 75580 48636 75620
rect 48676 75580 48718 75620
rect 48758 75580 48800 75620
rect 48472 75571 48840 75580
rect 63592 75620 63960 75629
rect 63632 75580 63674 75620
rect 63714 75580 63756 75620
rect 63796 75580 63838 75620
rect 63878 75580 63920 75620
rect 63592 75571 63960 75580
rect 78712 75620 79080 75629
rect 78752 75580 78794 75620
rect 78834 75580 78876 75620
rect 78916 75580 78958 75620
rect 78998 75580 79040 75620
rect 78712 75571 79080 75580
rect 93832 75620 94200 75629
rect 93872 75580 93914 75620
rect 93954 75580 93996 75620
rect 94036 75580 94078 75620
rect 94118 75580 94160 75620
rect 93832 75571 94200 75580
rect 652 75284 692 75293
rect 652 74705 692 75244
rect 844 75032 884 75041
rect 748 74992 844 75032
rect 651 74696 693 74705
rect 651 74656 652 74696
rect 692 74656 693 74696
rect 651 74647 693 74656
rect 651 72932 693 72941
rect 651 72892 652 72932
rect 692 72892 693 72932
rect 651 72883 693 72892
rect 652 72798 692 72883
rect 652 71504 692 71513
rect 652 71009 692 71464
rect 651 71000 693 71009
rect 651 70960 652 71000
rect 692 70960 693 71000
rect 651 70951 693 70960
rect 651 69236 693 69245
rect 651 69196 652 69236
rect 692 69196 693 69236
rect 651 69187 693 69196
rect 652 69102 692 69187
rect 652 67724 692 67733
rect 555 67472 597 67481
rect 555 67432 556 67472
rect 596 67432 597 67472
rect 555 67423 597 67432
rect 556 47321 596 67423
rect 652 67313 692 67684
rect 651 67304 693 67313
rect 651 67264 652 67304
rect 692 67264 693 67304
rect 651 67255 693 67264
rect 652 66212 692 66221
rect 652 65465 692 66172
rect 651 65456 693 65465
rect 651 65416 652 65456
rect 692 65416 693 65456
rect 651 65407 693 65416
rect 652 63860 692 63869
rect 652 63617 692 63820
rect 651 63608 693 63617
rect 651 63568 652 63608
rect 692 63568 693 63608
rect 651 63559 693 63568
rect 748 63029 788 74992
rect 844 74983 884 74992
rect 4352 74864 4720 74873
rect 4392 74824 4434 74864
rect 4474 74824 4516 74864
rect 4556 74824 4598 74864
rect 4638 74824 4680 74864
rect 4352 74815 4720 74824
rect 19472 74864 19840 74873
rect 19512 74824 19554 74864
rect 19594 74824 19636 74864
rect 19676 74824 19718 74864
rect 19758 74824 19800 74864
rect 19472 74815 19840 74824
rect 34592 74864 34960 74873
rect 34632 74824 34674 74864
rect 34714 74824 34756 74864
rect 34796 74824 34838 74864
rect 34878 74824 34920 74864
rect 34592 74815 34960 74824
rect 49712 74864 50080 74873
rect 49752 74824 49794 74864
rect 49834 74824 49876 74864
rect 49916 74824 49958 74864
rect 49998 74824 50040 74864
rect 49712 74815 50080 74824
rect 64832 74864 65200 74873
rect 64872 74824 64914 74864
rect 64954 74824 64996 74864
rect 65036 74824 65078 74864
rect 65118 74824 65160 74864
rect 64832 74815 65200 74824
rect 79952 74864 80320 74873
rect 79992 74824 80034 74864
rect 80074 74824 80116 74864
rect 80156 74824 80198 74864
rect 80238 74824 80280 74864
rect 79952 74815 80320 74824
rect 95072 74864 95440 74873
rect 95112 74824 95154 74864
rect 95194 74824 95236 74864
rect 95276 74824 95318 74864
rect 95358 74824 95400 74864
rect 95072 74815 95440 74824
rect 3112 74108 3480 74117
rect 3152 74068 3194 74108
rect 3234 74068 3276 74108
rect 3316 74068 3358 74108
rect 3398 74068 3440 74108
rect 3112 74059 3480 74068
rect 18232 74108 18600 74117
rect 18272 74068 18314 74108
rect 18354 74068 18396 74108
rect 18436 74068 18478 74108
rect 18518 74068 18560 74108
rect 18232 74059 18600 74068
rect 33352 74108 33720 74117
rect 33392 74068 33434 74108
rect 33474 74068 33516 74108
rect 33556 74068 33598 74108
rect 33638 74068 33680 74108
rect 33352 74059 33720 74068
rect 48472 74108 48840 74117
rect 48512 74068 48554 74108
rect 48594 74068 48636 74108
rect 48676 74068 48718 74108
rect 48758 74068 48800 74108
rect 48472 74059 48840 74068
rect 63592 74108 63960 74117
rect 63632 74068 63674 74108
rect 63714 74068 63756 74108
rect 63796 74068 63838 74108
rect 63878 74068 63920 74108
rect 63592 74059 63960 74068
rect 78712 74108 79080 74117
rect 78752 74068 78794 74108
rect 78834 74068 78876 74108
rect 78916 74068 78958 74108
rect 78998 74068 79040 74108
rect 78712 74059 79080 74068
rect 93832 74108 94200 74117
rect 93872 74068 93914 74108
rect 93954 74068 93996 74108
rect 94036 74068 94078 74108
rect 94118 74068 94160 74108
rect 93832 74059 94200 74068
rect 4352 73352 4720 73361
rect 4392 73312 4434 73352
rect 4474 73312 4516 73352
rect 4556 73312 4598 73352
rect 4638 73312 4680 73352
rect 4352 73303 4720 73312
rect 19472 73352 19840 73361
rect 19512 73312 19554 73352
rect 19594 73312 19636 73352
rect 19676 73312 19718 73352
rect 19758 73312 19800 73352
rect 19472 73303 19840 73312
rect 34592 73352 34960 73361
rect 34632 73312 34674 73352
rect 34714 73312 34756 73352
rect 34796 73312 34838 73352
rect 34878 73312 34920 73352
rect 34592 73303 34960 73312
rect 49712 73352 50080 73361
rect 49752 73312 49794 73352
rect 49834 73312 49876 73352
rect 49916 73312 49958 73352
rect 49998 73312 50040 73352
rect 49712 73303 50080 73312
rect 64832 73352 65200 73361
rect 64872 73312 64914 73352
rect 64954 73312 64996 73352
rect 65036 73312 65078 73352
rect 65118 73312 65160 73352
rect 64832 73303 65200 73312
rect 79952 73352 80320 73361
rect 79992 73312 80034 73352
rect 80074 73312 80116 73352
rect 80156 73312 80198 73352
rect 80238 73312 80280 73352
rect 79952 73303 80320 73312
rect 95072 73352 95440 73361
rect 95112 73312 95154 73352
rect 95194 73312 95236 73352
rect 95276 73312 95318 73352
rect 95358 73312 95400 73352
rect 95072 73303 95440 73312
rect 844 72764 884 72773
rect 884 72724 1076 72764
rect 844 72715 884 72724
rect 844 71504 884 71513
rect 884 71464 980 71504
rect 844 71455 884 71464
rect 843 68984 885 68993
rect 843 68944 844 68984
rect 884 68944 885 68984
rect 843 68935 885 68944
rect 844 68850 884 68935
rect 843 67472 885 67481
rect 843 67432 844 67472
rect 884 67432 885 67472
rect 843 67423 885 67432
rect 844 67338 884 67423
rect 843 65960 885 65969
rect 843 65920 844 65960
rect 884 65920 885 65960
rect 843 65911 885 65920
rect 844 65826 884 65911
rect 843 63692 885 63701
rect 843 63652 844 63692
rect 884 63652 885 63692
rect 843 63643 885 63652
rect 844 63558 884 63643
rect 747 63020 789 63029
rect 747 62980 748 63020
rect 788 62980 789 63020
rect 747 62971 789 62980
rect 652 62348 692 62357
rect 652 61769 692 62308
rect 843 62180 885 62189
rect 843 62140 844 62180
rect 884 62140 885 62180
rect 843 62131 885 62140
rect 844 62046 884 62131
rect 651 61760 693 61769
rect 651 61720 652 61760
rect 692 61720 693 61760
rect 651 61711 693 61720
rect 843 60332 885 60341
rect 843 60292 844 60332
rect 884 60292 885 60332
rect 843 60283 885 60292
rect 844 60198 884 60283
rect 652 60164 692 60173
rect 652 59921 692 60124
rect 651 59912 693 59921
rect 651 59872 652 59912
rect 692 59872 693 59912
rect 651 59863 693 59872
rect 652 58652 692 58661
rect 652 58073 692 58612
rect 844 58400 884 58409
rect 651 58064 693 58073
rect 651 58024 652 58064
rect 692 58024 693 58064
rect 651 58015 693 58024
rect 844 57149 884 58360
rect 843 57140 885 57149
rect 843 57100 844 57140
rect 884 57100 885 57140
rect 843 57091 885 57100
rect 651 56300 693 56309
rect 651 56260 652 56300
rect 692 56260 693 56300
rect 651 56251 693 56260
rect 652 56166 692 56251
rect 940 56216 980 71464
rect 1036 57989 1076 72724
rect 3112 72596 3480 72605
rect 3152 72556 3194 72596
rect 3234 72556 3276 72596
rect 3316 72556 3358 72596
rect 3398 72556 3440 72596
rect 3112 72547 3480 72556
rect 18232 72596 18600 72605
rect 18272 72556 18314 72596
rect 18354 72556 18396 72596
rect 18436 72556 18478 72596
rect 18518 72556 18560 72596
rect 18232 72547 18600 72556
rect 33352 72596 33720 72605
rect 33392 72556 33434 72596
rect 33474 72556 33516 72596
rect 33556 72556 33598 72596
rect 33638 72556 33680 72596
rect 33352 72547 33720 72556
rect 48472 72596 48840 72605
rect 48512 72556 48554 72596
rect 48594 72556 48636 72596
rect 48676 72556 48718 72596
rect 48758 72556 48800 72596
rect 48472 72547 48840 72556
rect 63592 72596 63960 72605
rect 63632 72556 63674 72596
rect 63714 72556 63756 72596
rect 63796 72556 63838 72596
rect 63878 72556 63920 72596
rect 63592 72547 63960 72556
rect 78712 72596 79080 72605
rect 78752 72556 78794 72596
rect 78834 72556 78876 72596
rect 78916 72556 78958 72596
rect 78998 72556 79040 72596
rect 78712 72547 79080 72556
rect 93832 72596 94200 72605
rect 93872 72556 93914 72596
rect 93954 72556 93996 72596
rect 94036 72556 94078 72596
rect 94118 72556 94160 72596
rect 93832 72547 94200 72556
rect 4352 71840 4720 71849
rect 4392 71800 4434 71840
rect 4474 71800 4516 71840
rect 4556 71800 4598 71840
rect 4638 71800 4680 71840
rect 4352 71791 4720 71800
rect 19472 71840 19840 71849
rect 19512 71800 19554 71840
rect 19594 71800 19636 71840
rect 19676 71800 19718 71840
rect 19758 71800 19800 71840
rect 19472 71791 19840 71800
rect 34592 71840 34960 71849
rect 34632 71800 34674 71840
rect 34714 71800 34756 71840
rect 34796 71800 34838 71840
rect 34878 71800 34920 71840
rect 34592 71791 34960 71800
rect 49712 71840 50080 71849
rect 49752 71800 49794 71840
rect 49834 71800 49876 71840
rect 49916 71800 49958 71840
rect 49998 71800 50040 71840
rect 49712 71791 50080 71800
rect 64832 71840 65200 71849
rect 64872 71800 64914 71840
rect 64954 71800 64996 71840
rect 65036 71800 65078 71840
rect 65118 71800 65160 71840
rect 64832 71791 65200 71800
rect 79952 71840 80320 71849
rect 79992 71800 80034 71840
rect 80074 71800 80116 71840
rect 80156 71800 80198 71840
rect 80238 71800 80280 71840
rect 79952 71791 80320 71800
rect 95072 71840 95440 71849
rect 95112 71800 95154 71840
rect 95194 71800 95236 71840
rect 95276 71800 95318 71840
rect 95358 71800 95400 71840
rect 95072 71791 95440 71800
rect 3112 71084 3480 71093
rect 3152 71044 3194 71084
rect 3234 71044 3276 71084
rect 3316 71044 3358 71084
rect 3398 71044 3440 71084
rect 3112 71035 3480 71044
rect 18232 71084 18600 71093
rect 18272 71044 18314 71084
rect 18354 71044 18396 71084
rect 18436 71044 18478 71084
rect 18518 71044 18560 71084
rect 18232 71035 18600 71044
rect 33352 71084 33720 71093
rect 33392 71044 33434 71084
rect 33474 71044 33516 71084
rect 33556 71044 33598 71084
rect 33638 71044 33680 71084
rect 33352 71035 33720 71044
rect 48472 71084 48840 71093
rect 48512 71044 48554 71084
rect 48594 71044 48636 71084
rect 48676 71044 48718 71084
rect 48758 71044 48800 71084
rect 48472 71035 48840 71044
rect 63592 71084 63960 71093
rect 63632 71044 63674 71084
rect 63714 71044 63756 71084
rect 63796 71044 63838 71084
rect 63878 71044 63920 71084
rect 63592 71035 63960 71044
rect 78712 71084 79080 71093
rect 78752 71044 78794 71084
rect 78834 71044 78876 71084
rect 78916 71044 78958 71084
rect 78998 71044 79040 71084
rect 78712 71035 79080 71044
rect 93832 71084 94200 71093
rect 93872 71044 93914 71084
rect 93954 71044 93996 71084
rect 94036 71044 94078 71084
rect 94118 71044 94160 71084
rect 93832 71035 94200 71044
rect 4352 70328 4720 70337
rect 4392 70288 4434 70328
rect 4474 70288 4516 70328
rect 4556 70288 4598 70328
rect 4638 70288 4680 70328
rect 4352 70279 4720 70288
rect 19472 70328 19840 70337
rect 19512 70288 19554 70328
rect 19594 70288 19636 70328
rect 19676 70288 19718 70328
rect 19758 70288 19800 70328
rect 19472 70279 19840 70288
rect 34592 70328 34960 70337
rect 34632 70288 34674 70328
rect 34714 70288 34756 70328
rect 34796 70288 34838 70328
rect 34878 70288 34920 70328
rect 34592 70279 34960 70288
rect 49712 70328 50080 70337
rect 49752 70288 49794 70328
rect 49834 70288 49876 70328
rect 49916 70288 49958 70328
rect 49998 70288 50040 70328
rect 49712 70279 50080 70288
rect 64832 70328 65200 70337
rect 64872 70288 64914 70328
rect 64954 70288 64996 70328
rect 65036 70288 65078 70328
rect 65118 70288 65160 70328
rect 64832 70279 65200 70288
rect 79952 70328 80320 70337
rect 79992 70288 80034 70328
rect 80074 70288 80116 70328
rect 80156 70288 80198 70328
rect 80238 70288 80280 70328
rect 79952 70279 80320 70288
rect 95072 70328 95440 70337
rect 95112 70288 95154 70328
rect 95194 70288 95236 70328
rect 95276 70288 95318 70328
rect 95358 70288 95400 70328
rect 95072 70279 95440 70288
rect 3112 69572 3480 69581
rect 3152 69532 3194 69572
rect 3234 69532 3276 69572
rect 3316 69532 3358 69572
rect 3398 69532 3440 69572
rect 3112 69523 3480 69532
rect 18232 69572 18600 69581
rect 18272 69532 18314 69572
rect 18354 69532 18396 69572
rect 18436 69532 18478 69572
rect 18518 69532 18560 69572
rect 18232 69523 18600 69532
rect 33352 69572 33720 69581
rect 33392 69532 33434 69572
rect 33474 69532 33516 69572
rect 33556 69532 33598 69572
rect 33638 69532 33680 69572
rect 33352 69523 33720 69532
rect 48472 69572 48840 69581
rect 48512 69532 48554 69572
rect 48594 69532 48636 69572
rect 48676 69532 48718 69572
rect 48758 69532 48800 69572
rect 48472 69523 48840 69532
rect 63592 69572 63960 69581
rect 63632 69532 63674 69572
rect 63714 69532 63756 69572
rect 63796 69532 63838 69572
rect 63878 69532 63920 69572
rect 63592 69523 63960 69532
rect 78712 69572 79080 69581
rect 78752 69532 78794 69572
rect 78834 69532 78876 69572
rect 78916 69532 78958 69572
rect 78998 69532 79040 69572
rect 78712 69523 79080 69532
rect 93832 69572 94200 69581
rect 93872 69532 93914 69572
rect 93954 69532 93996 69572
rect 94036 69532 94078 69572
rect 94118 69532 94160 69572
rect 93832 69523 94200 69532
rect 1227 68984 1269 68993
rect 1227 68944 1228 68984
rect 1268 68944 1269 68984
rect 1227 68935 1269 68944
rect 1131 65960 1173 65969
rect 1131 65920 1132 65960
rect 1172 65920 1173 65960
rect 1131 65911 1173 65920
rect 1035 57980 1077 57989
rect 1035 57940 1036 57980
rect 1076 57940 1077 57980
rect 1035 57931 1077 57940
rect 940 56176 1076 56216
rect 747 56132 789 56141
rect 747 56092 748 56132
rect 788 56092 789 56132
rect 747 56083 789 56092
rect 844 56132 884 56141
rect 884 56092 980 56132
rect 844 56083 884 56092
rect 652 54788 692 54797
rect 652 54377 692 54748
rect 651 54368 693 54377
rect 651 54328 652 54368
rect 692 54328 693 54368
rect 651 54319 693 54328
rect 651 52604 693 52613
rect 651 52564 652 52604
rect 692 52564 693 52604
rect 651 52555 693 52564
rect 652 52470 692 52555
rect 652 51092 692 51101
rect 748 51092 788 56083
rect 844 54620 884 54629
rect 844 52529 884 54580
rect 940 52697 980 56092
rect 1036 52865 1076 56176
rect 1035 52856 1077 52865
rect 1035 52816 1036 52856
rect 1076 52816 1077 52856
rect 1035 52807 1077 52816
rect 939 52688 981 52697
rect 939 52648 940 52688
rect 980 52648 981 52688
rect 939 52639 981 52648
rect 843 52520 885 52529
rect 843 52480 844 52520
rect 884 52480 885 52520
rect 843 52471 885 52480
rect 844 52352 884 52361
rect 884 52312 1076 52352
rect 844 52303 884 52312
rect 748 51052 980 51092
rect 652 50681 692 51052
rect 844 50840 884 50849
rect 651 50672 693 50681
rect 651 50632 652 50672
rect 692 50632 693 50672
rect 651 50623 693 50632
rect 652 49580 692 49589
rect 652 48833 692 49540
rect 844 49505 884 50800
rect 843 49496 885 49505
rect 843 49456 844 49496
rect 884 49456 885 49496
rect 843 49447 885 49456
rect 844 49328 884 49337
rect 651 48824 693 48833
rect 651 48784 652 48824
rect 692 48784 693 48824
rect 651 48775 693 48784
rect 747 47900 789 47909
rect 747 47860 748 47900
rect 788 47860 789 47900
rect 747 47851 789 47860
rect 555 47312 597 47321
rect 555 47272 556 47312
rect 596 47272 597 47312
rect 555 47263 597 47272
rect 652 47228 692 47237
rect 652 46985 692 47188
rect 651 46976 693 46985
rect 651 46936 652 46976
rect 692 46936 693 46976
rect 651 46927 693 46936
rect 652 45968 692 45977
rect 652 45137 692 45928
rect 651 45128 693 45137
rect 651 45088 652 45128
rect 692 45088 693 45128
rect 651 45079 693 45088
rect 651 43280 693 43289
rect 651 43240 652 43280
rect 692 43240 693 43280
rect 651 43231 693 43240
rect 652 43146 692 43231
rect 652 41768 692 41777
rect 652 41441 692 41728
rect 748 41600 788 47851
rect 844 47573 884 49288
rect 843 47564 885 47573
rect 843 47524 844 47564
rect 884 47524 885 47564
rect 843 47515 885 47524
rect 844 47060 884 47069
rect 844 45977 884 47020
rect 940 46640 980 51052
rect 1036 47489 1076 52312
rect 1035 47480 1077 47489
rect 1035 47440 1036 47480
rect 1076 47440 1077 47480
rect 1035 47431 1077 47440
rect 940 46600 1076 46640
rect 843 45968 885 45977
rect 843 45928 844 45968
rect 884 45928 885 45968
rect 843 45919 885 45928
rect 748 41560 980 41600
rect 651 41432 693 41441
rect 651 41392 652 41432
rect 692 41392 693 41432
rect 651 41383 693 41392
rect 652 39920 692 39929
rect 652 39593 692 39880
rect 651 39584 693 39593
rect 651 39544 652 39584
rect 692 39544 693 39584
rect 651 39535 693 39544
rect 652 38408 692 38417
rect 652 37745 692 38368
rect 651 37736 693 37745
rect 651 37696 652 37736
rect 692 37696 693 37736
rect 651 37687 693 37696
rect 651 35888 693 35897
rect 651 35848 652 35888
rect 692 35848 693 35888
rect 651 35839 693 35848
rect 652 35720 692 35839
rect 652 35671 692 35680
rect 652 34208 692 34217
rect 652 34049 692 34168
rect 651 34040 693 34049
rect 651 34000 652 34040
rect 692 34000 693 34040
rect 651 33991 693 34000
rect 652 32696 692 32705
rect 652 32201 692 32656
rect 651 32192 693 32201
rect 651 32152 652 32192
rect 692 32152 693 32192
rect 651 32143 693 32152
rect 652 30848 692 30857
rect 652 30353 692 30808
rect 651 30344 693 30353
rect 651 30304 652 30344
rect 692 30304 693 30344
rect 651 30295 693 30304
rect 652 29336 692 29345
rect 652 28505 692 29296
rect 651 28496 693 28505
rect 651 28456 652 28496
rect 692 28456 693 28496
rect 651 28447 693 28456
rect 651 26648 693 26657
rect 651 26608 652 26648
rect 692 26608 693 26648
rect 651 26599 693 26608
rect 652 26514 692 26599
rect 652 25136 692 25145
rect 652 24809 692 25096
rect 651 24800 693 24809
rect 651 24760 652 24800
rect 692 24760 693 24800
rect 651 24751 693 24760
rect 652 23288 692 23297
rect 652 22961 692 23248
rect 651 22952 693 22961
rect 651 22912 652 22952
rect 692 22912 693 22952
rect 651 22903 693 22912
rect 652 21776 692 21785
rect 652 21113 692 21736
rect 651 21104 693 21113
rect 651 21064 652 21104
rect 692 21064 693 21104
rect 651 21055 693 21064
rect 651 19256 693 19265
rect 651 19216 652 19256
rect 692 19216 693 19256
rect 651 19207 693 19216
rect 652 19088 692 19207
rect 652 19039 692 19048
rect 652 17576 692 17585
rect 652 17417 692 17536
rect 651 17408 693 17417
rect 651 17368 652 17408
rect 692 17368 693 17408
rect 651 17359 693 17368
rect 843 16316 885 16325
rect 843 16276 844 16316
rect 884 16276 885 16316
rect 843 16267 885 16276
rect 844 16182 884 16267
rect 652 16064 692 16073
rect 652 15569 692 16024
rect 651 15560 693 15569
rect 651 15520 652 15560
rect 692 15520 693 15560
rect 651 15511 693 15520
rect 940 15140 980 41560
rect 748 15100 980 15140
rect 651 13796 693 13805
rect 651 13756 652 13796
rect 692 13756 693 13796
rect 651 13747 693 13756
rect 652 13662 692 13747
rect 652 12284 692 12293
rect 652 11873 692 12244
rect 651 11864 693 11873
rect 651 11824 652 11864
rect 692 11824 693 11864
rect 651 11815 693 11824
rect 651 10016 693 10025
rect 651 9976 652 10016
rect 692 9976 693 10016
rect 651 9967 693 9976
rect 652 9882 692 9967
rect 652 8504 692 8513
rect 652 8177 692 8464
rect 651 8168 693 8177
rect 651 8128 652 8168
rect 692 8128 693 8168
rect 651 8119 693 8128
rect 652 6329 692 6414
rect 748 6404 788 15100
rect 844 13964 884 13973
rect 1036 13964 1076 46600
rect 1132 45809 1172 65911
rect 1228 51857 1268 68935
rect 4352 68816 4720 68825
rect 4392 68776 4434 68816
rect 4474 68776 4516 68816
rect 4556 68776 4598 68816
rect 4638 68776 4680 68816
rect 4352 68767 4720 68776
rect 19472 68816 19840 68825
rect 19512 68776 19554 68816
rect 19594 68776 19636 68816
rect 19676 68776 19718 68816
rect 19758 68776 19800 68816
rect 19472 68767 19840 68776
rect 34592 68816 34960 68825
rect 34632 68776 34674 68816
rect 34714 68776 34756 68816
rect 34796 68776 34838 68816
rect 34878 68776 34920 68816
rect 34592 68767 34960 68776
rect 49712 68816 50080 68825
rect 49752 68776 49794 68816
rect 49834 68776 49876 68816
rect 49916 68776 49958 68816
rect 49998 68776 50040 68816
rect 49712 68767 50080 68776
rect 64832 68816 65200 68825
rect 64872 68776 64914 68816
rect 64954 68776 64996 68816
rect 65036 68776 65078 68816
rect 65118 68776 65160 68816
rect 64832 68767 65200 68776
rect 79952 68816 80320 68825
rect 79992 68776 80034 68816
rect 80074 68776 80116 68816
rect 80156 68776 80198 68816
rect 80238 68776 80280 68816
rect 79952 68767 80320 68776
rect 95072 68816 95440 68825
rect 95112 68776 95154 68816
rect 95194 68776 95236 68816
rect 95276 68776 95318 68816
rect 95358 68776 95400 68816
rect 95072 68767 95440 68776
rect 3112 68060 3480 68069
rect 3152 68020 3194 68060
rect 3234 68020 3276 68060
rect 3316 68020 3358 68060
rect 3398 68020 3440 68060
rect 3112 68011 3480 68020
rect 18232 68060 18600 68069
rect 18272 68020 18314 68060
rect 18354 68020 18396 68060
rect 18436 68020 18478 68060
rect 18518 68020 18560 68060
rect 18232 68011 18600 68020
rect 33352 68060 33720 68069
rect 33392 68020 33434 68060
rect 33474 68020 33516 68060
rect 33556 68020 33598 68060
rect 33638 68020 33680 68060
rect 33352 68011 33720 68020
rect 48472 68060 48840 68069
rect 48512 68020 48554 68060
rect 48594 68020 48636 68060
rect 48676 68020 48718 68060
rect 48758 68020 48800 68060
rect 48472 68011 48840 68020
rect 63592 68060 63960 68069
rect 63632 68020 63674 68060
rect 63714 68020 63756 68060
rect 63796 68020 63838 68060
rect 63878 68020 63920 68060
rect 63592 68011 63960 68020
rect 78712 68060 79080 68069
rect 78752 68020 78794 68060
rect 78834 68020 78876 68060
rect 78916 68020 78958 68060
rect 78998 68020 79040 68060
rect 78712 68011 79080 68020
rect 93832 68060 94200 68069
rect 93872 68020 93914 68060
rect 93954 68020 93996 68060
rect 94036 68020 94078 68060
rect 94118 68020 94160 68060
rect 93832 68011 94200 68020
rect 4352 67304 4720 67313
rect 4392 67264 4434 67304
rect 4474 67264 4516 67304
rect 4556 67264 4598 67304
rect 4638 67264 4680 67304
rect 4352 67255 4720 67264
rect 19472 67304 19840 67313
rect 19512 67264 19554 67304
rect 19594 67264 19636 67304
rect 19676 67264 19718 67304
rect 19758 67264 19800 67304
rect 19472 67255 19840 67264
rect 34592 67304 34960 67313
rect 34632 67264 34674 67304
rect 34714 67264 34756 67304
rect 34796 67264 34838 67304
rect 34878 67264 34920 67304
rect 34592 67255 34960 67264
rect 49712 67304 50080 67313
rect 49752 67264 49794 67304
rect 49834 67264 49876 67304
rect 49916 67264 49958 67304
rect 49998 67264 50040 67304
rect 49712 67255 50080 67264
rect 64832 67304 65200 67313
rect 64872 67264 64914 67304
rect 64954 67264 64996 67304
rect 65036 67264 65078 67304
rect 65118 67264 65160 67304
rect 64832 67255 65200 67264
rect 79952 67304 80320 67313
rect 79992 67264 80034 67304
rect 80074 67264 80116 67304
rect 80156 67264 80198 67304
rect 80238 67264 80280 67304
rect 79952 67255 80320 67264
rect 95072 67304 95440 67313
rect 95112 67264 95154 67304
rect 95194 67264 95236 67304
rect 95276 67264 95318 67304
rect 95358 67264 95400 67304
rect 95072 67255 95440 67264
rect 3112 66548 3480 66557
rect 3152 66508 3194 66548
rect 3234 66508 3276 66548
rect 3316 66508 3358 66548
rect 3398 66508 3440 66548
rect 3112 66499 3480 66508
rect 18232 66548 18600 66557
rect 18272 66508 18314 66548
rect 18354 66508 18396 66548
rect 18436 66508 18478 66548
rect 18518 66508 18560 66548
rect 18232 66499 18600 66508
rect 33352 66548 33720 66557
rect 33392 66508 33434 66548
rect 33474 66508 33516 66548
rect 33556 66508 33598 66548
rect 33638 66508 33680 66548
rect 33352 66499 33720 66508
rect 48472 66548 48840 66557
rect 48512 66508 48554 66548
rect 48594 66508 48636 66548
rect 48676 66508 48718 66548
rect 48758 66508 48800 66548
rect 48472 66499 48840 66508
rect 63592 66548 63960 66557
rect 63632 66508 63674 66548
rect 63714 66508 63756 66548
rect 63796 66508 63838 66548
rect 63878 66508 63920 66548
rect 63592 66499 63960 66508
rect 78712 66548 79080 66557
rect 78752 66508 78794 66548
rect 78834 66508 78876 66548
rect 78916 66508 78958 66548
rect 78998 66508 79040 66548
rect 78712 66499 79080 66508
rect 93832 66548 94200 66557
rect 93872 66508 93914 66548
rect 93954 66508 93996 66548
rect 94036 66508 94078 66548
rect 94118 66508 94160 66548
rect 93832 66499 94200 66508
rect 4352 65792 4720 65801
rect 4392 65752 4434 65792
rect 4474 65752 4516 65792
rect 4556 65752 4598 65792
rect 4638 65752 4680 65792
rect 4352 65743 4720 65752
rect 19472 65792 19840 65801
rect 19512 65752 19554 65792
rect 19594 65752 19636 65792
rect 19676 65752 19718 65792
rect 19758 65752 19800 65792
rect 19472 65743 19840 65752
rect 34592 65792 34960 65801
rect 34632 65752 34674 65792
rect 34714 65752 34756 65792
rect 34796 65752 34838 65792
rect 34878 65752 34920 65792
rect 34592 65743 34960 65752
rect 49712 65792 50080 65801
rect 49752 65752 49794 65792
rect 49834 65752 49876 65792
rect 49916 65752 49958 65792
rect 49998 65752 50040 65792
rect 49712 65743 50080 65752
rect 64832 65792 65200 65801
rect 64872 65752 64914 65792
rect 64954 65752 64996 65792
rect 65036 65752 65078 65792
rect 65118 65752 65160 65792
rect 64832 65743 65200 65752
rect 79952 65792 80320 65801
rect 79992 65752 80034 65792
rect 80074 65752 80116 65792
rect 80156 65752 80198 65792
rect 80238 65752 80280 65792
rect 79952 65743 80320 65752
rect 95072 65792 95440 65801
rect 95112 65752 95154 65792
rect 95194 65752 95236 65792
rect 95276 65752 95318 65792
rect 95358 65752 95400 65792
rect 95072 65743 95440 65752
rect 3112 65036 3480 65045
rect 3152 64996 3194 65036
rect 3234 64996 3276 65036
rect 3316 64996 3358 65036
rect 3398 64996 3440 65036
rect 3112 64987 3480 64996
rect 18232 65036 18600 65045
rect 18272 64996 18314 65036
rect 18354 64996 18396 65036
rect 18436 64996 18478 65036
rect 18518 64996 18560 65036
rect 18232 64987 18600 64996
rect 33352 65036 33720 65045
rect 33392 64996 33434 65036
rect 33474 64996 33516 65036
rect 33556 64996 33598 65036
rect 33638 64996 33680 65036
rect 33352 64987 33720 64996
rect 48472 65036 48840 65045
rect 48512 64996 48554 65036
rect 48594 64996 48636 65036
rect 48676 64996 48718 65036
rect 48758 64996 48800 65036
rect 48472 64987 48840 64996
rect 63592 65036 63960 65045
rect 63632 64996 63674 65036
rect 63714 64996 63756 65036
rect 63796 64996 63838 65036
rect 63878 64996 63920 65036
rect 63592 64987 63960 64996
rect 78712 65036 79080 65045
rect 78752 64996 78794 65036
rect 78834 64996 78876 65036
rect 78916 64996 78958 65036
rect 78998 64996 79040 65036
rect 78712 64987 79080 64996
rect 93832 65036 94200 65045
rect 93872 64996 93914 65036
rect 93954 64996 93996 65036
rect 94036 64996 94078 65036
rect 94118 64996 94160 65036
rect 93832 64987 94200 64996
rect 4352 64280 4720 64289
rect 4392 64240 4434 64280
rect 4474 64240 4516 64280
rect 4556 64240 4598 64280
rect 4638 64240 4680 64280
rect 4352 64231 4720 64240
rect 19472 64280 19840 64289
rect 19512 64240 19554 64280
rect 19594 64240 19636 64280
rect 19676 64240 19718 64280
rect 19758 64240 19800 64280
rect 19472 64231 19840 64240
rect 34592 64280 34960 64289
rect 34632 64240 34674 64280
rect 34714 64240 34756 64280
rect 34796 64240 34838 64280
rect 34878 64240 34920 64280
rect 34592 64231 34960 64240
rect 49712 64280 50080 64289
rect 49752 64240 49794 64280
rect 49834 64240 49876 64280
rect 49916 64240 49958 64280
rect 49998 64240 50040 64280
rect 49712 64231 50080 64240
rect 64832 64280 65200 64289
rect 64872 64240 64914 64280
rect 64954 64240 64996 64280
rect 65036 64240 65078 64280
rect 65118 64240 65160 64280
rect 64832 64231 65200 64240
rect 79952 64280 80320 64289
rect 79992 64240 80034 64280
rect 80074 64240 80116 64280
rect 80156 64240 80198 64280
rect 80238 64240 80280 64280
rect 79952 64231 80320 64240
rect 95072 64280 95440 64289
rect 95112 64240 95154 64280
rect 95194 64240 95236 64280
rect 95276 64240 95318 64280
rect 95358 64240 95400 64280
rect 95072 64231 95440 64240
rect 13227 63692 13269 63701
rect 13227 63652 13228 63692
rect 13268 63652 13269 63692
rect 13227 63643 13269 63652
rect 3112 63524 3480 63533
rect 3152 63484 3194 63524
rect 3234 63484 3276 63524
rect 3316 63484 3358 63524
rect 3398 63484 3440 63524
rect 3112 63475 3480 63484
rect 6507 63020 6549 63029
rect 6507 62980 6508 63020
rect 6548 62980 6549 63020
rect 6507 62971 6549 62980
rect 4352 62768 4720 62777
rect 4392 62728 4434 62768
rect 4474 62728 4516 62768
rect 4556 62728 4598 62768
rect 4638 62728 4680 62768
rect 4352 62719 4720 62728
rect 3112 62012 3480 62021
rect 3152 61972 3194 62012
rect 3234 61972 3276 62012
rect 3316 61972 3358 62012
rect 3398 61972 3440 62012
rect 3112 61963 3480 61972
rect 4352 61256 4720 61265
rect 4392 61216 4434 61256
rect 4474 61216 4516 61256
rect 4556 61216 4598 61256
rect 4638 61216 4680 61256
rect 4352 61207 4720 61216
rect 6508 60920 6548 62971
rect 6508 60871 6548 60880
rect 6604 60920 6644 60929
rect 3112 60500 3480 60509
rect 3152 60460 3194 60500
rect 3234 60460 3276 60500
rect 3316 60460 3358 60500
rect 3398 60460 3440 60500
rect 3112 60451 3480 60460
rect 6604 60341 6644 60880
rect 6892 60836 6932 60845
rect 6603 60332 6645 60341
rect 6603 60292 6604 60332
rect 6644 60292 6645 60332
rect 6603 60283 6645 60292
rect 6796 60080 6836 60089
rect 6508 59912 6548 59921
rect 4352 59744 4720 59753
rect 4392 59704 4434 59744
rect 4474 59704 4516 59744
rect 4556 59704 4598 59744
rect 4638 59704 4680 59744
rect 4352 59695 4720 59704
rect 6508 59240 6548 59872
rect 6412 59200 6548 59240
rect 6796 59240 6836 60040
rect 6892 60080 6932 60796
rect 6892 60031 6932 60040
rect 6796 59200 7316 59240
rect 3112 58988 3480 58997
rect 3152 58948 3194 58988
rect 3234 58948 3276 58988
rect 3316 58948 3358 58988
rect 3398 58948 3440 58988
rect 3112 58939 3480 58948
rect 4352 58232 4720 58241
rect 4392 58192 4434 58232
rect 4474 58192 4516 58232
rect 4556 58192 4598 58232
rect 4638 58192 4680 58232
rect 4352 58183 4720 58192
rect 5835 57980 5877 57989
rect 5835 57940 5836 57980
rect 5876 57940 5877 57980
rect 5835 57931 5877 57940
rect 3112 57476 3480 57485
rect 3152 57436 3194 57476
rect 3234 57436 3276 57476
rect 3316 57436 3358 57476
rect 3398 57436 3440 57476
rect 3112 57427 3480 57436
rect 5836 57056 5876 57931
rect 6219 57896 6261 57905
rect 6219 57856 6220 57896
rect 6260 57856 6261 57896
rect 6219 57847 6261 57856
rect 6315 57896 6357 57905
rect 6315 57856 6316 57896
rect 6356 57856 6357 57896
rect 6315 57847 6357 57856
rect 6220 57149 6260 57847
rect 6316 57762 6356 57847
rect 6412 57224 6452 59200
rect 6508 57905 6548 57990
rect 6507 57896 6549 57905
rect 6507 57856 6508 57896
rect 6548 57856 6549 57896
rect 6507 57847 6549 57856
rect 6508 57644 6548 57653
rect 6548 57604 7124 57644
rect 6508 57595 6548 57604
rect 6412 57184 6836 57224
rect 6027 57140 6069 57149
rect 6219 57140 6261 57149
rect 6027 57100 6028 57140
rect 6068 57100 6071 57140
rect 6027 57091 6071 57100
rect 6219 57100 6220 57140
rect 6260 57100 6261 57140
rect 6219 57091 6261 57100
rect 6031 57079 6071 57091
rect 5836 56981 5876 57016
rect 5931 57056 5973 57065
rect 5931 57016 5932 57056
rect 5972 57016 5973 57056
rect 5931 57007 5973 57016
rect 6031 57008 6071 57039
rect 6220 57056 6260 57091
rect 5835 56972 5877 56981
rect 5835 56932 5836 56972
rect 5876 56932 5877 56972
rect 5835 56923 5877 56932
rect 5836 56921 5876 56923
rect 5932 56922 5972 57007
rect 6220 57005 6260 57016
rect 6507 57056 6549 57065
rect 6507 57016 6508 57056
rect 6548 57016 6549 57056
rect 6507 57007 6549 57016
rect 6508 56922 6548 57007
rect 6700 56888 6740 56897
rect 4352 56720 4720 56729
rect 4392 56680 4434 56720
rect 4474 56680 4516 56720
rect 4556 56680 4598 56720
rect 4638 56680 4680 56720
rect 4352 56671 4720 56680
rect 5643 56384 5685 56393
rect 5643 56344 5644 56384
rect 5684 56344 5685 56384
rect 5643 56335 5685 56344
rect 6603 56384 6645 56393
rect 6603 56344 6604 56384
rect 6644 56344 6645 56384
rect 6603 56335 6645 56344
rect 6700 56384 6740 56848
rect 6700 56335 6740 56344
rect 3112 55964 3480 55973
rect 3152 55924 3194 55964
rect 3234 55924 3276 55964
rect 3316 55924 3358 55964
rect 3398 55924 3440 55964
rect 3112 55915 3480 55924
rect 4352 55208 4720 55217
rect 4392 55168 4434 55208
rect 4474 55168 4516 55208
rect 4556 55168 4598 55208
rect 4638 55168 4680 55208
rect 4352 55159 4720 55168
rect 3112 54452 3480 54461
rect 3152 54412 3194 54452
rect 3234 54412 3276 54452
rect 3316 54412 3358 54452
rect 3398 54412 3440 54452
rect 3112 54403 3480 54412
rect 4352 53696 4720 53705
rect 4392 53656 4434 53696
rect 4474 53656 4516 53696
rect 4556 53656 4598 53696
rect 4638 53656 4680 53696
rect 4352 53647 4720 53656
rect 3112 52940 3480 52949
rect 3152 52900 3194 52940
rect 3234 52900 3276 52940
rect 3316 52900 3358 52940
rect 3398 52900 3440 52940
rect 3112 52891 3480 52900
rect 5644 52772 5684 56335
rect 6604 56250 6644 56335
rect 6796 56216 6836 57184
rect 6988 57056 7028 57065
rect 6988 56393 7028 57016
rect 7084 57056 7124 57604
rect 7084 57007 7124 57016
rect 7179 57056 7221 57065
rect 7179 57016 7180 57056
rect 7220 57016 7221 57056
rect 7179 57007 7221 57016
rect 7276 57056 7316 59200
rect 7276 57007 7316 57016
rect 7180 56922 7220 57007
rect 6987 56384 7029 56393
rect 6987 56344 6988 56384
rect 7028 56344 7029 56384
rect 6987 56335 7029 56344
rect 6796 56176 7124 56216
rect 6411 56132 6453 56141
rect 6411 56092 6412 56132
rect 6452 56092 6453 56132
rect 6411 56083 6453 56092
rect 6412 55998 6452 56083
rect 6412 53360 6452 53369
rect 6604 53360 6644 53369
rect 6452 53320 6548 53360
rect 6412 53311 6452 53320
rect 5835 53108 5877 53117
rect 5835 53068 5836 53108
rect 5876 53068 5877 53108
rect 5835 53059 5877 53068
rect 6411 53108 6453 53117
rect 6411 53068 6412 53108
rect 6452 53068 6453 53108
rect 6411 53059 6453 53068
rect 5644 52723 5684 52732
rect 5739 52604 5781 52613
rect 5739 52564 5740 52604
rect 5780 52564 5781 52604
rect 5739 52555 5781 52564
rect 2283 52520 2325 52529
rect 2283 52480 2284 52520
rect 2324 52480 2325 52520
rect 2283 52471 2325 52480
rect 4107 52520 4149 52529
rect 4107 52480 4108 52520
rect 4148 52480 4149 52520
rect 4107 52471 4149 52480
rect 5644 52520 5684 52529
rect 2187 52016 2229 52025
rect 2187 51976 2188 52016
rect 2228 51976 2229 52016
rect 2187 51967 2229 51976
rect 2188 51932 2228 51967
rect 2188 51881 2228 51892
rect 1227 51848 1269 51857
rect 1227 51808 1228 51848
rect 1268 51808 1269 51848
rect 1227 51799 1269 51808
rect 2091 51848 2133 51857
rect 2091 51808 2092 51848
rect 2132 51808 2133 51848
rect 2091 51799 2133 51808
rect 2284 51848 2324 52471
rect 3243 52016 3285 52025
rect 3243 51976 3244 52016
rect 3284 51976 3285 52016
rect 3243 51967 3285 51976
rect 2955 51932 2997 51941
rect 2955 51892 2956 51932
rect 2996 51892 2997 51932
rect 2955 51883 2997 51892
rect 2476 51848 2516 51857
rect 2324 51808 2476 51848
rect 2284 51799 2324 51808
rect 2476 51799 2516 51808
rect 2763 51848 2805 51857
rect 2763 51808 2764 51848
rect 2804 51808 2805 51848
rect 2763 51799 2805 51808
rect 2092 51714 2132 51799
rect 2764 51714 2804 51799
rect 2956 51798 2996 51883
rect 3244 51848 3284 51967
rect 3915 51932 3957 51941
rect 3915 51892 3916 51932
rect 3956 51892 3957 51932
rect 3915 51883 3957 51892
rect 3244 51799 3284 51808
rect 3435 51848 3477 51857
rect 3435 51808 3436 51848
rect 3476 51808 3477 51848
rect 3435 51799 3477 51808
rect 3916 51848 3956 51883
rect 3436 51714 3476 51799
rect 3916 51797 3956 51808
rect 4011 51848 4053 51857
rect 4011 51808 4012 51848
rect 4052 51808 4053 51848
rect 4011 51799 4053 51808
rect 4108 51848 4148 52471
rect 4352 52184 4720 52193
rect 4392 52144 4434 52184
rect 4474 52144 4516 52184
rect 4556 52144 4598 52184
rect 4638 52144 4680 52184
rect 4352 52135 4720 52144
rect 5547 52016 5589 52025
rect 5547 51976 5548 52016
rect 5588 51976 5589 52016
rect 5547 51967 5589 51976
rect 5644 52016 5684 52480
rect 5740 52520 5780 52555
rect 5740 52469 5780 52480
rect 5644 51967 5684 51976
rect 4108 51799 4148 51808
rect 5259 51848 5301 51857
rect 5259 51808 5260 51848
rect 5300 51808 5301 51848
rect 5259 51799 5301 51808
rect 5356 51848 5396 51857
rect 5451 51848 5493 51857
rect 5396 51808 5452 51848
rect 5492 51808 5493 51848
rect 5356 51799 5396 51808
rect 5451 51799 5493 51808
rect 5548 51848 5588 51967
rect 5548 51799 5588 51808
rect 5740 51848 5780 51857
rect 5836 51848 5876 53059
rect 6412 52974 6452 53059
rect 6508 52865 6548 53320
rect 6644 53320 6740 53360
rect 6604 53311 6644 53320
rect 6184 52856 6226 52865
rect 6184 52816 6185 52856
rect 6225 52816 6226 52856
rect 6184 52807 6226 52816
rect 6507 52856 6549 52865
rect 6507 52816 6508 52856
rect 6548 52816 6549 52856
rect 6507 52807 6549 52816
rect 6027 52688 6069 52697
rect 6027 52648 6028 52688
rect 6068 52648 6069 52688
rect 6027 52639 6069 52648
rect 5931 52520 5973 52529
rect 5931 52480 5932 52520
rect 5972 52480 5973 52520
rect 5931 52471 5973 52480
rect 6028 52520 6068 52639
rect 6185 52535 6225 52807
rect 6315 52604 6357 52613
rect 6315 52564 6316 52604
rect 6356 52564 6357 52604
rect 6315 52555 6357 52564
rect 6185 52486 6225 52495
rect 6028 52471 6068 52480
rect 5780 51808 5876 51848
rect 5740 51799 5780 51808
rect 4012 51714 4052 51799
rect 5260 51714 5300 51799
rect 5932 51773 5972 52471
rect 6219 52352 6261 52361
rect 6219 52312 6220 52352
rect 6260 52312 6261 52352
rect 6219 52303 6261 52312
rect 6220 51848 6260 52303
rect 6316 52016 6356 52555
rect 6508 52520 6548 52807
rect 6700 52697 6740 53320
rect 6699 52688 6741 52697
rect 6699 52648 6700 52688
rect 6740 52648 6741 52688
rect 6699 52639 6741 52648
rect 6604 52520 6644 52529
rect 6508 52480 6604 52520
rect 6604 52471 6644 52480
rect 6700 52520 6740 52639
rect 6700 52471 6740 52480
rect 6411 52352 6453 52361
rect 6411 52312 6412 52352
rect 6452 52312 6453 52352
rect 6411 52303 6453 52312
rect 6412 52218 6452 52303
rect 6316 51967 6356 51976
rect 5931 51764 5973 51773
rect 5931 51724 5932 51764
rect 5972 51724 5973 51764
rect 5931 51715 5973 51724
rect 6123 51764 6165 51773
rect 6123 51724 6124 51764
rect 6164 51724 6165 51764
rect 6123 51715 6165 51724
rect 2667 51680 2709 51689
rect 2667 51640 2668 51680
rect 2708 51640 2709 51680
rect 2667 51631 2709 51640
rect 2668 51008 2708 51631
rect 3340 51596 3380 51605
rect 2860 51556 3340 51596
rect 2764 51008 2804 51017
rect 2668 50968 2764 51008
rect 2764 50959 2804 50968
rect 2860 51008 2900 51556
rect 3340 51547 3380 51556
rect 3112 51428 3480 51437
rect 3152 51388 3194 51428
rect 3234 51388 3276 51428
rect 3316 51388 3358 51428
rect 3398 51388 3440 51428
rect 3112 51379 3480 51388
rect 2860 50959 2900 50968
rect 1899 50840 1941 50849
rect 1899 50800 1900 50840
rect 1940 50800 1941 50840
rect 1899 50791 1941 50800
rect 2475 50840 2517 50849
rect 2475 50800 2476 50840
rect 2516 50800 2517 50840
rect 2475 50791 2517 50800
rect 1131 45800 1173 45809
rect 1131 45760 1132 45800
rect 1172 45760 1173 45800
rect 1131 45751 1173 45760
rect 1131 44792 1173 44801
rect 1131 44752 1132 44792
rect 1172 44752 1173 44792
rect 1131 44743 1173 44752
rect 884 13924 1076 13964
rect 844 13915 884 13924
rect 843 12452 885 12461
rect 843 12412 844 12452
rect 884 12412 885 12452
rect 843 12403 885 12412
rect 844 12318 884 12403
rect 843 10268 885 10277
rect 843 10228 844 10268
rect 884 10228 885 10268
rect 843 10219 885 10228
rect 844 10134 884 10219
rect 843 8756 885 8765
rect 843 8716 844 8756
rect 884 8716 885 8756
rect 843 8707 885 8716
rect 844 8622 884 8707
rect 844 6404 884 6413
rect 748 6364 844 6404
rect 844 6355 884 6364
rect 651 6320 693 6329
rect 651 6280 652 6320
rect 692 6280 693 6320
rect 651 6271 693 6280
rect 843 4892 885 4901
rect 843 4852 844 4892
rect 884 4852 885 4892
rect 843 4843 885 4852
rect 844 4758 884 4843
rect 652 4724 692 4733
rect 652 4481 692 4684
rect 651 4472 693 4481
rect 651 4432 652 4472
rect 692 4432 693 4472
rect 651 4423 693 4432
rect 652 2792 692 2801
rect 652 2633 692 2752
rect 844 2708 884 2717
rect 1132 2708 1172 44743
rect 1900 12461 1940 50791
rect 2476 50706 2516 50791
rect 4352 50672 4720 50681
rect 4392 50632 4434 50672
rect 4474 50632 4516 50672
rect 4556 50632 4598 50672
rect 4638 50632 4680 50672
rect 4352 50623 4720 50632
rect 3112 49916 3480 49925
rect 3152 49876 3194 49916
rect 3234 49876 3276 49916
rect 3316 49876 3358 49916
rect 3398 49876 3440 49916
rect 3112 49867 3480 49876
rect 4352 49160 4720 49169
rect 4392 49120 4434 49160
rect 4474 49120 4516 49160
rect 4556 49120 4598 49160
rect 4638 49120 4680 49160
rect 4352 49111 4720 49120
rect 3112 48404 3480 48413
rect 3152 48364 3194 48404
rect 3234 48364 3276 48404
rect 3316 48364 3358 48404
rect 3398 48364 3440 48404
rect 3112 48355 3480 48364
rect 3915 47984 3957 47993
rect 3915 47944 3916 47984
rect 3956 47944 3957 47984
rect 3915 47935 3957 47944
rect 6124 47984 6164 51715
rect 6220 51689 6260 51808
rect 6411 51848 6453 51857
rect 6411 51808 6412 51848
rect 6452 51808 6453 51848
rect 6411 51799 6453 51808
rect 6795 51848 6837 51857
rect 6795 51808 6796 51848
rect 6836 51808 6837 51848
rect 6795 51799 6837 51808
rect 6892 51848 6932 51857
rect 6412 51714 6452 51799
rect 6796 51714 6836 51799
rect 6892 51689 6932 51808
rect 6219 51680 6261 51689
rect 6219 51640 6220 51680
rect 6260 51640 6261 51680
rect 6219 51631 6261 51640
rect 6891 51680 6933 51689
rect 6891 51640 6892 51680
rect 6932 51640 6933 51680
rect 6891 51631 6933 51640
rect 6700 51596 6740 51605
rect 6124 47935 6164 47944
rect 6219 47984 6261 47993
rect 6219 47944 6220 47984
rect 6260 47944 6261 47984
rect 6219 47935 6261 47944
rect 6316 47984 6356 47993
rect 1995 47480 2037 47489
rect 1995 47440 1996 47480
rect 2036 47440 2037 47480
rect 1995 47431 2037 47440
rect 2283 47480 2325 47489
rect 2283 47440 2284 47480
rect 2324 47440 2325 47480
rect 2283 47431 2325 47440
rect 3916 47480 3956 47935
rect 6220 47850 6260 47935
rect 4352 47648 4720 47657
rect 4392 47608 4434 47648
rect 4474 47608 4516 47648
rect 4556 47608 4598 47648
rect 4638 47608 4680 47648
rect 4352 47599 4720 47608
rect 3916 47431 3956 47440
rect 4011 47480 4053 47489
rect 4011 47440 4012 47480
rect 4052 47440 4053 47480
rect 4011 47431 4053 47440
rect 6316 47480 6356 47944
rect 6411 47984 6453 47993
rect 6411 47944 6412 47984
rect 6452 47944 6453 47984
rect 6411 47935 6453 47944
rect 6412 47850 6452 47935
rect 6316 47431 6356 47440
rect 1996 47346 2036 47431
rect 2284 47346 2324 47431
rect 2475 47396 2517 47405
rect 2475 47356 2476 47396
rect 2516 47356 2517 47396
rect 2475 47347 2517 47356
rect 2955 47396 2997 47405
rect 2955 47356 2956 47396
rect 2996 47356 2997 47396
rect 2955 47347 2997 47356
rect 2091 47312 2133 47321
rect 2091 47272 2092 47312
rect 2132 47272 2133 47312
rect 2091 47263 2133 47272
rect 2476 47312 2516 47347
rect 2092 47178 2132 47263
rect 2476 47228 2516 47272
rect 2763 47312 2805 47321
rect 2763 47272 2764 47312
rect 2804 47272 2805 47312
rect 2763 47263 2805 47272
rect 2476 47188 2612 47228
rect 2572 46472 2612 47188
rect 2668 46640 2708 46649
rect 2764 46640 2804 47263
rect 2956 47262 2996 47347
rect 3724 47312 3764 47321
rect 3244 47272 3724 47312
rect 3244 47060 3284 47272
rect 3724 47263 3764 47272
rect 3820 47312 3860 47321
rect 3820 47153 3860 47272
rect 4012 47312 4052 47431
rect 5835 47396 5877 47405
rect 5835 47356 5836 47396
rect 5876 47356 5877 47396
rect 5835 47347 5877 47356
rect 6603 47396 6645 47405
rect 6603 47356 6604 47396
rect 6644 47356 6645 47396
rect 6603 47347 6645 47356
rect 4012 47263 4052 47272
rect 5836 47312 5876 47347
rect 5836 47261 5876 47272
rect 5932 47312 5972 47323
rect 5932 47237 5972 47272
rect 6507 47312 6549 47321
rect 6507 47272 6508 47312
rect 6548 47272 6549 47312
rect 6507 47263 6549 47272
rect 6604 47312 6644 47347
rect 5931 47228 5973 47237
rect 5931 47188 5932 47228
rect 5972 47188 5973 47228
rect 5931 47179 5973 47188
rect 6508 47178 6548 47263
rect 6604 47261 6644 47272
rect 3819 47144 3861 47153
rect 3819 47104 3820 47144
rect 3860 47104 3861 47144
rect 3819 47095 3861 47104
rect 2860 47020 3284 47060
rect 5644 47060 5684 47069
rect 2860 46724 2900 47020
rect 3112 46892 3480 46901
rect 3152 46852 3194 46892
rect 3234 46852 3276 46892
rect 3316 46852 3358 46892
rect 3398 46852 3440 46892
rect 3112 46843 3480 46852
rect 2860 46675 2900 46684
rect 2708 46600 2804 46640
rect 2668 46591 2708 46600
rect 2668 46472 2708 46481
rect 2572 46432 2668 46472
rect 2668 46423 2708 46432
rect 4352 46136 4720 46145
rect 4392 46096 4434 46136
rect 4474 46096 4516 46136
rect 4556 46096 4598 46136
rect 4638 46096 4680 46136
rect 4352 46087 4720 46096
rect 3112 45380 3480 45389
rect 3152 45340 3194 45380
rect 3234 45340 3276 45380
rect 3316 45340 3358 45380
rect 3398 45340 3440 45380
rect 3112 45331 3480 45340
rect 4352 44624 4720 44633
rect 4392 44584 4434 44624
rect 4474 44584 4516 44624
rect 4556 44584 4598 44624
rect 4638 44584 4680 44624
rect 4352 44575 4720 44584
rect 3112 43868 3480 43877
rect 3152 43828 3194 43868
rect 3234 43828 3276 43868
rect 3316 43828 3358 43868
rect 3398 43828 3440 43868
rect 3112 43819 3480 43828
rect 4352 43112 4720 43121
rect 4392 43072 4434 43112
rect 4474 43072 4516 43112
rect 4556 43072 4598 43112
rect 4638 43072 4680 43112
rect 4352 43063 4720 43072
rect 3112 42356 3480 42365
rect 3152 42316 3194 42356
rect 3234 42316 3276 42356
rect 3316 42316 3358 42356
rect 3398 42316 3440 42356
rect 3112 42307 3480 42316
rect 4352 41600 4720 41609
rect 4392 41560 4434 41600
rect 4474 41560 4516 41600
rect 4556 41560 4598 41600
rect 4638 41560 4680 41600
rect 4352 41551 4720 41560
rect 3112 40844 3480 40853
rect 3152 40804 3194 40844
rect 3234 40804 3276 40844
rect 3316 40804 3358 40844
rect 3398 40804 3440 40844
rect 3112 40795 3480 40804
rect 4352 40088 4720 40097
rect 4392 40048 4434 40088
rect 4474 40048 4516 40088
rect 4556 40048 4598 40088
rect 4638 40048 4680 40088
rect 4352 40039 4720 40048
rect 3112 39332 3480 39341
rect 3152 39292 3194 39332
rect 3234 39292 3276 39332
rect 3316 39292 3358 39332
rect 3398 39292 3440 39332
rect 3112 39283 3480 39292
rect 4352 38576 4720 38585
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4352 38527 4720 38536
rect 3112 37820 3480 37829
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3112 37771 3480 37780
rect 4352 37064 4720 37073
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4352 37015 4720 37024
rect 3112 36308 3480 36317
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3112 36259 3480 36268
rect 4352 35552 4720 35561
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4352 35503 4720 35512
rect 3112 34796 3480 34805
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3112 34747 3480 34756
rect 4352 34040 4720 34049
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4352 33991 4720 34000
rect 3112 33284 3480 33293
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3112 33235 3480 33244
rect 4352 32528 4720 32537
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4352 32479 4720 32488
rect 3112 31772 3480 31781
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3112 31723 3480 31732
rect 4352 31016 4720 31025
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4352 30967 4720 30976
rect 3112 30260 3480 30269
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3112 30211 3480 30220
rect 4352 29504 4720 29513
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4352 29455 4720 29464
rect 3112 28748 3480 28757
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3112 28699 3480 28708
rect 4352 27992 4720 28001
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4352 27943 4720 27952
rect 3112 27236 3480 27245
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3112 27187 3480 27196
rect 4352 26480 4720 26489
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4352 26431 4720 26440
rect 3112 25724 3480 25733
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3112 25675 3480 25684
rect 4352 24968 4720 24977
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4352 24919 4720 24928
rect 3112 24212 3480 24221
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3112 24163 3480 24172
rect 4352 23456 4720 23465
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4352 23407 4720 23416
rect 3112 22700 3480 22709
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3112 22651 3480 22660
rect 4352 21944 4720 21953
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4352 21895 4720 21904
rect 3112 21188 3480 21197
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3112 21139 3480 21148
rect 4352 20432 4720 20441
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4352 20383 4720 20392
rect 3112 19676 3480 19685
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3112 19627 3480 19636
rect 4352 18920 4720 18929
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4352 18871 4720 18880
rect 3112 18164 3480 18173
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3112 18115 3480 18124
rect 4352 17408 4720 17417
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4352 17359 4720 17368
rect 3112 16652 3480 16661
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3112 16603 3480 16612
rect 4352 15896 4720 15905
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4352 15847 4720 15856
rect 3112 15140 3480 15149
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3112 15091 3480 15100
rect 4352 14384 4720 14393
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4352 14335 4720 14344
rect 3112 13628 3480 13637
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3112 13579 3480 13588
rect 4352 12872 4720 12881
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4352 12823 4720 12832
rect 1899 12452 1941 12461
rect 1899 12412 1900 12452
rect 1940 12412 1941 12452
rect 1899 12403 1941 12412
rect 3112 12116 3480 12125
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3112 12067 3480 12076
rect 4352 11360 4720 11369
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4352 11311 4720 11320
rect 3112 10604 3480 10613
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3112 10555 3480 10564
rect 4352 9848 4720 9857
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4352 9799 4720 9808
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 5644 8765 5684 47020
rect 6700 10277 6740 51556
rect 6796 47312 6836 47321
rect 6796 47069 6836 47272
rect 6988 47312 7028 47321
rect 6891 47228 6933 47237
rect 6891 47188 6892 47228
rect 6932 47188 6933 47228
rect 6891 47179 6933 47188
rect 6892 47094 6932 47179
rect 6988 47153 7028 47272
rect 6987 47144 7029 47153
rect 6987 47104 6988 47144
rect 7028 47104 7029 47144
rect 6987 47095 7029 47104
rect 6795 47060 6837 47069
rect 6795 47020 6796 47060
rect 6836 47020 6837 47060
rect 6795 47011 6837 47020
rect 7084 16325 7124 56176
rect 7851 49496 7893 49505
rect 7851 49456 7852 49496
rect 7892 49456 7893 49496
rect 7851 49447 7893 49456
rect 7563 47984 7605 47993
rect 7563 47944 7564 47984
rect 7604 47944 7605 47984
rect 7563 47935 7605 47944
rect 7372 47321 7412 47406
rect 7371 47312 7413 47321
rect 7371 47272 7372 47312
rect 7412 47272 7413 47312
rect 7371 47263 7413 47272
rect 7564 47312 7604 47935
rect 7564 47263 7604 47272
rect 7371 47144 7413 47153
rect 7371 47104 7372 47144
rect 7412 47104 7413 47144
rect 7371 47095 7413 47104
rect 7372 47010 7412 47095
rect 7563 47060 7605 47069
rect 7563 47020 7564 47060
rect 7604 47020 7605 47060
rect 7563 47011 7605 47020
rect 7564 45968 7604 47011
rect 7564 45919 7604 45928
rect 7852 45968 7892 49447
rect 9484 47984 9524 47993
rect 9387 47900 9429 47909
rect 9387 47860 9388 47900
rect 9428 47860 9429 47900
rect 9387 47851 9429 47860
rect 9388 47766 9428 47851
rect 9484 47321 9524 47944
rect 9867 47984 9909 47993
rect 9867 47944 9868 47984
rect 9908 47944 9909 47984
rect 9867 47935 9909 47944
rect 9868 47850 9908 47935
rect 13131 47564 13173 47573
rect 13131 47524 13132 47564
rect 13172 47524 13173 47564
rect 13131 47515 13173 47524
rect 13132 47480 13172 47515
rect 13132 47429 13172 47440
rect 13228 47321 13268 63643
rect 18232 63524 18600 63533
rect 18272 63484 18314 63524
rect 18354 63484 18396 63524
rect 18436 63484 18478 63524
rect 18518 63484 18560 63524
rect 18232 63475 18600 63484
rect 33352 63524 33720 63533
rect 33392 63484 33434 63524
rect 33474 63484 33516 63524
rect 33556 63484 33598 63524
rect 33638 63484 33680 63524
rect 33352 63475 33720 63484
rect 48472 63524 48840 63533
rect 48512 63484 48554 63524
rect 48594 63484 48636 63524
rect 48676 63484 48718 63524
rect 48758 63484 48800 63524
rect 48472 63475 48840 63484
rect 63592 63524 63960 63533
rect 63632 63484 63674 63524
rect 63714 63484 63756 63524
rect 63796 63484 63838 63524
rect 63878 63484 63920 63524
rect 63592 63475 63960 63484
rect 78712 63524 79080 63533
rect 78752 63484 78794 63524
rect 78834 63484 78876 63524
rect 78916 63484 78958 63524
rect 78998 63484 79040 63524
rect 78712 63475 79080 63484
rect 93832 63524 94200 63533
rect 93872 63484 93914 63524
rect 93954 63484 93996 63524
rect 94036 63484 94078 63524
rect 94118 63484 94160 63524
rect 93832 63475 94200 63484
rect 19472 62768 19840 62777
rect 19512 62728 19554 62768
rect 19594 62728 19636 62768
rect 19676 62728 19718 62768
rect 19758 62728 19800 62768
rect 19472 62719 19840 62728
rect 34592 62768 34960 62777
rect 34632 62728 34674 62768
rect 34714 62728 34756 62768
rect 34796 62728 34838 62768
rect 34878 62728 34920 62768
rect 34592 62719 34960 62728
rect 49712 62768 50080 62777
rect 49752 62728 49794 62768
rect 49834 62728 49876 62768
rect 49916 62728 49958 62768
rect 49998 62728 50040 62768
rect 49712 62719 50080 62728
rect 64832 62768 65200 62777
rect 64872 62728 64914 62768
rect 64954 62728 64996 62768
rect 65036 62728 65078 62768
rect 65118 62728 65160 62768
rect 64832 62719 65200 62728
rect 79952 62768 80320 62777
rect 79992 62728 80034 62768
rect 80074 62728 80116 62768
rect 80156 62728 80198 62768
rect 80238 62728 80280 62768
rect 79952 62719 80320 62728
rect 95072 62768 95440 62777
rect 95112 62728 95154 62768
rect 95194 62728 95236 62768
rect 95276 62728 95318 62768
rect 95358 62728 95400 62768
rect 95072 62719 95440 62728
rect 14187 62180 14229 62189
rect 14187 62140 14188 62180
rect 14228 62140 14229 62180
rect 14187 62131 14229 62140
rect 13803 47984 13845 47993
rect 13803 47944 13804 47984
rect 13844 47944 13845 47984
rect 13803 47935 13845 47944
rect 13611 47564 13653 47573
rect 13611 47524 13612 47564
rect 13652 47524 13653 47564
rect 13611 47515 13653 47524
rect 8043 47312 8085 47321
rect 8043 47272 8044 47312
rect 8084 47272 8085 47312
rect 8043 47263 8085 47272
rect 9483 47312 9525 47321
rect 9483 47272 9484 47312
rect 9524 47272 9525 47312
rect 9483 47263 9525 47272
rect 13227 47312 13269 47321
rect 13227 47272 13228 47312
rect 13268 47272 13269 47312
rect 13227 47263 13269 47272
rect 13612 47312 13652 47515
rect 13612 47263 13652 47272
rect 8044 45968 8084 47263
rect 13228 47178 13268 47263
rect 13420 47060 13460 47069
rect 13460 47020 13748 47060
rect 13420 47011 13460 47020
rect 13708 46556 13748 47020
rect 13804 46640 13844 47935
rect 14092 47396 14132 47407
rect 14092 47321 14132 47356
rect 13899 47312 13941 47321
rect 13899 47272 13900 47312
rect 13940 47272 13941 47312
rect 13899 47263 13941 47272
rect 14091 47312 14133 47321
rect 14091 47272 14092 47312
rect 14132 47272 14133 47312
rect 14091 47263 14133 47272
rect 13900 47178 13940 47263
rect 13804 46591 13844 46600
rect 13708 46507 13748 46516
rect 14091 46472 14133 46481
rect 14091 46432 14092 46472
rect 14132 46432 14133 46472
rect 14091 46423 14133 46432
rect 14092 46338 14132 46423
rect 14091 45968 14133 45977
rect 7892 45928 7988 45968
rect 7852 45919 7892 45928
rect 7755 45800 7797 45809
rect 7755 45760 7756 45800
rect 7796 45760 7797 45800
rect 7948 45800 7988 45928
rect 8044 45919 8084 45928
rect 8140 45928 8372 45968
rect 8140 45800 8180 45928
rect 7948 45760 8180 45800
rect 8235 45800 8277 45809
rect 8235 45760 8236 45800
rect 8276 45760 8277 45800
rect 7755 45751 7797 45760
rect 8235 45751 8277 45760
rect 8332 45800 8372 45928
rect 14091 45928 14092 45968
rect 14132 45928 14133 45968
rect 14091 45919 14133 45928
rect 14092 45834 14132 45919
rect 8332 45751 8372 45760
rect 14188 45800 14228 62131
rect 18232 62012 18600 62021
rect 18272 61972 18314 62012
rect 18354 61972 18396 62012
rect 18436 61972 18478 62012
rect 18518 61972 18560 62012
rect 18232 61963 18600 61972
rect 33352 62012 33720 62021
rect 33392 61972 33434 62012
rect 33474 61972 33516 62012
rect 33556 61972 33598 62012
rect 33638 61972 33680 62012
rect 33352 61963 33720 61972
rect 48472 62012 48840 62021
rect 48512 61972 48554 62012
rect 48594 61972 48636 62012
rect 48676 61972 48718 62012
rect 48758 61972 48800 62012
rect 48472 61963 48840 61972
rect 63592 62012 63960 62021
rect 63632 61972 63674 62012
rect 63714 61972 63756 62012
rect 63796 61972 63838 62012
rect 63878 61972 63920 62012
rect 63592 61963 63960 61972
rect 78712 62012 79080 62021
rect 78752 61972 78794 62012
rect 78834 61972 78876 62012
rect 78916 61972 78958 62012
rect 78998 61972 79040 62012
rect 78712 61963 79080 61972
rect 93832 62012 94200 62021
rect 93872 61972 93914 62012
rect 93954 61972 93996 62012
rect 94036 61972 94078 62012
rect 94118 61972 94160 62012
rect 93832 61963 94200 61972
rect 19472 61256 19840 61265
rect 19512 61216 19554 61256
rect 19594 61216 19636 61256
rect 19676 61216 19718 61256
rect 19758 61216 19800 61256
rect 19472 61207 19840 61216
rect 34592 61256 34960 61265
rect 34632 61216 34674 61256
rect 34714 61216 34756 61256
rect 34796 61216 34838 61256
rect 34878 61216 34920 61256
rect 34592 61207 34960 61216
rect 49712 61256 50080 61265
rect 49752 61216 49794 61256
rect 49834 61216 49876 61256
rect 49916 61216 49958 61256
rect 49998 61216 50040 61256
rect 49712 61207 50080 61216
rect 64832 61256 65200 61265
rect 64872 61216 64914 61256
rect 64954 61216 64996 61256
rect 65036 61216 65078 61256
rect 65118 61216 65160 61256
rect 64832 61207 65200 61216
rect 79952 61256 80320 61265
rect 79992 61216 80034 61256
rect 80074 61216 80116 61256
rect 80156 61216 80198 61256
rect 80238 61216 80280 61256
rect 79952 61207 80320 61216
rect 95072 61256 95440 61265
rect 95112 61216 95154 61256
rect 95194 61216 95236 61256
rect 95276 61216 95318 61256
rect 95358 61216 95400 61256
rect 95072 61207 95440 61216
rect 18232 60500 18600 60509
rect 18272 60460 18314 60500
rect 18354 60460 18396 60500
rect 18436 60460 18478 60500
rect 18518 60460 18560 60500
rect 18232 60451 18600 60460
rect 33352 60500 33720 60509
rect 33392 60460 33434 60500
rect 33474 60460 33516 60500
rect 33556 60460 33598 60500
rect 33638 60460 33680 60500
rect 33352 60451 33720 60460
rect 48472 60500 48840 60509
rect 48512 60460 48554 60500
rect 48594 60460 48636 60500
rect 48676 60460 48718 60500
rect 48758 60460 48800 60500
rect 48472 60451 48840 60460
rect 63592 60500 63960 60509
rect 63632 60460 63674 60500
rect 63714 60460 63756 60500
rect 63796 60460 63838 60500
rect 63878 60460 63920 60500
rect 63592 60451 63960 60460
rect 78712 60500 79080 60509
rect 78752 60460 78794 60500
rect 78834 60460 78876 60500
rect 78916 60460 78958 60500
rect 78998 60460 79040 60500
rect 78712 60451 79080 60460
rect 93832 60500 94200 60509
rect 93872 60460 93914 60500
rect 93954 60460 93996 60500
rect 94036 60460 94078 60500
rect 94118 60460 94160 60500
rect 93832 60451 94200 60460
rect 19472 59744 19840 59753
rect 19512 59704 19554 59744
rect 19594 59704 19636 59744
rect 19676 59704 19718 59744
rect 19758 59704 19800 59744
rect 19472 59695 19840 59704
rect 34592 59744 34960 59753
rect 34632 59704 34674 59744
rect 34714 59704 34756 59744
rect 34796 59704 34838 59744
rect 34878 59704 34920 59744
rect 34592 59695 34960 59704
rect 49712 59744 50080 59753
rect 49752 59704 49794 59744
rect 49834 59704 49876 59744
rect 49916 59704 49958 59744
rect 49998 59704 50040 59744
rect 49712 59695 50080 59704
rect 64832 59744 65200 59753
rect 64872 59704 64914 59744
rect 64954 59704 64996 59744
rect 65036 59704 65078 59744
rect 65118 59704 65160 59744
rect 64832 59695 65200 59704
rect 79952 59744 80320 59753
rect 79992 59704 80034 59744
rect 80074 59704 80116 59744
rect 80156 59704 80198 59744
rect 80238 59704 80280 59744
rect 79952 59695 80320 59704
rect 95072 59744 95440 59753
rect 95112 59704 95154 59744
rect 95194 59704 95236 59744
rect 95276 59704 95318 59744
rect 95358 59704 95400 59744
rect 95072 59695 95440 59704
rect 18232 58988 18600 58997
rect 18272 58948 18314 58988
rect 18354 58948 18396 58988
rect 18436 58948 18478 58988
rect 18518 58948 18560 58988
rect 18232 58939 18600 58948
rect 33352 58988 33720 58997
rect 33392 58948 33434 58988
rect 33474 58948 33516 58988
rect 33556 58948 33598 58988
rect 33638 58948 33680 58988
rect 33352 58939 33720 58948
rect 48472 58988 48840 58997
rect 48512 58948 48554 58988
rect 48594 58948 48636 58988
rect 48676 58948 48718 58988
rect 48758 58948 48800 58988
rect 48472 58939 48840 58948
rect 63592 58988 63960 58997
rect 63632 58948 63674 58988
rect 63714 58948 63756 58988
rect 63796 58948 63838 58988
rect 63878 58948 63920 58988
rect 63592 58939 63960 58948
rect 78712 58988 79080 58997
rect 78752 58948 78794 58988
rect 78834 58948 78876 58988
rect 78916 58948 78958 58988
rect 78998 58948 79040 58988
rect 78712 58939 79080 58948
rect 93832 58988 94200 58997
rect 93872 58948 93914 58988
rect 93954 58948 93996 58988
rect 94036 58948 94078 58988
rect 94118 58948 94160 58988
rect 93832 58939 94200 58948
rect 19472 58232 19840 58241
rect 19512 58192 19554 58232
rect 19594 58192 19636 58232
rect 19676 58192 19718 58232
rect 19758 58192 19800 58232
rect 19472 58183 19840 58192
rect 34592 58232 34960 58241
rect 34632 58192 34674 58232
rect 34714 58192 34756 58232
rect 34796 58192 34838 58232
rect 34878 58192 34920 58232
rect 34592 58183 34960 58192
rect 49712 58232 50080 58241
rect 49752 58192 49794 58232
rect 49834 58192 49876 58232
rect 49916 58192 49958 58232
rect 49998 58192 50040 58232
rect 49712 58183 50080 58192
rect 64832 58232 65200 58241
rect 64872 58192 64914 58232
rect 64954 58192 64996 58232
rect 65036 58192 65078 58232
rect 65118 58192 65160 58232
rect 64832 58183 65200 58192
rect 79952 58232 80320 58241
rect 79992 58192 80034 58232
rect 80074 58192 80116 58232
rect 80156 58192 80198 58232
rect 80238 58192 80280 58232
rect 79952 58183 80320 58192
rect 95072 58232 95440 58241
rect 95112 58192 95154 58232
rect 95194 58192 95236 58232
rect 95276 58192 95318 58232
rect 95358 58192 95400 58232
rect 95072 58183 95440 58192
rect 18232 57476 18600 57485
rect 18272 57436 18314 57476
rect 18354 57436 18396 57476
rect 18436 57436 18478 57476
rect 18518 57436 18560 57476
rect 18232 57427 18600 57436
rect 33352 57476 33720 57485
rect 33392 57436 33434 57476
rect 33474 57436 33516 57476
rect 33556 57436 33598 57476
rect 33638 57436 33680 57476
rect 33352 57427 33720 57436
rect 48472 57476 48840 57485
rect 48512 57436 48554 57476
rect 48594 57436 48636 57476
rect 48676 57436 48718 57476
rect 48758 57436 48800 57476
rect 48472 57427 48840 57436
rect 63592 57476 63960 57485
rect 63632 57436 63674 57476
rect 63714 57436 63756 57476
rect 63796 57436 63838 57476
rect 63878 57436 63920 57476
rect 63592 57427 63960 57436
rect 78712 57476 79080 57485
rect 78752 57436 78794 57476
rect 78834 57436 78876 57476
rect 78916 57436 78958 57476
rect 78998 57436 79040 57476
rect 78712 57427 79080 57436
rect 93832 57476 94200 57485
rect 93872 57436 93914 57476
rect 93954 57436 93996 57476
rect 94036 57436 94078 57476
rect 94118 57436 94160 57476
rect 93832 57427 94200 57436
rect 19472 56720 19840 56729
rect 19512 56680 19554 56720
rect 19594 56680 19636 56720
rect 19676 56680 19718 56720
rect 19758 56680 19800 56720
rect 19472 56671 19840 56680
rect 34592 56720 34960 56729
rect 34632 56680 34674 56720
rect 34714 56680 34756 56720
rect 34796 56680 34838 56720
rect 34878 56680 34920 56720
rect 34592 56671 34960 56680
rect 49712 56720 50080 56729
rect 49752 56680 49794 56720
rect 49834 56680 49876 56720
rect 49916 56680 49958 56720
rect 49998 56680 50040 56720
rect 49712 56671 50080 56680
rect 64832 56720 65200 56729
rect 64872 56680 64914 56720
rect 64954 56680 64996 56720
rect 65036 56680 65078 56720
rect 65118 56680 65160 56720
rect 64832 56671 65200 56680
rect 79952 56720 80320 56729
rect 79992 56680 80034 56720
rect 80074 56680 80116 56720
rect 80156 56680 80198 56720
rect 80238 56680 80280 56720
rect 79952 56671 80320 56680
rect 95072 56720 95440 56729
rect 95112 56680 95154 56720
rect 95194 56680 95236 56720
rect 95276 56680 95318 56720
rect 95358 56680 95400 56720
rect 95072 56671 95440 56680
rect 18232 55964 18600 55973
rect 18272 55924 18314 55964
rect 18354 55924 18396 55964
rect 18436 55924 18478 55964
rect 18518 55924 18560 55964
rect 18232 55915 18600 55924
rect 33352 55964 33720 55973
rect 33392 55924 33434 55964
rect 33474 55924 33516 55964
rect 33556 55924 33598 55964
rect 33638 55924 33680 55964
rect 33352 55915 33720 55924
rect 48472 55964 48840 55973
rect 48512 55924 48554 55964
rect 48594 55924 48636 55964
rect 48676 55924 48718 55964
rect 48758 55924 48800 55964
rect 48472 55915 48840 55924
rect 63592 55964 63960 55973
rect 63632 55924 63674 55964
rect 63714 55924 63756 55964
rect 63796 55924 63838 55964
rect 63878 55924 63920 55964
rect 63592 55915 63960 55924
rect 78712 55964 79080 55973
rect 78752 55924 78794 55964
rect 78834 55924 78876 55964
rect 78916 55924 78958 55964
rect 78998 55924 79040 55964
rect 78712 55915 79080 55924
rect 93832 55964 94200 55973
rect 93872 55924 93914 55964
rect 93954 55924 93996 55964
rect 94036 55924 94078 55964
rect 94118 55924 94160 55964
rect 93832 55915 94200 55924
rect 19472 55208 19840 55217
rect 19512 55168 19554 55208
rect 19594 55168 19636 55208
rect 19676 55168 19718 55208
rect 19758 55168 19800 55208
rect 19472 55159 19840 55168
rect 34592 55208 34960 55217
rect 34632 55168 34674 55208
rect 34714 55168 34756 55208
rect 34796 55168 34838 55208
rect 34878 55168 34920 55208
rect 34592 55159 34960 55168
rect 49712 55208 50080 55217
rect 49752 55168 49794 55208
rect 49834 55168 49876 55208
rect 49916 55168 49958 55208
rect 49998 55168 50040 55208
rect 49712 55159 50080 55168
rect 64832 55208 65200 55217
rect 64872 55168 64914 55208
rect 64954 55168 64996 55208
rect 65036 55168 65078 55208
rect 65118 55168 65160 55208
rect 64832 55159 65200 55168
rect 79952 55208 80320 55217
rect 79992 55168 80034 55208
rect 80074 55168 80116 55208
rect 80156 55168 80198 55208
rect 80238 55168 80280 55208
rect 79952 55159 80320 55168
rect 95072 55208 95440 55217
rect 95112 55168 95154 55208
rect 95194 55168 95236 55208
rect 95276 55168 95318 55208
rect 95358 55168 95400 55208
rect 95072 55159 95440 55168
rect 18232 54452 18600 54461
rect 18272 54412 18314 54452
rect 18354 54412 18396 54452
rect 18436 54412 18478 54452
rect 18518 54412 18560 54452
rect 18232 54403 18600 54412
rect 33352 54452 33720 54461
rect 33392 54412 33434 54452
rect 33474 54412 33516 54452
rect 33556 54412 33598 54452
rect 33638 54412 33680 54452
rect 33352 54403 33720 54412
rect 48472 54452 48840 54461
rect 48512 54412 48554 54452
rect 48594 54412 48636 54452
rect 48676 54412 48718 54452
rect 48758 54412 48800 54452
rect 48472 54403 48840 54412
rect 63592 54452 63960 54461
rect 63632 54412 63674 54452
rect 63714 54412 63756 54452
rect 63796 54412 63838 54452
rect 63878 54412 63920 54452
rect 63592 54403 63960 54412
rect 78712 54452 79080 54461
rect 78752 54412 78794 54452
rect 78834 54412 78876 54452
rect 78916 54412 78958 54452
rect 78998 54412 79040 54452
rect 78712 54403 79080 54412
rect 93832 54452 94200 54461
rect 93872 54412 93914 54452
rect 93954 54412 93996 54452
rect 94036 54412 94078 54452
rect 94118 54412 94160 54452
rect 93832 54403 94200 54412
rect 19472 53696 19840 53705
rect 19512 53656 19554 53696
rect 19594 53656 19636 53696
rect 19676 53656 19718 53696
rect 19758 53656 19800 53696
rect 19472 53647 19840 53656
rect 34592 53696 34960 53705
rect 34632 53656 34674 53696
rect 34714 53656 34756 53696
rect 34796 53656 34838 53696
rect 34878 53656 34920 53696
rect 34592 53647 34960 53656
rect 49712 53696 50080 53705
rect 49752 53656 49794 53696
rect 49834 53656 49876 53696
rect 49916 53656 49958 53696
rect 49998 53656 50040 53696
rect 49712 53647 50080 53656
rect 64832 53696 65200 53705
rect 64872 53656 64914 53696
rect 64954 53656 64996 53696
rect 65036 53656 65078 53696
rect 65118 53656 65160 53696
rect 64832 53647 65200 53656
rect 79952 53696 80320 53705
rect 79992 53656 80034 53696
rect 80074 53656 80116 53696
rect 80156 53656 80198 53696
rect 80238 53656 80280 53696
rect 79952 53647 80320 53656
rect 95072 53696 95440 53705
rect 95112 53656 95154 53696
rect 95194 53656 95236 53696
rect 95276 53656 95318 53696
rect 95358 53656 95400 53696
rect 95072 53647 95440 53656
rect 18232 52940 18600 52949
rect 18272 52900 18314 52940
rect 18354 52900 18396 52940
rect 18436 52900 18478 52940
rect 18518 52900 18560 52940
rect 18232 52891 18600 52900
rect 33352 52940 33720 52949
rect 33392 52900 33434 52940
rect 33474 52900 33516 52940
rect 33556 52900 33598 52940
rect 33638 52900 33680 52940
rect 33352 52891 33720 52900
rect 48472 52940 48840 52949
rect 48512 52900 48554 52940
rect 48594 52900 48636 52940
rect 48676 52900 48718 52940
rect 48758 52900 48800 52940
rect 48472 52891 48840 52900
rect 63592 52940 63960 52949
rect 63632 52900 63674 52940
rect 63714 52900 63756 52940
rect 63796 52900 63838 52940
rect 63878 52900 63920 52940
rect 63592 52891 63960 52900
rect 78712 52940 79080 52949
rect 78752 52900 78794 52940
rect 78834 52900 78876 52940
rect 78916 52900 78958 52940
rect 78998 52900 79040 52940
rect 78712 52891 79080 52900
rect 93832 52940 94200 52949
rect 93872 52900 93914 52940
rect 93954 52900 93996 52940
rect 94036 52900 94078 52940
rect 94118 52900 94160 52940
rect 93832 52891 94200 52900
rect 19472 52184 19840 52193
rect 19512 52144 19554 52184
rect 19594 52144 19636 52184
rect 19676 52144 19718 52184
rect 19758 52144 19800 52184
rect 19472 52135 19840 52144
rect 34592 52184 34960 52193
rect 34632 52144 34674 52184
rect 34714 52144 34756 52184
rect 34796 52144 34838 52184
rect 34878 52144 34920 52184
rect 34592 52135 34960 52144
rect 49712 52184 50080 52193
rect 49752 52144 49794 52184
rect 49834 52144 49876 52184
rect 49916 52144 49958 52184
rect 49998 52144 50040 52184
rect 49712 52135 50080 52144
rect 64832 52184 65200 52193
rect 64872 52144 64914 52184
rect 64954 52144 64996 52184
rect 65036 52144 65078 52184
rect 65118 52144 65160 52184
rect 64832 52135 65200 52144
rect 79952 52184 80320 52193
rect 79992 52144 80034 52184
rect 80074 52144 80116 52184
rect 80156 52144 80198 52184
rect 80238 52144 80280 52184
rect 79952 52135 80320 52144
rect 95072 52184 95440 52193
rect 95112 52144 95154 52184
rect 95194 52144 95236 52184
rect 95276 52144 95318 52184
rect 95358 52144 95400 52184
rect 95072 52135 95440 52144
rect 18232 51428 18600 51437
rect 18272 51388 18314 51428
rect 18354 51388 18396 51428
rect 18436 51388 18478 51428
rect 18518 51388 18560 51428
rect 18232 51379 18600 51388
rect 33352 51428 33720 51437
rect 33392 51388 33434 51428
rect 33474 51388 33516 51428
rect 33556 51388 33598 51428
rect 33638 51388 33680 51428
rect 33352 51379 33720 51388
rect 48472 51428 48840 51437
rect 48512 51388 48554 51428
rect 48594 51388 48636 51428
rect 48676 51388 48718 51428
rect 48758 51388 48800 51428
rect 48472 51379 48840 51388
rect 63592 51428 63960 51437
rect 63632 51388 63674 51428
rect 63714 51388 63756 51428
rect 63796 51388 63838 51428
rect 63878 51388 63920 51428
rect 63592 51379 63960 51388
rect 78712 51428 79080 51437
rect 78752 51388 78794 51428
rect 78834 51388 78876 51428
rect 78916 51388 78958 51428
rect 78998 51388 79040 51428
rect 78712 51379 79080 51388
rect 93832 51428 94200 51437
rect 93872 51388 93914 51428
rect 93954 51388 93996 51428
rect 94036 51388 94078 51428
rect 94118 51388 94160 51428
rect 93832 51379 94200 51388
rect 19472 50672 19840 50681
rect 19512 50632 19554 50672
rect 19594 50632 19636 50672
rect 19676 50632 19718 50672
rect 19758 50632 19800 50672
rect 19472 50623 19840 50632
rect 34592 50672 34960 50681
rect 34632 50632 34674 50672
rect 34714 50632 34756 50672
rect 34796 50632 34838 50672
rect 34878 50632 34920 50672
rect 34592 50623 34960 50632
rect 49712 50672 50080 50681
rect 49752 50632 49794 50672
rect 49834 50632 49876 50672
rect 49916 50632 49958 50672
rect 49998 50632 50040 50672
rect 49712 50623 50080 50632
rect 64832 50672 65200 50681
rect 64872 50632 64914 50672
rect 64954 50632 64996 50672
rect 65036 50632 65078 50672
rect 65118 50632 65160 50672
rect 64832 50623 65200 50632
rect 79952 50672 80320 50681
rect 79992 50632 80034 50672
rect 80074 50632 80116 50672
rect 80156 50632 80198 50672
rect 80238 50632 80280 50672
rect 79952 50623 80320 50632
rect 95072 50672 95440 50681
rect 95112 50632 95154 50672
rect 95194 50632 95236 50672
rect 95276 50632 95318 50672
rect 95358 50632 95400 50672
rect 95072 50623 95440 50632
rect 18232 49916 18600 49925
rect 18272 49876 18314 49916
rect 18354 49876 18396 49916
rect 18436 49876 18478 49916
rect 18518 49876 18560 49916
rect 18232 49867 18600 49876
rect 33352 49916 33720 49925
rect 33392 49876 33434 49916
rect 33474 49876 33516 49916
rect 33556 49876 33598 49916
rect 33638 49876 33680 49916
rect 33352 49867 33720 49876
rect 48472 49916 48840 49925
rect 48512 49876 48554 49916
rect 48594 49876 48636 49916
rect 48676 49876 48718 49916
rect 48758 49876 48800 49916
rect 48472 49867 48840 49876
rect 63592 49916 63960 49925
rect 63632 49876 63674 49916
rect 63714 49876 63756 49916
rect 63796 49876 63838 49916
rect 63878 49876 63920 49916
rect 63592 49867 63960 49876
rect 78712 49916 79080 49925
rect 78752 49876 78794 49916
rect 78834 49876 78876 49916
rect 78916 49876 78958 49916
rect 78998 49876 79040 49916
rect 78712 49867 79080 49876
rect 93832 49916 94200 49925
rect 93872 49876 93914 49916
rect 93954 49876 93996 49916
rect 94036 49876 94078 49916
rect 94118 49876 94160 49916
rect 93832 49867 94200 49876
rect 19472 49160 19840 49169
rect 19512 49120 19554 49160
rect 19594 49120 19636 49160
rect 19676 49120 19718 49160
rect 19758 49120 19800 49160
rect 19472 49111 19840 49120
rect 34592 49160 34960 49169
rect 34632 49120 34674 49160
rect 34714 49120 34756 49160
rect 34796 49120 34838 49160
rect 34878 49120 34920 49160
rect 34592 49111 34960 49120
rect 49712 49160 50080 49169
rect 49752 49120 49794 49160
rect 49834 49120 49876 49160
rect 49916 49120 49958 49160
rect 49998 49120 50040 49160
rect 49712 49111 50080 49120
rect 64832 49160 65200 49169
rect 64872 49120 64914 49160
rect 64954 49120 64996 49160
rect 65036 49120 65078 49160
rect 65118 49120 65160 49160
rect 64832 49111 65200 49120
rect 79952 49160 80320 49169
rect 79992 49120 80034 49160
rect 80074 49120 80116 49160
rect 80156 49120 80198 49160
rect 80238 49120 80280 49160
rect 79952 49111 80320 49120
rect 95072 49160 95440 49169
rect 95112 49120 95154 49160
rect 95194 49120 95236 49160
rect 95276 49120 95318 49160
rect 95358 49120 95400 49160
rect 95072 49111 95440 49120
rect 18232 48404 18600 48413
rect 18272 48364 18314 48404
rect 18354 48364 18396 48404
rect 18436 48364 18478 48404
rect 18518 48364 18560 48404
rect 18232 48355 18600 48364
rect 33352 48404 33720 48413
rect 33392 48364 33434 48404
rect 33474 48364 33516 48404
rect 33556 48364 33598 48404
rect 33638 48364 33680 48404
rect 33352 48355 33720 48364
rect 48472 48404 48840 48413
rect 48512 48364 48554 48404
rect 48594 48364 48636 48404
rect 48676 48364 48718 48404
rect 48758 48364 48800 48404
rect 48472 48355 48840 48364
rect 63592 48404 63960 48413
rect 63632 48364 63674 48404
rect 63714 48364 63756 48404
rect 63796 48364 63838 48404
rect 63878 48364 63920 48404
rect 63592 48355 63960 48364
rect 78712 48404 79080 48413
rect 78752 48364 78794 48404
rect 78834 48364 78876 48404
rect 78916 48364 78958 48404
rect 78998 48364 79040 48404
rect 78712 48355 79080 48364
rect 93832 48404 94200 48413
rect 93872 48364 93914 48404
rect 93954 48364 93996 48404
rect 94036 48364 94078 48404
rect 94118 48364 94160 48404
rect 93832 48355 94200 48364
rect 19472 47648 19840 47657
rect 19512 47608 19554 47648
rect 19594 47608 19636 47648
rect 19676 47608 19718 47648
rect 19758 47608 19800 47648
rect 19472 47599 19840 47608
rect 34592 47648 34960 47657
rect 34632 47608 34674 47648
rect 34714 47608 34756 47648
rect 34796 47608 34838 47648
rect 34878 47608 34920 47648
rect 34592 47599 34960 47608
rect 49712 47648 50080 47657
rect 49752 47608 49794 47648
rect 49834 47608 49876 47648
rect 49916 47608 49958 47648
rect 49998 47608 50040 47648
rect 49712 47599 50080 47608
rect 64832 47648 65200 47657
rect 64872 47608 64914 47648
rect 64954 47608 64996 47648
rect 65036 47608 65078 47648
rect 65118 47608 65160 47648
rect 64832 47599 65200 47608
rect 79952 47648 80320 47657
rect 79992 47608 80034 47648
rect 80074 47608 80116 47648
rect 80156 47608 80198 47648
rect 80238 47608 80280 47648
rect 79952 47599 80320 47608
rect 95072 47648 95440 47657
rect 95112 47608 95154 47648
rect 95194 47608 95236 47648
rect 95276 47608 95318 47648
rect 95358 47608 95400 47648
rect 95072 47599 95440 47608
rect 14476 47396 14516 47405
rect 14283 47312 14325 47321
rect 14283 47272 14284 47312
rect 14324 47272 14325 47312
rect 14283 47263 14325 47272
rect 14284 46556 14324 47263
rect 14284 46507 14324 46516
rect 14379 46472 14421 46481
rect 14379 46432 14380 46472
rect 14420 46432 14421 46472
rect 14379 46423 14421 46432
rect 14380 45968 14420 46423
rect 14380 45919 14420 45928
rect 7756 45666 7796 45751
rect 8236 45666 8276 45751
rect 14188 44960 14228 45760
rect 14188 44911 14228 44920
rect 14091 44792 14133 44801
rect 14091 44752 14092 44792
rect 14132 44752 14133 44792
rect 14091 44743 14133 44752
rect 14092 44658 14132 44743
rect 7083 16316 7125 16325
rect 7083 16276 7084 16316
rect 7124 16276 7125 16316
rect 7083 16267 7125 16276
rect 6699 10268 6741 10277
rect 6699 10228 6700 10268
rect 6740 10228 6741 10268
rect 6699 10219 6741 10228
rect 5643 8756 5685 8765
rect 5643 8716 5644 8756
rect 5684 8716 5685 8756
rect 5643 8707 5685 8716
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 14476 4901 14516 47356
rect 14571 47312 14613 47321
rect 14571 47272 14572 47312
rect 14612 47272 14613 47312
rect 14571 47263 14613 47272
rect 14956 47312 14996 47321
rect 14572 47178 14612 47263
rect 14956 46481 14996 47272
rect 18232 46892 18600 46901
rect 18272 46852 18314 46892
rect 18354 46852 18396 46892
rect 18436 46852 18478 46892
rect 18518 46852 18560 46892
rect 18232 46843 18600 46852
rect 33352 46892 33720 46901
rect 33392 46852 33434 46892
rect 33474 46852 33516 46892
rect 33556 46852 33598 46892
rect 33638 46852 33680 46892
rect 33352 46843 33720 46852
rect 48472 46892 48840 46901
rect 48512 46852 48554 46892
rect 48594 46852 48636 46892
rect 48676 46852 48718 46892
rect 48758 46852 48800 46892
rect 48472 46843 48840 46852
rect 63592 46892 63960 46901
rect 63632 46852 63674 46892
rect 63714 46852 63756 46892
rect 63796 46852 63838 46892
rect 63878 46852 63920 46892
rect 63592 46843 63960 46852
rect 78712 46892 79080 46901
rect 78752 46852 78794 46892
rect 78834 46852 78876 46892
rect 78916 46852 78958 46892
rect 78998 46852 79040 46892
rect 78712 46843 79080 46852
rect 93832 46892 94200 46901
rect 93872 46852 93914 46892
rect 93954 46852 93996 46892
rect 94036 46852 94078 46892
rect 94118 46852 94160 46892
rect 93832 46843 94200 46852
rect 14955 46472 14997 46481
rect 14955 46432 14956 46472
rect 14996 46432 14997 46472
rect 14955 46423 14997 46432
rect 19472 46136 19840 46145
rect 19512 46096 19554 46136
rect 19594 46096 19636 46136
rect 19676 46096 19718 46136
rect 19758 46096 19800 46136
rect 19472 46087 19840 46096
rect 34592 46136 34960 46145
rect 34632 46096 34674 46136
rect 34714 46096 34756 46136
rect 34796 46096 34838 46136
rect 34878 46096 34920 46136
rect 34592 46087 34960 46096
rect 49712 46136 50080 46145
rect 49752 46096 49794 46136
rect 49834 46096 49876 46136
rect 49916 46096 49958 46136
rect 49998 46096 50040 46136
rect 49712 46087 50080 46096
rect 64832 46136 65200 46145
rect 64872 46096 64914 46136
rect 64954 46096 64996 46136
rect 65036 46096 65078 46136
rect 65118 46096 65160 46136
rect 64832 46087 65200 46096
rect 79952 46136 80320 46145
rect 79992 46096 80034 46136
rect 80074 46096 80116 46136
rect 80156 46096 80198 46136
rect 80238 46096 80280 46136
rect 79952 46087 80320 46096
rect 95072 46136 95440 46145
rect 95112 46096 95154 46136
rect 95194 46096 95236 46136
rect 95276 46096 95318 46136
rect 95358 46096 95400 46136
rect 95072 46087 95440 46096
rect 14571 45968 14613 45977
rect 14571 45928 14572 45968
rect 14612 45928 14613 45968
rect 14571 45919 14613 45928
rect 14572 44960 14612 45919
rect 18232 45380 18600 45389
rect 18272 45340 18314 45380
rect 18354 45340 18396 45380
rect 18436 45340 18478 45380
rect 18518 45340 18560 45380
rect 18232 45331 18600 45340
rect 33352 45380 33720 45389
rect 33392 45340 33434 45380
rect 33474 45340 33516 45380
rect 33556 45340 33598 45380
rect 33638 45340 33680 45380
rect 33352 45331 33720 45340
rect 48472 45380 48840 45389
rect 48512 45340 48554 45380
rect 48594 45340 48636 45380
rect 48676 45340 48718 45380
rect 48758 45340 48800 45380
rect 48472 45331 48840 45340
rect 63592 45380 63960 45389
rect 63632 45340 63674 45380
rect 63714 45340 63756 45380
rect 63796 45340 63838 45380
rect 63878 45340 63920 45380
rect 63592 45331 63960 45340
rect 78712 45380 79080 45389
rect 78752 45340 78794 45380
rect 78834 45340 78876 45380
rect 78916 45340 78958 45380
rect 78998 45340 79040 45380
rect 78712 45331 79080 45340
rect 93832 45380 94200 45389
rect 93872 45340 93914 45380
rect 93954 45340 93996 45380
rect 94036 45340 94078 45380
rect 94118 45340 94160 45380
rect 93832 45331 94200 45340
rect 14572 44911 14612 44920
rect 19472 44624 19840 44633
rect 19512 44584 19554 44624
rect 19594 44584 19636 44624
rect 19676 44584 19718 44624
rect 19758 44584 19800 44624
rect 19472 44575 19840 44584
rect 34592 44624 34960 44633
rect 34632 44584 34674 44624
rect 34714 44584 34756 44624
rect 34796 44584 34838 44624
rect 34878 44584 34920 44624
rect 34592 44575 34960 44584
rect 49712 44624 50080 44633
rect 49752 44584 49794 44624
rect 49834 44584 49876 44624
rect 49916 44584 49958 44624
rect 49998 44584 50040 44624
rect 49712 44575 50080 44584
rect 64832 44624 65200 44633
rect 64872 44584 64914 44624
rect 64954 44584 64996 44624
rect 65036 44584 65078 44624
rect 65118 44584 65160 44624
rect 64832 44575 65200 44584
rect 79952 44624 80320 44633
rect 79992 44584 80034 44624
rect 80074 44584 80116 44624
rect 80156 44584 80198 44624
rect 80238 44584 80280 44624
rect 79952 44575 80320 44584
rect 95072 44624 95440 44633
rect 95112 44584 95154 44624
rect 95194 44584 95236 44624
rect 95276 44584 95318 44624
rect 95358 44584 95400 44624
rect 95072 44575 95440 44584
rect 18232 43868 18600 43877
rect 18272 43828 18314 43868
rect 18354 43828 18396 43868
rect 18436 43828 18478 43868
rect 18518 43828 18560 43868
rect 18232 43819 18600 43828
rect 33352 43868 33720 43877
rect 33392 43828 33434 43868
rect 33474 43828 33516 43868
rect 33556 43828 33598 43868
rect 33638 43828 33680 43868
rect 33352 43819 33720 43828
rect 48472 43868 48840 43877
rect 48512 43828 48554 43868
rect 48594 43828 48636 43868
rect 48676 43828 48718 43868
rect 48758 43828 48800 43868
rect 48472 43819 48840 43828
rect 63592 43868 63960 43877
rect 63632 43828 63674 43868
rect 63714 43828 63756 43868
rect 63796 43828 63838 43868
rect 63878 43828 63920 43868
rect 63592 43819 63960 43828
rect 78712 43868 79080 43877
rect 78752 43828 78794 43868
rect 78834 43828 78876 43868
rect 78916 43828 78958 43868
rect 78998 43828 79040 43868
rect 78712 43819 79080 43828
rect 93832 43868 94200 43877
rect 93872 43828 93914 43868
rect 93954 43828 93996 43868
rect 94036 43828 94078 43868
rect 94118 43828 94160 43868
rect 93832 43819 94200 43828
rect 19472 43112 19840 43121
rect 19512 43072 19554 43112
rect 19594 43072 19636 43112
rect 19676 43072 19718 43112
rect 19758 43072 19800 43112
rect 19472 43063 19840 43072
rect 34592 43112 34960 43121
rect 34632 43072 34674 43112
rect 34714 43072 34756 43112
rect 34796 43072 34838 43112
rect 34878 43072 34920 43112
rect 34592 43063 34960 43072
rect 49712 43112 50080 43121
rect 49752 43072 49794 43112
rect 49834 43072 49876 43112
rect 49916 43072 49958 43112
rect 49998 43072 50040 43112
rect 49712 43063 50080 43072
rect 64832 43112 65200 43121
rect 64872 43072 64914 43112
rect 64954 43072 64996 43112
rect 65036 43072 65078 43112
rect 65118 43072 65160 43112
rect 64832 43063 65200 43072
rect 79952 43112 80320 43121
rect 79992 43072 80034 43112
rect 80074 43072 80116 43112
rect 80156 43072 80198 43112
rect 80238 43072 80280 43112
rect 79952 43063 80320 43072
rect 95072 43112 95440 43121
rect 95112 43072 95154 43112
rect 95194 43072 95236 43112
rect 95276 43072 95318 43112
rect 95358 43072 95400 43112
rect 95072 43063 95440 43072
rect 18232 42356 18600 42365
rect 18272 42316 18314 42356
rect 18354 42316 18396 42356
rect 18436 42316 18478 42356
rect 18518 42316 18560 42356
rect 18232 42307 18600 42316
rect 33352 42356 33720 42365
rect 33392 42316 33434 42356
rect 33474 42316 33516 42356
rect 33556 42316 33598 42356
rect 33638 42316 33680 42356
rect 33352 42307 33720 42316
rect 48472 42356 48840 42365
rect 48512 42316 48554 42356
rect 48594 42316 48636 42356
rect 48676 42316 48718 42356
rect 48758 42316 48800 42356
rect 48472 42307 48840 42316
rect 63592 42356 63960 42365
rect 63632 42316 63674 42356
rect 63714 42316 63756 42356
rect 63796 42316 63838 42356
rect 63878 42316 63920 42356
rect 63592 42307 63960 42316
rect 78712 42356 79080 42365
rect 78752 42316 78794 42356
rect 78834 42316 78876 42356
rect 78916 42316 78958 42356
rect 78998 42316 79040 42356
rect 78712 42307 79080 42316
rect 93832 42356 94200 42365
rect 93872 42316 93914 42356
rect 93954 42316 93996 42356
rect 94036 42316 94078 42356
rect 94118 42316 94160 42356
rect 93832 42307 94200 42316
rect 19472 41600 19840 41609
rect 19512 41560 19554 41600
rect 19594 41560 19636 41600
rect 19676 41560 19718 41600
rect 19758 41560 19800 41600
rect 19472 41551 19840 41560
rect 34592 41600 34960 41609
rect 34632 41560 34674 41600
rect 34714 41560 34756 41600
rect 34796 41560 34838 41600
rect 34878 41560 34920 41600
rect 34592 41551 34960 41560
rect 49712 41600 50080 41609
rect 49752 41560 49794 41600
rect 49834 41560 49876 41600
rect 49916 41560 49958 41600
rect 49998 41560 50040 41600
rect 49712 41551 50080 41560
rect 64832 41600 65200 41609
rect 64872 41560 64914 41600
rect 64954 41560 64996 41600
rect 65036 41560 65078 41600
rect 65118 41560 65160 41600
rect 64832 41551 65200 41560
rect 79952 41600 80320 41609
rect 79992 41560 80034 41600
rect 80074 41560 80116 41600
rect 80156 41560 80198 41600
rect 80238 41560 80280 41600
rect 79952 41551 80320 41560
rect 95072 41600 95440 41609
rect 95112 41560 95154 41600
rect 95194 41560 95236 41600
rect 95276 41560 95318 41600
rect 95358 41560 95400 41600
rect 95072 41551 95440 41560
rect 18232 40844 18600 40853
rect 18272 40804 18314 40844
rect 18354 40804 18396 40844
rect 18436 40804 18478 40844
rect 18518 40804 18560 40844
rect 18232 40795 18600 40804
rect 33352 40844 33720 40853
rect 33392 40804 33434 40844
rect 33474 40804 33516 40844
rect 33556 40804 33598 40844
rect 33638 40804 33680 40844
rect 33352 40795 33720 40804
rect 48472 40844 48840 40853
rect 48512 40804 48554 40844
rect 48594 40804 48636 40844
rect 48676 40804 48718 40844
rect 48758 40804 48800 40844
rect 48472 40795 48840 40804
rect 63592 40844 63960 40853
rect 63632 40804 63674 40844
rect 63714 40804 63756 40844
rect 63796 40804 63838 40844
rect 63878 40804 63920 40844
rect 63592 40795 63960 40804
rect 78712 40844 79080 40853
rect 78752 40804 78794 40844
rect 78834 40804 78876 40844
rect 78916 40804 78958 40844
rect 78998 40804 79040 40844
rect 78712 40795 79080 40804
rect 93832 40844 94200 40853
rect 93872 40804 93914 40844
rect 93954 40804 93996 40844
rect 94036 40804 94078 40844
rect 94118 40804 94160 40844
rect 93832 40795 94200 40804
rect 19472 40088 19840 40097
rect 19512 40048 19554 40088
rect 19594 40048 19636 40088
rect 19676 40048 19718 40088
rect 19758 40048 19800 40088
rect 19472 40039 19840 40048
rect 34592 40088 34960 40097
rect 34632 40048 34674 40088
rect 34714 40048 34756 40088
rect 34796 40048 34838 40088
rect 34878 40048 34920 40088
rect 34592 40039 34960 40048
rect 49712 40088 50080 40097
rect 49752 40048 49794 40088
rect 49834 40048 49876 40088
rect 49916 40048 49958 40088
rect 49998 40048 50040 40088
rect 49712 40039 50080 40048
rect 64832 40088 65200 40097
rect 64872 40048 64914 40088
rect 64954 40048 64996 40088
rect 65036 40048 65078 40088
rect 65118 40048 65160 40088
rect 64832 40039 65200 40048
rect 79952 40088 80320 40097
rect 79992 40048 80034 40088
rect 80074 40048 80116 40088
rect 80156 40048 80198 40088
rect 80238 40048 80280 40088
rect 79952 40039 80320 40048
rect 95072 40088 95440 40097
rect 95112 40048 95154 40088
rect 95194 40048 95236 40088
rect 95276 40048 95318 40088
rect 95358 40048 95400 40088
rect 95072 40039 95440 40048
rect 18232 39332 18600 39341
rect 18272 39292 18314 39332
rect 18354 39292 18396 39332
rect 18436 39292 18478 39332
rect 18518 39292 18560 39332
rect 18232 39283 18600 39292
rect 33352 39332 33720 39341
rect 33392 39292 33434 39332
rect 33474 39292 33516 39332
rect 33556 39292 33598 39332
rect 33638 39292 33680 39332
rect 33352 39283 33720 39292
rect 48472 39332 48840 39341
rect 48512 39292 48554 39332
rect 48594 39292 48636 39332
rect 48676 39292 48718 39332
rect 48758 39292 48800 39332
rect 48472 39283 48840 39292
rect 63592 39332 63960 39341
rect 63632 39292 63674 39332
rect 63714 39292 63756 39332
rect 63796 39292 63838 39332
rect 63878 39292 63920 39332
rect 63592 39283 63960 39292
rect 78712 39332 79080 39341
rect 78752 39292 78794 39332
rect 78834 39292 78876 39332
rect 78916 39292 78958 39332
rect 78998 39292 79040 39332
rect 78712 39283 79080 39292
rect 93832 39332 94200 39341
rect 93872 39292 93914 39332
rect 93954 39292 93996 39332
rect 94036 39292 94078 39332
rect 94118 39292 94160 39332
rect 93832 39283 94200 39292
rect 19472 38576 19840 38585
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19472 38527 19840 38536
rect 34592 38576 34960 38585
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34592 38527 34960 38536
rect 49712 38576 50080 38585
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 49712 38527 50080 38536
rect 64832 38576 65200 38585
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 64832 38527 65200 38536
rect 79952 38576 80320 38585
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 79952 38527 80320 38536
rect 95072 38576 95440 38585
rect 95112 38536 95154 38576
rect 95194 38536 95236 38576
rect 95276 38536 95318 38576
rect 95358 38536 95400 38576
rect 95072 38527 95440 38536
rect 18232 37820 18600 37829
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18232 37771 18600 37780
rect 33352 37820 33720 37829
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33352 37771 33720 37780
rect 48472 37820 48840 37829
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48472 37771 48840 37780
rect 63592 37820 63960 37829
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63592 37771 63960 37780
rect 78712 37820 79080 37829
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 78712 37771 79080 37780
rect 93832 37820 94200 37829
rect 93872 37780 93914 37820
rect 93954 37780 93996 37820
rect 94036 37780 94078 37820
rect 94118 37780 94160 37820
rect 93832 37771 94200 37780
rect 19472 37064 19840 37073
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19472 37015 19840 37024
rect 34592 37064 34960 37073
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34592 37015 34960 37024
rect 49712 37064 50080 37073
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 49712 37015 50080 37024
rect 64832 37064 65200 37073
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 64832 37015 65200 37024
rect 79952 37064 80320 37073
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 79952 37015 80320 37024
rect 95072 37064 95440 37073
rect 95112 37024 95154 37064
rect 95194 37024 95236 37064
rect 95276 37024 95318 37064
rect 95358 37024 95400 37064
rect 95072 37015 95440 37024
rect 18232 36308 18600 36317
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18232 36259 18600 36268
rect 33352 36308 33720 36317
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33352 36259 33720 36268
rect 48472 36308 48840 36317
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48472 36259 48840 36268
rect 63592 36308 63960 36317
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63592 36259 63960 36268
rect 78712 36308 79080 36317
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 78712 36259 79080 36268
rect 93832 36308 94200 36317
rect 93872 36268 93914 36308
rect 93954 36268 93996 36308
rect 94036 36268 94078 36308
rect 94118 36268 94160 36308
rect 93832 36259 94200 36268
rect 19472 35552 19840 35561
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19472 35503 19840 35512
rect 34592 35552 34960 35561
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34592 35503 34960 35512
rect 49712 35552 50080 35561
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 49712 35503 50080 35512
rect 64832 35552 65200 35561
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 64832 35503 65200 35512
rect 79952 35552 80320 35561
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 79952 35503 80320 35512
rect 95072 35552 95440 35561
rect 95112 35512 95154 35552
rect 95194 35512 95236 35552
rect 95276 35512 95318 35552
rect 95358 35512 95400 35552
rect 95072 35503 95440 35512
rect 18232 34796 18600 34805
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18232 34747 18600 34756
rect 33352 34796 33720 34805
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33352 34747 33720 34756
rect 48472 34796 48840 34805
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48472 34747 48840 34756
rect 63592 34796 63960 34805
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63592 34747 63960 34756
rect 78712 34796 79080 34805
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 78712 34747 79080 34756
rect 93832 34796 94200 34805
rect 93872 34756 93914 34796
rect 93954 34756 93996 34796
rect 94036 34756 94078 34796
rect 94118 34756 94160 34796
rect 93832 34747 94200 34756
rect 19472 34040 19840 34049
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19472 33991 19840 34000
rect 34592 34040 34960 34049
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34592 33991 34960 34000
rect 49712 34040 50080 34049
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 49712 33991 50080 34000
rect 64832 34040 65200 34049
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 64832 33991 65200 34000
rect 79952 34040 80320 34049
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 79952 33991 80320 34000
rect 95072 34040 95440 34049
rect 95112 34000 95154 34040
rect 95194 34000 95236 34040
rect 95276 34000 95318 34040
rect 95358 34000 95400 34040
rect 95072 33991 95440 34000
rect 18232 33284 18600 33293
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18232 33235 18600 33244
rect 33352 33284 33720 33293
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33352 33235 33720 33244
rect 48472 33284 48840 33293
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48472 33235 48840 33244
rect 63592 33284 63960 33293
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63592 33235 63960 33244
rect 78712 33284 79080 33293
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 78712 33235 79080 33244
rect 93832 33284 94200 33293
rect 93872 33244 93914 33284
rect 93954 33244 93996 33284
rect 94036 33244 94078 33284
rect 94118 33244 94160 33284
rect 93832 33235 94200 33244
rect 19472 32528 19840 32537
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19472 32479 19840 32488
rect 34592 32528 34960 32537
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34592 32479 34960 32488
rect 49712 32528 50080 32537
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 49712 32479 50080 32488
rect 64832 32528 65200 32537
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 64832 32479 65200 32488
rect 79952 32528 80320 32537
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 79952 32479 80320 32488
rect 95072 32528 95440 32537
rect 95112 32488 95154 32528
rect 95194 32488 95236 32528
rect 95276 32488 95318 32528
rect 95358 32488 95400 32528
rect 95072 32479 95440 32488
rect 18232 31772 18600 31781
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18232 31723 18600 31732
rect 33352 31772 33720 31781
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33352 31723 33720 31732
rect 48472 31772 48840 31781
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48472 31723 48840 31732
rect 63592 31772 63960 31781
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63592 31723 63960 31732
rect 78712 31772 79080 31781
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 78712 31723 79080 31732
rect 93832 31772 94200 31781
rect 93872 31732 93914 31772
rect 93954 31732 93996 31772
rect 94036 31732 94078 31772
rect 94118 31732 94160 31772
rect 93832 31723 94200 31732
rect 19472 31016 19840 31025
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19472 30967 19840 30976
rect 34592 31016 34960 31025
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34592 30967 34960 30976
rect 49712 31016 50080 31025
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 49712 30967 50080 30976
rect 64832 31016 65200 31025
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 64832 30967 65200 30976
rect 79952 31016 80320 31025
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 79952 30967 80320 30976
rect 95072 31016 95440 31025
rect 95112 30976 95154 31016
rect 95194 30976 95236 31016
rect 95276 30976 95318 31016
rect 95358 30976 95400 31016
rect 95072 30967 95440 30976
rect 18232 30260 18600 30269
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18232 30211 18600 30220
rect 33352 30260 33720 30269
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33352 30211 33720 30220
rect 48472 30260 48840 30269
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48472 30211 48840 30220
rect 63592 30260 63960 30269
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63592 30211 63960 30220
rect 78712 30260 79080 30269
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 78712 30211 79080 30220
rect 93832 30260 94200 30269
rect 93872 30220 93914 30260
rect 93954 30220 93996 30260
rect 94036 30220 94078 30260
rect 94118 30220 94160 30260
rect 93832 30211 94200 30220
rect 19472 29504 19840 29513
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19472 29455 19840 29464
rect 34592 29504 34960 29513
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34592 29455 34960 29464
rect 49712 29504 50080 29513
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 49712 29455 50080 29464
rect 64832 29504 65200 29513
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 64832 29455 65200 29464
rect 79952 29504 80320 29513
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 79952 29455 80320 29464
rect 95072 29504 95440 29513
rect 95112 29464 95154 29504
rect 95194 29464 95236 29504
rect 95276 29464 95318 29504
rect 95358 29464 95400 29504
rect 95072 29455 95440 29464
rect 18232 28748 18600 28757
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18232 28699 18600 28708
rect 33352 28748 33720 28757
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33352 28699 33720 28708
rect 48472 28748 48840 28757
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48472 28699 48840 28708
rect 63592 28748 63960 28757
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63592 28699 63960 28708
rect 78712 28748 79080 28757
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 78712 28699 79080 28708
rect 93832 28748 94200 28757
rect 93872 28708 93914 28748
rect 93954 28708 93996 28748
rect 94036 28708 94078 28748
rect 94118 28708 94160 28748
rect 93832 28699 94200 28708
rect 19472 27992 19840 28001
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19472 27943 19840 27952
rect 34592 27992 34960 28001
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34592 27943 34960 27952
rect 49712 27992 50080 28001
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 49712 27943 50080 27952
rect 64832 27992 65200 28001
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 64832 27943 65200 27952
rect 79952 27992 80320 28001
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 79952 27943 80320 27952
rect 95072 27992 95440 28001
rect 95112 27952 95154 27992
rect 95194 27952 95236 27992
rect 95276 27952 95318 27992
rect 95358 27952 95400 27992
rect 95072 27943 95440 27952
rect 18232 27236 18600 27245
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18232 27187 18600 27196
rect 33352 27236 33720 27245
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33352 27187 33720 27196
rect 48472 27236 48840 27245
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48472 27187 48840 27196
rect 63592 27236 63960 27245
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63592 27187 63960 27196
rect 78712 27236 79080 27245
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 78712 27187 79080 27196
rect 93832 27236 94200 27245
rect 93872 27196 93914 27236
rect 93954 27196 93996 27236
rect 94036 27196 94078 27236
rect 94118 27196 94160 27236
rect 93832 27187 94200 27196
rect 19472 26480 19840 26489
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19472 26431 19840 26440
rect 34592 26480 34960 26489
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34592 26431 34960 26440
rect 49712 26480 50080 26489
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 49712 26431 50080 26440
rect 64832 26480 65200 26489
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 64832 26431 65200 26440
rect 79952 26480 80320 26489
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 79952 26431 80320 26440
rect 95072 26480 95440 26489
rect 95112 26440 95154 26480
rect 95194 26440 95236 26480
rect 95276 26440 95318 26480
rect 95358 26440 95400 26480
rect 95072 26431 95440 26440
rect 18232 25724 18600 25733
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18232 25675 18600 25684
rect 33352 25724 33720 25733
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33352 25675 33720 25684
rect 48472 25724 48840 25733
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48472 25675 48840 25684
rect 63592 25724 63960 25733
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63592 25675 63960 25684
rect 78712 25724 79080 25733
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 78712 25675 79080 25684
rect 93832 25724 94200 25733
rect 93872 25684 93914 25724
rect 93954 25684 93996 25724
rect 94036 25684 94078 25724
rect 94118 25684 94160 25724
rect 93832 25675 94200 25684
rect 19472 24968 19840 24977
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19472 24919 19840 24928
rect 34592 24968 34960 24977
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34592 24919 34960 24928
rect 49712 24968 50080 24977
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 49712 24919 50080 24928
rect 64832 24968 65200 24977
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 64832 24919 65200 24928
rect 79952 24968 80320 24977
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 79952 24919 80320 24928
rect 95072 24968 95440 24977
rect 95112 24928 95154 24968
rect 95194 24928 95236 24968
rect 95276 24928 95318 24968
rect 95358 24928 95400 24968
rect 95072 24919 95440 24928
rect 18232 24212 18600 24221
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18232 24163 18600 24172
rect 33352 24212 33720 24221
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33352 24163 33720 24172
rect 48472 24212 48840 24221
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48472 24163 48840 24172
rect 63592 24212 63960 24221
rect 63632 24172 63674 24212
rect 63714 24172 63756 24212
rect 63796 24172 63838 24212
rect 63878 24172 63920 24212
rect 63592 24163 63960 24172
rect 78712 24212 79080 24221
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 78712 24163 79080 24172
rect 93832 24212 94200 24221
rect 93872 24172 93914 24212
rect 93954 24172 93996 24212
rect 94036 24172 94078 24212
rect 94118 24172 94160 24212
rect 93832 24163 94200 24172
rect 19472 23456 19840 23465
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19472 23407 19840 23416
rect 34592 23456 34960 23465
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34592 23407 34960 23416
rect 49712 23456 50080 23465
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 49712 23407 50080 23416
rect 64832 23456 65200 23465
rect 64872 23416 64914 23456
rect 64954 23416 64996 23456
rect 65036 23416 65078 23456
rect 65118 23416 65160 23456
rect 64832 23407 65200 23416
rect 79952 23456 80320 23465
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 79952 23407 80320 23416
rect 95072 23456 95440 23465
rect 95112 23416 95154 23456
rect 95194 23416 95236 23456
rect 95276 23416 95318 23456
rect 95358 23416 95400 23456
rect 95072 23407 95440 23416
rect 18232 22700 18600 22709
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18232 22651 18600 22660
rect 33352 22700 33720 22709
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33352 22651 33720 22660
rect 48472 22700 48840 22709
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48472 22651 48840 22660
rect 63592 22700 63960 22709
rect 63632 22660 63674 22700
rect 63714 22660 63756 22700
rect 63796 22660 63838 22700
rect 63878 22660 63920 22700
rect 63592 22651 63960 22660
rect 78712 22700 79080 22709
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 78712 22651 79080 22660
rect 93832 22700 94200 22709
rect 93872 22660 93914 22700
rect 93954 22660 93996 22700
rect 94036 22660 94078 22700
rect 94118 22660 94160 22700
rect 93832 22651 94200 22660
rect 19472 21944 19840 21953
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19472 21895 19840 21904
rect 34592 21944 34960 21953
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34592 21895 34960 21904
rect 49712 21944 50080 21953
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 49712 21895 50080 21904
rect 64832 21944 65200 21953
rect 64872 21904 64914 21944
rect 64954 21904 64996 21944
rect 65036 21904 65078 21944
rect 65118 21904 65160 21944
rect 64832 21895 65200 21904
rect 79952 21944 80320 21953
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 79952 21895 80320 21904
rect 95072 21944 95440 21953
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95072 21895 95440 21904
rect 18232 21188 18600 21197
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18232 21139 18600 21148
rect 33352 21188 33720 21197
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33352 21139 33720 21148
rect 48472 21188 48840 21197
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48472 21139 48840 21148
rect 63592 21188 63960 21197
rect 63632 21148 63674 21188
rect 63714 21148 63756 21188
rect 63796 21148 63838 21188
rect 63878 21148 63920 21188
rect 63592 21139 63960 21148
rect 78712 21188 79080 21197
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 78712 21139 79080 21148
rect 93832 21188 94200 21197
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 93832 21139 94200 21148
rect 19472 20432 19840 20441
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19472 20383 19840 20392
rect 34592 20432 34960 20441
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34592 20383 34960 20392
rect 49712 20432 50080 20441
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 49712 20383 50080 20392
rect 64832 20432 65200 20441
rect 64872 20392 64914 20432
rect 64954 20392 64996 20432
rect 65036 20392 65078 20432
rect 65118 20392 65160 20432
rect 64832 20383 65200 20392
rect 79952 20432 80320 20441
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 79952 20383 80320 20392
rect 95072 20432 95440 20441
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95072 20383 95440 20392
rect 18232 19676 18600 19685
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18232 19627 18600 19636
rect 33352 19676 33720 19685
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33352 19627 33720 19636
rect 48472 19676 48840 19685
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48472 19627 48840 19636
rect 63592 19676 63960 19685
rect 63632 19636 63674 19676
rect 63714 19636 63756 19676
rect 63796 19636 63838 19676
rect 63878 19636 63920 19676
rect 63592 19627 63960 19636
rect 78712 19676 79080 19685
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 78712 19627 79080 19636
rect 93832 19676 94200 19685
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 93832 19627 94200 19636
rect 19472 18920 19840 18929
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19472 18871 19840 18880
rect 34592 18920 34960 18929
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34592 18871 34960 18880
rect 49712 18920 50080 18929
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 49712 18871 50080 18880
rect 64832 18920 65200 18929
rect 64872 18880 64914 18920
rect 64954 18880 64996 18920
rect 65036 18880 65078 18920
rect 65118 18880 65160 18920
rect 64832 18871 65200 18880
rect 79952 18920 80320 18929
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 79952 18871 80320 18880
rect 95072 18920 95440 18929
rect 95112 18880 95154 18920
rect 95194 18880 95236 18920
rect 95276 18880 95318 18920
rect 95358 18880 95400 18920
rect 95072 18871 95440 18880
rect 18232 18164 18600 18173
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18232 18115 18600 18124
rect 33352 18164 33720 18173
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33352 18115 33720 18124
rect 48472 18164 48840 18173
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48472 18115 48840 18124
rect 63592 18164 63960 18173
rect 63632 18124 63674 18164
rect 63714 18124 63756 18164
rect 63796 18124 63838 18164
rect 63878 18124 63920 18164
rect 63592 18115 63960 18124
rect 78712 18164 79080 18173
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 78712 18115 79080 18124
rect 93832 18164 94200 18173
rect 93872 18124 93914 18164
rect 93954 18124 93996 18164
rect 94036 18124 94078 18164
rect 94118 18124 94160 18164
rect 93832 18115 94200 18124
rect 19472 17408 19840 17417
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19472 17359 19840 17368
rect 34592 17408 34960 17417
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34592 17359 34960 17368
rect 49712 17408 50080 17417
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 49712 17359 50080 17368
rect 64832 17408 65200 17417
rect 64872 17368 64914 17408
rect 64954 17368 64996 17408
rect 65036 17368 65078 17408
rect 65118 17368 65160 17408
rect 64832 17359 65200 17368
rect 79952 17408 80320 17417
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 79952 17359 80320 17368
rect 95072 17408 95440 17417
rect 95112 17368 95154 17408
rect 95194 17368 95236 17408
rect 95276 17368 95318 17408
rect 95358 17368 95400 17408
rect 95072 17359 95440 17368
rect 18232 16652 18600 16661
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18232 16603 18600 16612
rect 33352 16652 33720 16661
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33352 16603 33720 16612
rect 48472 16652 48840 16661
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48472 16603 48840 16612
rect 63592 16652 63960 16661
rect 63632 16612 63674 16652
rect 63714 16612 63756 16652
rect 63796 16612 63838 16652
rect 63878 16612 63920 16652
rect 63592 16603 63960 16612
rect 78712 16652 79080 16661
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 78712 16603 79080 16612
rect 93832 16652 94200 16661
rect 93872 16612 93914 16652
rect 93954 16612 93996 16652
rect 94036 16612 94078 16652
rect 94118 16612 94160 16652
rect 93832 16603 94200 16612
rect 19472 15896 19840 15905
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19472 15847 19840 15856
rect 34592 15896 34960 15905
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34592 15847 34960 15856
rect 49712 15896 50080 15905
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 49712 15847 50080 15856
rect 64832 15896 65200 15905
rect 64872 15856 64914 15896
rect 64954 15856 64996 15896
rect 65036 15856 65078 15896
rect 65118 15856 65160 15896
rect 64832 15847 65200 15856
rect 79952 15896 80320 15905
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 79952 15847 80320 15856
rect 95072 15896 95440 15905
rect 95112 15856 95154 15896
rect 95194 15856 95236 15896
rect 95276 15856 95318 15896
rect 95358 15856 95400 15896
rect 95072 15847 95440 15856
rect 18232 15140 18600 15149
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18232 15091 18600 15100
rect 33352 15140 33720 15149
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 33352 15091 33720 15100
rect 48472 15140 48840 15149
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48472 15091 48840 15100
rect 63592 15140 63960 15149
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63592 15091 63960 15100
rect 78712 15140 79080 15149
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 78712 15091 79080 15100
rect 93832 15140 94200 15149
rect 93872 15100 93914 15140
rect 93954 15100 93996 15140
rect 94036 15100 94078 15140
rect 94118 15100 94160 15140
rect 93832 15091 94200 15100
rect 19472 14384 19840 14393
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19472 14335 19840 14344
rect 34592 14384 34960 14393
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34592 14335 34960 14344
rect 49712 14384 50080 14393
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 49712 14335 50080 14344
rect 64832 14384 65200 14393
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 64832 14335 65200 14344
rect 79952 14384 80320 14393
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 79952 14335 80320 14344
rect 95072 14384 95440 14393
rect 95112 14344 95154 14384
rect 95194 14344 95236 14384
rect 95276 14344 95318 14384
rect 95358 14344 95400 14384
rect 95072 14335 95440 14344
rect 18232 13628 18600 13637
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18232 13579 18600 13588
rect 33352 13628 33720 13637
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33352 13579 33720 13588
rect 48472 13628 48840 13637
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48472 13579 48840 13588
rect 63592 13628 63960 13637
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63592 13579 63960 13588
rect 78712 13628 79080 13637
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 78712 13579 79080 13588
rect 93832 13628 94200 13637
rect 93872 13588 93914 13628
rect 93954 13588 93996 13628
rect 94036 13588 94078 13628
rect 94118 13588 94160 13628
rect 93832 13579 94200 13588
rect 19472 12872 19840 12881
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19472 12823 19840 12832
rect 34592 12872 34960 12881
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34592 12823 34960 12832
rect 49712 12872 50080 12881
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 49712 12823 50080 12832
rect 64832 12872 65200 12881
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 64832 12823 65200 12832
rect 79952 12872 80320 12881
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 79952 12823 80320 12832
rect 95072 12872 95440 12881
rect 95112 12832 95154 12872
rect 95194 12832 95236 12872
rect 95276 12832 95318 12872
rect 95358 12832 95400 12872
rect 95072 12823 95440 12832
rect 18232 12116 18600 12125
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18232 12067 18600 12076
rect 33352 12116 33720 12125
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33352 12067 33720 12076
rect 48472 12116 48840 12125
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48472 12067 48840 12076
rect 63592 12116 63960 12125
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63592 12067 63960 12076
rect 78712 12116 79080 12125
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 78712 12067 79080 12076
rect 93832 12116 94200 12125
rect 93872 12076 93914 12116
rect 93954 12076 93996 12116
rect 94036 12076 94078 12116
rect 94118 12076 94160 12116
rect 93832 12067 94200 12076
rect 19472 11360 19840 11369
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19472 11311 19840 11320
rect 34592 11360 34960 11369
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34592 11311 34960 11320
rect 49712 11360 50080 11369
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 49712 11311 50080 11320
rect 64832 11360 65200 11369
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 64832 11311 65200 11320
rect 79952 11360 80320 11369
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 79952 11311 80320 11320
rect 95072 11360 95440 11369
rect 95112 11320 95154 11360
rect 95194 11320 95236 11360
rect 95276 11320 95318 11360
rect 95358 11320 95400 11360
rect 95072 11311 95440 11320
rect 18232 10604 18600 10613
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18232 10555 18600 10564
rect 33352 10604 33720 10613
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33352 10555 33720 10564
rect 48472 10604 48840 10613
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48472 10555 48840 10564
rect 63592 10604 63960 10613
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63592 10555 63960 10564
rect 78712 10604 79080 10613
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 78712 10555 79080 10564
rect 93832 10604 94200 10613
rect 93872 10564 93914 10604
rect 93954 10564 93996 10604
rect 94036 10564 94078 10604
rect 94118 10564 94160 10604
rect 93832 10555 94200 10564
rect 19472 9848 19840 9857
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19472 9799 19840 9808
rect 34592 9848 34960 9857
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34592 9799 34960 9808
rect 49712 9848 50080 9857
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 49712 9799 50080 9808
rect 64832 9848 65200 9857
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 64832 9799 65200 9808
rect 79952 9848 80320 9857
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 79952 9799 80320 9808
rect 95072 9848 95440 9857
rect 95112 9808 95154 9848
rect 95194 9808 95236 9848
rect 95276 9808 95318 9848
rect 95358 9808 95400 9848
rect 95072 9799 95440 9808
rect 18232 9092 18600 9101
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18232 9043 18600 9052
rect 33352 9092 33720 9101
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33352 9043 33720 9052
rect 48472 9092 48840 9101
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48472 9043 48840 9052
rect 63592 9092 63960 9101
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63592 9043 63960 9052
rect 78712 9092 79080 9101
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 78712 9043 79080 9052
rect 93832 9092 94200 9101
rect 93872 9052 93914 9092
rect 93954 9052 93996 9092
rect 94036 9052 94078 9092
rect 94118 9052 94160 9092
rect 93832 9043 94200 9052
rect 19472 8336 19840 8345
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19472 8287 19840 8296
rect 34592 8336 34960 8345
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34592 8287 34960 8296
rect 49712 8336 50080 8345
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 49712 8287 50080 8296
rect 64832 8336 65200 8345
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 64832 8287 65200 8296
rect 79952 8336 80320 8345
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 79952 8287 80320 8296
rect 95072 8336 95440 8345
rect 95112 8296 95154 8336
rect 95194 8296 95236 8336
rect 95276 8296 95318 8336
rect 95358 8296 95400 8336
rect 95072 8287 95440 8296
rect 18232 7580 18600 7589
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18232 7531 18600 7540
rect 33352 7580 33720 7589
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33352 7531 33720 7540
rect 48472 7580 48840 7589
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48472 7531 48840 7540
rect 63592 7580 63960 7589
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63592 7531 63960 7540
rect 78712 7580 79080 7589
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 78712 7531 79080 7540
rect 93832 7580 94200 7589
rect 93872 7540 93914 7580
rect 93954 7540 93996 7580
rect 94036 7540 94078 7580
rect 94118 7540 94160 7580
rect 93832 7531 94200 7540
rect 19472 6824 19840 6833
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19472 6775 19840 6784
rect 34592 6824 34960 6833
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34592 6775 34960 6784
rect 49712 6824 50080 6833
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 49712 6775 50080 6784
rect 64832 6824 65200 6833
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 64832 6775 65200 6784
rect 79952 6824 80320 6833
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 79952 6775 80320 6784
rect 95072 6824 95440 6833
rect 95112 6784 95154 6824
rect 95194 6784 95236 6824
rect 95276 6784 95318 6824
rect 95358 6784 95400 6824
rect 95072 6775 95440 6784
rect 18232 6068 18600 6077
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18232 6019 18600 6028
rect 33352 6068 33720 6077
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33352 6019 33720 6028
rect 48472 6068 48840 6077
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48472 6019 48840 6028
rect 63592 6068 63960 6077
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63592 6019 63960 6028
rect 78712 6068 79080 6077
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 78712 6019 79080 6028
rect 93832 6068 94200 6077
rect 93872 6028 93914 6068
rect 93954 6028 93996 6068
rect 94036 6028 94078 6068
rect 94118 6028 94160 6068
rect 93832 6019 94200 6028
rect 19472 5312 19840 5321
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19472 5263 19840 5272
rect 34592 5312 34960 5321
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34592 5263 34960 5272
rect 49712 5312 50080 5321
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 49712 5263 50080 5272
rect 64832 5312 65200 5321
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 64832 5263 65200 5272
rect 79952 5312 80320 5321
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 79952 5263 80320 5272
rect 95072 5312 95440 5321
rect 95112 5272 95154 5312
rect 95194 5272 95236 5312
rect 95276 5272 95318 5312
rect 95358 5272 95400 5312
rect 95072 5263 95440 5272
rect 14475 4892 14517 4901
rect 14475 4852 14476 4892
rect 14516 4852 14517 4892
rect 14475 4843 14517 4852
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 18232 4556 18600 4565
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18232 4507 18600 4516
rect 33352 4556 33720 4565
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33352 4507 33720 4516
rect 48472 4556 48840 4565
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48472 4507 48840 4516
rect 63592 4556 63960 4565
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63592 4507 63960 4516
rect 78712 4556 79080 4565
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 78712 4507 79080 4516
rect 93832 4556 94200 4565
rect 93872 4516 93914 4556
rect 93954 4516 93996 4556
rect 94036 4516 94078 4556
rect 94118 4516 94160 4556
rect 93832 4507 94200 4516
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 19472 3800 19840 3809
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19472 3751 19840 3760
rect 34592 3800 34960 3809
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34592 3751 34960 3760
rect 49712 3800 50080 3809
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 49712 3751 50080 3760
rect 64832 3800 65200 3809
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 64832 3751 65200 3760
rect 79952 3800 80320 3809
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 79952 3751 80320 3760
rect 95072 3800 95440 3809
rect 95112 3760 95154 3800
rect 95194 3760 95236 3800
rect 95276 3760 95318 3800
rect 95358 3760 95400 3800
rect 95072 3751 95440 3760
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 18232 3044 18600 3053
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18232 2995 18600 3004
rect 33352 3044 33720 3053
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33352 2995 33720 3004
rect 48472 3044 48840 3053
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48472 2995 48840 3004
rect 63592 3044 63960 3053
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63592 2995 63960 3004
rect 78712 3044 79080 3053
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 78712 2995 79080 3004
rect 93832 3044 94200 3053
rect 93872 3004 93914 3044
rect 93954 3004 93996 3044
rect 94036 3004 94078 3044
rect 94118 3004 94160 3044
rect 93832 2995 94200 3004
rect 884 2668 1172 2708
rect 844 2659 884 2668
rect 651 2624 693 2633
rect 651 2584 652 2624
rect 692 2584 693 2624
rect 651 2575 693 2584
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 19472 2288 19840 2297
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19472 2239 19840 2248
rect 34592 2288 34960 2297
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34592 2239 34960 2248
rect 49712 2288 50080 2297
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 49712 2239 50080 2248
rect 64832 2288 65200 2297
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 64832 2239 65200 2248
rect 79952 2288 80320 2297
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 79952 2239 80320 2248
rect 95072 2288 95440 2297
rect 95112 2248 95154 2288
rect 95194 2248 95236 2288
rect 95276 2248 95318 2288
rect 95358 2248 95400 2288
rect 95072 2239 95440 2248
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 18232 1532 18600 1541
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18232 1483 18600 1492
rect 33352 1532 33720 1541
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33352 1483 33720 1492
rect 48472 1532 48840 1541
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48472 1483 48840 1492
rect 63592 1532 63960 1541
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63592 1483 63960 1492
rect 78712 1532 79080 1541
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 78712 1483 79080 1492
rect 93832 1532 94200 1541
rect 93872 1492 93914 1532
rect 93954 1492 93996 1532
rect 94036 1492 94078 1532
rect 94118 1492 94160 1532
rect 93832 1483 94200 1492
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
rect 19472 776 19840 785
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19472 727 19840 736
rect 34592 776 34960 785
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34592 727 34960 736
rect 49712 776 50080 785
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 49712 727 50080 736
rect 64832 776 65200 785
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 64832 727 65200 736
rect 79952 776 80320 785
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 79952 727 80320 736
rect 95072 776 95440 785
rect 95112 736 95154 776
rect 95194 736 95236 776
rect 95276 736 95318 776
rect 95358 736 95400 776
rect 95072 727 95440 736
<< via2 >>
rect 3112 81628 3152 81668
rect 3194 81628 3234 81668
rect 3276 81628 3316 81668
rect 3358 81628 3398 81668
rect 3440 81628 3480 81668
rect 18232 81628 18272 81668
rect 18314 81628 18354 81668
rect 18396 81628 18436 81668
rect 18478 81628 18518 81668
rect 18560 81628 18600 81668
rect 33352 81628 33392 81668
rect 33434 81628 33474 81668
rect 33516 81628 33556 81668
rect 33598 81628 33638 81668
rect 33680 81628 33720 81668
rect 48472 81628 48512 81668
rect 48554 81628 48594 81668
rect 48636 81628 48676 81668
rect 48718 81628 48758 81668
rect 48800 81628 48840 81668
rect 63592 81628 63632 81668
rect 63674 81628 63714 81668
rect 63756 81628 63796 81668
rect 63838 81628 63878 81668
rect 63920 81628 63960 81668
rect 78712 81628 78752 81668
rect 78794 81628 78834 81668
rect 78876 81628 78916 81668
rect 78958 81628 78998 81668
rect 79040 81628 79080 81668
rect 93832 81628 93872 81668
rect 93914 81628 93954 81668
rect 93996 81628 94036 81668
rect 94078 81628 94118 81668
rect 94160 81628 94200 81668
rect 4352 80872 4392 80912
rect 4434 80872 4474 80912
rect 4516 80872 4556 80912
rect 4598 80872 4638 80912
rect 4680 80872 4720 80912
rect 19472 80872 19512 80912
rect 19554 80872 19594 80912
rect 19636 80872 19676 80912
rect 19718 80872 19758 80912
rect 19800 80872 19840 80912
rect 34592 80872 34632 80912
rect 34674 80872 34714 80912
rect 34756 80872 34796 80912
rect 34838 80872 34878 80912
rect 34920 80872 34960 80912
rect 49712 80872 49752 80912
rect 49794 80872 49834 80912
rect 49876 80872 49916 80912
rect 49958 80872 49998 80912
rect 50040 80872 50080 80912
rect 64832 80872 64872 80912
rect 64914 80872 64954 80912
rect 64996 80872 65036 80912
rect 65078 80872 65118 80912
rect 65160 80872 65200 80912
rect 79952 80872 79992 80912
rect 80034 80872 80074 80912
rect 80116 80872 80156 80912
rect 80198 80872 80238 80912
rect 80280 80872 80320 80912
rect 95072 80872 95112 80912
rect 95154 80872 95194 80912
rect 95236 80872 95276 80912
rect 95318 80872 95358 80912
rect 95400 80872 95440 80912
rect 3112 80116 3152 80156
rect 3194 80116 3234 80156
rect 3276 80116 3316 80156
rect 3358 80116 3398 80156
rect 3440 80116 3480 80156
rect 18232 80116 18272 80156
rect 18314 80116 18354 80156
rect 18396 80116 18436 80156
rect 18478 80116 18518 80156
rect 18560 80116 18600 80156
rect 33352 80116 33392 80156
rect 33434 80116 33474 80156
rect 33516 80116 33556 80156
rect 33598 80116 33638 80156
rect 33680 80116 33720 80156
rect 48472 80116 48512 80156
rect 48554 80116 48594 80156
rect 48636 80116 48676 80156
rect 48718 80116 48758 80156
rect 48800 80116 48840 80156
rect 63592 80116 63632 80156
rect 63674 80116 63714 80156
rect 63756 80116 63796 80156
rect 63838 80116 63878 80156
rect 63920 80116 63960 80156
rect 78712 80116 78752 80156
rect 78794 80116 78834 80156
rect 78876 80116 78916 80156
rect 78958 80116 78998 80156
rect 79040 80116 79080 80156
rect 93832 80116 93872 80156
rect 93914 80116 93954 80156
rect 93996 80116 94036 80156
rect 94078 80116 94118 80156
rect 94160 80116 94200 80156
rect 4352 79360 4392 79400
rect 4434 79360 4474 79400
rect 4516 79360 4556 79400
rect 4598 79360 4638 79400
rect 4680 79360 4720 79400
rect 19472 79360 19512 79400
rect 19554 79360 19594 79400
rect 19636 79360 19676 79400
rect 19718 79360 19758 79400
rect 19800 79360 19840 79400
rect 34592 79360 34632 79400
rect 34674 79360 34714 79400
rect 34756 79360 34796 79400
rect 34838 79360 34878 79400
rect 34920 79360 34960 79400
rect 49712 79360 49752 79400
rect 49794 79360 49834 79400
rect 49876 79360 49916 79400
rect 49958 79360 49998 79400
rect 50040 79360 50080 79400
rect 64832 79360 64872 79400
rect 64914 79360 64954 79400
rect 64996 79360 65036 79400
rect 65078 79360 65118 79400
rect 65160 79360 65200 79400
rect 79952 79360 79992 79400
rect 80034 79360 80074 79400
rect 80116 79360 80156 79400
rect 80198 79360 80238 79400
rect 80280 79360 80320 79400
rect 95072 79360 95112 79400
rect 95154 79360 95194 79400
rect 95236 79360 95276 79400
rect 95318 79360 95358 79400
rect 95400 79360 95440 79400
rect 3112 78604 3152 78644
rect 3194 78604 3234 78644
rect 3276 78604 3316 78644
rect 3358 78604 3398 78644
rect 3440 78604 3480 78644
rect 18232 78604 18272 78644
rect 18314 78604 18354 78644
rect 18396 78604 18436 78644
rect 18478 78604 18518 78644
rect 18560 78604 18600 78644
rect 33352 78604 33392 78644
rect 33434 78604 33474 78644
rect 33516 78604 33556 78644
rect 33598 78604 33638 78644
rect 33680 78604 33720 78644
rect 48472 78604 48512 78644
rect 48554 78604 48594 78644
rect 48636 78604 48676 78644
rect 48718 78604 48758 78644
rect 48800 78604 48840 78644
rect 63592 78604 63632 78644
rect 63674 78604 63714 78644
rect 63756 78604 63796 78644
rect 63838 78604 63878 78644
rect 63920 78604 63960 78644
rect 78712 78604 78752 78644
rect 78794 78604 78834 78644
rect 78876 78604 78916 78644
rect 78958 78604 78998 78644
rect 79040 78604 79080 78644
rect 93832 78604 93872 78644
rect 93914 78604 93954 78644
rect 93996 78604 94036 78644
rect 94078 78604 94118 78644
rect 94160 78604 94200 78644
rect 4352 77848 4392 77888
rect 4434 77848 4474 77888
rect 4516 77848 4556 77888
rect 4598 77848 4638 77888
rect 4680 77848 4720 77888
rect 19472 77848 19512 77888
rect 19554 77848 19594 77888
rect 19636 77848 19676 77888
rect 19718 77848 19758 77888
rect 19800 77848 19840 77888
rect 34592 77848 34632 77888
rect 34674 77848 34714 77888
rect 34756 77848 34796 77888
rect 34838 77848 34878 77888
rect 34920 77848 34960 77888
rect 49712 77848 49752 77888
rect 49794 77848 49834 77888
rect 49876 77848 49916 77888
rect 49958 77848 49998 77888
rect 50040 77848 50080 77888
rect 64832 77848 64872 77888
rect 64914 77848 64954 77888
rect 64996 77848 65036 77888
rect 65078 77848 65118 77888
rect 65160 77848 65200 77888
rect 79952 77848 79992 77888
rect 80034 77848 80074 77888
rect 80116 77848 80156 77888
rect 80198 77848 80238 77888
rect 80280 77848 80320 77888
rect 95072 77848 95112 77888
rect 95154 77848 95194 77888
rect 95236 77848 95276 77888
rect 95318 77848 95358 77888
rect 95400 77848 95440 77888
rect 3112 77092 3152 77132
rect 3194 77092 3234 77132
rect 3276 77092 3316 77132
rect 3358 77092 3398 77132
rect 3440 77092 3480 77132
rect 18232 77092 18272 77132
rect 18314 77092 18354 77132
rect 18396 77092 18436 77132
rect 18478 77092 18518 77132
rect 18560 77092 18600 77132
rect 33352 77092 33392 77132
rect 33434 77092 33474 77132
rect 33516 77092 33556 77132
rect 33598 77092 33638 77132
rect 33680 77092 33720 77132
rect 48472 77092 48512 77132
rect 48554 77092 48594 77132
rect 48636 77092 48676 77132
rect 48718 77092 48758 77132
rect 48800 77092 48840 77132
rect 63592 77092 63632 77132
rect 63674 77092 63714 77132
rect 63756 77092 63796 77132
rect 63838 77092 63878 77132
rect 63920 77092 63960 77132
rect 78712 77092 78752 77132
rect 78794 77092 78834 77132
rect 78876 77092 78916 77132
rect 78958 77092 78998 77132
rect 79040 77092 79080 77132
rect 93832 77092 93872 77132
rect 93914 77092 93954 77132
rect 93996 77092 94036 77132
rect 94078 77092 94118 77132
rect 94160 77092 94200 77132
rect 4352 76336 4392 76376
rect 4434 76336 4474 76376
rect 4516 76336 4556 76376
rect 4598 76336 4638 76376
rect 4680 76336 4720 76376
rect 19472 76336 19512 76376
rect 19554 76336 19594 76376
rect 19636 76336 19676 76376
rect 19718 76336 19758 76376
rect 19800 76336 19840 76376
rect 34592 76336 34632 76376
rect 34674 76336 34714 76376
rect 34756 76336 34796 76376
rect 34838 76336 34878 76376
rect 34920 76336 34960 76376
rect 49712 76336 49752 76376
rect 49794 76336 49834 76376
rect 49876 76336 49916 76376
rect 49958 76336 49998 76376
rect 50040 76336 50080 76376
rect 64832 76336 64872 76376
rect 64914 76336 64954 76376
rect 64996 76336 65036 76376
rect 65078 76336 65118 76376
rect 65160 76336 65200 76376
rect 79952 76336 79992 76376
rect 80034 76336 80074 76376
rect 80116 76336 80156 76376
rect 80198 76336 80238 76376
rect 80280 76336 80320 76376
rect 95072 76336 95112 76376
rect 95154 76336 95194 76376
rect 95236 76336 95276 76376
rect 95318 76336 95358 76376
rect 95400 76336 95440 76376
rect 3112 75580 3152 75620
rect 3194 75580 3234 75620
rect 3276 75580 3316 75620
rect 3358 75580 3398 75620
rect 3440 75580 3480 75620
rect 18232 75580 18272 75620
rect 18314 75580 18354 75620
rect 18396 75580 18436 75620
rect 18478 75580 18518 75620
rect 18560 75580 18600 75620
rect 33352 75580 33392 75620
rect 33434 75580 33474 75620
rect 33516 75580 33556 75620
rect 33598 75580 33638 75620
rect 33680 75580 33720 75620
rect 48472 75580 48512 75620
rect 48554 75580 48594 75620
rect 48636 75580 48676 75620
rect 48718 75580 48758 75620
rect 48800 75580 48840 75620
rect 63592 75580 63632 75620
rect 63674 75580 63714 75620
rect 63756 75580 63796 75620
rect 63838 75580 63878 75620
rect 63920 75580 63960 75620
rect 78712 75580 78752 75620
rect 78794 75580 78834 75620
rect 78876 75580 78916 75620
rect 78958 75580 78998 75620
rect 79040 75580 79080 75620
rect 93832 75580 93872 75620
rect 93914 75580 93954 75620
rect 93996 75580 94036 75620
rect 94078 75580 94118 75620
rect 94160 75580 94200 75620
rect 652 74656 692 74696
rect 652 72892 692 72932
rect 652 70960 692 71000
rect 652 69196 692 69236
rect 556 67432 596 67472
rect 652 67264 692 67304
rect 652 65416 692 65456
rect 652 63568 692 63608
rect 4352 74824 4392 74864
rect 4434 74824 4474 74864
rect 4516 74824 4556 74864
rect 4598 74824 4638 74864
rect 4680 74824 4720 74864
rect 19472 74824 19512 74864
rect 19554 74824 19594 74864
rect 19636 74824 19676 74864
rect 19718 74824 19758 74864
rect 19800 74824 19840 74864
rect 34592 74824 34632 74864
rect 34674 74824 34714 74864
rect 34756 74824 34796 74864
rect 34838 74824 34878 74864
rect 34920 74824 34960 74864
rect 49712 74824 49752 74864
rect 49794 74824 49834 74864
rect 49876 74824 49916 74864
rect 49958 74824 49998 74864
rect 50040 74824 50080 74864
rect 64832 74824 64872 74864
rect 64914 74824 64954 74864
rect 64996 74824 65036 74864
rect 65078 74824 65118 74864
rect 65160 74824 65200 74864
rect 79952 74824 79992 74864
rect 80034 74824 80074 74864
rect 80116 74824 80156 74864
rect 80198 74824 80238 74864
rect 80280 74824 80320 74864
rect 95072 74824 95112 74864
rect 95154 74824 95194 74864
rect 95236 74824 95276 74864
rect 95318 74824 95358 74864
rect 95400 74824 95440 74864
rect 3112 74068 3152 74108
rect 3194 74068 3234 74108
rect 3276 74068 3316 74108
rect 3358 74068 3398 74108
rect 3440 74068 3480 74108
rect 18232 74068 18272 74108
rect 18314 74068 18354 74108
rect 18396 74068 18436 74108
rect 18478 74068 18518 74108
rect 18560 74068 18600 74108
rect 33352 74068 33392 74108
rect 33434 74068 33474 74108
rect 33516 74068 33556 74108
rect 33598 74068 33638 74108
rect 33680 74068 33720 74108
rect 48472 74068 48512 74108
rect 48554 74068 48594 74108
rect 48636 74068 48676 74108
rect 48718 74068 48758 74108
rect 48800 74068 48840 74108
rect 63592 74068 63632 74108
rect 63674 74068 63714 74108
rect 63756 74068 63796 74108
rect 63838 74068 63878 74108
rect 63920 74068 63960 74108
rect 78712 74068 78752 74108
rect 78794 74068 78834 74108
rect 78876 74068 78916 74108
rect 78958 74068 78998 74108
rect 79040 74068 79080 74108
rect 93832 74068 93872 74108
rect 93914 74068 93954 74108
rect 93996 74068 94036 74108
rect 94078 74068 94118 74108
rect 94160 74068 94200 74108
rect 4352 73312 4392 73352
rect 4434 73312 4474 73352
rect 4516 73312 4556 73352
rect 4598 73312 4638 73352
rect 4680 73312 4720 73352
rect 19472 73312 19512 73352
rect 19554 73312 19594 73352
rect 19636 73312 19676 73352
rect 19718 73312 19758 73352
rect 19800 73312 19840 73352
rect 34592 73312 34632 73352
rect 34674 73312 34714 73352
rect 34756 73312 34796 73352
rect 34838 73312 34878 73352
rect 34920 73312 34960 73352
rect 49712 73312 49752 73352
rect 49794 73312 49834 73352
rect 49876 73312 49916 73352
rect 49958 73312 49998 73352
rect 50040 73312 50080 73352
rect 64832 73312 64872 73352
rect 64914 73312 64954 73352
rect 64996 73312 65036 73352
rect 65078 73312 65118 73352
rect 65160 73312 65200 73352
rect 79952 73312 79992 73352
rect 80034 73312 80074 73352
rect 80116 73312 80156 73352
rect 80198 73312 80238 73352
rect 80280 73312 80320 73352
rect 95072 73312 95112 73352
rect 95154 73312 95194 73352
rect 95236 73312 95276 73352
rect 95318 73312 95358 73352
rect 95400 73312 95440 73352
rect 844 68944 884 68984
rect 844 67432 884 67472
rect 844 65920 884 65960
rect 844 63652 884 63692
rect 748 62980 788 63020
rect 844 62140 884 62180
rect 652 61720 692 61760
rect 844 60292 884 60332
rect 652 59872 692 59912
rect 652 58024 692 58064
rect 844 57100 884 57140
rect 652 56260 692 56300
rect 3112 72556 3152 72596
rect 3194 72556 3234 72596
rect 3276 72556 3316 72596
rect 3358 72556 3398 72596
rect 3440 72556 3480 72596
rect 18232 72556 18272 72596
rect 18314 72556 18354 72596
rect 18396 72556 18436 72596
rect 18478 72556 18518 72596
rect 18560 72556 18600 72596
rect 33352 72556 33392 72596
rect 33434 72556 33474 72596
rect 33516 72556 33556 72596
rect 33598 72556 33638 72596
rect 33680 72556 33720 72596
rect 48472 72556 48512 72596
rect 48554 72556 48594 72596
rect 48636 72556 48676 72596
rect 48718 72556 48758 72596
rect 48800 72556 48840 72596
rect 63592 72556 63632 72596
rect 63674 72556 63714 72596
rect 63756 72556 63796 72596
rect 63838 72556 63878 72596
rect 63920 72556 63960 72596
rect 78712 72556 78752 72596
rect 78794 72556 78834 72596
rect 78876 72556 78916 72596
rect 78958 72556 78998 72596
rect 79040 72556 79080 72596
rect 93832 72556 93872 72596
rect 93914 72556 93954 72596
rect 93996 72556 94036 72596
rect 94078 72556 94118 72596
rect 94160 72556 94200 72596
rect 4352 71800 4392 71840
rect 4434 71800 4474 71840
rect 4516 71800 4556 71840
rect 4598 71800 4638 71840
rect 4680 71800 4720 71840
rect 19472 71800 19512 71840
rect 19554 71800 19594 71840
rect 19636 71800 19676 71840
rect 19718 71800 19758 71840
rect 19800 71800 19840 71840
rect 34592 71800 34632 71840
rect 34674 71800 34714 71840
rect 34756 71800 34796 71840
rect 34838 71800 34878 71840
rect 34920 71800 34960 71840
rect 49712 71800 49752 71840
rect 49794 71800 49834 71840
rect 49876 71800 49916 71840
rect 49958 71800 49998 71840
rect 50040 71800 50080 71840
rect 64832 71800 64872 71840
rect 64914 71800 64954 71840
rect 64996 71800 65036 71840
rect 65078 71800 65118 71840
rect 65160 71800 65200 71840
rect 79952 71800 79992 71840
rect 80034 71800 80074 71840
rect 80116 71800 80156 71840
rect 80198 71800 80238 71840
rect 80280 71800 80320 71840
rect 95072 71800 95112 71840
rect 95154 71800 95194 71840
rect 95236 71800 95276 71840
rect 95318 71800 95358 71840
rect 95400 71800 95440 71840
rect 3112 71044 3152 71084
rect 3194 71044 3234 71084
rect 3276 71044 3316 71084
rect 3358 71044 3398 71084
rect 3440 71044 3480 71084
rect 18232 71044 18272 71084
rect 18314 71044 18354 71084
rect 18396 71044 18436 71084
rect 18478 71044 18518 71084
rect 18560 71044 18600 71084
rect 33352 71044 33392 71084
rect 33434 71044 33474 71084
rect 33516 71044 33556 71084
rect 33598 71044 33638 71084
rect 33680 71044 33720 71084
rect 48472 71044 48512 71084
rect 48554 71044 48594 71084
rect 48636 71044 48676 71084
rect 48718 71044 48758 71084
rect 48800 71044 48840 71084
rect 63592 71044 63632 71084
rect 63674 71044 63714 71084
rect 63756 71044 63796 71084
rect 63838 71044 63878 71084
rect 63920 71044 63960 71084
rect 78712 71044 78752 71084
rect 78794 71044 78834 71084
rect 78876 71044 78916 71084
rect 78958 71044 78998 71084
rect 79040 71044 79080 71084
rect 93832 71044 93872 71084
rect 93914 71044 93954 71084
rect 93996 71044 94036 71084
rect 94078 71044 94118 71084
rect 94160 71044 94200 71084
rect 4352 70288 4392 70328
rect 4434 70288 4474 70328
rect 4516 70288 4556 70328
rect 4598 70288 4638 70328
rect 4680 70288 4720 70328
rect 19472 70288 19512 70328
rect 19554 70288 19594 70328
rect 19636 70288 19676 70328
rect 19718 70288 19758 70328
rect 19800 70288 19840 70328
rect 34592 70288 34632 70328
rect 34674 70288 34714 70328
rect 34756 70288 34796 70328
rect 34838 70288 34878 70328
rect 34920 70288 34960 70328
rect 49712 70288 49752 70328
rect 49794 70288 49834 70328
rect 49876 70288 49916 70328
rect 49958 70288 49998 70328
rect 50040 70288 50080 70328
rect 64832 70288 64872 70328
rect 64914 70288 64954 70328
rect 64996 70288 65036 70328
rect 65078 70288 65118 70328
rect 65160 70288 65200 70328
rect 79952 70288 79992 70328
rect 80034 70288 80074 70328
rect 80116 70288 80156 70328
rect 80198 70288 80238 70328
rect 80280 70288 80320 70328
rect 95072 70288 95112 70328
rect 95154 70288 95194 70328
rect 95236 70288 95276 70328
rect 95318 70288 95358 70328
rect 95400 70288 95440 70328
rect 3112 69532 3152 69572
rect 3194 69532 3234 69572
rect 3276 69532 3316 69572
rect 3358 69532 3398 69572
rect 3440 69532 3480 69572
rect 18232 69532 18272 69572
rect 18314 69532 18354 69572
rect 18396 69532 18436 69572
rect 18478 69532 18518 69572
rect 18560 69532 18600 69572
rect 33352 69532 33392 69572
rect 33434 69532 33474 69572
rect 33516 69532 33556 69572
rect 33598 69532 33638 69572
rect 33680 69532 33720 69572
rect 48472 69532 48512 69572
rect 48554 69532 48594 69572
rect 48636 69532 48676 69572
rect 48718 69532 48758 69572
rect 48800 69532 48840 69572
rect 63592 69532 63632 69572
rect 63674 69532 63714 69572
rect 63756 69532 63796 69572
rect 63838 69532 63878 69572
rect 63920 69532 63960 69572
rect 78712 69532 78752 69572
rect 78794 69532 78834 69572
rect 78876 69532 78916 69572
rect 78958 69532 78998 69572
rect 79040 69532 79080 69572
rect 93832 69532 93872 69572
rect 93914 69532 93954 69572
rect 93996 69532 94036 69572
rect 94078 69532 94118 69572
rect 94160 69532 94200 69572
rect 1228 68944 1268 68984
rect 1132 65920 1172 65960
rect 1036 57940 1076 57980
rect 748 56092 788 56132
rect 652 54328 692 54368
rect 652 52564 692 52604
rect 1036 52816 1076 52856
rect 940 52648 980 52688
rect 844 52480 884 52520
rect 652 50632 692 50672
rect 844 49456 884 49496
rect 652 48784 692 48824
rect 748 47860 788 47900
rect 556 47272 596 47312
rect 652 46936 692 46976
rect 652 45088 692 45128
rect 652 43240 692 43280
rect 844 47524 884 47564
rect 1036 47440 1076 47480
rect 844 45928 884 45968
rect 652 41392 692 41432
rect 652 39544 692 39584
rect 652 37696 692 37736
rect 652 35848 692 35888
rect 652 34000 692 34040
rect 652 32152 692 32192
rect 652 30304 692 30344
rect 652 28456 692 28496
rect 652 26608 692 26648
rect 652 24760 692 24800
rect 652 22912 692 22952
rect 652 21064 692 21104
rect 652 19216 692 19256
rect 652 17368 692 17408
rect 844 16276 884 16316
rect 652 15520 692 15560
rect 652 13756 692 13796
rect 652 11824 692 11864
rect 652 9976 692 10016
rect 652 8128 692 8168
rect 4352 68776 4392 68816
rect 4434 68776 4474 68816
rect 4516 68776 4556 68816
rect 4598 68776 4638 68816
rect 4680 68776 4720 68816
rect 19472 68776 19512 68816
rect 19554 68776 19594 68816
rect 19636 68776 19676 68816
rect 19718 68776 19758 68816
rect 19800 68776 19840 68816
rect 34592 68776 34632 68816
rect 34674 68776 34714 68816
rect 34756 68776 34796 68816
rect 34838 68776 34878 68816
rect 34920 68776 34960 68816
rect 49712 68776 49752 68816
rect 49794 68776 49834 68816
rect 49876 68776 49916 68816
rect 49958 68776 49998 68816
rect 50040 68776 50080 68816
rect 64832 68776 64872 68816
rect 64914 68776 64954 68816
rect 64996 68776 65036 68816
rect 65078 68776 65118 68816
rect 65160 68776 65200 68816
rect 79952 68776 79992 68816
rect 80034 68776 80074 68816
rect 80116 68776 80156 68816
rect 80198 68776 80238 68816
rect 80280 68776 80320 68816
rect 95072 68776 95112 68816
rect 95154 68776 95194 68816
rect 95236 68776 95276 68816
rect 95318 68776 95358 68816
rect 95400 68776 95440 68816
rect 3112 68020 3152 68060
rect 3194 68020 3234 68060
rect 3276 68020 3316 68060
rect 3358 68020 3398 68060
rect 3440 68020 3480 68060
rect 18232 68020 18272 68060
rect 18314 68020 18354 68060
rect 18396 68020 18436 68060
rect 18478 68020 18518 68060
rect 18560 68020 18600 68060
rect 33352 68020 33392 68060
rect 33434 68020 33474 68060
rect 33516 68020 33556 68060
rect 33598 68020 33638 68060
rect 33680 68020 33720 68060
rect 48472 68020 48512 68060
rect 48554 68020 48594 68060
rect 48636 68020 48676 68060
rect 48718 68020 48758 68060
rect 48800 68020 48840 68060
rect 63592 68020 63632 68060
rect 63674 68020 63714 68060
rect 63756 68020 63796 68060
rect 63838 68020 63878 68060
rect 63920 68020 63960 68060
rect 78712 68020 78752 68060
rect 78794 68020 78834 68060
rect 78876 68020 78916 68060
rect 78958 68020 78998 68060
rect 79040 68020 79080 68060
rect 93832 68020 93872 68060
rect 93914 68020 93954 68060
rect 93996 68020 94036 68060
rect 94078 68020 94118 68060
rect 94160 68020 94200 68060
rect 4352 67264 4392 67304
rect 4434 67264 4474 67304
rect 4516 67264 4556 67304
rect 4598 67264 4638 67304
rect 4680 67264 4720 67304
rect 19472 67264 19512 67304
rect 19554 67264 19594 67304
rect 19636 67264 19676 67304
rect 19718 67264 19758 67304
rect 19800 67264 19840 67304
rect 34592 67264 34632 67304
rect 34674 67264 34714 67304
rect 34756 67264 34796 67304
rect 34838 67264 34878 67304
rect 34920 67264 34960 67304
rect 49712 67264 49752 67304
rect 49794 67264 49834 67304
rect 49876 67264 49916 67304
rect 49958 67264 49998 67304
rect 50040 67264 50080 67304
rect 64832 67264 64872 67304
rect 64914 67264 64954 67304
rect 64996 67264 65036 67304
rect 65078 67264 65118 67304
rect 65160 67264 65200 67304
rect 79952 67264 79992 67304
rect 80034 67264 80074 67304
rect 80116 67264 80156 67304
rect 80198 67264 80238 67304
rect 80280 67264 80320 67304
rect 95072 67264 95112 67304
rect 95154 67264 95194 67304
rect 95236 67264 95276 67304
rect 95318 67264 95358 67304
rect 95400 67264 95440 67304
rect 3112 66508 3152 66548
rect 3194 66508 3234 66548
rect 3276 66508 3316 66548
rect 3358 66508 3398 66548
rect 3440 66508 3480 66548
rect 18232 66508 18272 66548
rect 18314 66508 18354 66548
rect 18396 66508 18436 66548
rect 18478 66508 18518 66548
rect 18560 66508 18600 66548
rect 33352 66508 33392 66548
rect 33434 66508 33474 66548
rect 33516 66508 33556 66548
rect 33598 66508 33638 66548
rect 33680 66508 33720 66548
rect 48472 66508 48512 66548
rect 48554 66508 48594 66548
rect 48636 66508 48676 66548
rect 48718 66508 48758 66548
rect 48800 66508 48840 66548
rect 63592 66508 63632 66548
rect 63674 66508 63714 66548
rect 63756 66508 63796 66548
rect 63838 66508 63878 66548
rect 63920 66508 63960 66548
rect 78712 66508 78752 66548
rect 78794 66508 78834 66548
rect 78876 66508 78916 66548
rect 78958 66508 78998 66548
rect 79040 66508 79080 66548
rect 93832 66508 93872 66548
rect 93914 66508 93954 66548
rect 93996 66508 94036 66548
rect 94078 66508 94118 66548
rect 94160 66508 94200 66548
rect 4352 65752 4392 65792
rect 4434 65752 4474 65792
rect 4516 65752 4556 65792
rect 4598 65752 4638 65792
rect 4680 65752 4720 65792
rect 19472 65752 19512 65792
rect 19554 65752 19594 65792
rect 19636 65752 19676 65792
rect 19718 65752 19758 65792
rect 19800 65752 19840 65792
rect 34592 65752 34632 65792
rect 34674 65752 34714 65792
rect 34756 65752 34796 65792
rect 34838 65752 34878 65792
rect 34920 65752 34960 65792
rect 49712 65752 49752 65792
rect 49794 65752 49834 65792
rect 49876 65752 49916 65792
rect 49958 65752 49998 65792
rect 50040 65752 50080 65792
rect 64832 65752 64872 65792
rect 64914 65752 64954 65792
rect 64996 65752 65036 65792
rect 65078 65752 65118 65792
rect 65160 65752 65200 65792
rect 79952 65752 79992 65792
rect 80034 65752 80074 65792
rect 80116 65752 80156 65792
rect 80198 65752 80238 65792
rect 80280 65752 80320 65792
rect 95072 65752 95112 65792
rect 95154 65752 95194 65792
rect 95236 65752 95276 65792
rect 95318 65752 95358 65792
rect 95400 65752 95440 65792
rect 3112 64996 3152 65036
rect 3194 64996 3234 65036
rect 3276 64996 3316 65036
rect 3358 64996 3398 65036
rect 3440 64996 3480 65036
rect 18232 64996 18272 65036
rect 18314 64996 18354 65036
rect 18396 64996 18436 65036
rect 18478 64996 18518 65036
rect 18560 64996 18600 65036
rect 33352 64996 33392 65036
rect 33434 64996 33474 65036
rect 33516 64996 33556 65036
rect 33598 64996 33638 65036
rect 33680 64996 33720 65036
rect 48472 64996 48512 65036
rect 48554 64996 48594 65036
rect 48636 64996 48676 65036
rect 48718 64996 48758 65036
rect 48800 64996 48840 65036
rect 63592 64996 63632 65036
rect 63674 64996 63714 65036
rect 63756 64996 63796 65036
rect 63838 64996 63878 65036
rect 63920 64996 63960 65036
rect 78712 64996 78752 65036
rect 78794 64996 78834 65036
rect 78876 64996 78916 65036
rect 78958 64996 78998 65036
rect 79040 64996 79080 65036
rect 93832 64996 93872 65036
rect 93914 64996 93954 65036
rect 93996 64996 94036 65036
rect 94078 64996 94118 65036
rect 94160 64996 94200 65036
rect 4352 64240 4392 64280
rect 4434 64240 4474 64280
rect 4516 64240 4556 64280
rect 4598 64240 4638 64280
rect 4680 64240 4720 64280
rect 19472 64240 19512 64280
rect 19554 64240 19594 64280
rect 19636 64240 19676 64280
rect 19718 64240 19758 64280
rect 19800 64240 19840 64280
rect 34592 64240 34632 64280
rect 34674 64240 34714 64280
rect 34756 64240 34796 64280
rect 34838 64240 34878 64280
rect 34920 64240 34960 64280
rect 49712 64240 49752 64280
rect 49794 64240 49834 64280
rect 49876 64240 49916 64280
rect 49958 64240 49998 64280
rect 50040 64240 50080 64280
rect 64832 64240 64872 64280
rect 64914 64240 64954 64280
rect 64996 64240 65036 64280
rect 65078 64240 65118 64280
rect 65160 64240 65200 64280
rect 79952 64240 79992 64280
rect 80034 64240 80074 64280
rect 80116 64240 80156 64280
rect 80198 64240 80238 64280
rect 80280 64240 80320 64280
rect 95072 64240 95112 64280
rect 95154 64240 95194 64280
rect 95236 64240 95276 64280
rect 95318 64240 95358 64280
rect 95400 64240 95440 64280
rect 13228 63652 13268 63692
rect 3112 63484 3152 63524
rect 3194 63484 3234 63524
rect 3276 63484 3316 63524
rect 3358 63484 3398 63524
rect 3440 63484 3480 63524
rect 6508 62980 6548 63020
rect 4352 62728 4392 62768
rect 4434 62728 4474 62768
rect 4516 62728 4556 62768
rect 4598 62728 4638 62768
rect 4680 62728 4720 62768
rect 3112 61972 3152 62012
rect 3194 61972 3234 62012
rect 3276 61972 3316 62012
rect 3358 61972 3398 62012
rect 3440 61972 3480 62012
rect 4352 61216 4392 61256
rect 4434 61216 4474 61256
rect 4516 61216 4556 61256
rect 4598 61216 4638 61256
rect 4680 61216 4720 61256
rect 3112 60460 3152 60500
rect 3194 60460 3234 60500
rect 3276 60460 3316 60500
rect 3358 60460 3398 60500
rect 3440 60460 3480 60500
rect 6604 60292 6644 60332
rect 4352 59704 4392 59744
rect 4434 59704 4474 59744
rect 4516 59704 4556 59744
rect 4598 59704 4638 59744
rect 4680 59704 4720 59744
rect 3112 58948 3152 58988
rect 3194 58948 3234 58988
rect 3276 58948 3316 58988
rect 3358 58948 3398 58988
rect 3440 58948 3480 58988
rect 4352 58192 4392 58232
rect 4434 58192 4474 58232
rect 4516 58192 4556 58232
rect 4598 58192 4638 58232
rect 4680 58192 4720 58232
rect 5836 57940 5876 57980
rect 3112 57436 3152 57476
rect 3194 57436 3234 57476
rect 3276 57436 3316 57476
rect 3358 57436 3398 57476
rect 3440 57436 3480 57476
rect 6220 57856 6260 57896
rect 6316 57856 6356 57896
rect 6508 57856 6548 57896
rect 6028 57100 6068 57140
rect 6220 57100 6260 57140
rect 5932 57016 5972 57056
rect 5836 56932 5876 56972
rect 6508 57016 6548 57056
rect 4352 56680 4392 56720
rect 4434 56680 4474 56720
rect 4516 56680 4556 56720
rect 4598 56680 4638 56720
rect 4680 56680 4720 56720
rect 5644 56344 5684 56384
rect 6604 56344 6644 56384
rect 3112 55924 3152 55964
rect 3194 55924 3234 55964
rect 3276 55924 3316 55964
rect 3358 55924 3398 55964
rect 3440 55924 3480 55964
rect 4352 55168 4392 55208
rect 4434 55168 4474 55208
rect 4516 55168 4556 55208
rect 4598 55168 4638 55208
rect 4680 55168 4720 55208
rect 3112 54412 3152 54452
rect 3194 54412 3234 54452
rect 3276 54412 3316 54452
rect 3358 54412 3398 54452
rect 3440 54412 3480 54452
rect 4352 53656 4392 53696
rect 4434 53656 4474 53696
rect 4516 53656 4556 53696
rect 4598 53656 4638 53696
rect 4680 53656 4720 53696
rect 3112 52900 3152 52940
rect 3194 52900 3234 52940
rect 3276 52900 3316 52940
rect 3358 52900 3398 52940
rect 3440 52900 3480 52940
rect 7180 57016 7220 57056
rect 6988 56344 7028 56384
rect 6412 56092 6452 56132
rect 5836 53068 5876 53108
rect 6412 53068 6452 53108
rect 5740 52564 5780 52604
rect 2284 52480 2324 52520
rect 4108 52480 4148 52520
rect 2188 51976 2228 52016
rect 1228 51808 1268 51848
rect 2092 51808 2132 51848
rect 3244 51976 3284 52016
rect 2956 51892 2996 51932
rect 2764 51808 2804 51848
rect 3916 51892 3956 51932
rect 3436 51808 3476 51848
rect 4012 51808 4052 51848
rect 4352 52144 4392 52184
rect 4434 52144 4474 52184
rect 4516 52144 4556 52184
rect 4598 52144 4638 52184
rect 4680 52144 4720 52184
rect 5548 51976 5588 52016
rect 5260 51808 5300 51848
rect 5452 51808 5492 51848
rect 6185 52816 6225 52856
rect 6508 52816 6548 52856
rect 6028 52648 6068 52688
rect 5932 52480 5972 52520
rect 6316 52564 6356 52604
rect 6220 52312 6260 52352
rect 6700 52648 6740 52688
rect 6412 52312 6452 52352
rect 5932 51724 5972 51764
rect 6124 51724 6164 51764
rect 2668 51640 2708 51680
rect 3112 51388 3152 51428
rect 3194 51388 3234 51428
rect 3276 51388 3316 51428
rect 3358 51388 3398 51428
rect 3440 51388 3480 51428
rect 1900 50800 1940 50840
rect 2476 50800 2516 50840
rect 1132 45760 1172 45800
rect 1132 44752 1172 44792
rect 844 12412 884 12452
rect 844 10228 884 10268
rect 844 8716 884 8756
rect 652 6280 692 6320
rect 844 4852 884 4892
rect 652 4432 692 4472
rect 4352 50632 4392 50672
rect 4434 50632 4474 50672
rect 4516 50632 4556 50672
rect 4598 50632 4638 50672
rect 4680 50632 4720 50672
rect 3112 49876 3152 49916
rect 3194 49876 3234 49916
rect 3276 49876 3316 49916
rect 3358 49876 3398 49916
rect 3440 49876 3480 49916
rect 4352 49120 4392 49160
rect 4434 49120 4474 49160
rect 4516 49120 4556 49160
rect 4598 49120 4638 49160
rect 4680 49120 4720 49160
rect 3112 48364 3152 48404
rect 3194 48364 3234 48404
rect 3276 48364 3316 48404
rect 3358 48364 3398 48404
rect 3440 48364 3480 48404
rect 3916 47944 3956 47984
rect 6412 51808 6452 51848
rect 6796 51808 6836 51848
rect 6220 51640 6260 51680
rect 6892 51640 6932 51680
rect 6220 47944 6260 47984
rect 1996 47440 2036 47480
rect 2284 47440 2324 47480
rect 4352 47608 4392 47648
rect 4434 47608 4474 47648
rect 4516 47608 4556 47648
rect 4598 47608 4638 47648
rect 4680 47608 4720 47648
rect 4012 47440 4052 47480
rect 6412 47944 6452 47984
rect 2476 47356 2516 47396
rect 2956 47356 2996 47396
rect 2092 47272 2132 47312
rect 2764 47272 2804 47312
rect 5836 47356 5876 47396
rect 6604 47356 6644 47396
rect 6508 47272 6548 47312
rect 5932 47188 5972 47228
rect 3820 47104 3860 47144
rect 3112 46852 3152 46892
rect 3194 46852 3234 46892
rect 3276 46852 3316 46892
rect 3358 46852 3398 46892
rect 3440 46852 3480 46892
rect 4352 46096 4392 46136
rect 4434 46096 4474 46136
rect 4516 46096 4556 46136
rect 4598 46096 4638 46136
rect 4680 46096 4720 46136
rect 3112 45340 3152 45380
rect 3194 45340 3234 45380
rect 3276 45340 3316 45380
rect 3358 45340 3398 45380
rect 3440 45340 3480 45380
rect 4352 44584 4392 44624
rect 4434 44584 4474 44624
rect 4516 44584 4556 44624
rect 4598 44584 4638 44624
rect 4680 44584 4720 44624
rect 3112 43828 3152 43868
rect 3194 43828 3234 43868
rect 3276 43828 3316 43868
rect 3358 43828 3398 43868
rect 3440 43828 3480 43868
rect 4352 43072 4392 43112
rect 4434 43072 4474 43112
rect 4516 43072 4556 43112
rect 4598 43072 4638 43112
rect 4680 43072 4720 43112
rect 3112 42316 3152 42356
rect 3194 42316 3234 42356
rect 3276 42316 3316 42356
rect 3358 42316 3398 42356
rect 3440 42316 3480 42356
rect 4352 41560 4392 41600
rect 4434 41560 4474 41600
rect 4516 41560 4556 41600
rect 4598 41560 4638 41600
rect 4680 41560 4720 41600
rect 3112 40804 3152 40844
rect 3194 40804 3234 40844
rect 3276 40804 3316 40844
rect 3358 40804 3398 40844
rect 3440 40804 3480 40844
rect 4352 40048 4392 40088
rect 4434 40048 4474 40088
rect 4516 40048 4556 40088
rect 4598 40048 4638 40088
rect 4680 40048 4720 40088
rect 3112 39292 3152 39332
rect 3194 39292 3234 39332
rect 3276 39292 3316 39332
rect 3358 39292 3398 39332
rect 3440 39292 3480 39332
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 1900 12412 1940 12452
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 6892 47188 6932 47228
rect 6988 47104 7028 47144
rect 6796 47020 6836 47060
rect 7852 49456 7892 49496
rect 7564 47944 7604 47984
rect 7372 47272 7412 47312
rect 7372 47104 7412 47144
rect 7564 47020 7604 47060
rect 9388 47860 9428 47900
rect 9868 47944 9908 47984
rect 13132 47524 13172 47564
rect 18232 63484 18272 63524
rect 18314 63484 18354 63524
rect 18396 63484 18436 63524
rect 18478 63484 18518 63524
rect 18560 63484 18600 63524
rect 33352 63484 33392 63524
rect 33434 63484 33474 63524
rect 33516 63484 33556 63524
rect 33598 63484 33638 63524
rect 33680 63484 33720 63524
rect 48472 63484 48512 63524
rect 48554 63484 48594 63524
rect 48636 63484 48676 63524
rect 48718 63484 48758 63524
rect 48800 63484 48840 63524
rect 63592 63484 63632 63524
rect 63674 63484 63714 63524
rect 63756 63484 63796 63524
rect 63838 63484 63878 63524
rect 63920 63484 63960 63524
rect 78712 63484 78752 63524
rect 78794 63484 78834 63524
rect 78876 63484 78916 63524
rect 78958 63484 78998 63524
rect 79040 63484 79080 63524
rect 93832 63484 93872 63524
rect 93914 63484 93954 63524
rect 93996 63484 94036 63524
rect 94078 63484 94118 63524
rect 94160 63484 94200 63524
rect 19472 62728 19512 62768
rect 19554 62728 19594 62768
rect 19636 62728 19676 62768
rect 19718 62728 19758 62768
rect 19800 62728 19840 62768
rect 34592 62728 34632 62768
rect 34674 62728 34714 62768
rect 34756 62728 34796 62768
rect 34838 62728 34878 62768
rect 34920 62728 34960 62768
rect 49712 62728 49752 62768
rect 49794 62728 49834 62768
rect 49876 62728 49916 62768
rect 49958 62728 49998 62768
rect 50040 62728 50080 62768
rect 64832 62728 64872 62768
rect 64914 62728 64954 62768
rect 64996 62728 65036 62768
rect 65078 62728 65118 62768
rect 65160 62728 65200 62768
rect 79952 62728 79992 62768
rect 80034 62728 80074 62768
rect 80116 62728 80156 62768
rect 80198 62728 80238 62768
rect 80280 62728 80320 62768
rect 95072 62728 95112 62768
rect 95154 62728 95194 62768
rect 95236 62728 95276 62768
rect 95318 62728 95358 62768
rect 95400 62728 95440 62768
rect 14188 62140 14228 62180
rect 13804 47944 13844 47984
rect 13612 47524 13652 47564
rect 8044 47272 8084 47312
rect 9484 47272 9524 47312
rect 13228 47272 13268 47312
rect 13900 47272 13940 47312
rect 14092 47272 14132 47312
rect 14092 46432 14132 46472
rect 7756 45760 7796 45800
rect 8236 45760 8276 45800
rect 14092 45928 14132 45968
rect 18232 61972 18272 62012
rect 18314 61972 18354 62012
rect 18396 61972 18436 62012
rect 18478 61972 18518 62012
rect 18560 61972 18600 62012
rect 33352 61972 33392 62012
rect 33434 61972 33474 62012
rect 33516 61972 33556 62012
rect 33598 61972 33638 62012
rect 33680 61972 33720 62012
rect 48472 61972 48512 62012
rect 48554 61972 48594 62012
rect 48636 61972 48676 62012
rect 48718 61972 48758 62012
rect 48800 61972 48840 62012
rect 63592 61972 63632 62012
rect 63674 61972 63714 62012
rect 63756 61972 63796 62012
rect 63838 61972 63878 62012
rect 63920 61972 63960 62012
rect 78712 61972 78752 62012
rect 78794 61972 78834 62012
rect 78876 61972 78916 62012
rect 78958 61972 78998 62012
rect 79040 61972 79080 62012
rect 93832 61972 93872 62012
rect 93914 61972 93954 62012
rect 93996 61972 94036 62012
rect 94078 61972 94118 62012
rect 94160 61972 94200 62012
rect 19472 61216 19512 61256
rect 19554 61216 19594 61256
rect 19636 61216 19676 61256
rect 19718 61216 19758 61256
rect 19800 61216 19840 61256
rect 34592 61216 34632 61256
rect 34674 61216 34714 61256
rect 34756 61216 34796 61256
rect 34838 61216 34878 61256
rect 34920 61216 34960 61256
rect 49712 61216 49752 61256
rect 49794 61216 49834 61256
rect 49876 61216 49916 61256
rect 49958 61216 49998 61256
rect 50040 61216 50080 61256
rect 64832 61216 64872 61256
rect 64914 61216 64954 61256
rect 64996 61216 65036 61256
rect 65078 61216 65118 61256
rect 65160 61216 65200 61256
rect 79952 61216 79992 61256
rect 80034 61216 80074 61256
rect 80116 61216 80156 61256
rect 80198 61216 80238 61256
rect 80280 61216 80320 61256
rect 95072 61216 95112 61256
rect 95154 61216 95194 61256
rect 95236 61216 95276 61256
rect 95318 61216 95358 61256
rect 95400 61216 95440 61256
rect 18232 60460 18272 60500
rect 18314 60460 18354 60500
rect 18396 60460 18436 60500
rect 18478 60460 18518 60500
rect 18560 60460 18600 60500
rect 33352 60460 33392 60500
rect 33434 60460 33474 60500
rect 33516 60460 33556 60500
rect 33598 60460 33638 60500
rect 33680 60460 33720 60500
rect 48472 60460 48512 60500
rect 48554 60460 48594 60500
rect 48636 60460 48676 60500
rect 48718 60460 48758 60500
rect 48800 60460 48840 60500
rect 63592 60460 63632 60500
rect 63674 60460 63714 60500
rect 63756 60460 63796 60500
rect 63838 60460 63878 60500
rect 63920 60460 63960 60500
rect 78712 60460 78752 60500
rect 78794 60460 78834 60500
rect 78876 60460 78916 60500
rect 78958 60460 78998 60500
rect 79040 60460 79080 60500
rect 93832 60460 93872 60500
rect 93914 60460 93954 60500
rect 93996 60460 94036 60500
rect 94078 60460 94118 60500
rect 94160 60460 94200 60500
rect 19472 59704 19512 59744
rect 19554 59704 19594 59744
rect 19636 59704 19676 59744
rect 19718 59704 19758 59744
rect 19800 59704 19840 59744
rect 34592 59704 34632 59744
rect 34674 59704 34714 59744
rect 34756 59704 34796 59744
rect 34838 59704 34878 59744
rect 34920 59704 34960 59744
rect 49712 59704 49752 59744
rect 49794 59704 49834 59744
rect 49876 59704 49916 59744
rect 49958 59704 49998 59744
rect 50040 59704 50080 59744
rect 64832 59704 64872 59744
rect 64914 59704 64954 59744
rect 64996 59704 65036 59744
rect 65078 59704 65118 59744
rect 65160 59704 65200 59744
rect 79952 59704 79992 59744
rect 80034 59704 80074 59744
rect 80116 59704 80156 59744
rect 80198 59704 80238 59744
rect 80280 59704 80320 59744
rect 95072 59704 95112 59744
rect 95154 59704 95194 59744
rect 95236 59704 95276 59744
rect 95318 59704 95358 59744
rect 95400 59704 95440 59744
rect 18232 58948 18272 58988
rect 18314 58948 18354 58988
rect 18396 58948 18436 58988
rect 18478 58948 18518 58988
rect 18560 58948 18600 58988
rect 33352 58948 33392 58988
rect 33434 58948 33474 58988
rect 33516 58948 33556 58988
rect 33598 58948 33638 58988
rect 33680 58948 33720 58988
rect 48472 58948 48512 58988
rect 48554 58948 48594 58988
rect 48636 58948 48676 58988
rect 48718 58948 48758 58988
rect 48800 58948 48840 58988
rect 63592 58948 63632 58988
rect 63674 58948 63714 58988
rect 63756 58948 63796 58988
rect 63838 58948 63878 58988
rect 63920 58948 63960 58988
rect 78712 58948 78752 58988
rect 78794 58948 78834 58988
rect 78876 58948 78916 58988
rect 78958 58948 78998 58988
rect 79040 58948 79080 58988
rect 93832 58948 93872 58988
rect 93914 58948 93954 58988
rect 93996 58948 94036 58988
rect 94078 58948 94118 58988
rect 94160 58948 94200 58988
rect 19472 58192 19512 58232
rect 19554 58192 19594 58232
rect 19636 58192 19676 58232
rect 19718 58192 19758 58232
rect 19800 58192 19840 58232
rect 34592 58192 34632 58232
rect 34674 58192 34714 58232
rect 34756 58192 34796 58232
rect 34838 58192 34878 58232
rect 34920 58192 34960 58232
rect 49712 58192 49752 58232
rect 49794 58192 49834 58232
rect 49876 58192 49916 58232
rect 49958 58192 49998 58232
rect 50040 58192 50080 58232
rect 64832 58192 64872 58232
rect 64914 58192 64954 58232
rect 64996 58192 65036 58232
rect 65078 58192 65118 58232
rect 65160 58192 65200 58232
rect 79952 58192 79992 58232
rect 80034 58192 80074 58232
rect 80116 58192 80156 58232
rect 80198 58192 80238 58232
rect 80280 58192 80320 58232
rect 95072 58192 95112 58232
rect 95154 58192 95194 58232
rect 95236 58192 95276 58232
rect 95318 58192 95358 58232
rect 95400 58192 95440 58232
rect 18232 57436 18272 57476
rect 18314 57436 18354 57476
rect 18396 57436 18436 57476
rect 18478 57436 18518 57476
rect 18560 57436 18600 57476
rect 33352 57436 33392 57476
rect 33434 57436 33474 57476
rect 33516 57436 33556 57476
rect 33598 57436 33638 57476
rect 33680 57436 33720 57476
rect 48472 57436 48512 57476
rect 48554 57436 48594 57476
rect 48636 57436 48676 57476
rect 48718 57436 48758 57476
rect 48800 57436 48840 57476
rect 63592 57436 63632 57476
rect 63674 57436 63714 57476
rect 63756 57436 63796 57476
rect 63838 57436 63878 57476
rect 63920 57436 63960 57476
rect 78712 57436 78752 57476
rect 78794 57436 78834 57476
rect 78876 57436 78916 57476
rect 78958 57436 78998 57476
rect 79040 57436 79080 57476
rect 93832 57436 93872 57476
rect 93914 57436 93954 57476
rect 93996 57436 94036 57476
rect 94078 57436 94118 57476
rect 94160 57436 94200 57476
rect 19472 56680 19512 56720
rect 19554 56680 19594 56720
rect 19636 56680 19676 56720
rect 19718 56680 19758 56720
rect 19800 56680 19840 56720
rect 34592 56680 34632 56720
rect 34674 56680 34714 56720
rect 34756 56680 34796 56720
rect 34838 56680 34878 56720
rect 34920 56680 34960 56720
rect 49712 56680 49752 56720
rect 49794 56680 49834 56720
rect 49876 56680 49916 56720
rect 49958 56680 49998 56720
rect 50040 56680 50080 56720
rect 64832 56680 64872 56720
rect 64914 56680 64954 56720
rect 64996 56680 65036 56720
rect 65078 56680 65118 56720
rect 65160 56680 65200 56720
rect 79952 56680 79992 56720
rect 80034 56680 80074 56720
rect 80116 56680 80156 56720
rect 80198 56680 80238 56720
rect 80280 56680 80320 56720
rect 95072 56680 95112 56720
rect 95154 56680 95194 56720
rect 95236 56680 95276 56720
rect 95318 56680 95358 56720
rect 95400 56680 95440 56720
rect 18232 55924 18272 55964
rect 18314 55924 18354 55964
rect 18396 55924 18436 55964
rect 18478 55924 18518 55964
rect 18560 55924 18600 55964
rect 33352 55924 33392 55964
rect 33434 55924 33474 55964
rect 33516 55924 33556 55964
rect 33598 55924 33638 55964
rect 33680 55924 33720 55964
rect 48472 55924 48512 55964
rect 48554 55924 48594 55964
rect 48636 55924 48676 55964
rect 48718 55924 48758 55964
rect 48800 55924 48840 55964
rect 63592 55924 63632 55964
rect 63674 55924 63714 55964
rect 63756 55924 63796 55964
rect 63838 55924 63878 55964
rect 63920 55924 63960 55964
rect 78712 55924 78752 55964
rect 78794 55924 78834 55964
rect 78876 55924 78916 55964
rect 78958 55924 78998 55964
rect 79040 55924 79080 55964
rect 93832 55924 93872 55964
rect 93914 55924 93954 55964
rect 93996 55924 94036 55964
rect 94078 55924 94118 55964
rect 94160 55924 94200 55964
rect 19472 55168 19512 55208
rect 19554 55168 19594 55208
rect 19636 55168 19676 55208
rect 19718 55168 19758 55208
rect 19800 55168 19840 55208
rect 34592 55168 34632 55208
rect 34674 55168 34714 55208
rect 34756 55168 34796 55208
rect 34838 55168 34878 55208
rect 34920 55168 34960 55208
rect 49712 55168 49752 55208
rect 49794 55168 49834 55208
rect 49876 55168 49916 55208
rect 49958 55168 49998 55208
rect 50040 55168 50080 55208
rect 64832 55168 64872 55208
rect 64914 55168 64954 55208
rect 64996 55168 65036 55208
rect 65078 55168 65118 55208
rect 65160 55168 65200 55208
rect 79952 55168 79992 55208
rect 80034 55168 80074 55208
rect 80116 55168 80156 55208
rect 80198 55168 80238 55208
rect 80280 55168 80320 55208
rect 95072 55168 95112 55208
rect 95154 55168 95194 55208
rect 95236 55168 95276 55208
rect 95318 55168 95358 55208
rect 95400 55168 95440 55208
rect 18232 54412 18272 54452
rect 18314 54412 18354 54452
rect 18396 54412 18436 54452
rect 18478 54412 18518 54452
rect 18560 54412 18600 54452
rect 33352 54412 33392 54452
rect 33434 54412 33474 54452
rect 33516 54412 33556 54452
rect 33598 54412 33638 54452
rect 33680 54412 33720 54452
rect 48472 54412 48512 54452
rect 48554 54412 48594 54452
rect 48636 54412 48676 54452
rect 48718 54412 48758 54452
rect 48800 54412 48840 54452
rect 63592 54412 63632 54452
rect 63674 54412 63714 54452
rect 63756 54412 63796 54452
rect 63838 54412 63878 54452
rect 63920 54412 63960 54452
rect 78712 54412 78752 54452
rect 78794 54412 78834 54452
rect 78876 54412 78916 54452
rect 78958 54412 78998 54452
rect 79040 54412 79080 54452
rect 93832 54412 93872 54452
rect 93914 54412 93954 54452
rect 93996 54412 94036 54452
rect 94078 54412 94118 54452
rect 94160 54412 94200 54452
rect 19472 53656 19512 53696
rect 19554 53656 19594 53696
rect 19636 53656 19676 53696
rect 19718 53656 19758 53696
rect 19800 53656 19840 53696
rect 34592 53656 34632 53696
rect 34674 53656 34714 53696
rect 34756 53656 34796 53696
rect 34838 53656 34878 53696
rect 34920 53656 34960 53696
rect 49712 53656 49752 53696
rect 49794 53656 49834 53696
rect 49876 53656 49916 53696
rect 49958 53656 49998 53696
rect 50040 53656 50080 53696
rect 64832 53656 64872 53696
rect 64914 53656 64954 53696
rect 64996 53656 65036 53696
rect 65078 53656 65118 53696
rect 65160 53656 65200 53696
rect 79952 53656 79992 53696
rect 80034 53656 80074 53696
rect 80116 53656 80156 53696
rect 80198 53656 80238 53696
rect 80280 53656 80320 53696
rect 95072 53656 95112 53696
rect 95154 53656 95194 53696
rect 95236 53656 95276 53696
rect 95318 53656 95358 53696
rect 95400 53656 95440 53696
rect 18232 52900 18272 52940
rect 18314 52900 18354 52940
rect 18396 52900 18436 52940
rect 18478 52900 18518 52940
rect 18560 52900 18600 52940
rect 33352 52900 33392 52940
rect 33434 52900 33474 52940
rect 33516 52900 33556 52940
rect 33598 52900 33638 52940
rect 33680 52900 33720 52940
rect 48472 52900 48512 52940
rect 48554 52900 48594 52940
rect 48636 52900 48676 52940
rect 48718 52900 48758 52940
rect 48800 52900 48840 52940
rect 63592 52900 63632 52940
rect 63674 52900 63714 52940
rect 63756 52900 63796 52940
rect 63838 52900 63878 52940
rect 63920 52900 63960 52940
rect 78712 52900 78752 52940
rect 78794 52900 78834 52940
rect 78876 52900 78916 52940
rect 78958 52900 78998 52940
rect 79040 52900 79080 52940
rect 93832 52900 93872 52940
rect 93914 52900 93954 52940
rect 93996 52900 94036 52940
rect 94078 52900 94118 52940
rect 94160 52900 94200 52940
rect 19472 52144 19512 52184
rect 19554 52144 19594 52184
rect 19636 52144 19676 52184
rect 19718 52144 19758 52184
rect 19800 52144 19840 52184
rect 34592 52144 34632 52184
rect 34674 52144 34714 52184
rect 34756 52144 34796 52184
rect 34838 52144 34878 52184
rect 34920 52144 34960 52184
rect 49712 52144 49752 52184
rect 49794 52144 49834 52184
rect 49876 52144 49916 52184
rect 49958 52144 49998 52184
rect 50040 52144 50080 52184
rect 64832 52144 64872 52184
rect 64914 52144 64954 52184
rect 64996 52144 65036 52184
rect 65078 52144 65118 52184
rect 65160 52144 65200 52184
rect 79952 52144 79992 52184
rect 80034 52144 80074 52184
rect 80116 52144 80156 52184
rect 80198 52144 80238 52184
rect 80280 52144 80320 52184
rect 95072 52144 95112 52184
rect 95154 52144 95194 52184
rect 95236 52144 95276 52184
rect 95318 52144 95358 52184
rect 95400 52144 95440 52184
rect 18232 51388 18272 51428
rect 18314 51388 18354 51428
rect 18396 51388 18436 51428
rect 18478 51388 18518 51428
rect 18560 51388 18600 51428
rect 33352 51388 33392 51428
rect 33434 51388 33474 51428
rect 33516 51388 33556 51428
rect 33598 51388 33638 51428
rect 33680 51388 33720 51428
rect 48472 51388 48512 51428
rect 48554 51388 48594 51428
rect 48636 51388 48676 51428
rect 48718 51388 48758 51428
rect 48800 51388 48840 51428
rect 63592 51388 63632 51428
rect 63674 51388 63714 51428
rect 63756 51388 63796 51428
rect 63838 51388 63878 51428
rect 63920 51388 63960 51428
rect 78712 51388 78752 51428
rect 78794 51388 78834 51428
rect 78876 51388 78916 51428
rect 78958 51388 78998 51428
rect 79040 51388 79080 51428
rect 93832 51388 93872 51428
rect 93914 51388 93954 51428
rect 93996 51388 94036 51428
rect 94078 51388 94118 51428
rect 94160 51388 94200 51428
rect 19472 50632 19512 50672
rect 19554 50632 19594 50672
rect 19636 50632 19676 50672
rect 19718 50632 19758 50672
rect 19800 50632 19840 50672
rect 34592 50632 34632 50672
rect 34674 50632 34714 50672
rect 34756 50632 34796 50672
rect 34838 50632 34878 50672
rect 34920 50632 34960 50672
rect 49712 50632 49752 50672
rect 49794 50632 49834 50672
rect 49876 50632 49916 50672
rect 49958 50632 49998 50672
rect 50040 50632 50080 50672
rect 64832 50632 64872 50672
rect 64914 50632 64954 50672
rect 64996 50632 65036 50672
rect 65078 50632 65118 50672
rect 65160 50632 65200 50672
rect 79952 50632 79992 50672
rect 80034 50632 80074 50672
rect 80116 50632 80156 50672
rect 80198 50632 80238 50672
rect 80280 50632 80320 50672
rect 95072 50632 95112 50672
rect 95154 50632 95194 50672
rect 95236 50632 95276 50672
rect 95318 50632 95358 50672
rect 95400 50632 95440 50672
rect 18232 49876 18272 49916
rect 18314 49876 18354 49916
rect 18396 49876 18436 49916
rect 18478 49876 18518 49916
rect 18560 49876 18600 49916
rect 33352 49876 33392 49916
rect 33434 49876 33474 49916
rect 33516 49876 33556 49916
rect 33598 49876 33638 49916
rect 33680 49876 33720 49916
rect 48472 49876 48512 49916
rect 48554 49876 48594 49916
rect 48636 49876 48676 49916
rect 48718 49876 48758 49916
rect 48800 49876 48840 49916
rect 63592 49876 63632 49916
rect 63674 49876 63714 49916
rect 63756 49876 63796 49916
rect 63838 49876 63878 49916
rect 63920 49876 63960 49916
rect 78712 49876 78752 49916
rect 78794 49876 78834 49916
rect 78876 49876 78916 49916
rect 78958 49876 78998 49916
rect 79040 49876 79080 49916
rect 93832 49876 93872 49916
rect 93914 49876 93954 49916
rect 93996 49876 94036 49916
rect 94078 49876 94118 49916
rect 94160 49876 94200 49916
rect 19472 49120 19512 49160
rect 19554 49120 19594 49160
rect 19636 49120 19676 49160
rect 19718 49120 19758 49160
rect 19800 49120 19840 49160
rect 34592 49120 34632 49160
rect 34674 49120 34714 49160
rect 34756 49120 34796 49160
rect 34838 49120 34878 49160
rect 34920 49120 34960 49160
rect 49712 49120 49752 49160
rect 49794 49120 49834 49160
rect 49876 49120 49916 49160
rect 49958 49120 49998 49160
rect 50040 49120 50080 49160
rect 64832 49120 64872 49160
rect 64914 49120 64954 49160
rect 64996 49120 65036 49160
rect 65078 49120 65118 49160
rect 65160 49120 65200 49160
rect 79952 49120 79992 49160
rect 80034 49120 80074 49160
rect 80116 49120 80156 49160
rect 80198 49120 80238 49160
rect 80280 49120 80320 49160
rect 95072 49120 95112 49160
rect 95154 49120 95194 49160
rect 95236 49120 95276 49160
rect 95318 49120 95358 49160
rect 95400 49120 95440 49160
rect 18232 48364 18272 48404
rect 18314 48364 18354 48404
rect 18396 48364 18436 48404
rect 18478 48364 18518 48404
rect 18560 48364 18600 48404
rect 33352 48364 33392 48404
rect 33434 48364 33474 48404
rect 33516 48364 33556 48404
rect 33598 48364 33638 48404
rect 33680 48364 33720 48404
rect 48472 48364 48512 48404
rect 48554 48364 48594 48404
rect 48636 48364 48676 48404
rect 48718 48364 48758 48404
rect 48800 48364 48840 48404
rect 63592 48364 63632 48404
rect 63674 48364 63714 48404
rect 63756 48364 63796 48404
rect 63838 48364 63878 48404
rect 63920 48364 63960 48404
rect 78712 48364 78752 48404
rect 78794 48364 78834 48404
rect 78876 48364 78916 48404
rect 78958 48364 78998 48404
rect 79040 48364 79080 48404
rect 93832 48364 93872 48404
rect 93914 48364 93954 48404
rect 93996 48364 94036 48404
rect 94078 48364 94118 48404
rect 94160 48364 94200 48404
rect 19472 47608 19512 47648
rect 19554 47608 19594 47648
rect 19636 47608 19676 47648
rect 19718 47608 19758 47648
rect 19800 47608 19840 47648
rect 34592 47608 34632 47648
rect 34674 47608 34714 47648
rect 34756 47608 34796 47648
rect 34838 47608 34878 47648
rect 34920 47608 34960 47648
rect 49712 47608 49752 47648
rect 49794 47608 49834 47648
rect 49876 47608 49916 47648
rect 49958 47608 49998 47648
rect 50040 47608 50080 47648
rect 64832 47608 64872 47648
rect 64914 47608 64954 47648
rect 64996 47608 65036 47648
rect 65078 47608 65118 47648
rect 65160 47608 65200 47648
rect 79952 47608 79992 47648
rect 80034 47608 80074 47648
rect 80116 47608 80156 47648
rect 80198 47608 80238 47648
rect 80280 47608 80320 47648
rect 95072 47608 95112 47648
rect 95154 47608 95194 47648
rect 95236 47608 95276 47648
rect 95318 47608 95358 47648
rect 95400 47608 95440 47648
rect 14284 47272 14324 47312
rect 14380 46432 14420 46472
rect 14092 44752 14132 44792
rect 7084 16276 7124 16316
rect 6700 10228 6740 10268
rect 5644 8716 5684 8756
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 14572 47272 14612 47312
rect 18232 46852 18272 46892
rect 18314 46852 18354 46892
rect 18396 46852 18436 46892
rect 18478 46852 18518 46892
rect 18560 46852 18600 46892
rect 33352 46852 33392 46892
rect 33434 46852 33474 46892
rect 33516 46852 33556 46892
rect 33598 46852 33638 46892
rect 33680 46852 33720 46892
rect 48472 46852 48512 46892
rect 48554 46852 48594 46892
rect 48636 46852 48676 46892
rect 48718 46852 48758 46892
rect 48800 46852 48840 46892
rect 63592 46852 63632 46892
rect 63674 46852 63714 46892
rect 63756 46852 63796 46892
rect 63838 46852 63878 46892
rect 63920 46852 63960 46892
rect 78712 46852 78752 46892
rect 78794 46852 78834 46892
rect 78876 46852 78916 46892
rect 78958 46852 78998 46892
rect 79040 46852 79080 46892
rect 93832 46852 93872 46892
rect 93914 46852 93954 46892
rect 93996 46852 94036 46892
rect 94078 46852 94118 46892
rect 94160 46852 94200 46892
rect 14956 46432 14996 46472
rect 19472 46096 19512 46136
rect 19554 46096 19594 46136
rect 19636 46096 19676 46136
rect 19718 46096 19758 46136
rect 19800 46096 19840 46136
rect 34592 46096 34632 46136
rect 34674 46096 34714 46136
rect 34756 46096 34796 46136
rect 34838 46096 34878 46136
rect 34920 46096 34960 46136
rect 49712 46096 49752 46136
rect 49794 46096 49834 46136
rect 49876 46096 49916 46136
rect 49958 46096 49998 46136
rect 50040 46096 50080 46136
rect 64832 46096 64872 46136
rect 64914 46096 64954 46136
rect 64996 46096 65036 46136
rect 65078 46096 65118 46136
rect 65160 46096 65200 46136
rect 79952 46096 79992 46136
rect 80034 46096 80074 46136
rect 80116 46096 80156 46136
rect 80198 46096 80238 46136
rect 80280 46096 80320 46136
rect 95072 46096 95112 46136
rect 95154 46096 95194 46136
rect 95236 46096 95276 46136
rect 95318 46096 95358 46136
rect 95400 46096 95440 46136
rect 14572 45928 14612 45968
rect 18232 45340 18272 45380
rect 18314 45340 18354 45380
rect 18396 45340 18436 45380
rect 18478 45340 18518 45380
rect 18560 45340 18600 45380
rect 33352 45340 33392 45380
rect 33434 45340 33474 45380
rect 33516 45340 33556 45380
rect 33598 45340 33638 45380
rect 33680 45340 33720 45380
rect 48472 45340 48512 45380
rect 48554 45340 48594 45380
rect 48636 45340 48676 45380
rect 48718 45340 48758 45380
rect 48800 45340 48840 45380
rect 63592 45340 63632 45380
rect 63674 45340 63714 45380
rect 63756 45340 63796 45380
rect 63838 45340 63878 45380
rect 63920 45340 63960 45380
rect 78712 45340 78752 45380
rect 78794 45340 78834 45380
rect 78876 45340 78916 45380
rect 78958 45340 78998 45380
rect 79040 45340 79080 45380
rect 93832 45340 93872 45380
rect 93914 45340 93954 45380
rect 93996 45340 94036 45380
rect 94078 45340 94118 45380
rect 94160 45340 94200 45380
rect 19472 44584 19512 44624
rect 19554 44584 19594 44624
rect 19636 44584 19676 44624
rect 19718 44584 19758 44624
rect 19800 44584 19840 44624
rect 34592 44584 34632 44624
rect 34674 44584 34714 44624
rect 34756 44584 34796 44624
rect 34838 44584 34878 44624
rect 34920 44584 34960 44624
rect 49712 44584 49752 44624
rect 49794 44584 49834 44624
rect 49876 44584 49916 44624
rect 49958 44584 49998 44624
rect 50040 44584 50080 44624
rect 64832 44584 64872 44624
rect 64914 44584 64954 44624
rect 64996 44584 65036 44624
rect 65078 44584 65118 44624
rect 65160 44584 65200 44624
rect 79952 44584 79992 44624
rect 80034 44584 80074 44624
rect 80116 44584 80156 44624
rect 80198 44584 80238 44624
rect 80280 44584 80320 44624
rect 95072 44584 95112 44624
rect 95154 44584 95194 44624
rect 95236 44584 95276 44624
rect 95318 44584 95358 44624
rect 95400 44584 95440 44624
rect 18232 43828 18272 43868
rect 18314 43828 18354 43868
rect 18396 43828 18436 43868
rect 18478 43828 18518 43868
rect 18560 43828 18600 43868
rect 33352 43828 33392 43868
rect 33434 43828 33474 43868
rect 33516 43828 33556 43868
rect 33598 43828 33638 43868
rect 33680 43828 33720 43868
rect 48472 43828 48512 43868
rect 48554 43828 48594 43868
rect 48636 43828 48676 43868
rect 48718 43828 48758 43868
rect 48800 43828 48840 43868
rect 63592 43828 63632 43868
rect 63674 43828 63714 43868
rect 63756 43828 63796 43868
rect 63838 43828 63878 43868
rect 63920 43828 63960 43868
rect 78712 43828 78752 43868
rect 78794 43828 78834 43868
rect 78876 43828 78916 43868
rect 78958 43828 78998 43868
rect 79040 43828 79080 43868
rect 93832 43828 93872 43868
rect 93914 43828 93954 43868
rect 93996 43828 94036 43868
rect 94078 43828 94118 43868
rect 94160 43828 94200 43868
rect 19472 43072 19512 43112
rect 19554 43072 19594 43112
rect 19636 43072 19676 43112
rect 19718 43072 19758 43112
rect 19800 43072 19840 43112
rect 34592 43072 34632 43112
rect 34674 43072 34714 43112
rect 34756 43072 34796 43112
rect 34838 43072 34878 43112
rect 34920 43072 34960 43112
rect 49712 43072 49752 43112
rect 49794 43072 49834 43112
rect 49876 43072 49916 43112
rect 49958 43072 49998 43112
rect 50040 43072 50080 43112
rect 64832 43072 64872 43112
rect 64914 43072 64954 43112
rect 64996 43072 65036 43112
rect 65078 43072 65118 43112
rect 65160 43072 65200 43112
rect 79952 43072 79992 43112
rect 80034 43072 80074 43112
rect 80116 43072 80156 43112
rect 80198 43072 80238 43112
rect 80280 43072 80320 43112
rect 95072 43072 95112 43112
rect 95154 43072 95194 43112
rect 95236 43072 95276 43112
rect 95318 43072 95358 43112
rect 95400 43072 95440 43112
rect 18232 42316 18272 42356
rect 18314 42316 18354 42356
rect 18396 42316 18436 42356
rect 18478 42316 18518 42356
rect 18560 42316 18600 42356
rect 33352 42316 33392 42356
rect 33434 42316 33474 42356
rect 33516 42316 33556 42356
rect 33598 42316 33638 42356
rect 33680 42316 33720 42356
rect 48472 42316 48512 42356
rect 48554 42316 48594 42356
rect 48636 42316 48676 42356
rect 48718 42316 48758 42356
rect 48800 42316 48840 42356
rect 63592 42316 63632 42356
rect 63674 42316 63714 42356
rect 63756 42316 63796 42356
rect 63838 42316 63878 42356
rect 63920 42316 63960 42356
rect 78712 42316 78752 42356
rect 78794 42316 78834 42356
rect 78876 42316 78916 42356
rect 78958 42316 78998 42356
rect 79040 42316 79080 42356
rect 93832 42316 93872 42356
rect 93914 42316 93954 42356
rect 93996 42316 94036 42356
rect 94078 42316 94118 42356
rect 94160 42316 94200 42356
rect 19472 41560 19512 41600
rect 19554 41560 19594 41600
rect 19636 41560 19676 41600
rect 19718 41560 19758 41600
rect 19800 41560 19840 41600
rect 34592 41560 34632 41600
rect 34674 41560 34714 41600
rect 34756 41560 34796 41600
rect 34838 41560 34878 41600
rect 34920 41560 34960 41600
rect 49712 41560 49752 41600
rect 49794 41560 49834 41600
rect 49876 41560 49916 41600
rect 49958 41560 49998 41600
rect 50040 41560 50080 41600
rect 64832 41560 64872 41600
rect 64914 41560 64954 41600
rect 64996 41560 65036 41600
rect 65078 41560 65118 41600
rect 65160 41560 65200 41600
rect 79952 41560 79992 41600
rect 80034 41560 80074 41600
rect 80116 41560 80156 41600
rect 80198 41560 80238 41600
rect 80280 41560 80320 41600
rect 95072 41560 95112 41600
rect 95154 41560 95194 41600
rect 95236 41560 95276 41600
rect 95318 41560 95358 41600
rect 95400 41560 95440 41600
rect 18232 40804 18272 40844
rect 18314 40804 18354 40844
rect 18396 40804 18436 40844
rect 18478 40804 18518 40844
rect 18560 40804 18600 40844
rect 33352 40804 33392 40844
rect 33434 40804 33474 40844
rect 33516 40804 33556 40844
rect 33598 40804 33638 40844
rect 33680 40804 33720 40844
rect 48472 40804 48512 40844
rect 48554 40804 48594 40844
rect 48636 40804 48676 40844
rect 48718 40804 48758 40844
rect 48800 40804 48840 40844
rect 63592 40804 63632 40844
rect 63674 40804 63714 40844
rect 63756 40804 63796 40844
rect 63838 40804 63878 40844
rect 63920 40804 63960 40844
rect 78712 40804 78752 40844
rect 78794 40804 78834 40844
rect 78876 40804 78916 40844
rect 78958 40804 78998 40844
rect 79040 40804 79080 40844
rect 93832 40804 93872 40844
rect 93914 40804 93954 40844
rect 93996 40804 94036 40844
rect 94078 40804 94118 40844
rect 94160 40804 94200 40844
rect 19472 40048 19512 40088
rect 19554 40048 19594 40088
rect 19636 40048 19676 40088
rect 19718 40048 19758 40088
rect 19800 40048 19840 40088
rect 34592 40048 34632 40088
rect 34674 40048 34714 40088
rect 34756 40048 34796 40088
rect 34838 40048 34878 40088
rect 34920 40048 34960 40088
rect 49712 40048 49752 40088
rect 49794 40048 49834 40088
rect 49876 40048 49916 40088
rect 49958 40048 49998 40088
rect 50040 40048 50080 40088
rect 64832 40048 64872 40088
rect 64914 40048 64954 40088
rect 64996 40048 65036 40088
rect 65078 40048 65118 40088
rect 65160 40048 65200 40088
rect 79952 40048 79992 40088
rect 80034 40048 80074 40088
rect 80116 40048 80156 40088
rect 80198 40048 80238 40088
rect 80280 40048 80320 40088
rect 95072 40048 95112 40088
rect 95154 40048 95194 40088
rect 95236 40048 95276 40088
rect 95318 40048 95358 40088
rect 95400 40048 95440 40088
rect 18232 39292 18272 39332
rect 18314 39292 18354 39332
rect 18396 39292 18436 39332
rect 18478 39292 18518 39332
rect 18560 39292 18600 39332
rect 33352 39292 33392 39332
rect 33434 39292 33474 39332
rect 33516 39292 33556 39332
rect 33598 39292 33638 39332
rect 33680 39292 33720 39332
rect 48472 39292 48512 39332
rect 48554 39292 48594 39332
rect 48636 39292 48676 39332
rect 48718 39292 48758 39332
rect 48800 39292 48840 39332
rect 63592 39292 63632 39332
rect 63674 39292 63714 39332
rect 63756 39292 63796 39332
rect 63838 39292 63878 39332
rect 63920 39292 63960 39332
rect 78712 39292 78752 39332
rect 78794 39292 78834 39332
rect 78876 39292 78916 39332
rect 78958 39292 78998 39332
rect 79040 39292 79080 39332
rect 93832 39292 93872 39332
rect 93914 39292 93954 39332
rect 93996 39292 94036 39332
rect 94078 39292 94118 39332
rect 94160 39292 94200 39332
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 95072 38536 95112 38576
rect 95154 38536 95194 38576
rect 95236 38536 95276 38576
rect 95318 38536 95358 38576
rect 95400 38536 95440 38576
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 93832 37780 93872 37820
rect 93914 37780 93954 37820
rect 93996 37780 94036 37820
rect 94078 37780 94118 37820
rect 94160 37780 94200 37820
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 95072 37024 95112 37064
rect 95154 37024 95194 37064
rect 95236 37024 95276 37064
rect 95318 37024 95358 37064
rect 95400 37024 95440 37064
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 93832 36268 93872 36308
rect 93914 36268 93954 36308
rect 93996 36268 94036 36308
rect 94078 36268 94118 36308
rect 94160 36268 94200 36308
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 95072 35512 95112 35552
rect 95154 35512 95194 35552
rect 95236 35512 95276 35552
rect 95318 35512 95358 35552
rect 95400 35512 95440 35552
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 93832 34756 93872 34796
rect 93914 34756 93954 34796
rect 93996 34756 94036 34796
rect 94078 34756 94118 34796
rect 94160 34756 94200 34796
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 95072 34000 95112 34040
rect 95154 34000 95194 34040
rect 95236 34000 95276 34040
rect 95318 34000 95358 34040
rect 95400 34000 95440 34040
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 93832 33244 93872 33284
rect 93914 33244 93954 33284
rect 93996 33244 94036 33284
rect 94078 33244 94118 33284
rect 94160 33244 94200 33284
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 95072 32488 95112 32528
rect 95154 32488 95194 32528
rect 95236 32488 95276 32528
rect 95318 32488 95358 32528
rect 95400 32488 95440 32528
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 93832 31732 93872 31772
rect 93914 31732 93954 31772
rect 93996 31732 94036 31772
rect 94078 31732 94118 31772
rect 94160 31732 94200 31772
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 95072 30976 95112 31016
rect 95154 30976 95194 31016
rect 95236 30976 95276 31016
rect 95318 30976 95358 31016
rect 95400 30976 95440 31016
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 93832 30220 93872 30260
rect 93914 30220 93954 30260
rect 93996 30220 94036 30260
rect 94078 30220 94118 30260
rect 94160 30220 94200 30260
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 95072 29464 95112 29504
rect 95154 29464 95194 29504
rect 95236 29464 95276 29504
rect 95318 29464 95358 29504
rect 95400 29464 95440 29504
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 93832 28708 93872 28748
rect 93914 28708 93954 28748
rect 93996 28708 94036 28748
rect 94078 28708 94118 28748
rect 94160 28708 94200 28748
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 95072 27952 95112 27992
rect 95154 27952 95194 27992
rect 95236 27952 95276 27992
rect 95318 27952 95358 27992
rect 95400 27952 95440 27992
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 93832 27196 93872 27236
rect 93914 27196 93954 27236
rect 93996 27196 94036 27236
rect 94078 27196 94118 27236
rect 94160 27196 94200 27236
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 95072 26440 95112 26480
rect 95154 26440 95194 26480
rect 95236 26440 95276 26480
rect 95318 26440 95358 26480
rect 95400 26440 95440 26480
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 93832 25684 93872 25724
rect 93914 25684 93954 25724
rect 93996 25684 94036 25724
rect 94078 25684 94118 25724
rect 94160 25684 94200 25724
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 95072 24928 95112 24968
rect 95154 24928 95194 24968
rect 95236 24928 95276 24968
rect 95318 24928 95358 24968
rect 95400 24928 95440 24968
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 63592 24172 63632 24212
rect 63674 24172 63714 24212
rect 63756 24172 63796 24212
rect 63838 24172 63878 24212
rect 63920 24172 63960 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 93832 24172 93872 24212
rect 93914 24172 93954 24212
rect 93996 24172 94036 24212
rect 94078 24172 94118 24212
rect 94160 24172 94200 24212
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 64832 23416 64872 23456
rect 64914 23416 64954 23456
rect 64996 23416 65036 23456
rect 65078 23416 65118 23456
rect 65160 23416 65200 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 95072 23416 95112 23456
rect 95154 23416 95194 23456
rect 95236 23416 95276 23456
rect 95318 23416 95358 23456
rect 95400 23416 95440 23456
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 63592 22660 63632 22700
rect 63674 22660 63714 22700
rect 63756 22660 63796 22700
rect 63838 22660 63878 22700
rect 63920 22660 63960 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 93832 22660 93872 22700
rect 93914 22660 93954 22700
rect 93996 22660 94036 22700
rect 94078 22660 94118 22700
rect 94160 22660 94200 22700
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 64832 21904 64872 21944
rect 64914 21904 64954 21944
rect 64996 21904 65036 21944
rect 65078 21904 65118 21944
rect 65160 21904 65200 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 63592 21148 63632 21188
rect 63674 21148 63714 21188
rect 63756 21148 63796 21188
rect 63838 21148 63878 21188
rect 63920 21148 63960 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 64832 20392 64872 20432
rect 64914 20392 64954 20432
rect 64996 20392 65036 20432
rect 65078 20392 65118 20432
rect 65160 20392 65200 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 63592 19636 63632 19676
rect 63674 19636 63714 19676
rect 63756 19636 63796 19676
rect 63838 19636 63878 19676
rect 63920 19636 63960 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 64832 18880 64872 18920
rect 64914 18880 64954 18920
rect 64996 18880 65036 18920
rect 65078 18880 65118 18920
rect 65160 18880 65200 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 95072 18880 95112 18920
rect 95154 18880 95194 18920
rect 95236 18880 95276 18920
rect 95318 18880 95358 18920
rect 95400 18880 95440 18920
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 63592 18124 63632 18164
rect 63674 18124 63714 18164
rect 63756 18124 63796 18164
rect 63838 18124 63878 18164
rect 63920 18124 63960 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 93832 18124 93872 18164
rect 93914 18124 93954 18164
rect 93996 18124 94036 18164
rect 94078 18124 94118 18164
rect 94160 18124 94200 18164
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 64832 17368 64872 17408
rect 64914 17368 64954 17408
rect 64996 17368 65036 17408
rect 65078 17368 65118 17408
rect 65160 17368 65200 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 95072 17368 95112 17408
rect 95154 17368 95194 17408
rect 95236 17368 95276 17408
rect 95318 17368 95358 17408
rect 95400 17368 95440 17408
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 63592 16612 63632 16652
rect 63674 16612 63714 16652
rect 63756 16612 63796 16652
rect 63838 16612 63878 16652
rect 63920 16612 63960 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 93832 16612 93872 16652
rect 93914 16612 93954 16652
rect 93996 16612 94036 16652
rect 94078 16612 94118 16652
rect 94160 16612 94200 16652
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 64832 15856 64872 15896
rect 64914 15856 64954 15896
rect 64996 15856 65036 15896
rect 65078 15856 65118 15896
rect 65160 15856 65200 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 95072 15856 95112 15896
rect 95154 15856 95194 15896
rect 95236 15856 95276 15896
rect 95318 15856 95358 15896
rect 95400 15856 95440 15896
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 93832 15100 93872 15140
rect 93914 15100 93954 15140
rect 93996 15100 94036 15140
rect 94078 15100 94118 15140
rect 94160 15100 94200 15140
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 95072 14344 95112 14384
rect 95154 14344 95194 14384
rect 95236 14344 95276 14384
rect 95318 14344 95358 14384
rect 95400 14344 95440 14384
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 93832 13588 93872 13628
rect 93914 13588 93954 13628
rect 93996 13588 94036 13628
rect 94078 13588 94118 13628
rect 94160 13588 94200 13628
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 95072 12832 95112 12872
rect 95154 12832 95194 12872
rect 95236 12832 95276 12872
rect 95318 12832 95358 12872
rect 95400 12832 95440 12872
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 93832 12076 93872 12116
rect 93914 12076 93954 12116
rect 93996 12076 94036 12116
rect 94078 12076 94118 12116
rect 94160 12076 94200 12116
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 95072 11320 95112 11360
rect 95154 11320 95194 11360
rect 95236 11320 95276 11360
rect 95318 11320 95358 11360
rect 95400 11320 95440 11360
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 93832 10564 93872 10604
rect 93914 10564 93954 10604
rect 93996 10564 94036 10604
rect 94078 10564 94118 10604
rect 94160 10564 94200 10604
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 95072 9808 95112 9848
rect 95154 9808 95194 9848
rect 95236 9808 95276 9848
rect 95318 9808 95358 9848
rect 95400 9808 95440 9848
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 93832 9052 93872 9092
rect 93914 9052 93954 9092
rect 93996 9052 94036 9092
rect 94078 9052 94118 9092
rect 94160 9052 94200 9092
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 95072 8296 95112 8336
rect 95154 8296 95194 8336
rect 95236 8296 95276 8336
rect 95318 8296 95358 8336
rect 95400 8296 95440 8336
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 93832 7540 93872 7580
rect 93914 7540 93954 7580
rect 93996 7540 94036 7580
rect 94078 7540 94118 7580
rect 94160 7540 94200 7580
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 95072 6784 95112 6824
rect 95154 6784 95194 6824
rect 95236 6784 95276 6824
rect 95318 6784 95358 6824
rect 95400 6784 95440 6824
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 93832 6028 93872 6068
rect 93914 6028 93954 6068
rect 93996 6028 94036 6068
rect 94078 6028 94118 6068
rect 94160 6028 94200 6068
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 95072 5272 95112 5312
rect 95154 5272 95194 5312
rect 95236 5272 95276 5312
rect 95318 5272 95358 5312
rect 95400 5272 95440 5312
rect 14476 4852 14516 4892
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 93832 4516 93872 4556
rect 93914 4516 93954 4556
rect 93996 4516 94036 4556
rect 94078 4516 94118 4556
rect 94160 4516 94200 4556
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 95072 3760 95112 3800
rect 95154 3760 95194 3800
rect 95236 3760 95276 3800
rect 95318 3760 95358 3800
rect 95400 3760 95440 3800
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 93832 3004 93872 3044
rect 93914 3004 93954 3044
rect 93996 3004 94036 3044
rect 94078 3004 94118 3044
rect 94160 3004 94200 3044
rect 652 2584 692 2624
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 95072 2248 95112 2288
rect 95154 2248 95194 2288
rect 95236 2248 95276 2288
rect 95318 2248 95358 2288
rect 95400 2248 95440 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 93832 1492 93872 1532
rect 93914 1492 93954 1532
rect 93996 1492 94036 1532
rect 94078 1492 94118 1532
rect 94160 1492 94200 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
rect 95072 736 95112 776
rect 95154 736 95194 776
rect 95236 736 95276 776
rect 95318 736 95358 776
rect 95400 736 95440 776
<< metal3 >>
rect 3103 81628 3112 81668
rect 3152 81628 3194 81668
rect 3234 81628 3276 81668
rect 3316 81628 3358 81668
rect 3398 81628 3440 81668
rect 3480 81628 3489 81668
rect 18223 81628 18232 81668
rect 18272 81628 18314 81668
rect 18354 81628 18396 81668
rect 18436 81628 18478 81668
rect 18518 81628 18560 81668
rect 18600 81628 18609 81668
rect 33343 81628 33352 81668
rect 33392 81628 33434 81668
rect 33474 81628 33516 81668
rect 33556 81628 33598 81668
rect 33638 81628 33680 81668
rect 33720 81628 33729 81668
rect 48463 81628 48472 81668
rect 48512 81628 48554 81668
rect 48594 81628 48636 81668
rect 48676 81628 48718 81668
rect 48758 81628 48800 81668
rect 48840 81628 48849 81668
rect 63583 81628 63592 81668
rect 63632 81628 63674 81668
rect 63714 81628 63756 81668
rect 63796 81628 63838 81668
rect 63878 81628 63920 81668
rect 63960 81628 63969 81668
rect 78703 81628 78712 81668
rect 78752 81628 78794 81668
rect 78834 81628 78876 81668
rect 78916 81628 78958 81668
rect 78998 81628 79040 81668
rect 79080 81628 79089 81668
rect 93823 81628 93832 81668
rect 93872 81628 93914 81668
rect 93954 81628 93996 81668
rect 94036 81628 94078 81668
rect 94118 81628 94160 81668
rect 94200 81628 94209 81668
rect 4343 80872 4352 80912
rect 4392 80872 4434 80912
rect 4474 80872 4516 80912
rect 4556 80872 4598 80912
rect 4638 80872 4680 80912
rect 4720 80872 4729 80912
rect 19463 80872 19472 80912
rect 19512 80872 19554 80912
rect 19594 80872 19636 80912
rect 19676 80872 19718 80912
rect 19758 80872 19800 80912
rect 19840 80872 19849 80912
rect 34583 80872 34592 80912
rect 34632 80872 34674 80912
rect 34714 80872 34756 80912
rect 34796 80872 34838 80912
rect 34878 80872 34920 80912
rect 34960 80872 34969 80912
rect 49703 80872 49712 80912
rect 49752 80872 49794 80912
rect 49834 80872 49876 80912
rect 49916 80872 49958 80912
rect 49998 80872 50040 80912
rect 50080 80872 50089 80912
rect 64823 80872 64832 80912
rect 64872 80872 64914 80912
rect 64954 80872 64996 80912
rect 65036 80872 65078 80912
rect 65118 80872 65160 80912
rect 65200 80872 65209 80912
rect 79943 80872 79952 80912
rect 79992 80872 80034 80912
rect 80074 80872 80116 80912
rect 80156 80872 80198 80912
rect 80238 80872 80280 80912
rect 80320 80872 80329 80912
rect 95063 80872 95072 80912
rect 95112 80872 95154 80912
rect 95194 80872 95236 80912
rect 95276 80872 95318 80912
rect 95358 80872 95400 80912
rect 95440 80872 95449 80912
rect 0 80180 80 80260
rect 3103 80116 3112 80156
rect 3152 80116 3194 80156
rect 3234 80116 3276 80156
rect 3316 80116 3358 80156
rect 3398 80116 3440 80156
rect 3480 80116 3489 80156
rect 18223 80116 18232 80156
rect 18272 80116 18314 80156
rect 18354 80116 18396 80156
rect 18436 80116 18478 80156
rect 18518 80116 18560 80156
rect 18600 80116 18609 80156
rect 33343 80116 33352 80156
rect 33392 80116 33434 80156
rect 33474 80116 33516 80156
rect 33556 80116 33598 80156
rect 33638 80116 33680 80156
rect 33720 80116 33729 80156
rect 48463 80116 48472 80156
rect 48512 80116 48554 80156
rect 48594 80116 48636 80156
rect 48676 80116 48718 80156
rect 48758 80116 48800 80156
rect 48840 80116 48849 80156
rect 63583 80116 63592 80156
rect 63632 80116 63674 80156
rect 63714 80116 63756 80156
rect 63796 80116 63838 80156
rect 63878 80116 63920 80156
rect 63960 80116 63969 80156
rect 78703 80116 78712 80156
rect 78752 80116 78794 80156
rect 78834 80116 78876 80156
rect 78916 80116 78958 80156
rect 78998 80116 79040 80156
rect 79080 80116 79089 80156
rect 93823 80116 93832 80156
rect 93872 80116 93914 80156
rect 93954 80116 93996 80156
rect 94036 80116 94078 80156
rect 94118 80116 94160 80156
rect 94200 80116 94209 80156
rect 4343 79360 4352 79400
rect 4392 79360 4434 79400
rect 4474 79360 4516 79400
rect 4556 79360 4598 79400
rect 4638 79360 4680 79400
rect 4720 79360 4729 79400
rect 19463 79360 19472 79400
rect 19512 79360 19554 79400
rect 19594 79360 19636 79400
rect 19676 79360 19718 79400
rect 19758 79360 19800 79400
rect 19840 79360 19849 79400
rect 34583 79360 34592 79400
rect 34632 79360 34674 79400
rect 34714 79360 34756 79400
rect 34796 79360 34838 79400
rect 34878 79360 34920 79400
rect 34960 79360 34969 79400
rect 49703 79360 49712 79400
rect 49752 79360 49794 79400
rect 49834 79360 49876 79400
rect 49916 79360 49958 79400
rect 49998 79360 50040 79400
rect 50080 79360 50089 79400
rect 64823 79360 64832 79400
rect 64872 79360 64914 79400
rect 64954 79360 64996 79400
rect 65036 79360 65078 79400
rect 65118 79360 65160 79400
rect 65200 79360 65209 79400
rect 79943 79360 79952 79400
rect 79992 79360 80034 79400
rect 80074 79360 80116 79400
rect 80156 79360 80198 79400
rect 80238 79360 80280 79400
rect 80320 79360 80329 79400
rect 95063 79360 95072 79400
rect 95112 79360 95154 79400
rect 95194 79360 95236 79400
rect 95276 79360 95318 79400
rect 95358 79360 95400 79400
rect 95440 79360 95449 79400
rect 3103 78604 3112 78644
rect 3152 78604 3194 78644
rect 3234 78604 3276 78644
rect 3316 78604 3358 78644
rect 3398 78604 3440 78644
rect 3480 78604 3489 78644
rect 18223 78604 18232 78644
rect 18272 78604 18314 78644
rect 18354 78604 18396 78644
rect 18436 78604 18478 78644
rect 18518 78604 18560 78644
rect 18600 78604 18609 78644
rect 33343 78604 33352 78644
rect 33392 78604 33434 78644
rect 33474 78604 33516 78644
rect 33556 78604 33598 78644
rect 33638 78604 33680 78644
rect 33720 78604 33729 78644
rect 48463 78604 48472 78644
rect 48512 78604 48554 78644
rect 48594 78604 48636 78644
rect 48676 78604 48718 78644
rect 48758 78604 48800 78644
rect 48840 78604 48849 78644
rect 63583 78604 63592 78644
rect 63632 78604 63674 78644
rect 63714 78604 63756 78644
rect 63796 78604 63838 78644
rect 63878 78604 63920 78644
rect 63960 78604 63969 78644
rect 78703 78604 78712 78644
rect 78752 78604 78794 78644
rect 78834 78604 78876 78644
rect 78916 78604 78958 78644
rect 78998 78604 79040 78644
rect 79080 78604 79089 78644
rect 93823 78604 93832 78644
rect 93872 78604 93914 78644
rect 93954 78604 93996 78644
rect 94036 78604 94078 78644
rect 94118 78604 94160 78644
rect 94200 78604 94209 78644
rect 0 78332 80 78412
rect 4343 77848 4352 77888
rect 4392 77848 4434 77888
rect 4474 77848 4516 77888
rect 4556 77848 4598 77888
rect 4638 77848 4680 77888
rect 4720 77848 4729 77888
rect 19463 77848 19472 77888
rect 19512 77848 19554 77888
rect 19594 77848 19636 77888
rect 19676 77848 19718 77888
rect 19758 77848 19800 77888
rect 19840 77848 19849 77888
rect 34583 77848 34592 77888
rect 34632 77848 34674 77888
rect 34714 77848 34756 77888
rect 34796 77848 34838 77888
rect 34878 77848 34920 77888
rect 34960 77848 34969 77888
rect 49703 77848 49712 77888
rect 49752 77848 49794 77888
rect 49834 77848 49876 77888
rect 49916 77848 49958 77888
rect 49998 77848 50040 77888
rect 50080 77848 50089 77888
rect 64823 77848 64832 77888
rect 64872 77848 64914 77888
rect 64954 77848 64996 77888
rect 65036 77848 65078 77888
rect 65118 77848 65160 77888
rect 65200 77848 65209 77888
rect 79943 77848 79952 77888
rect 79992 77848 80034 77888
rect 80074 77848 80116 77888
rect 80156 77848 80198 77888
rect 80238 77848 80280 77888
rect 80320 77848 80329 77888
rect 95063 77848 95072 77888
rect 95112 77848 95154 77888
rect 95194 77848 95236 77888
rect 95276 77848 95318 77888
rect 95358 77848 95400 77888
rect 95440 77848 95449 77888
rect 3103 77092 3112 77132
rect 3152 77092 3194 77132
rect 3234 77092 3276 77132
rect 3316 77092 3358 77132
rect 3398 77092 3440 77132
rect 3480 77092 3489 77132
rect 18223 77092 18232 77132
rect 18272 77092 18314 77132
rect 18354 77092 18396 77132
rect 18436 77092 18478 77132
rect 18518 77092 18560 77132
rect 18600 77092 18609 77132
rect 33343 77092 33352 77132
rect 33392 77092 33434 77132
rect 33474 77092 33516 77132
rect 33556 77092 33598 77132
rect 33638 77092 33680 77132
rect 33720 77092 33729 77132
rect 48463 77092 48472 77132
rect 48512 77092 48554 77132
rect 48594 77092 48636 77132
rect 48676 77092 48718 77132
rect 48758 77092 48800 77132
rect 48840 77092 48849 77132
rect 63583 77092 63592 77132
rect 63632 77092 63674 77132
rect 63714 77092 63756 77132
rect 63796 77092 63838 77132
rect 63878 77092 63920 77132
rect 63960 77092 63969 77132
rect 78703 77092 78712 77132
rect 78752 77092 78794 77132
rect 78834 77092 78876 77132
rect 78916 77092 78958 77132
rect 78998 77092 79040 77132
rect 79080 77092 79089 77132
rect 93823 77092 93832 77132
rect 93872 77092 93914 77132
rect 93954 77092 93996 77132
rect 94036 77092 94078 77132
rect 94118 77092 94160 77132
rect 94200 77092 94209 77132
rect 0 76484 80 76564
rect 4343 76336 4352 76376
rect 4392 76336 4434 76376
rect 4474 76336 4516 76376
rect 4556 76336 4598 76376
rect 4638 76336 4680 76376
rect 4720 76336 4729 76376
rect 19463 76336 19472 76376
rect 19512 76336 19554 76376
rect 19594 76336 19636 76376
rect 19676 76336 19718 76376
rect 19758 76336 19800 76376
rect 19840 76336 19849 76376
rect 34583 76336 34592 76376
rect 34632 76336 34674 76376
rect 34714 76336 34756 76376
rect 34796 76336 34838 76376
rect 34878 76336 34920 76376
rect 34960 76336 34969 76376
rect 49703 76336 49712 76376
rect 49752 76336 49794 76376
rect 49834 76336 49876 76376
rect 49916 76336 49958 76376
rect 49998 76336 50040 76376
rect 50080 76336 50089 76376
rect 64823 76336 64832 76376
rect 64872 76336 64914 76376
rect 64954 76336 64996 76376
rect 65036 76336 65078 76376
rect 65118 76336 65160 76376
rect 65200 76336 65209 76376
rect 79943 76336 79952 76376
rect 79992 76336 80034 76376
rect 80074 76336 80116 76376
rect 80156 76336 80198 76376
rect 80238 76336 80280 76376
rect 80320 76336 80329 76376
rect 95063 76336 95072 76376
rect 95112 76336 95154 76376
rect 95194 76336 95236 76376
rect 95276 76336 95318 76376
rect 95358 76336 95400 76376
rect 95440 76336 95449 76376
rect 3103 75580 3112 75620
rect 3152 75580 3194 75620
rect 3234 75580 3276 75620
rect 3316 75580 3358 75620
rect 3398 75580 3440 75620
rect 3480 75580 3489 75620
rect 18223 75580 18232 75620
rect 18272 75580 18314 75620
rect 18354 75580 18396 75620
rect 18436 75580 18478 75620
rect 18518 75580 18560 75620
rect 18600 75580 18609 75620
rect 33343 75580 33352 75620
rect 33392 75580 33434 75620
rect 33474 75580 33516 75620
rect 33556 75580 33598 75620
rect 33638 75580 33680 75620
rect 33720 75580 33729 75620
rect 48463 75580 48472 75620
rect 48512 75580 48554 75620
rect 48594 75580 48636 75620
rect 48676 75580 48718 75620
rect 48758 75580 48800 75620
rect 48840 75580 48849 75620
rect 63583 75580 63592 75620
rect 63632 75580 63674 75620
rect 63714 75580 63756 75620
rect 63796 75580 63838 75620
rect 63878 75580 63920 75620
rect 63960 75580 63969 75620
rect 78703 75580 78712 75620
rect 78752 75580 78794 75620
rect 78834 75580 78876 75620
rect 78916 75580 78958 75620
rect 78998 75580 79040 75620
rect 79080 75580 79089 75620
rect 93823 75580 93832 75620
rect 93872 75580 93914 75620
rect 93954 75580 93996 75620
rect 94036 75580 94078 75620
rect 94118 75580 94160 75620
rect 94200 75580 94209 75620
rect 4343 74824 4352 74864
rect 4392 74824 4434 74864
rect 4474 74824 4516 74864
rect 4556 74824 4598 74864
rect 4638 74824 4680 74864
rect 4720 74824 4729 74864
rect 19463 74824 19472 74864
rect 19512 74824 19554 74864
rect 19594 74824 19636 74864
rect 19676 74824 19718 74864
rect 19758 74824 19800 74864
rect 19840 74824 19849 74864
rect 34583 74824 34592 74864
rect 34632 74824 34674 74864
rect 34714 74824 34756 74864
rect 34796 74824 34838 74864
rect 34878 74824 34920 74864
rect 34960 74824 34969 74864
rect 49703 74824 49712 74864
rect 49752 74824 49794 74864
rect 49834 74824 49876 74864
rect 49916 74824 49958 74864
rect 49998 74824 50040 74864
rect 50080 74824 50089 74864
rect 64823 74824 64832 74864
rect 64872 74824 64914 74864
rect 64954 74824 64996 74864
rect 65036 74824 65078 74864
rect 65118 74824 65160 74864
rect 65200 74824 65209 74864
rect 79943 74824 79952 74864
rect 79992 74824 80034 74864
rect 80074 74824 80116 74864
rect 80156 74824 80198 74864
rect 80238 74824 80280 74864
rect 80320 74824 80329 74864
rect 95063 74824 95072 74864
rect 95112 74824 95154 74864
rect 95194 74824 95236 74864
rect 95276 74824 95318 74864
rect 95358 74824 95400 74864
rect 95440 74824 95449 74864
rect 0 74696 80 74716
rect 0 74656 652 74696
rect 692 74656 701 74696
rect 0 74636 80 74656
rect 3103 74068 3112 74108
rect 3152 74068 3194 74108
rect 3234 74068 3276 74108
rect 3316 74068 3358 74108
rect 3398 74068 3440 74108
rect 3480 74068 3489 74108
rect 18223 74068 18232 74108
rect 18272 74068 18314 74108
rect 18354 74068 18396 74108
rect 18436 74068 18478 74108
rect 18518 74068 18560 74108
rect 18600 74068 18609 74108
rect 33343 74068 33352 74108
rect 33392 74068 33434 74108
rect 33474 74068 33516 74108
rect 33556 74068 33598 74108
rect 33638 74068 33680 74108
rect 33720 74068 33729 74108
rect 48463 74068 48472 74108
rect 48512 74068 48554 74108
rect 48594 74068 48636 74108
rect 48676 74068 48718 74108
rect 48758 74068 48800 74108
rect 48840 74068 48849 74108
rect 63583 74068 63592 74108
rect 63632 74068 63674 74108
rect 63714 74068 63756 74108
rect 63796 74068 63838 74108
rect 63878 74068 63920 74108
rect 63960 74068 63969 74108
rect 78703 74068 78712 74108
rect 78752 74068 78794 74108
rect 78834 74068 78876 74108
rect 78916 74068 78958 74108
rect 78998 74068 79040 74108
rect 79080 74068 79089 74108
rect 93823 74068 93832 74108
rect 93872 74068 93914 74108
rect 93954 74068 93996 74108
rect 94036 74068 94078 74108
rect 94118 74068 94160 74108
rect 94200 74068 94209 74108
rect 4343 73312 4352 73352
rect 4392 73312 4434 73352
rect 4474 73312 4516 73352
rect 4556 73312 4598 73352
rect 4638 73312 4680 73352
rect 4720 73312 4729 73352
rect 19463 73312 19472 73352
rect 19512 73312 19554 73352
rect 19594 73312 19636 73352
rect 19676 73312 19718 73352
rect 19758 73312 19800 73352
rect 19840 73312 19849 73352
rect 34583 73312 34592 73352
rect 34632 73312 34674 73352
rect 34714 73312 34756 73352
rect 34796 73312 34838 73352
rect 34878 73312 34920 73352
rect 34960 73312 34969 73352
rect 49703 73312 49712 73352
rect 49752 73312 49794 73352
rect 49834 73312 49876 73352
rect 49916 73312 49958 73352
rect 49998 73312 50040 73352
rect 50080 73312 50089 73352
rect 64823 73312 64832 73352
rect 64872 73312 64914 73352
rect 64954 73312 64996 73352
rect 65036 73312 65078 73352
rect 65118 73312 65160 73352
rect 65200 73312 65209 73352
rect 79943 73312 79952 73352
rect 79992 73312 80034 73352
rect 80074 73312 80116 73352
rect 80156 73312 80198 73352
rect 80238 73312 80280 73352
rect 80320 73312 80329 73352
rect 95063 73312 95072 73352
rect 95112 73312 95154 73352
rect 95194 73312 95236 73352
rect 95276 73312 95318 73352
rect 95358 73312 95400 73352
rect 95440 73312 95449 73352
rect 643 72892 652 72932
rect 692 72892 701 72932
rect 0 72848 80 72868
rect 652 72848 692 72892
rect 0 72808 692 72848
rect 0 72788 80 72808
rect 3103 72556 3112 72596
rect 3152 72556 3194 72596
rect 3234 72556 3276 72596
rect 3316 72556 3358 72596
rect 3398 72556 3440 72596
rect 3480 72556 3489 72596
rect 18223 72556 18232 72596
rect 18272 72556 18314 72596
rect 18354 72556 18396 72596
rect 18436 72556 18478 72596
rect 18518 72556 18560 72596
rect 18600 72556 18609 72596
rect 33343 72556 33352 72596
rect 33392 72556 33434 72596
rect 33474 72556 33516 72596
rect 33556 72556 33598 72596
rect 33638 72556 33680 72596
rect 33720 72556 33729 72596
rect 48463 72556 48472 72596
rect 48512 72556 48554 72596
rect 48594 72556 48636 72596
rect 48676 72556 48718 72596
rect 48758 72556 48800 72596
rect 48840 72556 48849 72596
rect 63583 72556 63592 72596
rect 63632 72556 63674 72596
rect 63714 72556 63756 72596
rect 63796 72556 63838 72596
rect 63878 72556 63920 72596
rect 63960 72556 63969 72596
rect 78703 72556 78712 72596
rect 78752 72556 78794 72596
rect 78834 72556 78876 72596
rect 78916 72556 78958 72596
rect 78998 72556 79040 72596
rect 79080 72556 79089 72596
rect 93823 72556 93832 72596
rect 93872 72556 93914 72596
rect 93954 72556 93996 72596
rect 94036 72556 94078 72596
rect 94118 72556 94160 72596
rect 94200 72556 94209 72596
rect 4343 71800 4352 71840
rect 4392 71800 4434 71840
rect 4474 71800 4516 71840
rect 4556 71800 4598 71840
rect 4638 71800 4680 71840
rect 4720 71800 4729 71840
rect 19463 71800 19472 71840
rect 19512 71800 19554 71840
rect 19594 71800 19636 71840
rect 19676 71800 19718 71840
rect 19758 71800 19800 71840
rect 19840 71800 19849 71840
rect 34583 71800 34592 71840
rect 34632 71800 34674 71840
rect 34714 71800 34756 71840
rect 34796 71800 34838 71840
rect 34878 71800 34920 71840
rect 34960 71800 34969 71840
rect 49703 71800 49712 71840
rect 49752 71800 49794 71840
rect 49834 71800 49876 71840
rect 49916 71800 49958 71840
rect 49998 71800 50040 71840
rect 50080 71800 50089 71840
rect 64823 71800 64832 71840
rect 64872 71800 64914 71840
rect 64954 71800 64996 71840
rect 65036 71800 65078 71840
rect 65118 71800 65160 71840
rect 65200 71800 65209 71840
rect 79943 71800 79952 71840
rect 79992 71800 80034 71840
rect 80074 71800 80116 71840
rect 80156 71800 80198 71840
rect 80238 71800 80280 71840
rect 80320 71800 80329 71840
rect 95063 71800 95072 71840
rect 95112 71800 95154 71840
rect 95194 71800 95236 71840
rect 95276 71800 95318 71840
rect 95358 71800 95400 71840
rect 95440 71800 95449 71840
rect 3103 71044 3112 71084
rect 3152 71044 3194 71084
rect 3234 71044 3276 71084
rect 3316 71044 3358 71084
rect 3398 71044 3440 71084
rect 3480 71044 3489 71084
rect 18223 71044 18232 71084
rect 18272 71044 18314 71084
rect 18354 71044 18396 71084
rect 18436 71044 18478 71084
rect 18518 71044 18560 71084
rect 18600 71044 18609 71084
rect 33343 71044 33352 71084
rect 33392 71044 33434 71084
rect 33474 71044 33516 71084
rect 33556 71044 33598 71084
rect 33638 71044 33680 71084
rect 33720 71044 33729 71084
rect 48463 71044 48472 71084
rect 48512 71044 48554 71084
rect 48594 71044 48636 71084
rect 48676 71044 48718 71084
rect 48758 71044 48800 71084
rect 48840 71044 48849 71084
rect 63583 71044 63592 71084
rect 63632 71044 63674 71084
rect 63714 71044 63756 71084
rect 63796 71044 63838 71084
rect 63878 71044 63920 71084
rect 63960 71044 63969 71084
rect 78703 71044 78712 71084
rect 78752 71044 78794 71084
rect 78834 71044 78876 71084
rect 78916 71044 78958 71084
rect 78998 71044 79040 71084
rect 79080 71044 79089 71084
rect 93823 71044 93832 71084
rect 93872 71044 93914 71084
rect 93954 71044 93996 71084
rect 94036 71044 94078 71084
rect 94118 71044 94160 71084
rect 94200 71044 94209 71084
rect 0 71000 80 71020
rect 0 70960 652 71000
rect 692 70960 701 71000
rect 0 70940 80 70960
rect 4343 70288 4352 70328
rect 4392 70288 4434 70328
rect 4474 70288 4516 70328
rect 4556 70288 4598 70328
rect 4638 70288 4680 70328
rect 4720 70288 4729 70328
rect 19463 70288 19472 70328
rect 19512 70288 19554 70328
rect 19594 70288 19636 70328
rect 19676 70288 19718 70328
rect 19758 70288 19800 70328
rect 19840 70288 19849 70328
rect 34583 70288 34592 70328
rect 34632 70288 34674 70328
rect 34714 70288 34756 70328
rect 34796 70288 34838 70328
rect 34878 70288 34920 70328
rect 34960 70288 34969 70328
rect 49703 70288 49712 70328
rect 49752 70288 49794 70328
rect 49834 70288 49876 70328
rect 49916 70288 49958 70328
rect 49998 70288 50040 70328
rect 50080 70288 50089 70328
rect 64823 70288 64832 70328
rect 64872 70288 64914 70328
rect 64954 70288 64996 70328
rect 65036 70288 65078 70328
rect 65118 70288 65160 70328
rect 65200 70288 65209 70328
rect 79943 70288 79952 70328
rect 79992 70288 80034 70328
rect 80074 70288 80116 70328
rect 80156 70288 80198 70328
rect 80238 70288 80280 70328
rect 80320 70288 80329 70328
rect 95063 70288 95072 70328
rect 95112 70288 95154 70328
rect 95194 70288 95236 70328
rect 95276 70288 95318 70328
rect 95358 70288 95400 70328
rect 95440 70288 95449 70328
rect 3103 69532 3112 69572
rect 3152 69532 3194 69572
rect 3234 69532 3276 69572
rect 3316 69532 3358 69572
rect 3398 69532 3440 69572
rect 3480 69532 3489 69572
rect 18223 69532 18232 69572
rect 18272 69532 18314 69572
rect 18354 69532 18396 69572
rect 18436 69532 18478 69572
rect 18518 69532 18560 69572
rect 18600 69532 18609 69572
rect 33343 69532 33352 69572
rect 33392 69532 33434 69572
rect 33474 69532 33516 69572
rect 33556 69532 33598 69572
rect 33638 69532 33680 69572
rect 33720 69532 33729 69572
rect 48463 69532 48472 69572
rect 48512 69532 48554 69572
rect 48594 69532 48636 69572
rect 48676 69532 48718 69572
rect 48758 69532 48800 69572
rect 48840 69532 48849 69572
rect 63583 69532 63592 69572
rect 63632 69532 63674 69572
rect 63714 69532 63756 69572
rect 63796 69532 63838 69572
rect 63878 69532 63920 69572
rect 63960 69532 63969 69572
rect 78703 69532 78712 69572
rect 78752 69532 78794 69572
rect 78834 69532 78876 69572
rect 78916 69532 78958 69572
rect 78998 69532 79040 69572
rect 79080 69532 79089 69572
rect 93823 69532 93832 69572
rect 93872 69532 93914 69572
rect 93954 69532 93996 69572
rect 94036 69532 94078 69572
rect 94118 69532 94160 69572
rect 94200 69532 94209 69572
rect 643 69196 652 69236
rect 692 69196 701 69236
rect 0 69152 80 69172
rect 652 69152 692 69196
rect 0 69112 692 69152
rect 0 69092 80 69112
rect 835 68944 844 68984
rect 884 68944 1228 68984
rect 1268 68944 1277 68984
rect 4343 68776 4352 68816
rect 4392 68776 4434 68816
rect 4474 68776 4516 68816
rect 4556 68776 4598 68816
rect 4638 68776 4680 68816
rect 4720 68776 4729 68816
rect 19463 68776 19472 68816
rect 19512 68776 19554 68816
rect 19594 68776 19636 68816
rect 19676 68776 19718 68816
rect 19758 68776 19800 68816
rect 19840 68776 19849 68816
rect 34583 68776 34592 68816
rect 34632 68776 34674 68816
rect 34714 68776 34756 68816
rect 34796 68776 34838 68816
rect 34878 68776 34920 68816
rect 34960 68776 34969 68816
rect 49703 68776 49712 68816
rect 49752 68776 49794 68816
rect 49834 68776 49876 68816
rect 49916 68776 49958 68816
rect 49998 68776 50040 68816
rect 50080 68776 50089 68816
rect 64823 68776 64832 68816
rect 64872 68776 64914 68816
rect 64954 68776 64996 68816
rect 65036 68776 65078 68816
rect 65118 68776 65160 68816
rect 65200 68776 65209 68816
rect 79943 68776 79952 68816
rect 79992 68776 80034 68816
rect 80074 68776 80116 68816
rect 80156 68776 80198 68816
rect 80238 68776 80280 68816
rect 80320 68776 80329 68816
rect 95063 68776 95072 68816
rect 95112 68776 95154 68816
rect 95194 68776 95236 68816
rect 95276 68776 95318 68816
rect 95358 68776 95400 68816
rect 95440 68776 95449 68816
rect 3103 68020 3112 68060
rect 3152 68020 3194 68060
rect 3234 68020 3276 68060
rect 3316 68020 3358 68060
rect 3398 68020 3440 68060
rect 3480 68020 3489 68060
rect 18223 68020 18232 68060
rect 18272 68020 18314 68060
rect 18354 68020 18396 68060
rect 18436 68020 18478 68060
rect 18518 68020 18560 68060
rect 18600 68020 18609 68060
rect 33343 68020 33352 68060
rect 33392 68020 33434 68060
rect 33474 68020 33516 68060
rect 33556 68020 33598 68060
rect 33638 68020 33680 68060
rect 33720 68020 33729 68060
rect 48463 68020 48472 68060
rect 48512 68020 48554 68060
rect 48594 68020 48636 68060
rect 48676 68020 48718 68060
rect 48758 68020 48800 68060
rect 48840 68020 48849 68060
rect 63583 68020 63592 68060
rect 63632 68020 63674 68060
rect 63714 68020 63756 68060
rect 63796 68020 63838 68060
rect 63878 68020 63920 68060
rect 63960 68020 63969 68060
rect 78703 68020 78712 68060
rect 78752 68020 78794 68060
rect 78834 68020 78876 68060
rect 78916 68020 78958 68060
rect 78998 68020 79040 68060
rect 79080 68020 79089 68060
rect 93823 68020 93832 68060
rect 93872 68020 93914 68060
rect 93954 68020 93996 68060
rect 94036 68020 94078 68060
rect 94118 68020 94160 68060
rect 94200 68020 94209 68060
rect 547 67432 556 67472
rect 596 67432 844 67472
rect 884 67432 893 67472
rect 0 67304 80 67324
rect 0 67264 652 67304
rect 692 67264 701 67304
rect 4343 67264 4352 67304
rect 4392 67264 4434 67304
rect 4474 67264 4516 67304
rect 4556 67264 4598 67304
rect 4638 67264 4680 67304
rect 4720 67264 4729 67304
rect 19463 67264 19472 67304
rect 19512 67264 19554 67304
rect 19594 67264 19636 67304
rect 19676 67264 19718 67304
rect 19758 67264 19800 67304
rect 19840 67264 19849 67304
rect 34583 67264 34592 67304
rect 34632 67264 34674 67304
rect 34714 67264 34756 67304
rect 34796 67264 34838 67304
rect 34878 67264 34920 67304
rect 34960 67264 34969 67304
rect 49703 67264 49712 67304
rect 49752 67264 49794 67304
rect 49834 67264 49876 67304
rect 49916 67264 49958 67304
rect 49998 67264 50040 67304
rect 50080 67264 50089 67304
rect 64823 67264 64832 67304
rect 64872 67264 64914 67304
rect 64954 67264 64996 67304
rect 65036 67264 65078 67304
rect 65118 67264 65160 67304
rect 65200 67264 65209 67304
rect 79943 67264 79952 67304
rect 79992 67264 80034 67304
rect 80074 67264 80116 67304
rect 80156 67264 80198 67304
rect 80238 67264 80280 67304
rect 80320 67264 80329 67304
rect 95063 67264 95072 67304
rect 95112 67264 95154 67304
rect 95194 67264 95236 67304
rect 95276 67264 95318 67304
rect 95358 67264 95400 67304
rect 95440 67264 95449 67304
rect 0 67244 80 67264
rect 3103 66508 3112 66548
rect 3152 66508 3194 66548
rect 3234 66508 3276 66548
rect 3316 66508 3358 66548
rect 3398 66508 3440 66548
rect 3480 66508 3489 66548
rect 18223 66508 18232 66548
rect 18272 66508 18314 66548
rect 18354 66508 18396 66548
rect 18436 66508 18478 66548
rect 18518 66508 18560 66548
rect 18600 66508 18609 66548
rect 33343 66508 33352 66548
rect 33392 66508 33434 66548
rect 33474 66508 33516 66548
rect 33556 66508 33598 66548
rect 33638 66508 33680 66548
rect 33720 66508 33729 66548
rect 48463 66508 48472 66548
rect 48512 66508 48554 66548
rect 48594 66508 48636 66548
rect 48676 66508 48718 66548
rect 48758 66508 48800 66548
rect 48840 66508 48849 66548
rect 63583 66508 63592 66548
rect 63632 66508 63674 66548
rect 63714 66508 63756 66548
rect 63796 66508 63838 66548
rect 63878 66508 63920 66548
rect 63960 66508 63969 66548
rect 78703 66508 78712 66548
rect 78752 66508 78794 66548
rect 78834 66508 78876 66548
rect 78916 66508 78958 66548
rect 78998 66508 79040 66548
rect 79080 66508 79089 66548
rect 93823 66508 93832 66548
rect 93872 66508 93914 66548
rect 93954 66508 93996 66548
rect 94036 66508 94078 66548
rect 94118 66508 94160 66548
rect 94200 66508 94209 66548
rect 835 65920 844 65960
rect 884 65920 1132 65960
rect 1172 65920 1181 65960
rect 4343 65752 4352 65792
rect 4392 65752 4434 65792
rect 4474 65752 4516 65792
rect 4556 65752 4598 65792
rect 4638 65752 4680 65792
rect 4720 65752 4729 65792
rect 19463 65752 19472 65792
rect 19512 65752 19554 65792
rect 19594 65752 19636 65792
rect 19676 65752 19718 65792
rect 19758 65752 19800 65792
rect 19840 65752 19849 65792
rect 34583 65752 34592 65792
rect 34632 65752 34674 65792
rect 34714 65752 34756 65792
rect 34796 65752 34838 65792
rect 34878 65752 34920 65792
rect 34960 65752 34969 65792
rect 49703 65752 49712 65792
rect 49752 65752 49794 65792
rect 49834 65752 49876 65792
rect 49916 65752 49958 65792
rect 49998 65752 50040 65792
rect 50080 65752 50089 65792
rect 64823 65752 64832 65792
rect 64872 65752 64914 65792
rect 64954 65752 64996 65792
rect 65036 65752 65078 65792
rect 65118 65752 65160 65792
rect 65200 65752 65209 65792
rect 79943 65752 79952 65792
rect 79992 65752 80034 65792
rect 80074 65752 80116 65792
rect 80156 65752 80198 65792
rect 80238 65752 80280 65792
rect 80320 65752 80329 65792
rect 95063 65752 95072 65792
rect 95112 65752 95154 65792
rect 95194 65752 95236 65792
rect 95276 65752 95318 65792
rect 95358 65752 95400 65792
rect 95440 65752 95449 65792
rect 0 65456 80 65476
rect 0 65416 652 65456
rect 692 65416 701 65456
rect 0 65396 80 65416
rect 3103 64996 3112 65036
rect 3152 64996 3194 65036
rect 3234 64996 3276 65036
rect 3316 64996 3358 65036
rect 3398 64996 3440 65036
rect 3480 64996 3489 65036
rect 18223 64996 18232 65036
rect 18272 64996 18314 65036
rect 18354 64996 18396 65036
rect 18436 64996 18478 65036
rect 18518 64996 18560 65036
rect 18600 64996 18609 65036
rect 33343 64996 33352 65036
rect 33392 64996 33434 65036
rect 33474 64996 33516 65036
rect 33556 64996 33598 65036
rect 33638 64996 33680 65036
rect 33720 64996 33729 65036
rect 48463 64996 48472 65036
rect 48512 64996 48554 65036
rect 48594 64996 48636 65036
rect 48676 64996 48718 65036
rect 48758 64996 48800 65036
rect 48840 64996 48849 65036
rect 63583 64996 63592 65036
rect 63632 64996 63674 65036
rect 63714 64996 63756 65036
rect 63796 64996 63838 65036
rect 63878 64996 63920 65036
rect 63960 64996 63969 65036
rect 78703 64996 78712 65036
rect 78752 64996 78794 65036
rect 78834 64996 78876 65036
rect 78916 64996 78958 65036
rect 78998 64996 79040 65036
rect 79080 64996 79089 65036
rect 93823 64996 93832 65036
rect 93872 64996 93914 65036
rect 93954 64996 93996 65036
rect 94036 64996 94078 65036
rect 94118 64996 94160 65036
rect 94200 64996 94209 65036
rect 4343 64240 4352 64280
rect 4392 64240 4434 64280
rect 4474 64240 4516 64280
rect 4556 64240 4598 64280
rect 4638 64240 4680 64280
rect 4720 64240 4729 64280
rect 19463 64240 19472 64280
rect 19512 64240 19554 64280
rect 19594 64240 19636 64280
rect 19676 64240 19718 64280
rect 19758 64240 19800 64280
rect 19840 64240 19849 64280
rect 34583 64240 34592 64280
rect 34632 64240 34674 64280
rect 34714 64240 34756 64280
rect 34796 64240 34838 64280
rect 34878 64240 34920 64280
rect 34960 64240 34969 64280
rect 49703 64240 49712 64280
rect 49752 64240 49794 64280
rect 49834 64240 49876 64280
rect 49916 64240 49958 64280
rect 49998 64240 50040 64280
rect 50080 64240 50089 64280
rect 64823 64240 64832 64280
rect 64872 64240 64914 64280
rect 64954 64240 64996 64280
rect 65036 64240 65078 64280
rect 65118 64240 65160 64280
rect 65200 64240 65209 64280
rect 79943 64240 79952 64280
rect 79992 64240 80034 64280
rect 80074 64240 80116 64280
rect 80156 64240 80198 64280
rect 80238 64240 80280 64280
rect 80320 64240 80329 64280
rect 95063 64240 95072 64280
rect 95112 64240 95154 64280
rect 95194 64240 95236 64280
rect 95276 64240 95318 64280
rect 95358 64240 95400 64280
rect 95440 64240 95449 64280
rect 835 63652 844 63692
rect 884 63652 13228 63692
rect 13268 63652 13277 63692
rect 0 63608 80 63628
rect 0 63568 652 63608
rect 692 63568 701 63608
rect 0 63548 80 63568
rect 3103 63484 3112 63524
rect 3152 63484 3194 63524
rect 3234 63484 3276 63524
rect 3316 63484 3358 63524
rect 3398 63484 3440 63524
rect 3480 63484 3489 63524
rect 18223 63484 18232 63524
rect 18272 63484 18314 63524
rect 18354 63484 18396 63524
rect 18436 63484 18478 63524
rect 18518 63484 18560 63524
rect 18600 63484 18609 63524
rect 33343 63484 33352 63524
rect 33392 63484 33434 63524
rect 33474 63484 33516 63524
rect 33556 63484 33598 63524
rect 33638 63484 33680 63524
rect 33720 63484 33729 63524
rect 48463 63484 48472 63524
rect 48512 63484 48554 63524
rect 48594 63484 48636 63524
rect 48676 63484 48718 63524
rect 48758 63484 48800 63524
rect 48840 63484 48849 63524
rect 63583 63484 63592 63524
rect 63632 63484 63674 63524
rect 63714 63484 63756 63524
rect 63796 63484 63838 63524
rect 63878 63484 63920 63524
rect 63960 63484 63969 63524
rect 78703 63484 78712 63524
rect 78752 63484 78794 63524
rect 78834 63484 78876 63524
rect 78916 63484 78958 63524
rect 78998 63484 79040 63524
rect 79080 63484 79089 63524
rect 93823 63484 93832 63524
rect 93872 63484 93914 63524
rect 93954 63484 93996 63524
rect 94036 63484 94078 63524
rect 94118 63484 94160 63524
rect 94200 63484 94209 63524
rect 739 62980 748 63020
rect 788 62980 6508 63020
rect 6548 62980 6557 63020
rect 4343 62728 4352 62768
rect 4392 62728 4434 62768
rect 4474 62728 4516 62768
rect 4556 62728 4598 62768
rect 4638 62728 4680 62768
rect 4720 62728 4729 62768
rect 19463 62728 19472 62768
rect 19512 62728 19554 62768
rect 19594 62728 19636 62768
rect 19676 62728 19718 62768
rect 19758 62728 19800 62768
rect 19840 62728 19849 62768
rect 34583 62728 34592 62768
rect 34632 62728 34674 62768
rect 34714 62728 34756 62768
rect 34796 62728 34838 62768
rect 34878 62728 34920 62768
rect 34960 62728 34969 62768
rect 49703 62728 49712 62768
rect 49752 62728 49794 62768
rect 49834 62728 49876 62768
rect 49916 62728 49958 62768
rect 49998 62728 50040 62768
rect 50080 62728 50089 62768
rect 64823 62728 64832 62768
rect 64872 62728 64914 62768
rect 64954 62728 64996 62768
rect 65036 62728 65078 62768
rect 65118 62728 65160 62768
rect 65200 62728 65209 62768
rect 79943 62728 79952 62768
rect 79992 62728 80034 62768
rect 80074 62728 80116 62768
rect 80156 62728 80198 62768
rect 80238 62728 80280 62768
rect 80320 62728 80329 62768
rect 95063 62728 95072 62768
rect 95112 62728 95154 62768
rect 95194 62728 95236 62768
rect 95276 62728 95318 62768
rect 95358 62728 95400 62768
rect 95440 62728 95449 62768
rect 835 62140 844 62180
rect 884 62140 14188 62180
rect 14228 62140 14237 62180
rect 3103 61972 3112 62012
rect 3152 61972 3194 62012
rect 3234 61972 3276 62012
rect 3316 61972 3358 62012
rect 3398 61972 3440 62012
rect 3480 61972 3489 62012
rect 18223 61972 18232 62012
rect 18272 61972 18314 62012
rect 18354 61972 18396 62012
rect 18436 61972 18478 62012
rect 18518 61972 18560 62012
rect 18600 61972 18609 62012
rect 33343 61972 33352 62012
rect 33392 61972 33434 62012
rect 33474 61972 33516 62012
rect 33556 61972 33598 62012
rect 33638 61972 33680 62012
rect 33720 61972 33729 62012
rect 48463 61972 48472 62012
rect 48512 61972 48554 62012
rect 48594 61972 48636 62012
rect 48676 61972 48718 62012
rect 48758 61972 48800 62012
rect 48840 61972 48849 62012
rect 63583 61972 63592 62012
rect 63632 61972 63674 62012
rect 63714 61972 63756 62012
rect 63796 61972 63838 62012
rect 63878 61972 63920 62012
rect 63960 61972 63969 62012
rect 78703 61972 78712 62012
rect 78752 61972 78794 62012
rect 78834 61972 78876 62012
rect 78916 61972 78958 62012
rect 78998 61972 79040 62012
rect 79080 61972 79089 62012
rect 93823 61972 93832 62012
rect 93872 61972 93914 62012
rect 93954 61972 93996 62012
rect 94036 61972 94078 62012
rect 94118 61972 94160 62012
rect 94200 61972 94209 62012
rect 0 61760 80 61780
rect 0 61720 652 61760
rect 692 61720 701 61760
rect 0 61700 80 61720
rect 4343 61216 4352 61256
rect 4392 61216 4434 61256
rect 4474 61216 4516 61256
rect 4556 61216 4598 61256
rect 4638 61216 4680 61256
rect 4720 61216 4729 61256
rect 19463 61216 19472 61256
rect 19512 61216 19554 61256
rect 19594 61216 19636 61256
rect 19676 61216 19718 61256
rect 19758 61216 19800 61256
rect 19840 61216 19849 61256
rect 34583 61216 34592 61256
rect 34632 61216 34674 61256
rect 34714 61216 34756 61256
rect 34796 61216 34838 61256
rect 34878 61216 34920 61256
rect 34960 61216 34969 61256
rect 49703 61216 49712 61256
rect 49752 61216 49794 61256
rect 49834 61216 49876 61256
rect 49916 61216 49958 61256
rect 49998 61216 50040 61256
rect 50080 61216 50089 61256
rect 64823 61216 64832 61256
rect 64872 61216 64914 61256
rect 64954 61216 64996 61256
rect 65036 61216 65078 61256
rect 65118 61216 65160 61256
rect 65200 61216 65209 61256
rect 79943 61216 79952 61256
rect 79992 61216 80034 61256
rect 80074 61216 80116 61256
rect 80156 61216 80198 61256
rect 80238 61216 80280 61256
rect 80320 61216 80329 61256
rect 95063 61216 95072 61256
rect 95112 61216 95154 61256
rect 95194 61216 95236 61256
rect 95276 61216 95318 61256
rect 95358 61216 95400 61256
rect 95440 61216 95449 61256
rect 3103 60460 3112 60500
rect 3152 60460 3194 60500
rect 3234 60460 3276 60500
rect 3316 60460 3358 60500
rect 3398 60460 3440 60500
rect 3480 60460 3489 60500
rect 18223 60460 18232 60500
rect 18272 60460 18314 60500
rect 18354 60460 18396 60500
rect 18436 60460 18478 60500
rect 18518 60460 18560 60500
rect 18600 60460 18609 60500
rect 33343 60460 33352 60500
rect 33392 60460 33434 60500
rect 33474 60460 33516 60500
rect 33556 60460 33598 60500
rect 33638 60460 33680 60500
rect 33720 60460 33729 60500
rect 48463 60460 48472 60500
rect 48512 60460 48554 60500
rect 48594 60460 48636 60500
rect 48676 60460 48718 60500
rect 48758 60460 48800 60500
rect 48840 60460 48849 60500
rect 63583 60460 63592 60500
rect 63632 60460 63674 60500
rect 63714 60460 63756 60500
rect 63796 60460 63838 60500
rect 63878 60460 63920 60500
rect 63960 60460 63969 60500
rect 78703 60460 78712 60500
rect 78752 60460 78794 60500
rect 78834 60460 78876 60500
rect 78916 60460 78958 60500
rect 78998 60460 79040 60500
rect 79080 60460 79089 60500
rect 93823 60460 93832 60500
rect 93872 60460 93914 60500
rect 93954 60460 93996 60500
rect 94036 60460 94078 60500
rect 94118 60460 94160 60500
rect 94200 60460 94209 60500
rect 835 60292 844 60332
rect 884 60292 6604 60332
rect 6644 60292 6653 60332
rect 0 59912 80 59932
rect 0 59872 652 59912
rect 692 59872 701 59912
rect 0 59852 80 59872
rect 4343 59704 4352 59744
rect 4392 59704 4434 59744
rect 4474 59704 4516 59744
rect 4556 59704 4598 59744
rect 4638 59704 4680 59744
rect 4720 59704 4729 59744
rect 19463 59704 19472 59744
rect 19512 59704 19554 59744
rect 19594 59704 19636 59744
rect 19676 59704 19718 59744
rect 19758 59704 19800 59744
rect 19840 59704 19849 59744
rect 34583 59704 34592 59744
rect 34632 59704 34674 59744
rect 34714 59704 34756 59744
rect 34796 59704 34838 59744
rect 34878 59704 34920 59744
rect 34960 59704 34969 59744
rect 49703 59704 49712 59744
rect 49752 59704 49794 59744
rect 49834 59704 49876 59744
rect 49916 59704 49958 59744
rect 49998 59704 50040 59744
rect 50080 59704 50089 59744
rect 64823 59704 64832 59744
rect 64872 59704 64914 59744
rect 64954 59704 64996 59744
rect 65036 59704 65078 59744
rect 65118 59704 65160 59744
rect 65200 59704 65209 59744
rect 79943 59704 79952 59744
rect 79992 59704 80034 59744
rect 80074 59704 80116 59744
rect 80156 59704 80198 59744
rect 80238 59704 80280 59744
rect 80320 59704 80329 59744
rect 95063 59704 95072 59744
rect 95112 59704 95154 59744
rect 95194 59704 95236 59744
rect 95276 59704 95318 59744
rect 95358 59704 95400 59744
rect 95440 59704 95449 59744
rect 3103 58948 3112 58988
rect 3152 58948 3194 58988
rect 3234 58948 3276 58988
rect 3316 58948 3358 58988
rect 3398 58948 3440 58988
rect 3480 58948 3489 58988
rect 18223 58948 18232 58988
rect 18272 58948 18314 58988
rect 18354 58948 18396 58988
rect 18436 58948 18478 58988
rect 18518 58948 18560 58988
rect 18600 58948 18609 58988
rect 33343 58948 33352 58988
rect 33392 58948 33434 58988
rect 33474 58948 33516 58988
rect 33556 58948 33598 58988
rect 33638 58948 33680 58988
rect 33720 58948 33729 58988
rect 48463 58948 48472 58988
rect 48512 58948 48554 58988
rect 48594 58948 48636 58988
rect 48676 58948 48718 58988
rect 48758 58948 48800 58988
rect 48840 58948 48849 58988
rect 63583 58948 63592 58988
rect 63632 58948 63674 58988
rect 63714 58948 63756 58988
rect 63796 58948 63838 58988
rect 63878 58948 63920 58988
rect 63960 58948 63969 58988
rect 78703 58948 78712 58988
rect 78752 58948 78794 58988
rect 78834 58948 78876 58988
rect 78916 58948 78958 58988
rect 78998 58948 79040 58988
rect 79080 58948 79089 58988
rect 93823 58948 93832 58988
rect 93872 58948 93914 58988
rect 93954 58948 93996 58988
rect 94036 58948 94078 58988
rect 94118 58948 94160 58988
rect 94200 58948 94209 58988
rect 4343 58192 4352 58232
rect 4392 58192 4434 58232
rect 4474 58192 4516 58232
rect 4556 58192 4598 58232
rect 4638 58192 4680 58232
rect 4720 58192 4729 58232
rect 19463 58192 19472 58232
rect 19512 58192 19554 58232
rect 19594 58192 19636 58232
rect 19676 58192 19718 58232
rect 19758 58192 19800 58232
rect 19840 58192 19849 58232
rect 34583 58192 34592 58232
rect 34632 58192 34674 58232
rect 34714 58192 34756 58232
rect 34796 58192 34838 58232
rect 34878 58192 34920 58232
rect 34960 58192 34969 58232
rect 49703 58192 49712 58232
rect 49752 58192 49794 58232
rect 49834 58192 49876 58232
rect 49916 58192 49958 58232
rect 49998 58192 50040 58232
rect 50080 58192 50089 58232
rect 64823 58192 64832 58232
rect 64872 58192 64914 58232
rect 64954 58192 64996 58232
rect 65036 58192 65078 58232
rect 65118 58192 65160 58232
rect 65200 58192 65209 58232
rect 79943 58192 79952 58232
rect 79992 58192 80034 58232
rect 80074 58192 80116 58232
rect 80156 58192 80198 58232
rect 80238 58192 80280 58232
rect 80320 58192 80329 58232
rect 95063 58192 95072 58232
rect 95112 58192 95154 58232
rect 95194 58192 95236 58232
rect 95276 58192 95318 58232
rect 95358 58192 95400 58232
rect 95440 58192 95449 58232
rect 0 58064 80 58084
rect 0 58024 652 58064
rect 692 58024 701 58064
rect 0 58004 80 58024
rect 1027 57940 1036 57980
rect 1076 57940 5836 57980
rect 5876 57940 6548 57980
rect 6508 57896 6548 57940
rect 6192 57856 6220 57896
rect 6260 57856 6316 57896
rect 6356 57856 6384 57896
rect 6499 57856 6508 57896
rect 6548 57856 6557 57896
rect 3103 57436 3112 57476
rect 3152 57436 3194 57476
rect 3234 57436 3276 57476
rect 3316 57436 3358 57476
rect 3398 57436 3440 57476
rect 3480 57436 3489 57476
rect 18223 57436 18232 57476
rect 18272 57436 18314 57476
rect 18354 57436 18396 57476
rect 18436 57436 18478 57476
rect 18518 57436 18560 57476
rect 18600 57436 18609 57476
rect 33343 57436 33352 57476
rect 33392 57436 33434 57476
rect 33474 57436 33516 57476
rect 33556 57436 33598 57476
rect 33638 57436 33680 57476
rect 33720 57436 33729 57476
rect 48463 57436 48472 57476
rect 48512 57436 48554 57476
rect 48594 57436 48636 57476
rect 48676 57436 48718 57476
rect 48758 57436 48800 57476
rect 48840 57436 48849 57476
rect 63583 57436 63592 57476
rect 63632 57436 63674 57476
rect 63714 57436 63756 57476
rect 63796 57436 63838 57476
rect 63878 57436 63920 57476
rect 63960 57436 63969 57476
rect 78703 57436 78712 57476
rect 78752 57436 78794 57476
rect 78834 57436 78876 57476
rect 78916 57436 78958 57476
rect 78998 57436 79040 57476
rect 79080 57436 79089 57476
rect 93823 57436 93832 57476
rect 93872 57436 93914 57476
rect 93954 57436 93996 57476
rect 94036 57436 94078 57476
rect 94118 57436 94160 57476
rect 94200 57436 94209 57476
rect 835 57100 844 57140
rect 884 57100 6028 57140
rect 6068 57100 6220 57140
rect 6260 57100 6269 57140
rect 6412 57100 7220 57140
rect 6412 57056 6452 57100
rect 7180 57056 7220 57100
rect 5923 57016 5932 57056
rect 5972 57016 6452 57056
rect 6499 57016 6508 57056
rect 6548 57016 6557 57056
rect 7171 57016 7180 57056
rect 7220 57016 7229 57056
rect 6508 56972 6548 57016
rect 5827 56932 5836 56972
rect 5876 56932 6548 56972
rect 4343 56680 4352 56720
rect 4392 56680 4434 56720
rect 4474 56680 4516 56720
rect 4556 56680 4598 56720
rect 4638 56680 4680 56720
rect 4720 56680 4729 56720
rect 19463 56680 19472 56720
rect 19512 56680 19554 56720
rect 19594 56680 19636 56720
rect 19676 56680 19718 56720
rect 19758 56680 19800 56720
rect 19840 56680 19849 56720
rect 34583 56680 34592 56720
rect 34632 56680 34674 56720
rect 34714 56680 34756 56720
rect 34796 56680 34838 56720
rect 34878 56680 34920 56720
rect 34960 56680 34969 56720
rect 49703 56680 49712 56720
rect 49752 56680 49794 56720
rect 49834 56680 49876 56720
rect 49916 56680 49958 56720
rect 49998 56680 50040 56720
rect 50080 56680 50089 56720
rect 64823 56680 64832 56720
rect 64872 56680 64914 56720
rect 64954 56680 64996 56720
rect 65036 56680 65078 56720
rect 65118 56680 65160 56720
rect 65200 56680 65209 56720
rect 79943 56680 79952 56720
rect 79992 56680 80034 56720
rect 80074 56680 80116 56720
rect 80156 56680 80198 56720
rect 80238 56680 80280 56720
rect 80320 56680 80329 56720
rect 95063 56680 95072 56720
rect 95112 56680 95154 56720
rect 95194 56680 95236 56720
rect 95276 56680 95318 56720
rect 95358 56680 95400 56720
rect 95440 56680 95449 56720
rect 5635 56344 5644 56384
rect 5684 56344 6604 56384
rect 6644 56344 6988 56384
rect 7028 56344 7037 56384
rect 643 56260 652 56300
rect 692 56260 701 56300
rect 0 56216 80 56236
rect 652 56216 692 56260
rect 0 56176 692 56216
rect 0 56156 80 56176
rect 739 56092 748 56132
rect 788 56092 6412 56132
rect 6452 56092 6461 56132
rect 3103 55924 3112 55964
rect 3152 55924 3194 55964
rect 3234 55924 3276 55964
rect 3316 55924 3358 55964
rect 3398 55924 3440 55964
rect 3480 55924 3489 55964
rect 18223 55924 18232 55964
rect 18272 55924 18314 55964
rect 18354 55924 18396 55964
rect 18436 55924 18478 55964
rect 18518 55924 18560 55964
rect 18600 55924 18609 55964
rect 33343 55924 33352 55964
rect 33392 55924 33434 55964
rect 33474 55924 33516 55964
rect 33556 55924 33598 55964
rect 33638 55924 33680 55964
rect 33720 55924 33729 55964
rect 48463 55924 48472 55964
rect 48512 55924 48554 55964
rect 48594 55924 48636 55964
rect 48676 55924 48718 55964
rect 48758 55924 48800 55964
rect 48840 55924 48849 55964
rect 63583 55924 63592 55964
rect 63632 55924 63674 55964
rect 63714 55924 63756 55964
rect 63796 55924 63838 55964
rect 63878 55924 63920 55964
rect 63960 55924 63969 55964
rect 78703 55924 78712 55964
rect 78752 55924 78794 55964
rect 78834 55924 78876 55964
rect 78916 55924 78958 55964
rect 78998 55924 79040 55964
rect 79080 55924 79089 55964
rect 93823 55924 93832 55964
rect 93872 55924 93914 55964
rect 93954 55924 93996 55964
rect 94036 55924 94078 55964
rect 94118 55924 94160 55964
rect 94200 55924 94209 55964
rect 4343 55168 4352 55208
rect 4392 55168 4434 55208
rect 4474 55168 4516 55208
rect 4556 55168 4598 55208
rect 4638 55168 4680 55208
rect 4720 55168 4729 55208
rect 19463 55168 19472 55208
rect 19512 55168 19554 55208
rect 19594 55168 19636 55208
rect 19676 55168 19718 55208
rect 19758 55168 19800 55208
rect 19840 55168 19849 55208
rect 34583 55168 34592 55208
rect 34632 55168 34674 55208
rect 34714 55168 34756 55208
rect 34796 55168 34838 55208
rect 34878 55168 34920 55208
rect 34960 55168 34969 55208
rect 49703 55168 49712 55208
rect 49752 55168 49794 55208
rect 49834 55168 49876 55208
rect 49916 55168 49958 55208
rect 49998 55168 50040 55208
rect 50080 55168 50089 55208
rect 64823 55168 64832 55208
rect 64872 55168 64914 55208
rect 64954 55168 64996 55208
rect 65036 55168 65078 55208
rect 65118 55168 65160 55208
rect 65200 55168 65209 55208
rect 79943 55168 79952 55208
rect 79992 55168 80034 55208
rect 80074 55168 80116 55208
rect 80156 55168 80198 55208
rect 80238 55168 80280 55208
rect 80320 55168 80329 55208
rect 95063 55168 95072 55208
rect 95112 55168 95154 55208
rect 95194 55168 95236 55208
rect 95276 55168 95318 55208
rect 95358 55168 95400 55208
rect 95440 55168 95449 55208
rect 3103 54412 3112 54452
rect 3152 54412 3194 54452
rect 3234 54412 3276 54452
rect 3316 54412 3358 54452
rect 3398 54412 3440 54452
rect 3480 54412 3489 54452
rect 18223 54412 18232 54452
rect 18272 54412 18314 54452
rect 18354 54412 18396 54452
rect 18436 54412 18478 54452
rect 18518 54412 18560 54452
rect 18600 54412 18609 54452
rect 33343 54412 33352 54452
rect 33392 54412 33434 54452
rect 33474 54412 33516 54452
rect 33556 54412 33598 54452
rect 33638 54412 33680 54452
rect 33720 54412 33729 54452
rect 48463 54412 48472 54452
rect 48512 54412 48554 54452
rect 48594 54412 48636 54452
rect 48676 54412 48718 54452
rect 48758 54412 48800 54452
rect 48840 54412 48849 54452
rect 63583 54412 63592 54452
rect 63632 54412 63674 54452
rect 63714 54412 63756 54452
rect 63796 54412 63838 54452
rect 63878 54412 63920 54452
rect 63960 54412 63969 54452
rect 78703 54412 78712 54452
rect 78752 54412 78794 54452
rect 78834 54412 78876 54452
rect 78916 54412 78958 54452
rect 78998 54412 79040 54452
rect 79080 54412 79089 54452
rect 93823 54412 93832 54452
rect 93872 54412 93914 54452
rect 93954 54412 93996 54452
rect 94036 54412 94078 54452
rect 94118 54412 94160 54452
rect 94200 54412 94209 54452
rect 0 54368 80 54388
rect 0 54328 652 54368
rect 692 54328 701 54368
rect 0 54308 80 54328
rect 4343 53656 4352 53696
rect 4392 53656 4434 53696
rect 4474 53656 4516 53696
rect 4556 53656 4598 53696
rect 4638 53656 4680 53696
rect 4720 53656 4729 53696
rect 19463 53656 19472 53696
rect 19512 53656 19554 53696
rect 19594 53656 19636 53696
rect 19676 53656 19718 53696
rect 19758 53656 19800 53696
rect 19840 53656 19849 53696
rect 34583 53656 34592 53696
rect 34632 53656 34674 53696
rect 34714 53656 34756 53696
rect 34796 53656 34838 53696
rect 34878 53656 34920 53696
rect 34960 53656 34969 53696
rect 49703 53656 49712 53696
rect 49752 53656 49794 53696
rect 49834 53656 49876 53696
rect 49916 53656 49958 53696
rect 49998 53656 50040 53696
rect 50080 53656 50089 53696
rect 64823 53656 64832 53696
rect 64872 53656 64914 53696
rect 64954 53656 64996 53696
rect 65036 53656 65078 53696
rect 65118 53656 65160 53696
rect 65200 53656 65209 53696
rect 79943 53656 79952 53696
rect 79992 53656 80034 53696
rect 80074 53656 80116 53696
rect 80156 53656 80198 53696
rect 80238 53656 80280 53696
rect 80320 53656 80329 53696
rect 95063 53656 95072 53696
rect 95112 53656 95154 53696
rect 95194 53656 95236 53696
rect 95276 53656 95318 53696
rect 95358 53656 95400 53696
rect 95440 53656 95449 53696
rect 5827 53068 5836 53108
rect 5876 53068 6412 53108
rect 6452 53068 6461 53108
rect 3103 52900 3112 52940
rect 3152 52900 3194 52940
rect 3234 52900 3276 52940
rect 3316 52900 3358 52940
rect 3398 52900 3440 52940
rect 3480 52900 3489 52940
rect 18223 52900 18232 52940
rect 18272 52900 18314 52940
rect 18354 52900 18396 52940
rect 18436 52900 18478 52940
rect 18518 52900 18560 52940
rect 18600 52900 18609 52940
rect 33343 52900 33352 52940
rect 33392 52900 33434 52940
rect 33474 52900 33516 52940
rect 33556 52900 33598 52940
rect 33638 52900 33680 52940
rect 33720 52900 33729 52940
rect 48463 52900 48472 52940
rect 48512 52900 48554 52940
rect 48594 52900 48636 52940
rect 48676 52900 48718 52940
rect 48758 52900 48800 52940
rect 48840 52900 48849 52940
rect 63583 52900 63592 52940
rect 63632 52900 63674 52940
rect 63714 52900 63756 52940
rect 63796 52900 63838 52940
rect 63878 52900 63920 52940
rect 63960 52900 63969 52940
rect 78703 52900 78712 52940
rect 78752 52900 78794 52940
rect 78834 52900 78876 52940
rect 78916 52900 78958 52940
rect 78998 52900 79040 52940
rect 79080 52900 79089 52940
rect 93823 52900 93832 52940
rect 93872 52900 93914 52940
rect 93954 52900 93996 52940
rect 94036 52900 94078 52940
rect 94118 52900 94160 52940
rect 94200 52900 94209 52940
rect 1027 52816 1036 52856
rect 1076 52816 6185 52856
rect 6225 52816 6508 52856
rect 6548 52816 6557 52856
rect 931 52648 940 52688
rect 980 52648 6028 52688
rect 6068 52648 6700 52688
rect 6740 52648 6749 52688
rect 643 52564 652 52604
rect 692 52564 701 52604
rect 5731 52564 5740 52604
rect 5780 52564 6316 52604
rect 6356 52564 6365 52604
rect 0 52520 80 52540
rect 652 52520 692 52564
rect 0 52480 692 52520
rect 835 52480 844 52520
rect 884 52480 2284 52520
rect 2324 52480 2333 52520
rect 4099 52480 4108 52520
rect 4148 52480 5932 52520
rect 5972 52480 5981 52520
rect 0 52460 80 52480
rect 6211 52312 6220 52352
rect 6260 52312 6412 52352
rect 6452 52312 6461 52352
rect 4343 52144 4352 52184
rect 4392 52144 4434 52184
rect 4474 52144 4516 52184
rect 4556 52144 4598 52184
rect 4638 52144 4680 52184
rect 4720 52144 4729 52184
rect 19463 52144 19472 52184
rect 19512 52144 19554 52184
rect 19594 52144 19636 52184
rect 19676 52144 19718 52184
rect 19758 52144 19800 52184
rect 19840 52144 19849 52184
rect 34583 52144 34592 52184
rect 34632 52144 34674 52184
rect 34714 52144 34756 52184
rect 34796 52144 34838 52184
rect 34878 52144 34920 52184
rect 34960 52144 34969 52184
rect 49703 52144 49712 52184
rect 49752 52144 49794 52184
rect 49834 52144 49876 52184
rect 49916 52144 49958 52184
rect 49998 52144 50040 52184
rect 50080 52144 50089 52184
rect 64823 52144 64832 52184
rect 64872 52144 64914 52184
rect 64954 52144 64996 52184
rect 65036 52144 65078 52184
rect 65118 52144 65160 52184
rect 65200 52144 65209 52184
rect 79943 52144 79952 52184
rect 79992 52144 80034 52184
rect 80074 52144 80116 52184
rect 80156 52144 80198 52184
rect 80238 52144 80280 52184
rect 80320 52144 80329 52184
rect 95063 52144 95072 52184
rect 95112 52144 95154 52184
rect 95194 52144 95236 52184
rect 95276 52144 95318 52184
rect 95358 52144 95400 52184
rect 95440 52144 95449 52184
rect 2179 51976 2188 52016
rect 2228 51976 3244 52016
rect 3284 51976 5548 52016
rect 5588 51976 5597 52016
rect 2947 51892 2956 51932
rect 2996 51892 3916 51932
rect 3956 51892 5300 51932
rect 5260 51848 5300 51892
rect 1219 51808 1228 51848
rect 1268 51808 2092 51848
rect 2132 51808 2764 51848
rect 2804 51808 2813 51848
rect 3427 51808 3436 51848
rect 3476 51808 4012 51848
rect 4052 51808 4061 51848
rect 5251 51808 5260 51848
rect 5300 51808 5309 51848
rect 5443 51808 5452 51848
rect 5492 51808 6412 51848
rect 6452 51808 6796 51848
rect 6836 51808 6845 51848
rect 5923 51724 5932 51764
rect 5972 51724 6124 51764
rect 6164 51724 6932 51764
rect 6892 51680 6932 51724
rect 2659 51640 2668 51680
rect 2708 51640 6220 51680
rect 6260 51640 6269 51680
rect 6883 51640 6892 51680
rect 6932 51640 6941 51680
rect 3103 51388 3112 51428
rect 3152 51388 3194 51428
rect 3234 51388 3276 51428
rect 3316 51388 3358 51428
rect 3398 51388 3440 51428
rect 3480 51388 3489 51428
rect 18223 51388 18232 51428
rect 18272 51388 18314 51428
rect 18354 51388 18396 51428
rect 18436 51388 18478 51428
rect 18518 51388 18560 51428
rect 18600 51388 18609 51428
rect 33343 51388 33352 51428
rect 33392 51388 33434 51428
rect 33474 51388 33516 51428
rect 33556 51388 33598 51428
rect 33638 51388 33680 51428
rect 33720 51388 33729 51428
rect 48463 51388 48472 51428
rect 48512 51388 48554 51428
rect 48594 51388 48636 51428
rect 48676 51388 48718 51428
rect 48758 51388 48800 51428
rect 48840 51388 48849 51428
rect 63583 51388 63592 51428
rect 63632 51388 63674 51428
rect 63714 51388 63756 51428
rect 63796 51388 63838 51428
rect 63878 51388 63920 51428
rect 63960 51388 63969 51428
rect 78703 51388 78712 51428
rect 78752 51388 78794 51428
rect 78834 51388 78876 51428
rect 78916 51388 78958 51428
rect 78998 51388 79040 51428
rect 79080 51388 79089 51428
rect 93823 51388 93832 51428
rect 93872 51388 93914 51428
rect 93954 51388 93996 51428
rect 94036 51388 94078 51428
rect 94118 51388 94160 51428
rect 94200 51388 94209 51428
rect 1891 50800 1900 50840
rect 1940 50800 2476 50840
rect 2516 50800 2525 50840
rect 0 50672 80 50692
rect 0 50632 652 50672
rect 692 50632 701 50672
rect 4343 50632 4352 50672
rect 4392 50632 4434 50672
rect 4474 50632 4516 50672
rect 4556 50632 4598 50672
rect 4638 50632 4680 50672
rect 4720 50632 4729 50672
rect 19463 50632 19472 50672
rect 19512 50632 19554 50672
rect 19594 50632 19636 50672
rect 19676 50632 19718 50672
rect 19758 50632 19800 50672
rect 19840 50632 19849 50672
rect 34583 50632 34592 50672
rect 34632 50632 34674 50672
rect 34714 50632 34756 50672
rect 34796 50632 34838 50672
rect 34878 50632 34920 50672
rect 34960 50632 34969 50672
rect 49703 50632 49712 50672
rect 49752 50632 49794 50672
rect 49834 50632 49876 50672
rect 49916 50632 49958 50672
rect 49998 50632 50040 50672
rect 50080 50632 50089 50672
rect 64823 50632 64832 50672
rect 64872 50632 64914 50672
rect 64954 50632 64996 50672
rect 65036 50632 65078 50672
rect 65118 50632 65160 50672
rect 65200 50632 65209 50672
rect 79943 50632 79952 50672
rect 79992 50632 80034 50672
rect 80074 50632 80116 50672
rect 80156 50632 80198 50672
rect 80238 50632 80280 50672
rect 80320 50632 80329 50672
rect 95063 50632 95072 50672
rect 95112 50632 95154 50672
rect 95194 50632 95236 50672
rect 95276 50632 95318 50672
rect 95358 50632 95400 50672
rect 95440 50632 95449 50672
rect 0 50612 80 50632
rect 3103 49876 3112 49916
rect 3152 49876 3194 49916
rect 3234 49876 3276 49916
rect 3316 49876 3358 49916
rect 3398 49876 3440 49916
rect 3480 49876 3489 49916
rect 18223 49876 18232 49916
rect 18272 49876 18314 49916
rect 18354 49876 18396 49916
rect 18436 49876 18478 49916
rect 18518 49876 18560 49916
rect 18600 49876 18609 49916
rect 33343 49876 33352 49916
rect 33392 49876 33434 49916
rect 33474 49876 33516 49916
rect 33556 49876 33598 49916
rect 33638 49876 33680 49916
rect 33720 49876 33729 49916
rect 48463 49876 48472 49916
rect 48512 49876 48554 49916
rect 48594 49876 48636 49916
rect 48676 49876 48718 49916
rect 48758 49876 48800 49916
rect 48840 49876 48849 49916
rect 63583 49876 63592 49916
rect 63632 49876 63674 49916
rect 63714 49876 63756 49916
rect 63796 49876 63838 49916
rect 63878 49876 63920 49916
rect 63960 49876 63969 49916
rect 78703 49876 78712 49916
rect 78752 49876 78794 49916
rect 78834 49876 78876 49916
rect 78916 49876 78958 49916
rect 78998 49876 79040 49916
rect 79080 49876 79089 49916
rect 93823 49876 93832 49916
rect 93872 49876 93914 49916
rect 93954 49876 93996 49916
rect 94036 49876 94078 49916
rect 94118 49876 94160 49916
rect 94200 49876 94209 49916
rect 835 49456 844 49496
rect 884 49456 7852 49496
rect 7892 49456 7901 49496
rect 4343 49120 4352 49160
rect 4392 49120 4434 49160
rect 4474 49120 4516 49160
rect 4556 49120 4598 49160
rect 4638 49120 4680 49160
rect 4720 49120 4729 49160
rect 19463 49120 19472 49160
rect 19512 49120 19554 49160
rect 19594 49120 19636 49160
rect 19676 49120 19718 49160
rect 19758 49120 19800 49160
rect 19840 49120 19849 49160
rect 34583 49120 34592 49160
rect 34632 49120 34674 49160
rect 34714 49120 34756 49160
rect 34796 49120 34838 49160
rect 34878 49120 34920 49160
rect 34960 49120 34969 49160
rect 49703 49120 49712 49160
rect 49752 49120 49794 49160
rect 49834 49120 49876 49160
rect 49916 49120 49958 49160
rect 49998 49120 50040 49160
rect 50080 49120 50089 49160
rect 64823 49120 64832 49160
rect 64872 49120 64914 49160
rect 64954 49120 64996 49160
rect 65036 49120 65078 49160
rect 65118 49120 65160 49160
rect 65200 49120 65209 49160
rect 79943 49120 79952 49160
rect 79992 49120 80034 49160
rect 80074 49120 80116 49160
rect 80156 49120 80198 49160
rect 80238 49120 80280 49160
rect 80320 49120 80329 49160
rect 95063 49120 95072 49160
rect 95112 49120 95154 49160
rect 95194 49120 95236 49160
rect 95276 49120 95318 49160
rect 95358 49120 95400 49160
rect 95440 49120 95449 49160
rect 0 48824 80 48844
rect 0 48784 652 48824
rect 692 48784 701 48824
rect 0 48764 80 48784
rect 3103 48364 3112 48404
rect 3152 48364 3194 48404
rect 3234 48364 3276 48404
rect 3316 48364 3358 48404
rect 3398 48364 3440 48404
rect 3480 48364 3489 48404
rect 18223 48364 18232 48404
rect 18272 48364 18314 48404
rect 18354 48364 18396 48404
rect 18436 48364 18478 48404
rect 18518 48364 18560 48404
rect 18600 48364 18609 48404
rect 33343 48364 33352 48404
rect 33392 48364 33434 48404
rect 33474 48364 33516 48404
rect 33556 48364 33598 48404
rect 33638 48364 33680 48404
rect 33720 48364 33729 48404
rect 48463 48364 48472 48404
rect 48512 48364 48554 48404
rect 48594 48364 48636 48404
rect 48676 48364 48718 48404
rect 48758 48364 48800 48404
rect 48840 48364 48849 48404
rect 63583 48364 63592 48404
rect 63632 48364 63674 48404
rect 63714 48364 63756 48404
rect 63796 48364 63838 48404
rect 63878 48364 63920 48404
rect 63960 48364 63969 48404
rect 78703 48364 78712 48404
rect 78752 48364 78794 48404
rect 78834 48364 78876 48404
rect 78916 48364 78958 48404
rect 78998 48364 79040 48404
rect 79080 48364 79089 48404
rect 93823 48364 93832 48404
rect 93872 48364 93914 48404
rect 93954 48364 93996 48404
rect 94036 48364 94078 48404
rect 94118 48364 94160 48404
rect 94200 48364 94209 48404
rect 3907 47944 3916 47984
rect 3956 47944 6220 47984
rect 6260 47944 6269 47984
rect 6403 47944 6412 47984
rect 6452 47944 7564 47984
rect 7604 47944 9868 47984
rect 9908 47944 13804 47984
rect 13844 47944 13853 47984
rect 739 47860 748 47900
rect 788 47860 9388 47900
rect 9428 47860 9437 47900
rect 4343 47608 4352 47648
rect 4392 47608 4434 47648
rect 4474 47608 4516 47648
rect 4556 47608 4598 47648
rect 4638 47608 4680 47648
rect 4720 47608 4729 47648
rect 19463 47608 19472 47648
rect 19512 47608 19554 47648
rect 19594 47608 19636 47648
rect 19676 47608 19718 47648
rect 19758 47608 19800 47648
rect 19840 47608 19849 47648
rect 34583 47608 34592 47648
rect 34632 47608 34674 47648
rect 34714 47608 34756 47648
rect 34796 47608 34838 47648
rect 34878 47608 34920 47648
rect 34960 47608 34969 47648
rect 49703 47608 49712 47648
rect 49752 47608 49794 47648
rect 49834 47608 49876 47648
rect 49916 47608 49958 47648
rect 49998 47608 50040 47648
rect 50080 47608 50089 47648
rect 64823 47608 64832 47648
rect 64872 47608 64914 47648
rect 64954 47608 64996 47648
rect 65036 47608 65078 47648
rect 65118 47608 65160 47648
rect 65200 47608 65209 47648
rect 79943 47608 79952 47648
rect 79992 47608 80034 47648
rect 80074 47608 80116 47648
rect 80156 47608 80198 47648
rect 80238 47608 80280 47648
rect 80320 47608 80329 47648
rect 95063 47608 95072 47648
rect 95112 47608 95154 47648
rect 95194 47608 95236 47648
rect 95276 47608 95318 47648
rect 95358 47608 95400 47648
rect 95440 47608 95449 47648
rect 835 47524 844 47564
rect 884 47524 13132 47564
rect 13172 47524 13612 47564
rect 13652 47524 13661 47564
rect 1027 47440 1036 47480
rect 1076 47440 1996 47480
rect 2036 47440 2045 47480
rect 2275 47440 2284 47480
rect 2324 47440 4012 47480
rect 4052 47440 4061 47480
rect 1996 47396 2036 47440
rect 1996 47356 2476 47396
rect 2516 47356 2525 47396
rect 2947 47356 2956 47396
rect 2996 47356 5836 47396
rect 5876 47356 5885 47396
rect 6595 47356 6604 47396
rect 6644 47356 6653 47396
rect 5836 47312 5876 47356
rect 6604 47312 6644 47356
rect 547 47272 556 47312
rect 596 47272 2092 47312
rect 2132 47272 2764 47312
rect 2804 47272 2813 47312
rect 5836 47272 6508 47312
rect 6548 47272 6557 47312
rect 6604 47272 7372 47312
rect 7412 47272 8044 47312
rect 8084 47272 9484 47312
rect 9524 47272 9533 47312
rect 13219 47272 13228 47312
rect 13268 47272 13900 47312
rect 13940 47272 13949 47312
rect 14083 47272 14092 47312
rect 14132 47272 14284 47312
rect 14324 47272 14572 47312
rect 14612 47272 14621 47312
rect 5923 47188 5932 47228
rect 5972 47188 6892 47228
rect 6932 47188 6941 47228
rect 3811 47104 3820 47144
rect 3860 47104 6320 47144
rect 6979 47104 6988 47144
rect 7028 47104 7372 47144
rect 7412 47104 7421 47144
rect 6280 47060 6320 47104
rect 6280 47020 6796 47060
rect 6836 47020 7564 47060
rect 7604 47020 7613 47060
rect 0 46976 80 46996
rect 0 46936 652 46976
rect 692 46936 701 46976
rect 0 46916 80 46936
rect 3103 46852 3112 46892
rect 3152 46852 3194 46892
rect 3234 46852 3276 46892
rect 3316 46852 3358 46892
rect 3398 46852 3440 46892
rect 3480 46852 3489 46892
rect 18223 46852 18232 46892
rect 18272 46852 18314 46892
rect 18354 46852 18396 46892
rect 18436 46852 18478 46892
rect 18518 46852 18560 46892
rect 18600 46852 18609 46892
rect 33343 46852 33352 46892
rect 33392 46852 33434 46892
rect 33474 46852 33516 46892
rect 33556 46852 33598 46892
rect 33638 46852 33680 46892
rect 33720 46852 33729 46892
rect 48463 46852 48472 46892
rect 48512 46852 48554 46892
rect 48594 46852 48636 46892
rect 48676 46852 48718 46892
rect 48758 46852 48800 46892
rect 48840 46852 48849 46892
rect 63583 46852 63592 46892
rect 63632 46852 63674 46892
rect 63714 46852 63756 46892
rect 63796 46852 63838 46892
rect 63878 46852 63920 46892
rect 63960 46852 63969 46892
rect 78703 46852 78712 46892
rect 78752 46852 78794 46892
rect 78834 46852 78876 46892
rect 78916 46852 78958 46892
rect 78998 46852 79040 46892
rect 79080 46852 79089 46892
rect 93823 46852 93832 46892
rect 93872 46852 93914 46892
rect 93954 46852 93996 46892
rect 94036 46852 94078 46892
rect 94118 46852 94160 46892
rect 94200 46852 94209 46892
rect 14083 46432 14092 46472
rect 14132 46432 14380 46472
rect 14420 46432 14956 46472
rect 14996 46432 15005 46472
rect 4343 46096 4352 46136
rect 4392 46096 4434 46136
rect 4474 46096 4516 46136
rect 4556 46096 4598 46136
rect 4638 46096 4680 46136
rect 4720 46096 4729 46136
rect 19463 46096 19472 46136
rect 19512 46096 19554 46136
rect 19594 46096 19636 46136
rect 19676 46096 19718 46136
rect 19758 46096 19800 46136
rect 19840 46096 19849 46136
rect 34583 46096 34592 46136
rect 34632 46096 34674 46136
rect 34714 46096 34756 46136
rect 34796 46096 34838 46136
rect 34878 46096 34920 46136
rect 34960 46096 34969 46136
rect 49703 46096 49712 46136
rect 49752 46096 49794 46136
rect 49834 46096 49876 46136
rect 49916 46096 49958 46136
rect 49998 46096 50040 46136
rect 50080 46096 50089 46136
rect 64823 46096 64832 46136
rect 64872 46096 64914 46136
rect 64954 46096 64996 46136
rect 65036 46096 65078 46136
rect 65118 46096 65160 46136
rect 65200 46096 65209 46136
rect 79943 46096 79952 46136
rect 79992 46096 80034 46136
rect 80074 46096 80116 46136
rect 80156 46096 80198 46136
rect 80238 46096 80280 46136
rect 80320 46096 80329 46136
rect 95063 46096 95072 46136
rect 95112 46096 95154 46136
rect 95194 46096 95236 46136
rect 95276 46096 95318 46136
rect 95358 46096 95400 46136
rect 95440 46096 95449 46136
rect 835 45928 844 45968
rect 884 45928 14092 45968
rect 14132 45928 14572 45968
rect 14612 45928 14621 45968
rect 1123 45760 1132 45800
rect 1172 45760 7756 45800
rect 7796 45760 8236 45800
rect 8276 45760 8285 45800
rect 3103 45340 3112 45380
rect 3152 45340 3194 45380
rect 3234 45340 3276 45380
rect 3316 45340 3358 45380
rect 3398 45340 3440 45380
rect 3480 45340 3489 45380
rect 18223 45340 18232 45380
rect 18272 45340 18314 45380
rect 18354 45340 18396 45380
rect 18436 45340 18478 45380
rect 18518 45340 18560 45380
rect 18600 45340 18609 45380
rect 33343 45340 33352 45380
rect 33392 45340 33434 45380
rect 33474 45340 33516 45380
rect 33556 45340 33598 45380
rect 33638 45340 33680 45380
rect 33720 45340 33729 45380
rect 48463 45340 48472 45380
rect 48512 45340 48554 45380
rect 48594 45340 48636 45380
rect 48676 45340 48718 45380
rect 48758 45340 48800 45380
rect 48840 45340 48849 45380
rect 63583 45340 63592 45380
rect 63632 45340 63674 45380
rect 63714 45340 63756 45380
rect 63796 45340 63838 45380
rect 63878 45340 63920 45380
rect 63960 45340 63969 45380
rect 78703 45340 78712 45380
rect 78752 45340 78794 45380
rect 78834 45340 78876 45380
rect 78916 45340 78958 45380
rect 78998 45340 79040 45380
rect 79080 45340 79089 45380
rect 93823 45340 93832 45380
rect 93872 45340 93914 45380
rect 93954 45340 93996 45380
rect 94036 45340 94078 45380
rect 94118 45340 94160 45380
rect 94200 45340 94209 45380
rect 0 45128 80 45148
rect 0 45088 652 45128
rect 692 45088 701 45128
rect 0 45068 80 45088
rect 1123 44752 1132 44792
rect 1172 44752 14092 44792
rect 14132 44752 14141 44792
rect 4343 44584 4352 44624
rect 4392 44584 4434 44624
rect 4474 44584 4516 44624
rect 4556 44584 4598 44624
rect 4638 44584 4680 44624
rect 4720 44584 4729 44624
rect 19463 44584 19472 44624
rect 19512 44584 19554 44624
rect 19594 44584 19636 44624
rect 19676 44584 19718 44624
rect 19758 44584 19800 44624
rect 19840 44584 19849 44624
rect 34583 44584 34592 44624
rect 34632 44584 34674 44624
rect 34714 44584 34756 44624
rect 34796 44584 34838 44624
rect 34878 44584 34920 44624
rect 34960 44584 34969 44624
rect 49703 44584 49712 44624
rect 49752 44584 49794 44624
rect 49834 44584 49876 44624
rect 49916 44584 49958 44624
rect 49998 44584 50040 44624
rect 50080 44584 50089 44624
rect 64823 44584 64832 44624
rect 64872 44584 64914 44624
rect 64954 44584 64996 44624
rect 65036 44584 65078 44624
rect 65118 44584 65160 44624
rect 65200 44584 65209 44624
rect 79943 44584 79952 44624
rect 79992 44584 80034 44624
rect 80074 44584 80116 44624
rect 80156 44584 80198 44624
rect 80238 44584 80280 44624
rect 80320 44584 80329 44624
rect 95063 44584 95072 44624
rect 95112 44584 95154 44624
rect 95194 44584 95236 44624
rect 95276 44584 95318 44624
rect 95358 44584 95400 44624
rect 95440 44584 95449 44624
rect 3103 43828 3112 43868
rect 3152 43828 3194 43868
rect 3234 43828 3276 43868
rect 3316 43828 3358 43868
rect 3398 43828 3440 43868
rect 3480 43828 3489 43868
rect 18223 43828 18232 43868
rect 18272 43828 18314 43868
rect 18354 43828 18396 43868
rect 18436 43828 18478 43868
rect 18518 43828 18560 43868
rect 18600 43828 18609 43868
rect 33343 43828 33352 43868
rect 33392 43828 33434 43868
rect 33474 43828 33516 43868
rect 33556 43828 33598 43868
rect 33638 43828 33680 43868
rect 33720 43828 33729 43868
rect 48463 43828 48472 43868
rect 48512 43828 48554 43868
rect 48594 43828 48636 43868
rect 48676 43828 48718 43868
rect 48758 43828 48800 43868
rect 48840 43828 48849 43868
rect 63583 43828 63592 43868
rect 63632 43828 63674 43868
rect 63714 43828 63756 43868
rect 63796 43828 63838 43868
rect 63878 43828 63920 43868
rect 63960 43828 63969 43868
rect 78703 43828 78712 43868
rect 78752 43828 78794 43868
rect 78834 43828 78876 43868
rect 78916 43828 78958 43868
rect 78998 43828 79040 43868
rect 79080 43828 79089 43868
rect 93823 43828 93832 43868
rect 93872 43828 93914 43868
rect 93954 43828 93996 43868
rect 94036 43828 94078 43868
rect 94118 43828 94160 43868
rect 94200 43828 94209 43868
rect 0 43280 80 43300
rect 0 43240 652 43280
rect 692 43240 701 43280
rect 0 43220 80 43240
rect 4343 43072 4352 43112
rect 4392 43072 4434 43112
rect 4474 43072 4516 43112
rect 4556 43072 4598 43112
rect 4638 43072 4680 43112
rect 4720 43072 4729 43112
rect 19463 43072 19472 43112
rect 19512 43072 19554 43112
rect 19594 43072 19636 43112
rect 19676 43072 19718 43112
rect 19758 43072 19800 43112
rect 19840 43072 19849 43112
rect 34583 43072 34592 43112
rect 34632 43072 34674 43112
rect 34714 43072 34756 43112
rect 34796 43072 34838 43112
rect 34878 43072 34920 43112
rect 34960 43072 34969 43112
rect 49703 43072 49712 43112
rect 49752 43072 49794 43112
rect 49834 43072 49876 43112
rect 49916 43072 49958 43112
rect 49998 43072 50040 43112
rect 50080 43072 50089 43112
rect 64823 43072 64832 43112
rect 64872 43072 64914 43112
rect 64954 43072 64996 43112
rect 65036 43072 65078 43112
rect 65118 43072 65160 43112
rect 65200 43072 65209 43112
rect 79943 43072 79952 43112
rect 79992 43072 80034 43112
rect 80074 43072 80116 43112
rect 80156 43072 80198 43112
rect 80238 43072 80280 43112
rect 80320 43072 80329 43112
rect 95063 43072 95072 43112
rect 95112 43072 95154 43112
rect 95194 43072 95236 43112
rect 95276 43072 95318 43112
rect 95358 43072 95400 43112
rect 95440 43072 95449 43112
rect 3103 42316 3112 42356
rect 3152 42316 3194 42356
rect 3234 42316 3276 42356
rect 3316 42316 3358 42356
rect 3398 42316 3440 42356
rect 3480 42316 3489 42356
rect 18223 42316 18232 42356
rect 18272 42316 18314 42356
rect 18354 42316 18396 42356
rect 18436 42316 18478 42356
rect 18518 42316 18560 42356
rect 18600 42316 18609 42356
rect 33343 42316 33352 42356
rect 33392 42316 33434 42356
rect 33474 42316 33516 42356
rect 33556 42316 33598 42356
rect 33638 42316 33680 42356
rect 33720 42316 33729 42356
rect 48463 42316 48472 42356
rect 48512 42316 48554 42356
rect 48594 42316 48636 42356
rect 48676 42316 48718 42356
rect 48758 42316 48800 42356
rect 48840 42316 48849 42356
rect 63583 42316 63592 42356
rect 63632 42316 63674 42356
rect 63714 42316 63756 42356
rect 63796 42316 63838 42356
rect 63878 42316 63920 42356
rect 63960 42316 63969 42356
rect 78703 42316 78712 42356
rect 78752 42316 78794 42356
rect 78834 42316 78876 42356
rect 78916 42316 78958 42356
rect 78998 42316 79040 42356
rect 79080 42316 79089 42356
rect 93823 42316 93832 42356
rect 93872 42316 93914 42356
rect 93954 42316 93996 42356
rect 94036 42316 94078 42356
rect 94118 42316 94160 42356
rect 94200 42316 94209 42356
rect 4343 41560 4352 41600
rect 4392 41560 4434 41600
rect 4474 41560 4516 41600
rect 4556 41560 4598 41600
rect 4638 41560 4680 41600
rect 4720 41560 4729 41600
rect 19463 41560 19472 41600
rect 19512 41560 19554 41600
rect 19594 41560 19636 41600
rect 19676 41560 19718 41600
rect 19758 41560 19800 41600
rect 19840 41560 19849 41600
rect 34583 41560 34592 41600
rect 34632 41560 34674 41600
rect 34714 41560 34756 41600
rect 34796 41560 34838 41600
rect 34878 41560 34920 41600
rect 34960 41560 34969 41600
rect 49703 41560 49712 41600
rect 49752 41560 49794 41600
rect 49834 41560 49876 41600
rect 49916 41560 49958 41600
rect 49998 41560 50040 41600
rect 50080 41560 50089 41600
rect 64823 41560 64832 41600
rect 64872 41560 64914 41600
rect 64954 41560 64996 41600
rect 65036 41560 65078 41600
rect 65118 41560 65160 41600
rect 65200 41560 65209 41600
rect 79943 41560 79952 41600
rect 79992 41560 80034 41600
rect 80074 41560 80116 41600
rect 80156 41560 80198 41600
rect 80238 41560 80280 41600
rect 80320 41560 80329 41600
rect 95063 41560 95072 41600
rect 95112 41560 95154 41600
rect 95194 41560 95236 41600
rect 95276 41560 95318 41600
rect 95358 41560 95400 41600
rect 95440 41560 95449 41600
rect 0 41432 80 41452
rect 0 41392 652 41432
rect 692 41392 701 41432
rect 0 41372 80 41392
rect 3103 40804 3112 40844
rect 3152 40804 3194 40844
rect 3234 40804 3276 40844
rect 3316 40804 3358 40844
rect 3398 40804 3440 40844
rect 3480 40804 3489 40844
rect 18223 40804 18232 40844
rect 18272 40804 18314 40844
rect 18354 40804 18396 40844
rect 18436 40804 18478 40844
rect 18518 40804 18560 40844
rect 18600 40804 18609 40844
rect 33343 40804 33352 40844
rect 33392 40804 33434 40844
rect 33474 40804 33516 40844
rect 33556 40804 33598 40844
rect 33638 40804 33680 40844
rect 33720 40804 33729 40844
rect 48463 40804 48472 40844
rect 48512 40804 48554 40844
rect 48594 40804 48636 40844
rect 48676 40804 48718 40844
rect 48758 40804 48800 40844
rect 48840 40804 48849 40844
rect 63583 40804 63592 40844
rect 63632 40804 63674 40844
rect 63714 40804 63756 40844
rect 63796 40804 63838 40844
rect 63878 40804 63920 40844
rect 63960 40804 63969 40844
rect 78703 40804 78712 40844
rect 78752 40804 78794 40844
rect 78834 40804 78876 40844
rect 78916 40804 78958 40844
rect 78998 40804 79040 40844
rect 79080 40804 79089 40844
rect 93823 40804 93832 40844
rect 93872 40804 93914 40844
rect 93954 40804 93996 40844
rect 94036 40804 94078 40844
rect 94118 40804 94160 40844
rect 94200 40804 94209 40844
rect 4343 40048 4352 40088
rect 4392 40048 4434 40088
rect 4474 40048 4516 40088
rect 4556 40048 4598 40088
rect 4638 40048 4680 40088
rect 4720 40048 4729 40088
rect 19463 40048 19472 40088
rect 19512 40048 19554 40088
rect 19594 40048 19636 40088
rect 19676 40048 19718 40088
rect 19758 40048 19800 40088
rect 19840 40048 19849 40088
rect 34583 40048 34592 40088
rect 34632 40048 34674 40088
rect 34714 40048 34756 40088
rect 34796 40048 34838 40088
rect 34878 40048 34920 40088
rect 34960 40048 34969 40088
rect 49703 40048 49712 40088
rect 49752 40048 49794 40088
rect 49834 40048 49876 40088
rect 49916 40048 49958 40088
rect 49998 40048 50040 40088
rect 50080 40048 50089 40088
rect 64823 40048 64832 40088
rect 64872 40048 64914 40088
rect 64954 40048 64996 40088
rect 65036 40048 65078 40088
rect 65118 40048 65160 40088
rect 65200 40048 65209 40088
rect 79943 40048 79952 40088
rect 79992 40048 80034 40088
rect 80074 40048 80116 40088
rect 80156 40048 80198 40088
rect 80238 40048 80280 40088
rect 80320 40048 80329 40088
rect 95063 40048 95072 40088
rect 95112 40048 95154 40088
rect 95194 40048 95236 40088
rect 95276 40048 95318 40088
rect 95358 40048 95400 40088
rect 95440 40048 95449 40088
rect 0 39584 80 39604
rect 0 39544 652 39584
rect 692 39544 701 39584
rect 0 39524 80 39544
rect 3103 39292 3112 39332
rect 3152 39292 3194 39332
rect 3234 39292 3276 39332
rect 3316 39292 3358 39332
rect 3398 39292 3440 39332
rect 3480 39292 3489 39332
rect 18223 39292 18232 39332
rect 18272 39292 18314 39332
rect 18354 39292 18396 39332
rect 18436 39292 18478 39332
rect 18518 39292 18560 39332
rect 18600 39292 18609 39332
rect 33343 39292 33352 39332
rect 33392 39292 33434 39332
rect 33474 39292 33516 39332
rect 33556 39292 33598 39332
rect 33638 39292 33680 39332
rect 33720 39292 33729 39332
rect 48463 39292 48472 39332
rect 48512 39292 48554 39332
rect 48594 39292 48636 39332
rect 48676 39292 48718 39332
rect 48758 39292 48800 39332
rect 48840 39292 48849 39332
rect 63583 39292 63592 39332
rect 63632 39292 63674 39332
rect 63714 39292 63756 39332
rect 63796 39292 63838 39332
rect 63878 39292 63920 39332
rect 63960 39292 63969 39332
rect 78703 39292 78712 39332
rect 78752 39292 78794 39332
rect 78834 39292 78876 39332
rect 78916 39292 78958 39332
rect 78998 39292 79040 39332
rect 79080 39292 79089 39332
rect 93823 39292 93832 39332
rect 93872 39292 93914 39332
rect 93954 39292 93996 39332
rect 94036 39292 94078 39332
rect 94118 39292 94160 39332
rect 94200 39292 94209 39332
rect 4343 38536 4352 38576
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4720 38536 4729 38576
rect 19463 38536 19472 38576
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19840 38536 19849 38576
rect 34583 38536 34592 38576
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34960 38536 34969 38576
rect 49703 38536 49712 38576
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 50080 38536 50089 38576
rect 64823 38536 64832 38576
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 65200 38536 65209 38576
rect 79943 38536 79952 38576
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 80320 38536 80329 38576
rect 95063 38536 95072 38576
rect 95112 38536 95154 38576
rect 95194 38536 95236 38576
rect 95276 38536 95318 38576
rect 95358 38536 95400 38576
rect 95440 38536 95449 38576
rect 3103 37780 3112 37820
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3480 37780 3489 37820
rect 18223 37780 18232 37820
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18600 37780 18609 37820
rect 33343 37780 33352 37820
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33720 37780 33729 37820
rect 48463 37780 48472 37820
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48840 37780 48849 37820
rect 63583 37780 63592 37820
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63960 37780 63969 37820
rect 78703 37780 78712 37820
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 79080 37780 79089 37820
rect 93823 37780 93832 37820
rect 93872 37780 93914 37820
rect 93954 37780 93996 37820
rect 94036 37780 94078 37820
rect 94118 37780 94160 37820
rect 94200 37780 94209 37820
rect 0 37736 80 37756
rect 0 37696 652 37736
rect 692 37696 701 37736
rect 0 37676 80 37696
rect 4343 37024 4352 37064
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4720 37024 4729 37064
rect 19463 37024 19472 37064
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19840 37024 19849 37064
rect 34583 37024 34592 37064
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34960 37024 34969 37064
rect 49703 37024 49712 37064
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 50080 37024 50089 37064
rect 64823 37024 64832 37064
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 65200 37024 65209 37064
rect 79943 37024 79952 37064
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 80320 37024 80329 37064
rect 95063 37024 95072 37064
rect 95112 37024 95154 37064
rect 95194 37024 95236 37064
rect 95276 37024 95318 37064
rect 95358 37024 95400 37064
rect 95440 37024 95449 37064
rect 3103 36268 3112 36308
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3480 36268 3489 36308
rect 18223 36268 18232 36308
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18600 36268 18609 36308
rect 33343 36268 33352 36308
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33720 36268 33729 36308
rect 48463 36268 48472 36308
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48840 36268 48849 36308
rect 63583 36268 63592 36308
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63960 36268 63969 36308
rect 78703 36268 78712 36308
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 79080 36268 79089 36308
rect 93823 36268 93832 36308
rect 93872 36268 93914 36308
rect 93954 36268 93996 36308
rect 94036 36268 94078 36308
rect 94118 36268 94160 36308
rect 94200 36268 94209 36308
rect 0 35888 80 35908
rect 0 35848 652 35888
rect 692 35848 701 35888
rect 0 35828 80 35848
rect 4343 35512 4352 35552
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4720 35512 4729 35552
rect 19463 35512 19472 35552
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19840 35512 19849 35552
rect 34583 35512 34592 35552
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34960 35512 34969 35552
rect 49703 35512 49712 35552
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 50080 35512 50089 35552
rect 64823 35512 64832 35552
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 65200 35512 65209 35552
rect 79943 35512 79952 35552
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 80320 35512 80329 35552
rect 95063 35512 95072 35552
rect 95112 35512 95154 35552
rect 95194 35512 95236 35552
rect 95276 35512 95318 35552
rect 95358 35512 95400 35552
rect 95440 35512 95449 35552
rect 3103 34756 3112 34796
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3480 34756 3489 34796
rect 18223 34756 18232 34796
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18600 34756 18609 34796
rect 33343 34756 33352 34796
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33720 34756 33729 34796
rect 48463 34756 48472 34796
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48840 34756 48849 34796
rect 63583 34756 63592 34796
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63960 34756 63969 34796
rect 78703 34756 78712 34796
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 79080 34756 79089 34796
rect 93823 34756 93832 34796
rect 93872 34756 93914 34796
rect 93954 34756 93996 34796
rect 94036 34756 94078 34796
rect 94118 34756 94160 34796
rect 94200 34756 94209 34796
rect 0 34040 80 34060
rect 0 34000 652 34040
rect 692 34000 701 34040
rect 4343 34000 4352 34040
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4720 34000 4729 34040
rect 19463 34000 19472 34040
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19840 34000 19849 34040
rect 34583 34000 34592 34040
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34960 34000 34969 34040
rect 49703 34000 49712 34040
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 50080 34000 50089 34040
rect 64823 34000 64832 34040
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 65200 34000 65209 34040
rect 79943 34000 79952 34040
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 80320 34000 80329 34040
rect 95063 34000 95072 34040
rect 95112 34000 95154 34040
rect 95194 34000 95236 34040
rect 95276 34000 95318 34040
rect 95358 34000 95400 34040
rect 95440 34000 95449 34040
rect 0 33980 80 34000
rect 3103 33244 3112 33284
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3480 33244 3489 33284
rect 18223 33244 18232 33284
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18600 33244 18609 33284
rect 33343 33244 33352 33284
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33720 33244 33729 33284
rect 48463 33244 48472 33284
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48840 33244 48849 33284
rect 63583 33244 63592 33284
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63960 33244 63969 33284
rect 78703 33244 78712 33284
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 79080 33244 79089 33284
rect 93823 33244 93832 33284
rect 93872 33244 93914 33284
rect 93954 33244 93996 33284
rect 94036 33244 94078 33284
rect 94118 33244 94160 33284
rect 94200 33244 94209 33284
rect 4343 32488 4352 32528
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4720 32488 4729 32528
rect 19463 32488 19472 32528
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19840 32488 19849 32528
rect 34583 32488 34592 32528
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34960 32488 34969 32528
rect 49703 32488 49712 32528
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 50080 32488 50089 32528
rect 64823 32488 64832 32528
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 65200 32488 65209 32528
rect 79943 32488 79952 32528
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 80320 32488 80329 32528
rect 95063 32488 95072 32528
rect 95112 32488 95154 32528
rect 95194 32488 95236 32528
rect 95276 32488 95318 32528
rect 95358 32488 95400 32528
rect 95440 32488 95449 32528
rect 0 32192 80 32212
rect 0 32152 652 32192
rect 692 32152 701 32192
rect 0 32132 80 32152
rect 3103 31732 3112 31772
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3480 31732 3489 31772
rect 18223 31732 18232 31772
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18600 31732 18609 31772
rect 33343 31732 33352 31772
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33720 31732 33729 31772
rect 48463 31732 48472 31772
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48840 31732 48849 31772
rect 63583 31732 63592 31772
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63960 31732 63969 31772
rect 78703 31732 78712 31772
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 79080 31732 79089 31772
rect 93823 31732 93832 31772
rect 93872 31732 93914 31772
rect 93954 31732 93996 31772
rect 94036 31732 94078 31772
rect 94118 31732 94160 31772
rect 94200 31732 94209 31772
rect 4343 30976 4352 31016
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4720 30976 4729 31016
rect 19463 30976 19472 31016
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19840 30976 19849 31016
rect 34583 30976 34592 31016
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34960 30976 34969 31016
rect 49703 30976 49712 31016
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 50080 30976 50089 31016
rect 64823 30976 64832 31016
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 65200 30976 65209 31016
rect 79943 30976 79952 31016
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 80320 30976 80329 31016
rect 95063 30976 95072 31016
rect 95112 30976 95154 31016
rect 95194 30976 95236 31016
rect 95276 30976 95318 31016
rect 95358 30976 95400 31016
rect 95440 30976 95449 31016
rect 0 30344 80 30364
rect 0 30304 652 30344
rect 692 30304 701 30344
rect 0 30284 80 30304
rect 3103 30220 3112 30260
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3480 30220 3489 30260
rect 18223 30220 18232 30260
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18600 30220 18609 30260
rect 33343 30220 33352 30260
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33720 30220 33729 30260
rect 48463 30220 48472 30260
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48840 30220 48849 30260
rect 63583 30220 63592 30260
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63960 30220 63969 30260
rect 78703 30220 78712 30260
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 79080 30220 79089 30260
rect 93823 30220 93832 30260
rect 93872 30220 93914 30260
rect 93954 30220 93996 30260
rect 94036 30220 94078 30260
rect 94118 30220 94160 30260
rect 94200 30220 94209 30260
rect 4343 29464 4352 29504
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4720 29464 4729 29504
rect 19463 29464 19472 29504
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19840 29464 19849 29504
rect 34583 29464 34592 29504
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34960 29464 34969 29504
rect 49703 29464 49712 29504
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 50080 29464 50089 29504
rect 64823 29464 64832 29504
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 65200 29464 65209 29504
rect 79943 29464 79952 29504
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 80320 29464 80329 29504
rect 95063 29464 95072 29504
rect 95112 29464 95154 29504
rect 95194 29464 95236 29504
rect 95276 29464 95318 29504
rect 95358 29464 95400 29504
rect 95440 29464 95449 29504
rect 3103 28708 3112 28748
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3480 28708 3489 28748
rect 18223 28708 18232 28748
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18600 28708 18609 28748
rect 33343 28708 33352 28748
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33720 28708 33729 28748
rect 48463 28708 48472 28748
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48840 28708 48849 28748
rect 63583 28708 63592 28748
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63960 28708 63969 28748
rect 78703 28708 78712 28748
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 79080 28708 79089 28748
rect 93823 28708 93832 28748
rect 93872 28708 93914 28748
rect 93954 28708 93996 28748
rect 94036 28708 94078 28748
rect 94118 28708 94160 28748
rect 94200 28708 94209 28748
rect 0 28496 80 28516
rect 0 28456 652 28496
rect 692 28456 701 28496
rect 0 28436 80 28456
rect 4343 27952 4352 27992
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4720 27952 4729 27992
rect 19463 27952 19472 27992
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19840 27952 19849 27992
rect 34583 27952 34592 27992
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34960 27952 34969 27992
rect 49703 27952 49712 27992
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 50080 27952 50089 27992
rect 64823 27952 64832 27992
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 65200 27952 65209 27992
rect 79943 27952 79952 27992
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 80320 27952 80329 27992
rect 95063 27952 95072 27992
rect 95112 27952 95154 27992
rect 95194 27952 95236 27992
rect 95276 27952 95318 27992
rect 95358 27952 95400 27992
rect 95440 27952 95449 27992
rect 3103 27196 3112 27236
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3480 27196 3489 27236
rect 18223 27196 18232 27236
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18600 27196 18609 27236
rect 33343 27196 33352 27236
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33720 27196 33729 27236
rect 48463 27196 48472 27236
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48840 27196 48849 27236
rect 63583 27196 63592 27236
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63960 27196 63969 27236
rect 78703 27196 78712 27236
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 79080 27196 79089 27236
rect 93823 27196 93832 27236
rect 93872 27196 93914 27236
rect 93954 27196 93996 27236
rect 94036 27196 94078 27236
rect 94118 27196 94160 27236
rect 94200 27196 94209 27236
rect 0 26648 80 26668
rect 0 26608 652 26648
rect 692 26608 701 26648
rect 0 26588 80 26608
rect 4343 26440 4352 26480
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4720 26440 4729 26480
rect 19463 26440 19472 26480
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19840 26440 19849 26480
rect 34583 26440 34592 26480
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34960 26440 34969 26480
rect 49703 26440 49712 26480
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 50080 26440 50089 26480
rect 64823 26440 64832 26480
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 65200 26440 65209 26480
rect 79943 26440 79952 26480
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 80320 26440 80329 26480
rect 95063 26440 95072 26480
rect 95112 26440 95154 26480
rect 95194 26440 95236 26480
rect 95276 26440 95318 26480
rect 95358 26440 95400 26480
rect 95440 26440 95449 26480
rect 3103 25684 3112 25724
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3480 25684 3489 25724
rect 18223 25684 18232 25724
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18600 25684 18609 25724
rect 33343 25684 33352 25724
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33720 25684 33729 25724
rect 48463 25684 48472 25724
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48840 25684 48849 25724
rect 63583 25684 63592 25724
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63960 25684 63969 25724
rect 78703 25684 78712 25724
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 79080 25684 79089 25724
rect 93823 25684 93832 25724
rect 93872 25684 93914 25724
rect 93954 25684 93996 25724
rect 94036 25684 94078 25724
rect 94118 25684 94160 25724
rect 94200 25684 94209 25724
rect 4343 24928 4352 24968
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4720 24928 4729 24968
rect 19463 24928 19472 24968
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19840 24928 19849 24968
rect 34583 24928 34592 24968
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34960 24928 34969 24968
rect 49703 24928 49712 24968
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 50080 24928 50089 24968
rect 64823 24928 64832 24968
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 65200 24928 65209 24968
rect 79943 24928 79952 24968
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 80320 24928 80329 24968
rect 95063 24928 95072 24968
rect 95112 24928 95154 24968
rect 95194 24928 95236 24968
rect 95276 24928 95318 24968
rect 95358 24928 95400 24968
rect 95440 24928 95449 24968
rect 0 24800 80 24820
rect 0 24760 652 24800
rect 692 24760 701 24800
rect 0 24740 80 24760
rect 3103 24172 3112 24212
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3480 24172 3489 24212
rect 18223 24172 18232 24212
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18600 24172 18609 24212
rect 33343 24172 33352 24212
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33720 24172 33729 24212
rect 48463 24172 48472 24212
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48840 24172 48849 24212
rect 63583 24172 63592 24212
rect 63632 24172 63674 24212
rect 63714 24172 63756 24212
rect 63796 24172 63838 24212
rect 63878 24172 63920 24212
rect 63960 24172 63969 24212
rect 78703 24172 78712 24212
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 79080 24172 79089 24212
rect 93823 24172 93832 24212
rect 93872 24172 93914 24212
rect 93954 24172 93996 24212
rect 94036 24172 94078 24212
rect 94118 24172 94160 24212
rect 94200 24172 94209 24212
rect 4343 23416 4352 23456
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4720 23416 4729 23456
rect 19463 23416 19472 23456
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19840 23416 19849 23456
rect 34583 23416 34592 23456
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34960 23416 34969 23456
rect 49703 23416 49712 23456
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 50080 23416 50089 23456
rect 64823 23416 64832 23456
rect 64872 23416 64914 23456
rect 64954 23416 64996 23456
rect 65036 23416 65078 23456
rect 65118 23416 65160 23456
rect 65200 23416 65209 23456
rect 79943 23416 79952 23456
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 80320 23416 80329 23456
rect 95063 23416 95072 23456
rect 95112 23416 95154 23456
rect 95194 23416 95236 23456
rect 95276 23416 95318 23456
rect 95358 23416 95400 23456
rect 95440 23416 95449 23456
rect 0 22952 80 22972
rect 0 22912 652 22952
rect 692 22912 701 22952
rect 0 22892 80 22912
rect 3103 22660 3112 22700
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3480 22660 3489 22700
rect 18223 22660 18232 22700
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18600 22660 18609 22700
rect 33343 22660 33352 22700
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33720 22660 33729 22700
rect 48463 22660 48472 22700
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48840 22660 48849 22700
rect 63583 22660 63592 22700
rect 63632 22660 63674 22700
rect 63714 22660 63756 22700
rect 63796 22660 63838 22700
rect 63878 22660 63920 22700
rect 63960 22660 63969 22700
rect 78703 22660 78712 22700
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 79080 22660 79089 22700
rect 93823 22660 93832 22700
rect 93872 22660 93914 22700
rect 93954 22660 93996 22700
rect 94036 22660 94078 22700
rect 94118 22660 94160 22700
rect 94200 22660 94209 22700
rect 4343 21904 4352 21944
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4720 21904 4729 21944
rect 19463 21904 19472 21944
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19840 21904 19849 21944
rect 34583 21904 34592 21944
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34960 21904 34969 21944
rect 49703 21904 49712 21944
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 50080 21904 50089 21944
rect 64823 21904 64832 21944
rect 64872 21904 64914 21944
rect 64954 21904 64996 21944
rect 65036 21904 65078 21944
rect 65118 21904 65160 21944
rect 65200 21904 65209 21944
rect 79943 21904 79952 21944
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 80320 21904 80329 21944
rect 95063 21904 95072 21944
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95440 21904 95449 21944
rect 3103 21148 3112 21188
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3480 21148 3489 21188
rect 18223 21148 18232 21188
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18600 21148 18609 21188
rect 33343 21148 33352 21188
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33720 21148 33729 21188
rect 48463 21148 48472 21188
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48840 21148 48849 21188
rect 63583 21148 63592 21188
rect 63632 21148 63674 21188
rect 63714 21148 63756 21188
rect 63796 21148 63838 21188
rect 63878 21148 63920 21188
rect 63960 21148 63969 21188
rect 78703 21148 78712 21188
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 79080 21148 79089 21188
rect 93823 21148 93832 21188
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 94200 21148 94209 21188
rect 0 21104 80 21124
rect 0 21064 652 21104
rect 692 21064 701 21104
rect 0 21044 80 21064
rect 4343 20392 4352 20432
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4720 20392 4729 20432
rect 19463 20392 19472 20432
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19840 20392 19849 20432
rect 34583 20392 34592 20432
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34960 20392 34969 20432
rect 49703 20392 49712 20432
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 50080 20392 50089 20432
rect 64823 20392 64832 20432
rect 64872 20392 64914 20432
rect 64954 20392 64996 20432
rect 65036 20392 65078 20432
rect 65118 20392 65160 20432
rect 65200 20392 65209 20432
rect 79943 20392 79952 20432
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 80320 20392 80329 20432
rect 95063 20392 95072 20432
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95440 20392 95449 20432
rect 3103 19636 3112 19676
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3480 19636 3489 19676
rect 18223 19636 18232 19676
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18600 19636 18609 19676
rect 33343 19636 33352 19676
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33720 19636 33729 19676
rect 48463 19636 48472 19676
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48840 19636 48849 19676
rect 63583 19636 63592 19676
rect 63632 19636 63674 19676
rect 63714 19636 63756 19676
rect 63796 19636 63838 19676
rect 63878 19636 63920 19676
rect 63960 19636 63969 19676
rect 78703 19636 78712 19676
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 79080 19636 79089 19676
rect 93823 19636 93832 19676
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 94200 19636 94209 19676
rect 0 19256 80 19276
rect 0 19216 652 19256
rect 692 19216 701 19256
rect 0 19196 80 19216
rect 4343 18880 4352 18920
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4720 18880 4729 18920
rect 19463 18880 19472 18920
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19840 18880 19849 18920
rect 34583 18880 34592 18920
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34960 18880 34969 18920
rect 49703 18880 49712 18920
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 50080 18880 50089 18920
rect 64823 18880 64832 18920
rect 64872 18880 64914 18920
rect 64954 18880 64996 18920
rect 65036 18880 65078 18920
rect 65118 18880 65160 18920
rect 65200 18880 65209 18920
rect 79943 18880 79952 18920
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 80320 18880 80329 18920
rect 95063 18880 95072 18920
rect 95112 18880 95154 18920
rect 95194 18880 95236 18920
rect 95276 18880 95318 18920
rect 95358 18880 95400 18920
rect 95440 18880 95449 18920
rect 3103 18124 3112 18164
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3480 18124 3489 18164
rect 18223 18124 18232 18164
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18600 18124 18609 18164
rect 33343 18124 33352 18164
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33720 18124 33729 18164
rect 48463 18124 48472 18164
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48840 18124 48849 18164
rect 63583 18124 63592 18164
rect 63632 18124 63674 18164
rect 63714 18124 63756 18164
rect 63796 18124 63838 18164
rect 63878 18124 63920 18164
rect 63960 18124 63969 18164
rect 78703 18124 78712 18164
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 79080 18124 79089 18164
rect 93823 18124 93832 18164
rect 93872 18124 93914 18164
rect 93954 18124 93996 18164
rect 94036 18124 94078 18164
rect 94118 18124 94160 18164
rect 94200 18124 94209 18164
rect 0 17408 80 17428
rect 0 17368 652 17408
rect 692 17368 701 17408
rect 4343 17368 4352 17408
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4720 17368 4729 17408
rect 19463 17368 19472 17408
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19840 17368 19849 17408
rect 34583 17368 34592 17408
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34960 17368 34969 17408
rect 49703 17368 49712 17408
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 50080 17368 50089 17408
rect 64823 17368 64832 17408
rect 64872 17368 64914 17408
rect 64954 17368 64996 17408
rect 65036 17368 65078 17408
rect 65118 17368 65160 17408
rect 65200 17368 65209 17408
rect 79943 17368 79952 17408
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 80320 17368 80329 17408
rect 95063 17368 95072 17408
rect 95112 17368 95154 17408
rect 95194 17368 95236 17408
rect 95276 17368 95318 17408
rect 95358 17368 95400 17408
rect 95440 17368 95449 17408
rect 0 17348 80 17368
rect 3103 16612 3112 16652
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3480 16612 3489 16652
rect 18223 16612 18232 16652
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18600 16612 18609 16652
rect 33343 16612 33352 16652
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33720 16612 33729 16652
rect 48463 16612 48472 16652
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48840 16612 48849 16652
rect 63583 16612 63592 16652
rect 63632 16612 63674 16652
rect 63714 16612 63756 16652
rect 63796 16612 63838 16652
rect 63878 16612 63920 16652
rect 63960 16612 63969 16652
rect 78703 16612 78712 16652
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 79080 16612 79089 16652
rect 93823 16612 93832 16652
rect 93872 16612 93914 16652
rect 93954 16612 93996 16652
rect 94036 16612 94078 16652
rect 94118 16612 94160 16652
rect 94200 16612 94209 16652
rect 835 16276 844 16316
rect 884 16276 7084 16316
rect 7124 16276 7133 16316
rect 4343 15856 4352 15896
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4720 15856 4729 15896
rect 19463 15856 19472 15896
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19840 15856 19849 15896
rect 34583 15856 34592 15896
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34960 15856 34969 15896
rect 49703 15856 49712 15896
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 50080 15856 50089 15896
rect 64823 15856 64832 15896
rect 64872 15856 64914 15896
rect 64954 15856 64996 15896
rect 65036 15856 65078 15896
rect 65118 15856 65160 15896
rect 65200 15856 65209 15896
rect 79943 15856 79952 15896
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 80320 15856 80329 15896
rect 95063 15856 95072 15896
rect 95112 15856 95154 15896
rect 95194 15856 95236 15896
rect 95276 15856 95318 15896
rect 95358 15856 95400 15896
rect 95440 15856 95449 15896
rect 0 15560 80 15580
rect 0 15520 652 15560
rect 692 15520 701 15560
rect 0 15500 80 15520
rect 3103 15100 3112 15140
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3480 15100 3489 15140
rect 18223 15100 18232 15140
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18600 15100 18609 15140
rect 33343 15100 33352 15140
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 33720 15100 33729 15140
rect 48463 15100 48472 15140
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48840 15100 48849 15140
rect 63583 15100 63592 15140
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63960 15100 63969 15140
rect 78703 15100 78712 15140
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 79080 15100 79089 15140
rect 93823 15100 93832 15140
rect 93872 15100 93914 15140
rect 93954 15100 93996 15140
rect 94036 15100 94078 15140
rect 94118 15100 94160 15140
rect 94200 15100 94209 15140
rect 4343 14344 4352 14384
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4720 14344 4729 14384
rect 19463 14344 19472 14384
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19840 14344 19849 14384
rect 34583 14344 34592 14384
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34960 14344 34969 14384
rect 49703 14344 49712 14384
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 50080 14344 50089 14384
rect 64823 14344 64832 14384
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 65200 14344 65209 14384
rect 79943 14344 79952 14384
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 80320 14344 80329 14384
rect 95063 14344 95072 14384
rect 95112 14344 95154 14384
rect 95194 14344 95236 14384
rect 95276 14344 95318 14384
rect 95358 14344 95400 14384
rect 95440 14344 95449 14384
rect 643 13756 652 13796
rect 692 13756 701 13796
rect 0 13712 80 13732
rect 652 13712 692 13756
rect 0 13672 692 13712
rect 0 13652 80 13672
rect 3103 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 3489 13628
rect 18223 13588 18232 13628
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18600 13588 18609 13628
rect 33343 13588 33352 13628
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33720 13588 33729 13628
rect 48463 13588 48472 13628
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48840 13588 48849 13628
rect 63583 13588 63592 13628
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63960 13588 63969 13628
rect 78703 13588 78712 13628
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 79080 13588 79089 13628
rect 93823 13588 93832 13628
rect 93872 13588 93914 13628
rect 93954 13588 93996 13628
rect 94036 13588 94078 13628
rect 94118 13588 94160 13628
rect 94200 13588 94209 13628
rect 4343 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 4729 12872
rect 19463 12832 19472 12872
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19840 12832 19849 12872
rect 34583 12832 34592 12872
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34960 12832 34969 12872
rect 49703 12832 49712 12872
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 50080 12832 50089 12872
rect 64823 12832 64832 12872
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 65200 12832 65209 12872
rect 79943 12832 79952 12872
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 80320 12832 80329 12872
rect 95063 12832 95072 12872
rect 95112 12832 95154 12872
rect 95194 12832 95236 12872
rect 95276 12832 95318 12872
rect 95358 12832 95400 12872
rect 95440 12832 95449 12872
rect 835 12412 844 12452
rect 884 12412 1900 12452
rect 1940 12412 1949 12452
rect 3103 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 3489 12116
rect 18223 12076 18232 12116
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18600 12076 18609 12116
rect 33343 12076 33352 12116
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33720 12076 33729 12116
rect 48463 12076 48472 12116
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48840 12076 48849 12116
rect 63583 12076 63592 12116
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63960 12076 63969 12116
rect 78703 12076 78712 12116
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 79080 12076 79089 12116
rect 93823 12076 93832 12116
rect 93872 12076 93914 12116
rect 93954 12076 93996 12116
rect 94036 12076 94078 12116
rect 94118 12076 94160 12116
rect 94200 12076 94209 12116
rect 0 11864 80 11884
rect 0 11824 652 11864
rect 692 11824 701 11864
rect 0 11804 80 11824
rect 4343 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 4729 11360
rect 19463 11320 19472 11360
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19840 11320 19849 11360
rect 34583 11320 34592 11360
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34960 11320 34969 11360
rect 49703 11320 49712 11360
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 50080 11320 50089 11360
rect 64823 11320 64832 11360
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 65200 11320 65209 11360
rect 79943 11320 79952 11360
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 80320 11320 80329 11360
rect 95063 11320 95072 11360
rect 95112 11320 95154 11360
rect 95194 11320 95236 11360
rect 95276 11320 95318 11360
rect 95358 11320 95400 11360
rect 95440 11320 95449 11360
rect 3103 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 3489 10604
rect 18223 10564 18232 10604
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18600 10564 18609 10604
rect 33343 10564 33352 10604
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33720 10564 33729 10604
rect 48463 10564 48472 10604
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48840 10564 48849 10604
rect 63583 10564 63592 10604
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63960 10564 63969 10604
rect 78703 10564 78712 10604
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 79080 10564 79089 10604
rect 93823 10564 93832 10604
rect 93872 10564 93914 10604
rect 93954 10564 93996 10604
rect 94036 10564 94078 10604
rect 94118 10564 94160 10604
rect 94200 10564 94209 10604
rect 835 10228 844 10268
rect 884 10228 6700 10268
rect 6740 10228 6749 10268
rect 0 10016 80 10036
rect 0 9976 652 10016
rect 692 9976 701 10016
rect 0 9956 80 9976
rect 4343 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 4729 9848
rect 19463 9808 19472 9848
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19840 9808 19849 9848
rect 34583 9808 34592 9848
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34960 9808 34969 9848
rect 49703 9808 49712 9848
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 50080 9808 50089 9848
rect 64823 9808 64832 9848
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 65200 9808 65209 9848
rect 79943 9808 79952 9848
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 80320 9808 80329 9848
rect 95063 9808 95072 9848
rect 95112 9808 95154 9848
rect 95194 9808 95236 9848
rect 95276 9808 95318 9848
rect 95358 9808 95400 9848
rect 95440 9808 95449 9848
rect 3103 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 3489 9092
rect 18223 9052 18232 9092
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18600 9052 18609 9092
rect 33343 9052 33352 9092
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33720 9052 33729 9092
rect 48463 9052 48472 9092
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48840 9052 48849 9092
rect 63583 9052 63592 9092
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63960 9052 63969 9092
rect 78703 9052 78712 9092
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 79080 9052 79089 9092
rect 93823 9052 93832 9092
rect 93872 9052 93914 9092
rect 93954 9052 93996 9092
rect 94036 9052 94078 9092
rect 94118 9052 94160 9092
rect 94200 9052 94209 9092
rect 835 8716 844 8756
rect 884 8716 5644 8756
rect 5684 8716 5693 8756
rect 4343 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 4729 8336
rect 19463 8296 19472 8336
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19840 8296 19849 8336
rect 34583 8296 34592 8336
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34960 8296 34969 8336
rect 49703 8296 49712 8336
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 50080 8296 50089 8336
rect 64823 8296 64832 8336
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 65200 8296 65209 8336
rect 79943 8296 79952 8336
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 80320 8296 80329 8336
rect 95063 8296 95072 8336
rect 95112 8296 95154 8336
rect 95194 8296 95236 8336
rect 95276 8296 95318 8336
rect 95358 8296 95400 8336
rect 95440 8296 95449 8336
rect 0 8168 80 8188
rect 0 8128 652 8168
rect 692 8128 701 8168
rect 0 8108 80 8128
rect 3103 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 3489 7580
rect 18223 7540 18232 7580
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18600 7540 18609 7580
rect 33343 7540 33352 7580
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33720 7540 33729 7580
rect 48463 7540 48472 7580
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48840 7540 48849 7580
rect 63583 7540 63592 7580
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63960 7540 63969 7580
rect 78703 7540 78712 7580
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 79080 7540 79089 7580
rect 93823 7540 93832 7580
rect 93872 7540 93914 7580
rect 93954 7540 93996 7580
rect 94036 7540 94078 7580
rect 94118 7540 94160 7580
rect 94200 7540 94209 7580
rect 4343 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 4729 6824
rect 19463 6784 19472 6824
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19840 6784 19849 6824
rect 34583 6784 34592 6824
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34960 6784 34969 6824
rect 49703 6784 49712 6824
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 50080 6784 50089 6824
rect 64823 6784 64832 6824
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 65200 6784 65209 6824
rect 79943 6784 79952 6824
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 80320 6784 80329 6824
rect 95063 6784 95072 6824
rect 95112 6784 95154 6824
rect 95194 6784 95236 6824
rect 95276 6784 95318 6824
rect 95358 6784 95400 6824
rect 95440 6784 95449 6824
rect 0 6320 80 6340
rect 0 6280 652 6320
rect 692 6280 701 6320
rect 0 6260 80 6280
rect 3103 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 3489 6068
rect 18223 6028 18232 6068
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18600 6028 18609 6068
rect 33343 6028 33352 6068
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33720 6028 33729 6068
rect 48463 6028 48472 6068
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48840 6028 48849 6068
rect 63583 6028 63592 6068
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63960 6028 63969 6068
rect 78703 6028 78712 6068
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 79080 6028 79089 6068
rect 93823 6028 93832 6068
rect 93872 6028 93914 6068
rect 93954 6028 93996 6068
rect 94036 6028 94078 6068
rect 94118 6028 94160 6068
rect 94200 6028 94209 6068
rect 4343 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 4729 5312
rect 19463 5272 19472 5312
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19840 5272 19849 5312
rect 34583 5272 34592 5312
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34960 5272 34969 5312
rect 49703 5272 49712 5312
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 50080 5272 50089 5312
rect 64823 5272 64832 5312
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 65200 5272 65209 5312
rect 79943 5272 79952 5312
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 80320 5272 80329 5312
rect 95063 5272 95072 5312
rect 95112 5272 95154 5312
rect 95194 5272 95236 5312
rect 95276 5272 95318 5312
rect 95358 5272 95400 5312
rect 95440 5272 95449 5312
rect 835 4852 844 4892
rect 884 4852 14476 4892
rect 14516 4852 14525 4892
rect 3103 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 3489 4556
rect 18223 4516 18232 4556
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18600 4516 18609 4556
rect 33343 4516 33352 4556
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33720 4516 33729 4556
rect 48463 4516 48472 4556
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48840 4516 48849 4556
rect 63583 4516 63592 4556
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63960 4516 63969 4556
rect 78703 4516 78712 4556
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 79080 4516 79089 4556
rect 93823 4516 93832 4556
rect 93872 4516 93914 4556
rect 93954 4516 93996 4556
rect 94036 4516 94078 4556
rect 94118 4516 94160 4556
rect 94200 4516 94209 4556
rect 0 4472 80 4492
rect 0 4432 652 4472
rect 692 4432 701 4472
rect 0 4412 80 4432
rect 4343 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 4729 3800
rect 19463 3760 19472 3800
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19840 3760 19849 3800
rect 34583 3760 34592 3800
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34960 3760 34969 3800
rect 49703 3760 49712 3800
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 50080 3760 50089 3800
rect 64823 3760 64832 3800
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 65200 3760 65209 3800
rect 79943 3760 79952 3800
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 80320 3760 80329 3800
rect 95063 3760 95072 3800
rect 95112 3760 95154 3800
rect 95194 3760 95236 3800
rect 95276 3760 95318 3800
rect 95358 3760 95400 3800
rect 95440 3760 95449 3800
rect 3103 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 3489 3044
rect 18223 3004 18232 3044
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18600 3004 18609 3044
rect 33343 3004 33352 3044
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33720 3004 33729 3044
rect 48463 3004 48472 3044
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48840 3004 48849 3044
rect 63583 3004 63592 3044
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63960 3004 63969 3044
rect 78703 3004 78712 3044
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 79080 3004 79089 3044
rect 93823 3004 93832 3044
rect 93872 3004 93914 3044
rect 93954 3004 93996 3044
rect 94036 3004 94078 3044
rect 94118 3004 94160 3044
rect 94200 3004 94209 3044
rect 0 2624 80 2644
rect 0 2584 652 2624
rect 692 2584 701 2624
rect 0 2564 80 2584
rect 4343 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 4729 2288
rect 19463 2248 19472 2288
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19840 2248 19849 2288
rect 34583 2248 34592 2288
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34960 2248 34969 2288
rect 49703 2248 49712 2288
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 50080 2248 50089 2288
rect 64823 2248 64832 2288
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 65200 2248 65209 2288
rect 79943 2248 79952 2288
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 80320 2248 80329 2288
rect 95063 2248 95072 2288
rect 95112 2248 95154 2288
rect 95194 2248 95236 2288
rect 95276 2248 95318 2288
rect 95358 2248 95400 2288
rect 95440 2248 95449 2288
rect 3103 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 3489 1532
rect 18223 1492 18232 1532
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18600 1492 18609 1532
rect 33343 1492 33352 1532
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33720 1492 33729 1532
rect 48463 1492 48472 1532
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48840 1492 48849 1532
rect 63583 1492 63592 1532
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63960 1492 63969 1532
rect 78703 1492 78712 1532
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 79080 1492 79089 1532
rect 93823 1492 93832 1532
rect 93872 1492 93914 1532
rect 93954 1492 93996 1532
rect 94036 1492 94078 1532
rect 94118 1492 94160 1532
rect 94200 1492 94209 1532
rect 4343 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 4729 776
rect 19463 736 19472 776
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19840 736 19849 776
rect 34583 736 34592 776
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34960 736 34969 776
rect 49703 736 49712 776
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 50080 736 50089 776
rect 64823 736 64832 776
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 65200 736 65209 776
rect 79943 736 79952 776
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 80320 736 80329 776
rect 95063 736 95072 776
rect 95112 736 95154 776
rect 95194 736 95236 776
rect 95276 736 95318 776
rect 95358 736 95400 776
rect 95440 736 95449 776
<< via3 >>
rect 3112 81628 3152 81668
rect 3194 81628 3234 81668
rect 3276 81628 3316 81668
rect 3358 81628 3398 81668
rect 3440 81628 3480 81668
rect 18232 81628 18272 81668
rect 18314 81628 18354 81668
rect 18396 81628 18436 81668
rect 18478 81628 18518 81668
rect 18560 81628 18600 81668
rect 33352 81628 33392 81668
rect 33434 81628 33474 81668
rect 33516 81628 33556 81668
rect 33598 81628 33638 81668
rect 33680 81628 33720 81668
rect 48472 81628 48512 81668
rect 48554 81628 48594 81668
rect 48636 81628 48676 81668
rect 48718 81628 48758 81668
rect 48800 81628 48840 81668
rect 63592 81628 63632 81668
rect 63674 81628 63714 81668
rect 63756 81628 63796 81668
rect 63838 81628 63878 81668
rect 63920 81628 63960 81668
rect 78712 81628 78752 81668
rect 78794 81628 78834 81668
rect 78876 81628 78916 81668
rect 78958 81628 78998 81668
rect 79040 81628 79080 81668
rect 93832 81628 93872 81668
rect 93914 81628 93954 81668
rect 93996 81628 94036 81668
rect 94078 81628 94118 81668
rect 94160 81628 94200 81668
rect 4352 80872 4392 80912
rect 4434 80872 4474 80912
rect 4516 80872 4556 80912
rect 4598 80872 4638 80912
rect 4680 80872 4720 80912
rect 19472 80872 19512 80912
rect 19554 80872 19594 80912
rect 19636 80872 19676 80912
rect 19718 80872 19758 80912
rect 19800 80872 19840 80912
rect 34592 80872 34632 80912
rect 34674 80872 34714 80912
rect 34756 80872 34796 80912
rect 34838 80872 34878 80912
rect 34920 80872 34960 80912
rect 49712 80872 49752 80912
rect 49794 80872 49834 80912
rect 49876 80872 49916 80912
rect 49958 80872 49998 80912
rect 50040 80872 50080 80912
rect 64832 80872 64872 80912
rect 64914 80872 64954 80912
rect 64996 80872 65036 80912
rect 65078 80872 65118 80912
rect 65160 80872 65200 80912
rect 79952 80872 79992 80912
rect 80034 80872 80074 80912
rect 80116 80872 80156 80912
rect 80198 80872 80238 80912
rect 80280 80872 80320 80912
rect 95072 80872 95112 80912
rect 95154 80872 95194 80912
rect 95236 80872 95276 80912
rect 95318 80872 95358 80912
rect 95400 80872 95440 80912
rect 3112 80116 3152 80156
rect 3194 80116 3234 80156
rect 3276 80116 3316 80156
rect 3358 80116 3398 80156
rect 3440 80116 3480 80156
rect 18232 80116 18272 80156
rect 18314 80116 18354 80156
rect 18396 80116 18436 80156
rect 18478 80116 18518 80156
rect 18560 80116 18600 80156
rect 33352 80116 33392 80156
rect 33434 80116 33474 80156
rect 33516 80116 33556 80156
rect 33598 80116 33638 80156
rect 33680 80116 33720 80156
rect 48472 80116 48512 80156
rect 48554 80116 48594 80156
rect 48636 80116 48676 80156
rect 48718 80116 48758 80156
rect 48800 80116 48840 80156
rect 63592 80116 63632 80156
rect 63674 80116 63714 80156
rect 63756 80116 63796 80156
rect 63838 80116 63878 80156
rect 63920 80116 63960 80156
rect 78712 80116 78752 80156
rect 78794 80116 78834 80156
rect 78876 80116 78916 80156
rect 78958 80116 78998 80156
rect 79040 80116 79080 80156
rect 93832 80116 93872 80156
rect 93914 80116 93954 80156
rect 93996 80116 94036 80156
rect 94078 80116 94118 80156
rect 94160 80116 94200 80156
rect 4352 79360 4392 79400
rect 4434 79360 4474 79400
rect 4516 79360 4556 79400
rect 4598 79360 4638 79400
rect 4680 79360 4720 79400
rect 19472 79360 19512 79400
rect 19554 79360 19594 79400
rect 19636 79360 19676 79400
rect 19718 79360 19758 79400
rect 19800 79360 19840 79400
rect 34592 79360 34632 79400
rect 34674 79360 34714 79400
rect 34756 79360 34796 79400
rect 34838 79360 34878 79400
rect 34920 79360 34960 79400
rect 49712 79360 49752 79400
rect 49794 79360 49834 79400
rect 49876 79360 49916 79400
rect 49958 79360 49998 79400
rect 50040 79360 50080 79400
rect 64832 79360 64872 79400
rect 64914 79360 64954 79400
rect 64996 79360 65036 79400
rect 65078 79360 65118 79400
rect 65160 79360 65200 79400
rect 79952 79360 79992 79400
rect 80034 79360 80074 79400
rect 80116 79360 80156 79400
rect 80198 79360 80238 79400
rect 80280 79360 80320 79400
rect 95072 79360 95112 79400
rect 95154 79360 95194 79400
rect 95236 79360 95276 79400
rect 95318 79360 95358 79400
rect 95400 79360 95440 79400
rect 3112 78604 3152 78644
rect 3194 78604 3234 78644
rect 3276 78604 3316 78644
rect 3358 78604 3398 78644
rect 3440 78604 3480 78644
rect 18232 78604 18272 78644
rect 18314 78604 18354 78644
rect 18396 78604 18436 78644
rect 18478 78604 18518 78644
rect 18560 78604 18600 78644
rect 33352 78604 33392 78644
rect 33434 78604 33474 78644
rect 33516 78604 33556 78644
rect 33598 78604 33638 78644
rect 33680 78604 33720 78644
rect 48472 78604 48512 78644
rect 48554 78604 48594 78644
rect 48636 78604 48676 78644
rect 48718 78604 48758 78644
rect 48800 78604 48840 78644
rect 63592 78604 63632 78644
rect 63674 78604 63714 78644
rect 63756 78604 63796 78644
rect 63838 78604 63878 78644
rect 63920 78604 63960 78644
rect 78712 78604 78752 78644
rect 78794 78604 78834 78644
rect 78876 78604 78916 78644
rect 78958 78604 78998 78644
rect 79040 78604 79080 78644
rect 93832 78604 93872 78644
rect 93914 78604 93954 78644
rect 93996 78604 94036 78644
rect 94078 78604 94118 78644
rect 94160 78604 94200 78644
rect 4352 77848 4392 77888
rect 4434 77848 4474 77888
rect 4516 77848 4556 77888
rect 4598 77848 4638 77888
rect 4680 77848 4720 77888
rect 19472 77848 19512 77888
rect 19554 77848 19594 77888
rect 19636 77848 19676 77888
rect 19718 77848 19758 77888
rect 19800 77848 19840 77888
rect 34592 77848 34632 77888
rect 34674 77848 34714 77888
rect 34756 77848 34796 77888
rect 34838 77848 34878 77888
rect 34920 77848 34960 77888
rect 49712 77848 49752 77888
rect 49794 77848 49834 77888
rect 49876 77848 49916 77888
rect 49958 77848 49998 77888
rect 50040 77848 50080 77888
rect 64832 77848 64872 77888
rect 64914 77848 64954 77888
rect 64996 77848 65036 77888
rect 65078 77848 65118 77888
rect 65160 77848 65200 77888
rect 79952 77848 79992 77888
rect 80034 77848 80074 77888
rect 80116 77848 80156 77888
rect 80198 77848 80238 77888
rect 80280 77848 80320 77888
rect 95072 77848 95112 77888
rect 95154 77848 95194 77888
rect 95236 77848 95276 77888
rect 95318 77848 95358 77888
rect 95400 77848 95440 77888
rect 3112 77092 3152 77132
rect 3194 77092 3234 77132
rect 3276 77092 3316 77132
rect 3358 77092 3398 77132
rect 3440 77092 3480 77132
rect 18232 77092 18272 77132
rect 18314 77092 18354 77132
rect 18396 77092 18436 77132
rect 18478 77092 18518 77132
rect 18560 77092 18600 77132
rect 33352 77092 33392 77132
rect 33434 77092 33474 77132
rect 33516 77092 33556 77132
rect 33598 77092 33638 77132
rect 33680 77092 33720 77132
rect 48472 77092 48512 77132
rect 48554 77092 48594 77132
rect 48636 77092 48676 77132
rect 48718 77092 48758 77132
rect 48800 77092 48840 77132
rect 63592 77092 63632 77132
rect 63674 77092 63714 77132
rect 63756 77092 63796 77132
rect 63838 77092 63878 77132
rect 63920 77092 63960 77132
rect 78712 77092 78752 77132
rect 78794 77092 78834 77132
rect 78876 77092 78916 77132
rect 78958 77092 78998 77132
rect 79040 77092 79080 77132
rect 93832 77092 93872 77132
rect 93914 77092 93954 77132
rect 93996 77092 94036 77132
rect 94078 77092 94118 77132
rect 94160 77092 94200 77132
rect 4352 76336 4392 76376
rect 4434 76336 4474 76376
rect 4516 76336 4556 76376
rect 4598 76336 4638 76376
rect 4680 76336 4720 76376
rect 19472 76336 19512 76376
rect 19554 76336 19594 76376
rect 19636 76336 19676 76376
rect 19718 76336 19758 76376
rect 19800 76336 19840 76376
rect 34592 76336 34632 76376
rect 34674 76336 34714 76376
rect 34756 76336 34796 76376
rect 34838 76336 34878 76376
rect 34920 76336 34960 76376
rect 49712 76336 49752 76376
rect 49794 76336 49834 76376
rect 49876 76336 49916 76376
rect 49958 76336 49998 76376
rect 50040 76336 50080 76376
rect 64832 76336 64872 76376
rect 64914 76336 64954 76376
rect 64996 76336 65036 76376
rect 65078 76336 65118 76376
rect 65160 76336 65200 76376
rect 79952 76336 79992 76376
rect 80034 76336 80074 76376
rect 80116 76336 80156 76376
rect 80198 76336 80238 76376
rect 80280 76336 80320 76376
rect 95072 76336 95112 76376
rect 95154 76336 95194 76376
rect 95236 76336 95276 76376
rect 95318 76336 95358 76376
rect 95400 76336 95440 76376
rect 3112 75580 3152 75620
rect 3194 75580 3234 75620
rect 3276 75580 3316 75620
rect 3358 75580 3398 75620
rect 3440 75580 3480 75620
rect 18232 75580 18272 75620
rect 18314 75580 18354 75620
rect 18396 75580 18436 75620
rect 18478 75580 18518 75620
rect 18560 75580 18600 75620
rect 33352 75580 33392 75620
rect 33434 75580 33474 75620
rect 33516 75580 33556 75620
rect 33598 75580 33638 75620
rect 33680 75580 33720 75620
rect 48472 75580 48512 75620
rect 48554 75580 48594 75620
rect 48636 75580 48676 75620
rect 48718 75580 48758 75620
rect 48800 75580 48840 75620
rect 63592 75580 63632 75620
rect 63674 75580 63714 75620
rect 63756 75580 63796 75620
rect 63838 75580 63878 75620
rect 63920 75580 63960 75620
rect 78712 75580 78752 75620
rect 78794 75580 78834 75620
rect 78876 75580 78916 75620
rect 78958 75580 78998 75620
rect 79040 75580 79080 75620
rect 93832 75580 93872 75620
rect 93914 75580 93954 75620
rect 93996 75580 94036 75620
rect 94078 75580 94118 75620
rect 94160 75580 94200 75620
rect 4352 74824 4392 74864
rect 4434 74824 4474 74864
rect 4516 74824 4556 74864
rect 4598 74824 4638 74864
rect 4680 74824 4720 74864
rect 19472 74824 19512 74864
rect 19554 74824 19594 74864
rect 19636 74824 19676 74864
rect 19718 74824 19758 74864
rect 19800 74824 19840 74864
rect 34592 74824 34632 74864
rect 34674 74824 34714 74864
rect 34756 74824 34796 74864
rect 34838 74824 34878 74864
rect 34920 74824 34960 74864
rect 49712 74824 49752 74864
rect 49794 74824 49834 74864
rect 49876 74824 49916 74864
rect 49958 74824 49998 74864
rect 50040 74824 50080 74864
rect 64832 74824 64872 74864
rect 64914 74824 64954 74864
rect 64996 74824 65036 74864
rect 65078 74824 65118 74864
rect 65160 74824 65200 74864
rect 79952 74824 79992 74864
rect 80034 74824 80074 74864
rect 80116 74824 80156 74864
rect 80198 74824 80238 74864
rect 80280 74824 80320 74864
rect 95072 74824 95112 74864
rect 95154 74824 95194 74864
rect 95236 74824 95276 74864
rect 95318 74824 95358 74864
rect 95400 74824 95440 74864
rect 3112 74068 3152 74108
rect 3194 74068 3234 74108
rect 3276 74068 3316 74108
rect 3358 74068 3398 74108
rect 3440 74068 3480 74108
rect 18232 74068 18272 74108
rect 18314 74068 18354 74108
rect 18396 74068 18436 74108
rect 18478 74068 18518 74108
rect 18560 74068 18600 74108
rect 33352 74068 33392 74108
rect 33434 74068 33474 74108
rect 33516 74068 33556 74108
rect 33598 74068 33638 74108
rect 33680 74068 33720 74108
rect 48472 74068 48512 74108
rect 48554 74068 48594 74108
rect 48636 74068 48676 74108
rect 48718 74068 48758 74108
rect 48800 74068 48840 74108
rect 63592 74068 63632 74108
rect 63674 74068 63714 74108
rect 63756 74068 63796 74108
rect 63838 74068 63878 74108
rect 63920 74068 63960 74108
rect 78712 74068 78752 74108
rect 78794 74068 78834 74108
rect 78876 74068 78916 74108
rect 78958 74068 78998 74108
rect 79040 74068 79080 74108
rect 93832 74068 93872 74108
rect 93914 74068 93954 74108
rect 93996 74068 94036 74108
rect 94078 74068 94118 74108
rect 94160 74068 94200 74108
rect 4352 73312 4392 73352
rect 4434 73312 4474 73352
rect 4516 73312 4556 73352
rect 4598 73312 4638 73352
rect 4680 73312 4720 73352
rect 19472 73312 19512 73352
rect 19554 73312 19594 73352
rect 19636 73312 19676 73352
rect 19718 73312 19758 73352
rect 19800 73312 19840 73352
rect 34592 73312 34632 73352
rect 34674 73312 34714 73352
rect 34756 73312 34796 73352
rect 34838 73312 34878 73352
rect 34920 73312 34960 73352
rect 49712 73312 49752 73352
rect 49794 73312 49834 73352
rect 49876 73312 49916 73352
rect 49958 73312 49998 73352
rect 50040 73312 50080 73352
rect 64832 73312 64872 73352
rect 64914 73312 64954 73352
rect 64996 73312 65036 73352
rect 65078 73312 65118 73352
rect 65160 73312 65200 73352
rect 79952 73312 79992 73352
rect 80034 73312 80074 73352
rect 80116 73312 80156 73352
rect 80198 73312 80238 73352
rect 80280 73312 80320 73352
rect 95072 73312 95112 73352
rect 95154 73312 95194 73352
rect 95236 73312 95276 73352
rect 95318 73312 95358 73352
rect 95400 73312 95440 73352
rect 3112 72556 3152 72596
rect 3194 72556 3234 72596
rect 3276 72556 3316 72596
rect 3358 72556 3398 72596
rect 3440 72556 3480 72596
rect 18232 72556 18272 72596
rect 18314 72556 18354 72596
rect 18396 72556 18436 72596
rect 18478 72556 18518 72596
rect 18560 72556 18600 72596
rect 33352 72556 33392 72596
rect 33434 72556 33474 72596
rect 33516 72556 33556 72596
rect 33598 72556 33638 72596
rect 33680 72556 33720 72596
rect 48472 72556 48512 72596
rect 48554 72556 48594 72596
rect 48636 72556 48676 72596
rect 48718 72556 48758 72596
rect 48800 72556 48840 72596
rect 63592 72556 63632 72596
rect 63674 72556 63714 72596
rect 63756 72556 63796 72596
rect 63838 72556 63878 72596
rect 63920 72556 63960 72596
rect 78712 72556 78752 72596
rect 78794 72556 78834 72596
rect 78876 72556 78916 72596
rect 78958 72556 78998 72596
rect 79040 72556 79080 72596
rect 93832 72556 93872 72596
rect 93914 72556 93954 72596
rect 93996 72556 94036 72596
rect 94078 72556 94118 72596
rect 94160 72556 94200 72596
rect 4352 71800 4392 71840
rect 4434 71800 4474 71840
rect 4516 71800 4556 71840
rect 4598 71800 4638 71840
rect 4680 71800 4720 71840
rect 19472 71800 19512 71840
rect 19554 71800 19594 71840
rect 19636 71800 19676 71840
rect 19718 71800 19758 71840
rect 19800 71800 19840 71840
rect 34592 71800 34632 71840
rect 34674 71800 34714 71840
rect 34756 71800 34796 71840
rect 34838 71800 34878 71840
rect 34920 71800 34960 71840
rect 49712 71800 49752 71840
rect 49794 71800 49834 71840
rect 49876 71800 49916 71840
rect 49958 71800 49998 71840
rect 50040 71800 50080 71840
rect 64832 71800 64872 71840
rect 64914 71800 64954 71840
rect 64996 71800 65036 71840
rect 65078 71800 65118 71840
rect 65160 71800 65200 71840
rect 79952 71800 79992 71840
rect 80034 71800 80074 71840
rect 80116 71800 80156 71840
rect 80198 71800 80238 71840
rect 80280 71800 80320 71840
rect 95072 71800 95112 71840
rect 95154 71800 95194 71840
rect 95236 71800 95276 71840
rect 95318 71800 95358 71840
rect 95400 71800 95440 71840
rect 3112 71044 3152 71084
rect 3194 71044 3234 71084
rect 3276 71044 3316 71084
rect 3358 71044 3398 71084
rect 3440 71044 3480 71084
rect 18232 71044 18272 71084
rect 18314 71044 18354 71084
rect 18396 71044 18436 71084
rect 18478 71044 18518 71084
rect 18560 71044 18600 71084
rect 33352 71044 33392 71084
rect 33434 71044 33474 71084
rect 33516 71044 33556 71084
rect 33598 71044 33638 71084
rect 33680 71044 33720 71084
rect 48472 71044 48512 71084
rect 48554 71044 48594 71084
rect 48636 71044 48676 71084
rect 48718 71044 48758 71084
rect 48800 71044 48840 71084
rect 63592 71044 63632 71084
rect 63674 71044 63714 71084
rect 63756 71044 63796 71084
rect 63838 71044 63878 71084
rect 63920 71044 63960 71084
rect 78712 71044 78752 71084
rect 78794 71044 78834 71084
rect 78876 71044 78916 71084
rect 78958 71044 78998 71084
rect 79040 71044 79080 71084
rect 93832 71044 93872 71084
rect 93914 71044 93954 71084
rect 93996 71044 94036 71084
rect 94078 71044 94118 71084
rect 94160 71044 94200 71084
rect 4352 70288 4392 70328
rect 4434 70288 4474 70328
rect 4516 70288 4556 70328
rect 4598 70288 4638 70328
rect 4680 70288 4720 70328
rect 19472 70288 19512 70328
rect 19554 70288 19594 70328
rect 19636 70288 19676 70328
rect 19718 70288 19758 70328
rect 19800 70288 19840 70328
rect 34592 70288 34632 70328
rect 34674 70288 34714 70328
rect 34756 70288 34796 70328
rect 34838 70288 34878 70328
rect 34920 70288 34960 70328
rect 49712 70288 49752 70328
rect 49794 70288 49834 70328
rect 49876 70288 49916 70328
rect 49958 70288 49998 70328
rect 50040 70288 50080 70328
rect 64832 70288 64872 70328
rect 64914 70288 64954 70328
rect 64996 70288 65036 70328
rect 65078 70288 65118 70328
rect 65160 70288 65200 70328
rect 79952 70288 79992 70328
rect 80034 70288 80074 70328
rect 80116 70288 80156 70328
rect 80198 70288 80238 70328
rect 80280 70288 80320 70328
rect 95072 70288 95112 70328
rect 95154 70288 95194 70328
rect 95236 70288 95276 70328
rect 95318 70288 95358 70328
rect 95400 70288 95440 70328
rect 3112 69532 3152 69572
rect 3194 69532 3234 69572
rect 3276 69532 3316 69572
rect 3358 69532 3398 69572
rect 3440 69532 3480 69572
rect 18232 69532 18272 69572
rect 18314 69532 18354 69572
rect 18396 69532 18436 69572
rect 18478 69532 18518 69572
rect 18560 69532 18600 69572
rect 33352 69532 33392 69572
rect 33434 69532 33474 69572
rect 33516 69532 33556 69572
rect 33598 69532 33638 69572
rect 33680 69532 33720 69572
rect 48472 69532 48512 69572
rect 48554 69532 48594 69572
rect 48636 69532 48676 69572
rect 48718 69532 48758 69572
rect 48800 69532 48840 69572
rect 63592 69532 63632 69572
rect 63674 69532 63714 69572
rect 63756 69532 63796 69572
rect 63838 69532 63878 69572
rect 63920 69532 63960 69572
rect 78712 69532 78752 69572
rect 78794 69532 78834 69572
rect 78876 69532 78916 69572
rect 78958 69532 78998 69572
rect 79040 69532 79080 69572
rect 93832 69532 93872 69572
rect 93914 69532 93954 69572
rect 93996 69532 94036 69572
rect 94078 69532 94118 69572
rect 94160 69532 94200 69572
rect 4352 68776 4392 68816
rect 4434 68776 4474 68816
rect 4516 68776 4556 68816
rect 4598 68776 4638 68816
rect 4680 68776 4720 68816
rect 19472 68776 19512 68816
rect 19554 68776 19594 68816
rect 19636 68776 19676 68816
rect 19718 68776 19758 68816
rect 19800 68776 19840 68816
rect 34592 68776 34632 68816
rect 34674 68776 34714 68816
rect 34756 68776 34796 68816
rect 34838 68776 34878 68816
rect 34920 68776 34960 68816
rect 49712 68776 49752 68816
rect 49794 68776 49834 68816
rect 49876 68776 49916 68816
rect 49958 68776 49998 68816
rect 50040 68776 50080 68816
rect 64832 68776 64872 68816
rect 64914 68776 64954 68816
rect 64996 68776 65036 68816
rect 65078 68776 65118 68816
rect 65160 68776 65200 68816
rect 79952 68776 79992 68816
rect 80034 68776 80074 68816
rect 80116 68776 80156 68816
rect 80198 68776 80238 68816
rect 80280 68776 80320 68816
rect 95072 68776 95112 68816
rect 95154 68776 95194 68816
rect 95236 68776 95276 68816
rect 95318 68776 95358 68816
rect 95400 68776 95440 68816
rect 3112 68020 3152 68060
rect 3194 68020 3234 68060
rect 3276 68020 3316 68060
rect 3358 68020 3398 68060
rect 3440 68020 3480 68060
rect 18232 68020 18272 68060
rect 18314 68020 18354 68060
rect 18396 68020 18436 68060
rect 18478 68020 18518 68060
rect 18560 68020 18600 68060
rect 33352 68020 33392 68060
rect 33434 68020 33474 68060
rect 33516 68020 33556 68060
rect 33598 68020 33638 68060
rect 33680 68020 33720 68060
rect 48472 68020 48512 68060
rect 48554 68020 48594 68060
rect 48636 68020 48676 68060
rect 48718 68020 48758 68060
rect 48800 68020 48840 68060
rect 63592 68020 63632 68060
rect 63674 68020 63714 68060
rect 63756 68020 63796 68060
rect 63838 68020 63878 68060
rect 63920 68020 63960 68060
rect 78712 68020 78752 68060
rect 78794 68020 78834 68060
rect 78876 68020 78916 68060
rect 78958 68020 78998 68060
rect 79040 68020 79080 68060
rect 93832 68020 93872 68060
rect 93914 68020 93954 68060
rect 93996 68020 94036 68060
rect 94078 68020 94118 68060
rect 94160 68020 94200 68060
rect 4352 67264 4392 67304
rect 4434 67264 4474 67304
rect 4516 67264 4556 67304
rect 4598 67264 4638 67304
rect 4680 67264 4720 67304
rect 19472 67264 19512 67304
rect 19554 67264 19594 67304
rect 19636 67264 19676 67304
rect 19718 67264 19758 67304
rect 19800 67264 19840 67304
rect 34592 67264 34632 67304
rect 34674 67264 34714 67304
rect 34756 67264 34796 67304
rect 34838 67264 34878 67304
rect 34920 67264 34960 67304
rect 49712 67264 49752 67304
rect 49794 67264 49834 67304
rect 49876 67264 49916 67304
rect 49958 67264 49998 67304
rect 50040 67264 50080 67304
rect 64832 67264 64872 67304
rect 64914 67264 64954 67304
rect 64996 67264 65036 67304
rect 65078 67264 65118 67304
rect 65160 67264 65200 67304
rect 79952 67264 79992 67304
rect 80034 67264 80074 67304
rect 80116 67264 80156 67304
rect 80198 67264 80238 67304
rect 80280 67264 80320 67304
rect 95072 67264 95112 67304
rect 95154 67264 95194 67304
rect 95236 67264 95276 67304
rect 95318 67264 95358 67304
rect 95400 67264 95440 67304
rect 3112 66508 3152 66548
rect 3194 66508 3234 66548
rect 3276 66508 3316 66548
rect 3358 66508 3398 66548
rect 3440 66508 3480 66548
rect 18232 66508 18272 66548
rect 18314 66508 18354 66548
rect 18396 66508 18436 66548
rect 18478 66508 18518 66548
rect 18560 66508 18600 66548
rect 33352 66508 33392 66548
rect 33434 66508 33474 66548
rect 33516 66508 33556 66548
rect 33598 66508 33638 66548
rect 33680 66508 33720 66548
rect 48472 66508 48512 66548
rect 48554 66508 48594 66548
rect 48636 66508 48676 66548
rect 48718 66508 48758 66548
rect 48800 66508 48840 66548
rect 63592 66508 63632 66548
rect 63674 66508 63714 66548
rect 63756 66508 63796 66548
rect 63838 66508 63878 66548
rect 63920 66508 63960 66548
rect 78712 66508 78752 66548
rect 78794 66508 78834 66548
rect 78876 66508 78916 66548
rect 78958 66508 78998 66548
rect 79040 66508 79080 66548
rect 93832 66508 93872 66548
rect 93914 66508 93954 66548
rect 93996 66508 94036 66548
rect 94078 66508 94118 66548
rect 94160 66508 94200 66548
rect 4352 65752 4392 65792
rect 4434 65752 4474 65792
rect 4516 65752 4556 65792
rect 4598 65752 4638 65792
rect 4680 65752 4720 65792
rect 19472 65752 19512 65792
rect 19554 65752 19594 65792
rect 19636 65752 19676 65792
rect 19718 65752 19758 65792
rect 19800 65752 19840 65792
rect 34592 65752 34632 65792
rect 34674 65752 34714 65792
rect 34756 65752 34796 65792
rect 34838 65752 34878 65792
rect 34920 65752 34960 65792
rect 49712 65752 49752 65792
rect 49794 65752 49834 65792
rect 49876 65752 49916 65792
rect 49958 65752 49998 65792
rect 50040 65752 50080 65792
rect 64832 65752 64872 65792
rect 64914 65752 64954 65792
rect 64996 65752 65036 65792
rect 65078 65752 65118 65792
rect 65160 65752 65200 65792
rect 79952 65752 79992 65792
rect 80034 65752 80074 65792
rect 80116 65752 80156 65792
rect 80198 65752 80238 65792
rect 80280 65752 80320 65792
rect 95072 65752 95112 65792
rect 95154 65752 95194 65792
rect 95236 65752 95276 65792
rect 95318 65752 95358 65792
rect 95400 65752 95440 65792
rect 3112 64996 3152 65036
rect 3194 64996 3234 65036
rect 3276 64996 3316 65036
rect 3358 64996 3398 65036
rect 3440 64996 3480 65036
rect 18232 64996 18272 65036
rect 18314 64996 18354 65036
rect 18396 64996 18436 65036
rect 18478 64996 18518 65036
rect 18560 64996 18600 65036
rect 33352 64996 33392 65036
rect 33434 64996 33474 65036
rect 33516 64996 33556 65036
rect 33598 64996 33638 65036
rect 33680 64996 33720 65036
rect 48472 64996 48512 65036
rect 48554 64996 48594 65036
rect 48636 64996 48676 65036
rect 48718 64996 48758 65036
rect 48800 64996 48840 65036
rect 63592 64996 63632 65036
rect 63674 64996 63714 65036
rect 63756 64996 63796 65036
rect 63838 64996 63878 65036
rect 63920 64996 63960 65036
rect 78712 64996 78752 65036
rect 78794 64996 78834 65036
rect 78876 64996 78916 65036
rect 78958 64996 78998 65036
rect 79040 64996 79080 65036
rect 93832 64996 93872 65036
rect 93914 64996 93954 65036
rect 93996 64996 94036 65036
rect 94078 64996 94118 65036
rect 94160 64996 94200 65036
rect 4352 64240 4392 64280
rect 4434 64240 4474 64280
rect 4516 64240 4556 64280
rect 4598 64240 4638 64280
rect 4680 64240 4720 64280
rect 19472 64240 19512 64280
rect 19554 64240 19594 64280
rect 19636 64240 19676 64280
rect 19718 64240 19758 64280
rect 19800 64240 19840 64280
rect 34592 64240 34632 64280
rect 34674 64240 34714 64280
rect 34756 64240 34796 64280
rect 34838 64240 34878 64280
rect 34920 64240 34960 64280
rect 49712 64240 49752 64280
rect 49794 64240 49834 64280
rect 49876 64240 49916 64280
rect 49958 64240 49998 64280
rect 50040 64240 50080 64280
rect 64832 64240 64872 64280
rect 64914 64240 64954 64280
rect 64996 64240 65036 64280
rect 65078 64240 65118 64280
rect 65160 64240 65200 64280
rect 79952 64240 79992 64280
rect 80034 64240 80074 64280
rect 80116 64240 80156 64280
rect 80198 64240 80238 64280
rect 80280 64240 80320 64280
rect 95072 64240 95112 64280
rect 95154 64240 95194 64280
rect 95236 64240 95276 64280
rect 95318 64240 95358 64280
rect 95400 64240 95440 64280
rect 3112 63484 3152 63524
rect 3194 63484 3234 63524
rect 3276 63484 3316 63524
rect 3358 63484 3398 63524
rect 3440 63484 3480 63524
rect 18232 63484 18272 63524
rect 18314 63484 18354 63524
rect 18396 63484 18436 63524
rect 18478 63484 18518 63524
rect 18560 63484 18600 63524
rect 33352 63484 33392 63524
rect 33434 63484 33474 63524
rect 33516 63484 33556 63524
rect 33598 63484 33638 63524
rect 33680 63484 33720 63524
rect 48472 63484 48512 63524
rect 48554 63484 48594 63524
rect 48636 63484 48676 63524
rect 48718 63484 48758 63524
rect 48800 63484 48840 63524
rect 63592 63484 63632 63524
rect 63674 63484 63714 63524
rect 63756 63484 63796 63524
rect 63838 63484 63878 63524
rect 63920 63484 63960 63524
rect 78712 63484 78752 63524
rect 78794 63484 78834 63524
rect 78876 63484 78916 63524
rect 78958 63484 78998 63524
rect 79040 63484 79080 63524
rect 93832 63484 93872 63524
rect 93914 63484 93954 63524
rect 93996 63484 94036 63524
rect 94078 63484 94118 63524
rect 94160 63484 94200 63524
rect 4352 62728 4392 62768
rect 4434 62728 4474 62768
rect 4516 62728 4556 62768
rect 4598 62728 4638 62768
rect 4680 62728 4720 62768
rect 19472 62728 19512 62768
rect 19554 62728 19594 62768
rect 19636 62728 19676 62768
rect 19718 62728 19758 62768
rect 19800 62728 19840 62768
rect 34592 62728 34632 62768
rect 34674 62728 34714 62768
rect 34756 62728 34796 62768
rect 34838 62728 34878 62768
rect 34920 62728 34960 62768
rect 49712 62728 49752 62768
rect 49794 62728 49834 62768
rect 49876 62728 49916 62768
rect 49958 62728 49998 62768
rect 50040 62728 50080 62768
rect 64832 62728 64872 62768
rect 64914 62728 64954 62768
rect 64996 62728 65036 62768
rect 65078 62728 65118 62768
rect 65160 62728 65200 62768
rect 79952 62728 79992 62768
rect 80034 62728 80074 62768
rect 80116 62728 80156 62768
rect 80198 62728 80238 62768
rect 80280 62728 80320 62768
rect 95072 62728 95112 62768
rect 95154 62728 95194 62768
rect 95236 62728 95276 62768
rect 95318 62728 95358 62768
rect 95400 62728 95440 62768
rect 3112 61972 3152 62012
rect 3194 61972 3234 62012
rect 3276 61972 3316 62012
rect 3358 61972 3398 62012
rect 3440 61972 3480 62012
rect 18232 61972 18272 62012
rect 18314 61972 18354 62012
rect 18396 61972 18436 62012
rect 18478 61972 18518 62012
rect 18560 61972 18600 62012
rect 33352 61972 33392 62012
rect 33434 61972 33474 62012
rect 33516 61972 33556 62012
rect 33598 61972 33638 62012
rect 33680 61972 33720 62012
rect 48472 61972 48512 62012
rect 48554 61972 48594 62012
rect 48636 61972 48676 62012
rect 48718 61972 48758 62012
rect 48800 61972 48840 62012
rect 63592 61972 63632 62012
rect 63674 61972 63714 62012
rect 63756 61972 63796 62012
rect 63838 61972 63878 62012
rect 63920 61972 63960 62012
rect 78712 61972 78752 62012
rect 78794 61972 78834 62012
rect 78876 61972 78916 62012
rect 78958 61972 78998 62012
rect 79040 61972 79080 62012
rect 93832 61972 93872 62012
rect 93914 61972 93954 62012
rect 93996 61972 94036 62012
rect 94078 61972 94118 62012
rect 94160 61972 94200 62012
rect 4352 61216 4392 61256
rect 4434 61216 4474 61256
rect 4516 61216 4556 61256
rect 4598 61216 4638 61256
rect 4680 61216 4720 61256
rect 19472 61216 19512 61256
rect 19554 61216 19594 61256
rect 19636 61216 19676 61256
rect 19718 61216 19758 61256
rect 19800 61216 19840 61256
rect 34592 61216 34632 61256
rect 34674 61216 34714 61256
rect 34756 61216 34796 61256
rect 34838 61216 34878 61256
rect 34920 61216 34960 61256
rect 49712 61216 49752 61256
rect 49794 61216 49834 61256
rect 49876 61216 49916 61256
rect 49958 61216 49998 61256
rect 50040 61216 50080 61256
rect 64832 61216 64872 61256
rect 64914 61216 64954 61256
rect 64996 61216 65036 61256
rect 65078 61216 65118 61256
rect 65160 61216 65200 61256
rect 79952 61216 79992 61256
rect 80034 61216 80074 61256
rect 80116 61216 80156 61256
rect 80198 61216 80238 61256
rect 80280 61216 80320 61256
rect 95072 61216 95112 61256
rect 95154 61216 95194 61256
rect 95236 61216 95276 61256
rect 95318 61216 95358 61256
rect 95400 61216 95440 61256
rect 3112 60460 3152 60500
rect 3194 60460 3234 60500
rect 3276 60460 3316 60500
rect 3358 60460 3398 60500
rect 3440 60460 3480 60500
rect 18232 60460 18272 60500
rect 18314 60460 18354 60500
rect 18396 60460 18436 60500
rect 18478 60460 18518 60500
rect 18560 60460 18600 60500
rect 33352 60460 33392 60500
rect 33434 60460 33474 60500
rect 33516 60460 33556 60500
rect 33598 60460 33638 60500
rect 33680 60460 33720 60500
rect 48472 60460 48512 60500
rect 48554 60460 48594 60500
rect 48636 60460 48676 60500
rect 48718 60460 48758 60500
rect 48800 60460 48840 60500
rect 63592 60460 63632 60500
rect 63674 60460 63714 60500
rect 63756 60460 63796 60500
rect 63838 60460 63878 60500
rect 63920 60460 63960 60500
rect 78712 60460 78752 60500
rect 78794 60460 78834 60500
rect 78876 60460 78916 60500
rect 78958 60460 78998 60500
rect 79040 60460 79080 60500
rect 93832 60460 93872 60500
rect 93914 60460 93954 60500
rect 93996 60460 94036 60500
rect 94078 60460 94118 60500
rect 94160 60460 94200 60500
rect 4352 59704 4392 59744
rect 4434 59704 4474 59744
rect 4516 59704 4556 59744
rect 4598 59704 4638 59744
rect 4680 59704 4720 59744
rect 19472 59704 19512 59744
rect 19554 59704 19594 59744
rect 19636 59704 19676 59744
rect 19718 59704 19758 59744
rect 19800 59704 19840 59744
rect 34592 59704 34632 59744
rect 34674 59704 34714 59744
rect 34756 59704 34796 59744
rect 34838 59704 34878 59744
rect 34920 59704 34960 59744
rect 49712 59704 49752 59744
rect 49794 59704 49834 59744
rect 49876 59704 49916 59744
rect 49958 59704 49998 59744
rect 50040 59704 50080 59744
rect 64832 59704 64872 59744
rect 64914 59704 64954 59744
rect 64996 59704 65036 59744
rect 65078 59704 65118 59744
rect 65160 59704 65200 59744
rect 79952 59704 79992 59744
rect 80034 59704 80074 59744
rect 80116 59704 80156 59744
rect 80198 59704 80238 59744
rect 80280 59704 80320 59744
rect 95072 59704 95112 59744
rect 95154 59704 95194 59744
rect 95236 59704 95276 59744
rect 95318 59704 95358 59744
rect 95400 59704 95440 59744
rect 3112 58948 3152 58988
rect 3194 58948 3234 58988
rect 3276 58948 3316 58988
rect 3358 58948 3398 58988
rect 3440 58948 3480 58988
rect 18232 58948 18272 58988
rect 18314 58948 18354 58988
rect 18396 58948 18436 58988
rect 18478 58948 18518 58988
rect 18560 58948 18600 58988
rect 33352 58948 33392 58988
rect 33434 58948 33474 58988
rect 33516 58948 33556 58988
rect 33598 58948 33638 58988
rect 33680 58948 33720 58988
rect 48472 58948 48512 58988
rect 48554 58948 48594 58988
rect 48636 58948 48676 58988
rect 48718 58948 48758 58988
rect 48800 58948 48840 58988
rect 63592 58948 63632 58988
rect 63674 58948 63714 58988
rect 63756 58948 63796 58988
rect 63838 58948 63878 58988
rect 63920 58948 63960 58988
rect 78712 58948 78752 58988
rect 78794 58948 78834 58988
rect 78876 58948 78916 58988
rect 78958 58948 78998 58988
rect 79040 58948 79080 58988
rect 93832 58948 93872 58988
rect 93914 58948 93954 58988
rect 93996 58948 94036 58988
rect 94078 58948 94118 58988
rect 94160 58948 94200 58988
rect 4352 58192 4392 58232
rect 4434 58192 4474 58232
rect 4516 58192 4556 58232
rect 4598 58192 4638 58232
rect 4680 58192 4720 58232
rect 19472 58192 19512 58232
rect 19554 58192 19594 58232
rect 19636 58192 19676 58232
rect 19718 58192 19758 58232
rect 19800 58192 19840 58232
rect 34592 58192 34632 58232
rect 34674 58192 34714 58232
rect 34756 58192 34796 58232
rect 34838 58192 34878 58232
rect 34920 58192 34960 58232
rect 49712 58192 49752 58232
rect 49794 58192 49834 58232
rect 49876 58192 49916 58232
rect 49958 58192 49998 58232
rect 50040 58192 50080 58232
rect 64832 58192 64872 58232
rect 64914 58192 64954 58232
rect 64996 58192 65036 58232
rect 65078 58192 65118 58232
rect 65160 58192 65200 58232
rect 79952 58192 79992 58232
rect 80034 58192 80074 58232
rect 80116 58192 80156 58232
rect 80198 58192 80238 58232
rect 80280 58192 80320 58232
rect 95072 58192 95112 58232
rect 95154 58192 95194 58232
rect 95236 58192 95276 58232
rect 95318 58192 95358 58232
rect 95400 58192 95440 58232
rect 3112 57436 3152 57476
rect 3194 57436 3234 57476
rect 3276 57436 3316 57476
rect 3358 57436 3398 57476
rect 3440 57436 3480 57476
rect 18232 57436 18272 57476
rect 18314 57436 18354 57476
rect 18396 57436 18436 57476
rect 18478 57436 18518 57476
rect 18560 57436 18600 57476
rect 33352 57436 33392 57476
rect 33434 57436 33474 57476
rect 33516 57436 33556 57476
rect 33598 57436 33638 57476
rect 33680 57436 33720 57476
rect 48472 57436 48512 57476
rect 48554 57436 48594 57476
rect 48636 57436 48676 57476
rect 48718 57436 48758 57476
rect 48800 57436 48840 57476
rect 63592 57436 63632 57476
rect 63674 57436 63714 57476
rect 63756 57436 63796 57476
rect 63838 57436 63878 57476
rect 63920 57436 63960 57476
rect 78712 57436 78752 57476
rect 78794 57436 78834 57476
rect 78876 57436 78916 57476
rect 78958 57436 78998 57476
rect 79040 57436 79080 57476
rect 93832 57436 93872 57476
rect 93914 57436 93954 57476
rect 93996 57436 94036 57476
rect 94078 57436 94118 57476
rect 94160 57436 94200 57476
rect 4352 56680 4392 56720
rect 4434 56680 4474 56720
rect 4516 56680 4556 56720
rect 4598 56680 4638 56720
rect 4680 56680 4720 56720
rect 19472 56680 19512 56720
rect 19554 56680 19594 56720
rect 19636 56680 19676 56720
rect 19718 56680 19758 56720
rect 19800 56680 19840 56720
rect 34592 56680 34632 56720
rect 34674 56680 34714 56720
rect 34756 56680 34796 56720
rect 34838 56680 34878 56720
rect 34920 56680 34960 56720
rect 49712 56680 49752 56720
rect 49794 56680 49834 56720
rect 49876 56680 49916 56720
rect 49958 56680 49998 56720
rect 50040 56680 50080 56720
rect 64832 56680 64872 56720
rect 64914 56680 64954 56720
rect 64996 56680 65036 56720
rect 65078 56680 65118 56720
rect 65160 56680 65200 56720
rect 79952 56680 79992 56720
rect 80034 56680 80074 56720
rect 80116 56680 80156 56720
rect 80198 56680 80238 56720
rect 80280 56680 80320 56720
rect 95072 56680 95112 56720
rect 95154 56680 95194 56720
rect 95236 56680 95276 56720
rect 95318 56680 95358 56720
rect 95400 56680 95440 56720
rect 3112 55924 3152 55964
rect 3194 55924 3234 55964
rect 3276 55924 3316 55964
rect 3358 55924 3398 55964
rect 3440 55924 3480 55964
rect 18232 55924 18272 55964
rect 18314 55924 18354 55964
rect 18396 55924 18436 55964
rect 18478 55924 18518 55964
rect 18560 55924 18600 55964
rect 33352 55924 33392 55964
rect 33434 55924 33474 55964
rect 33516 55924 33556 55964
rect 33598 55924 33638 55964
rect 33680 55924 33720 55964
rect 48472 55924 48512 55964
rect 48554 55924 48594 55964
rect 48636 55924 48676 55964
rect 48718 55924 48758 55964
rect 48800 55924 48840 55964
rect 63592 55924 63632 55964
rect 63674 55924 63714 55964
rect 63756 55924 63796 55964
rect 63838 55924 63878 55964
rect 63920 55924 63960 55964
rect 78712 55924 78752 55964
rect 78794 55924 78834 55964
rect 78876 55924 78916 55964
rect 78958 55924 78998 55964
rect 79040 55924 79080 55964
rect 93832 55924 93872 55964
rect 93914 55924 93954 55964
rect 93996 55924 94036 55964
rect 94078 55924 94118 55964
rect 94160 55924 94200 55964
rect 4352 55168 4392 55208
rect 4434 55168 4474 55208
rect 4516 55168 4556 55208
rect 4598 55168 4638 55208
rect 4680 55168 4720 55208
rect 19472 55168 19512 55208
rect 19554 55168 19594 55208
rect 19636 55168 19676 55208
rect 19718 55168 19758 55208
rect 19800 55168 19840 55208
rect 34592 55168 34632 55208
rect 34674 55168 34714 55208
rect 34756 55168 34796 55208
rect 34838 55168 34878 55208
rect 34920 55168 34960 55208
rect 49712 55168 49752 55208
rect 49794 55168 49834 55208
rect 49876 55168 49916 55208
rect 49958 55168 49998 55208
rect 50040 55168 50080 55208
rect 64832 55168 64872 55208
rect 64914 55168 64954 55208
rect 64996 55168 65036 55208
rect 65078 55168 65118 55208
rect 65160 55168 65200 55208
rect 79952 55168 79992 55208
rect 80034 55168 80074 55208
rect 80116 55168 80156 55208
rect 80198 55168 80238 55208
rect 80280 55168 80320 55208
rect 95072 55168 95112 55208
rect 95154 55168 95194 55208
rect 95236 55168 95276 55208
rect 95318 55168 95358 55208
rect 95400 55168 95440 55208
rect 3112 54412 3152 54452
rect 3194 54412 3234 54452
rect 3276 54412 3316 54452
rect 3358 54412 3398 54452
rect 3440 54412 3480 54452
rect 18232 54412 18272 54452
rect 18314 54412 18354 54452
rect 18396 54412 18436 54452
rect 18478 54412 18518 54452
rect 18560 54412 18600 54452
rect 33352 54412 33392 54452
rect 33434 54412 33474 54452
rect 33516 54412 33556 54452
rect 33598 54412 33638 54452
rect 33680 54412 33720 54452
rect 48472 54412 48512 54452
rect 48554 54412 48594 54452
rect 48636 54412 48676 54452
rect 48718 54412 48758 54452
rect 48800 54412 48840 54452
rect 63592 54412 63632 54452
rect 63674 54412 63714 54452
rect 63756 54412 63796 54452
rect 63838 54412 63878 54452
rect 63920 54412 63960 54452
rect 78712 54412 78752 54452
rect 78794 54412 78834 54452
rect 78876 54412 78916 54452
rect 78958 54412 78998 54452
rect 79040 54412 79080 54452
rect 93832 54412 93872 54452
rect 93914 54412 93954 54452
rect 93996 54412 94036 54452
rect 94078 54412 94118 54452
rect 94160 54412 94200 54452
rect 4352 53656 4392 53696
rect 4434 53656 4474 53696
rect 4516 53656 4556 53696
rect 4598 53656 4638 53696
rect 4680 53656 4720 53696
rect 19472 53656 19512 53696
rect 19554 53656 19594 53696
rect 19636 53656 19676 53696
rect 19718 53656 19758 53696
rect 19800 53656 19840 53696
rect 34592 53656 34632 53696
rect 34674 53656 34714 53696
rect 34756 53656 34796 53696
rect 34838 53656 34878 53696
rect 34920 53656 34960 53696
rect 49712 53656 49752 53696
rect 49794 53656 49834 53696
rect 49876 53656 49916 53696
rect 49958 53656 49998 53696
rect 50040 53656 50080 53696
rect 64832 53656 64872 53696
rect 64914 53656 64954 53696
rect 64996 53656 65036 53696
rect 65078 53656 65118 53696
rect 65160 53656 65200 53696
rect 79952 53656 79992 53696
rect 80034 53656 80074 53696
rect 80116 53656 80156 53696
rect 80198 53656 80238 53696
rect 80280 53656 80320 53696
rect 95072 53656 95112 53696
rect 95154 53656 95194 53696
rect 95236 53656 95276 53696
rect 95318 53656 95358 53696
rect 95400 53656 95440 53696
rect 3112 52900 3152 52940
rect 3194 52900 3234 52940
rect 3276 52900 3316 52940
rect 3358 52900 3398 52940
rect 3440 52900 3480 52940
rect 18232 52900 18272 52940
rect 18314 52900 18354 52940
rect 18396 52900 18436 52940
rect 18478 52900 18518 52940
rect 18560 52900 18600 52940
rect 33352 52900 33392 52940
rect 33434 52900 33474 52940
rect 33516 52900 33556 52940
rect 33598 52900 33638 52940
rect 33680 52900 33720 52940
rect 48472 52900 48512 52940
rect 48554 52900 48594 52940
rect 48636 52900 48676 52940
rect 48718 52900 48758 52940
rect 48800 52900 48840 52940
rect 63592 52900 63632 52940
rect 63674 52900 63714 52940
rect 63756 52900 63796 52940
rect 63838 52900 63878 52940
rect 63920 52900 63960 52940
rect 78712 52900 78752 52940
rect 78794 52900 78834 52940
rect 78876 52900 78916 52940
rect 78958 52900 78998 52940
rect 79040 52900 79080 52940
rect 93832 52900 93872 52940
rect 93914 52900 93954 52940
rect 93996 52900 94036 52940
rect 94078 52900 94118 52940
rect 94160 52900 94200 52940
rect 4352 52144 4392 52184
rect 4434 52144 4474 52184
rect 4516 52144 4556 52184
rect 4598 52144 4638 52184
rect 4680 52144 4720 52184
rect 19472 52144 19512 52184
rect 19554 52144 19594 52184
rect 19636 52144 19676 52184
rect 19718 52144 19758 52184
rect 19800 52144 19840 52184
rect 34592 52144 34632 52184
rect 34674 52144 34714 52184
rect 34756 52144 34796 52184
rect 34838 52144 34878 52184
rect 34920 52144 34960 52184
rect 49712 52144 49752 52184
rect 49794 52144 49834 52184
rect 49876 52144 49916 52184
rect 49958 52144 49998 52184
rect 50040 52144 50080 52184
rect 64832 52144 64872 52184
rect 64914 52144 64954 52184
rect 64996 52144 65036 52184
rect 65078 52144 65118 52184
rect 65160 52144 65200 52184
rect 79952 52144 79992 52184
rect 80034 52144 80074 52184
rect 80116 52144 80156 52184
rect 80198 52144 80238 52184
rect 80280 52144 80320 52184
rect 95072 52144 95112 52184
rect 95154 52144 95194 52184
rect 95236 52144 95276 52184
rect 95318 52144 95358 52184
rect 95400 52144 95440 52184
rect 3112 51388 3152 51428
rect 3194 51388 3234 51428
rect 3276 51388 3316 51428
rect 3358 51388 3398 51428
rect 3440 51388 3480 51428
rect 18232 51388 18272 51428
rect 18314 51388 18354 51428
rect 18396 51388 18436 51428
rect 18478 51388 18518 51428
rect 18560 51388 18600 51428
rect 33352 51388 33392 51428
rect 33434 51388 33474 51428
rect 33516 51388 33556 51428
rect 33598 51388 33638 51428
rect 33680 51388 33720 51428
rect 48472 51388 48512 51428
rect 48554 51388 48594 51428
rect 48636 51388 48676 51428
rect 48718 51388 48758 51428
rect 48800 51388 48840 51428
rect 63592 51388 63632 51428
rect 63674 51388 63714 51428
rect 63756 51388 63796 51428
rect 63838 51388 63878 51428
rect 63920 51388 63960 51428
rect 78712 51388 78752 51428
rect 78794 51388 78834 51428
rect 78876 51388 78916 51428
rect 78958 51388 78998 51428
rect 79040 51388 79080 51428
rect 93832 51388 93872 51428
rect 93914 51388 93954 51428
rect 93996 51388 94036 51428
rect 94078 51388 94118 51428
rect 94160 51388 94200 51428
rect 4352 50632 4392 50672
rect 4434 50632 4474 50672
rect 4516 50632 4556 50672
rect 4598 50632 4638 50672
rect 4680 50632 4720 50672
rect 19472 50632 19512 50672
rect 19554 50632 19594 50672
rect 19636 50632 19676 50672
rect 19718 50632 19758 50672
rect 19800 50632 19840 50672
rect 34592 50632 34632 50672
rect 34674 50632 34714 50672
rect 34756 50632 34796 50672
rect 34838 50632 34878 50672
rect 34920 50632 34960 50672
rect 49712 50632 49752 50672
rect 49794 50632 49834 50672
rect 49876 50632 49916 50672
rect 49958 50632 49998 50672
rect 50040 50632 50080 50672
rect 64832 50632 64872 50672
rect 64914 50632 64954 50672
rect 64996 50632 65036 50672
rect 65078 50632 65118 50672
rect 65160 50632 65200 50672
rect 79952 50632 79992 50672
rect 80034 50632 80074 50672
rect 80116 50632 80156 50672
rect 80198 50632 80238 50672
rect 80280 50632 80320 50672
rect 95072 50632 95112 50672
rect 95154 50632 95194 50672
rect 95236 50632 95276 50672
rect 95318 50632 95358 50672
rect 95400 50632 95440 50672
rect 3112 49876 3152 49916
rect 3194 49876 3234 49916
rect 3276 49876 3316 49916
rect 3358 49876 3398 49916
rect 3440 49876 3480 49916
rect 18232 49876 18272 49916
rect 18314 49876 18354 49916
rect 18396 49876 18436 49916
rect 18478 49876 18518 49916
rect 18560 49876 18600 49916
rect 33352 49876 33392 49916
rect 33434 49876 33474 49916
rect 33516 49876 33556 49916
rect 33598 49876 33638 49916
rect 33680 49876 33720 49916
rect 48472 49876 48512 49916
rect 48554 49876 48594 49916
rect 48636 49876 48676 49916
rect 48718 49876 48758 49916
rect 48800 49876 48840 49916
rect 63592 49876 63632 49916
rect 63674 49876 63714 49916
rect 63756 49876 63796 49916
rect 63838 49876 63878 49916
rect 63920 49876 63960 49916
rect 78712 49876 78752 49916
rect 78794 49876 78834 49916
rect 78876 49876 78916 49916
rect 78958 49876 78998 49916
rect 79040 49876 79080 49916
rect 93832 49876 93872 49916
rect 93914 49876 93954 49916
rect 93996 49876 94036 49916
rect 94078 49876 94118 49916
rect 94160 49876 94200 49916
rect 4352 49120 4392 49160
rect 4434 49120 4474 49160
rect 4516 49120 4556 49160
rect 4598 49120 4638 49160
rect 4680 49120 4720 49160
rect 19472 49120 19512 49160
rect 19554 49120 19594 49160
rect 19636 49120 19676 49160
rect 19718 49120 19758 49160
rect 19800 49120 19840 49160
rect 34592 49120 34632 49160
rect 34674 49120 34714 49160
rect 34756 49120 34796 49160
rect 34838 49120 34878 49160
rect 34920 49120 34960 49160
rect 49712 49120 49752 49160
rect 49794 49120 49834 49160
rect 49876 49120 49916 49160
rect 49958 49120 49998 49160
rect 50040 49120 50080 49160
rect 64832 49120 64872 49160
rect 64914 49120 64954 49160
rect 64996 49120 65036 49160
rect 65078 49120 65118 49160
rect 65160 49120 65200 49160
rect 79952 49120 79992 49160
rect 80034 49120 80074 49160
rect 80116 49120 80156 49160
rect 80198 49120 80238 49160
rect 80280 49120 80320 49160
rect 95072 49120 95112 49160
rect 95154 49120 95194 49160
rect 95236 49120 95276 49160
rect 95318 49120 95358 49160
rect 95400 49120 95440 49160
rect 3112 48364 3152 48404
rect 3194 48364 3234 48404
rect 3276 48364 3316 48404
rect 3358 48364 3398 48404
rect 3440 48364 3480 48404
rect 18232 48364 18272 48404
rect 18314 48364 18354 48404
rect 18396 48364 18436 48404
rect 18478 48364 18518 48404
rect 18560 48364 18600 48404
rect 33352 48364 33392 48404
rect 33434 48364 33474 48404
rect 33516 48364 33556 48404
rect 33598 48364 33638 48404
rect 33680 48364 33720 48404
rect 48472 48364 48512 48404
rect 48554 48364 48594 48404
rect 48636 48364 48676 48404
rect 48718 48364 48758 48404
rect 48800 48364 48840 48404
rect 63592 48364 63632 48404
rect 63674 48364 63714 48404
rect 63756 48364 63796 48404
rect 63838 48364 63878 48404
rect 63920 48364 63960 48404
rect 78712 48364 78752 48404
rect 78794 48364 78834 48404
rect 78876 48364 78916 48404
rect 78958 48364 78998 48404
rect 79040 48364 79080 48404
rect 93832 48364 93872 48404
rect 93914 48364 93954 48404
rect 93996 48364 94036 48404
rect 94078 48364 94118 48404
rect 94160 48364 94200 48404
rect 4352 47608 4392 47648
rect 4434 47608 4474 47648
rect 4516 47608 4556 47648
rect 4598 47608 4638 47648
rect 4680 47608 4720 47648
rect 19472 47608 19512 47648
rect 19554 47608 19594 47648
rect 19636 47608 19676 47648
rect 19718 47608 19758 47648
rect 19800 47608 19840 47648
rect 34592 47608 34632 47648
rect 34674 47608 34714 47648
rect 34756 47608 34796 47648
rect 34838 47608 34878 47648
rect 34920 47608 34960 47648
rect 49712 47608 49752 47648
rect 49794 47608 49834 47648
rect 49876 47608 49916 47648
rect 49958 47608 49998 47648
rect 50040 47608 50080 47648
rect 64832 47608 64872 47648
rect 64914 47608 64954 47648
rect 64996 47608 65036 47648
rect 65078 47608 65118 47648
rect 65160 47608 65200 47648
rect 79952 47608 79992 47648
rect 80034 47608 80074 47648
rect 80116 47608 80156 47648
rect 80198 47608 80238 47648
rect 80280 47608 80320 47648
rect 95072 47608 95112 47648
rect 95154 47608 95194 47648
rect 95236 47608 95276 47648
rect 95318 47608 95358 47648
rect 95400 47608 95440 47648
rect 3112 46852 3152 46892
rect 3194 46852 3234 46892
rect 3276 46852 3316 46892
rect 3358 46852 3398 46892
rect 3440 46852 3480 46892
rect 18232 46852 18272 46892
rect 18314 46852 18354 46892
rect 18396 46852 18436 46892
rect 18478 46852 18518 46892
rect 18560 46852 18600 46892
rect 33352 46852 33392 46892
rect 33434 46852 33474 46892
rect 33516 46852 33556 46892
rect 33598 46852 33638 46892
rect 33680 46852 33720 46892
rect 48472 46852 48512 46892
rect 48554 46852 48594 46892
rect 48636 46852 48676 46892
rect 48718 46852 48758 46892
rect 48800 46852 48840 46892
rect 63592 46852 63632 46892
rect 63674 46852 63714 46892
rect 63756 46852 63796 46892
rect 63838 46852 63878 46892
rect 63920 46852 63960 46892
rect 78712 46852 78752 46892
rect 78794 46852 78834 46892
rect 78876 46852 78916 46892
rect 78958 46852 78998 46892
rect 79040 46852 79080 46892
rect 93832 46852 93872 46892
rect 93914 46852 93954 46892
rect 93996 46852 94036 46892
rect 94078 46852 94118 46892
rect 94160 46852 94200 46892
rect 4352 46096 4392 46136
rect 4434 46096 4474 46136
rect 4516 46096 4556 46136
rect 4598 46096 4638 46136
rect 4680 46096 4720 46136
rect 19472 46096 19512 46136
rect 19554 46096 19594 46136
rect 19636 46096 19676 46136
rect 19718 46096 19758 46136
rect 19800 46096 19840 46136
rect 34592 46096 34632 46136
rect 34674 46096 34714 46136
rect 34756 46096 34796 46136
rect 34838 46096 34878 46136
rect 34920 46096 34960 46136
rect 49712 46096 49752 46136
rect 49794 46096 49834 46136
rect 49876 46096 49916 46136
rect 49958 46096 49998 46136
rect 50040 46096 50080 46136
rect 64832 46096 64872 46136
rect 64914 46096 64954 46136
rect 64996 46096 65036 46136
rect 65078 46096 65118 46136
rect 65160 46096 65200 46136
rect 79952 46096 79992 46136
rect 80034 46096 80074 46136
rect 80116 46096 80156 46136
rect 80198 46096 80238 46136
rect 80280 46096 80320 46136
rect 95072 46096 95112 46136
rect 95154 46096 95194 46136
rect 95236 46096 95276 46136
rect 95318 46096 95358 46136
rect 95400 46096 95440 46136
rect 3112 45340 3152 45380
rect 3194 45340 3234 45380
rect 3276 45340 3316 45380
rect 3358 45340 3398 45380
rect 3440 45340 3480 45380
rect 18232 45340 18272 45380
rect 18314 45340 18354 45380
rect 18396 45340 18436 45380
rect 18478 45340 18518 45380
rect 18560 45340 18600 45380
rect 33352 45340 33392 45380
rect 33434 45340 33474 45380
rect 33516 45340 33556 45380
rect 33598 45340 33638 45380
rect 33680 45340 33720 45380
rect 48472 45340 48512 45380
rect 48554 45340 48594 45380
rect 48636 45340 48676 45380
rect 48718 45340 48758 45380
rect 48800 45340 48840 45380
rect 63592 45340 63632 45380
rect 63674 45340 63714 45380
rect 63756 45340 63796 45380
rect 63838 45340 63878 45380
rect 63920 45340 63960 45380
rect 78712 45340 78752 45380
rect 78794 45340 78834 45380
rect 78876 45340 78916 45380
rect 78958 45340 78998 45380
rect 79040 45340 79080 45380
rect 93832 45340 93872 45380
rect 93914 45340 93954 45380
rect 93996 45340 94036 45380
rect 94078 45340 94118 45380
rect 94160 45340 94200 45380
rect 4352 44584 4392 44624
rect 4434 44584 4474 44624
rect 4516 44584 4556 44624
rect 4598 44584 4638 44624
rect 4680 44584 4720 44624
rect 19472 44584 19512 44624
rect 19554 44584 19594 44624
rect 19636 44584 19676 44624
rect 19718 44584 19758 44624
rect 19800 44584 19840 44624
rect 34592 44584 34632 44624
rect 34674 44584 34714 44624
rect 34756 44584 34796 44624
rect 34838 44584 34878 44624
rect 34920 44584 34960 44624
rect 49712 44584 49752 44624
rect 49794 44584 49834 44624
rect 49876 44584 49916 44624
rect 49958 44584 49998 44624
rect 50040 44584 50080 44624
rect 64832 44584 64872 44624
rect 64914 44584 64954 44624
rect 64996 44584 65036 44624
rect 65078 44584 65118 44624
rect 65160 44584 65200 44624
rect 79952 44584 79992 44624
rect 80034 44584 80074 44624
rect 80116 44584 80156 44624
rect 80198 44584 80238 44624
rect 80280 44584 80320 44624
rect 95072 44584 95112 44624
rect 95154 44584 95194 44624
rect 95236 44584 95276 44624
rect 95318 44584 95358 44624
rect 95400 44584 95440 44624
rect 3112 43828 3152 43868
rect 3194 43828 3234 43868
rect 3276 43828 3316 43868
rect 3358 43828 3398 43868
rect 3440 43828 3480 43868
rect 18232 43828 18272 43868
rect 18314 43828 18354 43868
rect 18396 43828 18436 43868
rect 18478 43828 18518 43868
rect 18560 43828 18600 43868
rect 33352 43828 33392 43868
rect 33434 43828 33474 43868
rect 33516 43828 33556 43868
rect 33598 43828 33638 43868
rect 33680 43828 33720 43868
rect 48472 43828 48512 43868
rect 48554 43828 48594 43868
rect 48636 43828 48676 43868
rect 48718 43828 48758 43868
rect 48800 43828 48840 43868
rect 63592 43828 63632 43868
rect 63674 43828 63714 43868
rect 63756 43828 63796 43868
rect 63838 43828 63878 43868
rect 63920 43828 63960 43868
rect 78712 43828 78752 43868
rect 78794 43828 78834 43868
rect 78876 43828 78916 43868
rect 78958 43828 78998 43868
rect 79040 43828 79080 43868
rect 93832 43828 93872 43868
rect 93914 43828 93954 43868
rect 93996 43828 94036 43868
rect 94078 43828 94118 43868
rect 94160 43828 94200 43868
rect 4352 43072 4392 43112
rect 4434 43072 4474 43112
rect 4516 43072 4556 43112
rect 4598 43072 4638 43112
rect 4680 43072 4720 43112
rect 19472 43072 19512 43112
rect 19554 43072 19594 43112
rect 19636 43072 19676 43112
rect 19718 43072 19758 43112
rect 19800 43072 19840 43112
rect 34592 43072 34632 43112
rect 34674 43072 34714 43112
rect 34756 43072 34796 43112
rect 34838 43072 34878 43112
rect 34920 43072 34960 43112
rect 49712 43072 49752 43112
rect 49794 43072 49834 43112
rect 49876 43072 49916 43112
rect 49958 43072 49998 43112
rect 50040 43072 50080 43112
rect 64832 43072 64872 43112
rect 64914 43072 64954 43112
rect 64996 43072 65036 43112
rect 65078 43072 65118 43112
rect 65160 43072 65200 43112
rect 79952 43072 79992 43112
rect 80034 43072 80074 43112
rect 80116 43072 80156 43112
rect 80198 43072 80238 43112
rect 80280 43072 80320 43112
rect 95072 43072 95112 43112
rect 95154 43072 95194 43112
rect 95236 43072 95276 43112
rect 95318 43072 95358 43112
rect 95400 43072 95440 43112
rect 3112 42316 3152 42356
rect 3194 42316 3234 42356
rect 3276 42316 3316 42356
rect 3358 42316 3398 42356
rect 3440 42316 3480 42356
rect 18232 42316 18272 42356
rect 18314 42316 18354 42356
rect 18396 42316 18436 42356
rect 18478 42316 18518 42356
rect 18560 42316 18600 42356
rect 33352 42316 33392 42356
rect 33434 42316 33474 42356
rect 33516 42316 33556 42356
rect 33598 42316 33638 42356
rect 33680 42316 33720 42356
rect 48472 42316 48512 42356
rect 48554 42316 48594 42356
rect 48636 42316 48676 42356
rect 48718 42316 48758 42356
rect 48800 42316 48840 42356
rect 63592 42316 63632 42356
rect 63674 42316 63714 42356
rect 63756 42316 63796 42356
rect 63838 42316 63878 42356
rect 63920 42316 63960 42356
rect 78712 42316 78752 42356
rect 78794 42316 78834 42356
rect 78876 42316 78916 42356
rect 78958 42316 78998 42356
rect 79040 42316 79080 42356
rect 93832 42316 93872 42356
rect 93914 42316 93954 42356
rect 93996 42316 94036 42356
rect 94078 42316 94118 42356
rect 94160 42316 94200 42356
rect 4352 41560 4392 41600
rect 4434 41560 4474 41600
rect 4516 41560 4556 41600
rect 4598 41560 4638 41600
rect 4680 41560 4720 41600
rect 19472 41560 19512 41600
rect 19554 41560 19594 41600
rect 19636 41560 19676 41600
rect 19718 41560 19758 41600
rect 19800 41560 19840 41600
rect 34592 41560 34632 41600
rect 34674 41560 34714 41600
rect 34756 41560 34796 41600
rect 34838 41560 34878 41600
rect 34920 41560 34960 41600
rect 49712 41560 49752 41600
rect 49794 41560 49834 41600
rect 49876 41560 49916 41600
rect 49958 41560 49998 41600
rect 50040 41560 50080 41600
rect 64832 41560 64872 41600
rect 64914 41560 64954 41600
rect 64996 41560 65036 41600
rect 65078 41560 65118 41600
rect 65160 41560 65200 41600
rect 79952 41560 79992 41600
rect 80034 41560 80074 41600
rect 80116 41560 80156 41600
rect 80198 41560 80238 41600
rect 80280 41560 80320 41600
rect 95072 41560 95112 41600
rect 95154 41560 95194 41600
rect 95236 41560 95276 41600
rect 95318 41560 95358 41600
rect 95400 41560 95440 41600
rect 3112 40804 3152 40844
rect 3194 40804 3234 40844
rect 3276 40804 3316 40844
rect 3358 40804 3398 40844
rect 3440 40804 3480 40844
rect 18232 40804 18272 40844
rect 18314 40804 18354 40844
rect 18396 40804 18436 40844
rect 18478 40804 18518 40844
rect 18560 40804 18600 40844
rect 33352 40804 33392 40844
rect 33434 40804 33474 40844
rect 33516 40804 33556 40844
rect 33598 40804 33638 40844
rect 33680 40804 33720 40844
rect 48472 40804 48512 40844
rect 48554 40804 48594 40844
rect 48636 40804 48676 40844
rect 48718 40804 48758 40844
rect 48800 40804 48840 40844
rect 63592 40804 63632 40844
rect 63674 40804 63714 40844
rect 63756 40804 63796 40844
rect 63838 40804 63878 40844
rect 63920 40804 63960 40844
rect 78712 40804 78752 40844
rect 78794 40804 78834 40844
rect 78876 40804 78916 40844
rect 78958 40804 78998 40844
rect 79040 40804 79080 40844
rect 93832 40804 93872 40844
rect 93914 40804 93954 40844
rect 93996 40804 94036 40844
rect 94078 40804 94118 40844
rect 94160 40804 94200 40844
rect 4352 40048 4392 40088
rect 4434 40048 4474 40088
rect 4516 40048 4556 40088
rect 4598 40048 4638 40088
rect 4680 40048 4720 40088
rect 19472 40048 19512 40088
rect 19554 40048 19594 40088
rect 19636 40048 19676 40088
rect 19718 40048 19758 40088
rect 19800 40048 19840 40088
rect 34592 40048 34632 40088
rect 34674 40048 34714 40088
rect 34756 40048 34796 40088
rect 34838 40048 34878 40088
rect 34920 40048 34960 40088
rect 49712 40048 49752 40088
rect 49794 40048 49834 40088
rect 49876 40048 49916 40088
rect 49958 40048 49998 40088
rect 50040 40048 50080 40088
rect 64832 40048 64872 40088
rect 64914 40048 64954 40088
rect 64996 40048 65036 40088
rect 65078 40048 65118 40088
rect 65160 40048 65200 40088
rect 79952 40048 79992 40088
rect 80034 40048 80074 40088
rect 80116 40048 80156 40088
rect 80198 40048 80238 40088
rect 80280 40048 80320 40088
rect 95072 40048 95112 40088
rect 95154 40048 95194 40088
rect 95236 40048 95276 40088
rect 95318 40048 95358 40088
rect 95400 40048 95440 40088
rect 3112 39292 3152 39332
rect 3194 39292 3234 39332
rect 3276 39292 3316 39332
rect 3358 39292 3398 39332
rect 3440 39292 3480 39332
rect 18232 39292 18272 39332
rect 18314 39292 18354 39332
rect 18396 39292 18436 39332
rect 18478 39292 18518 39332
rect 18560 39292 18600 39332
rect 33352 39292 33392 39332
rect 33434 39292 33474 39332
rect 33516 39292 33556 39332
rect 33598 39292 33638 39332
rect 33680 39292 33720 39332
rect 48472 39292 48512 39332
rect 48554 39292 48594 39332
rect 48636 39292 48676 39332
rect 48718 39292 48758 39332
rect 48800 39292 48840 39332
rect 63592 39292 63632 39332
rect 63674 39292 63714 39332
rect 63756 39292 63796 39332
rect 63838 39292 63878 39332
rect 63920 39292 63960 39332
rect 78712 39292 78752 39332
rect 78794 39292 78834 39332
rect 78876 39292 78916 39332
rect 78958 39292 78998 39332
rect 79040 39292 79080 39332
rect 93832 39292 93872 39332
rect 93914 39292 93954 39332
rect 93996 39292 94036 39332
rect 94078 39292 94118 39332
rect 94160 39292 94200 39332
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 95072 38536 95112 38576
rect 95154 38536 95194 38576
rect 95236 38536 95276 38576
rect 95318 38536 95358 38576
rect 95400 38536 95440 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 93832 37780 93872 37820
rect 93914 37780 93954 37820
rect 93996 37780 94036 37820
rect 94078 37780 94118 37820
rect 94160 37780 94200 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 95072 37024 95112 37064
rect 95154 37024 95194 37064
rect 95236 37024 95276 37064
rect 95318 37024 95358 37064
rect 95400 37024 95440 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 93832 36268 93872 36308
rect 93914 36268 93954 36308
rect 93996 36268 94036 36308
rect 94078 36268 94118 36308
rect 94160 36268 94200 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 95072 35512 95112 35552
rect 95154 35512 95194 35552
rect 95236 35512 95276 35552
rect 95318 35512 95358 35552
rect 95400 35512 95440 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 93832 34756 93872 34796
rect 93914 34756 93954 34796
rect 93996 34756 94036 34796
rect 94078 34756 94118 34796
rect 94160 34756 94200 34796
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 95072 34000 95112 34040
rect 95154 34000 95194 34040
rect 95236 34000 95276 34040
rect 95318 34000 95358 34040
rect 95400 34000 95440 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 93832 33244 93872 33284
rect 93914 33244 93954 33284
rect 93996 33244 94036 33284
rect 94078 33244 94118 33284
rect 94160 33244 94200 33284
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 95072 32488 95112 32528
rect 95154 32488 95194 32528
rect 95236 32488 95276 32528
rect 95318 32488 95358 32528
rect 95400 32488 95440 32528
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 93832 31732 93872 31772
rect 93914 31732 93954 31772
rect 93996 31732 94036 31772
rect 94078 31732 94118 31772
rect 94160 31732 94200 31772
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 95072 30976 95112 31016
rect 95154 30976 95194 31016
rect 95236 30976 95276 31016
rect 95318 30976 95358 31016
rect 95400 30976 95440 31016
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 93832 30220 93872 30260
rect 93914 30220 93954 30260
rect 93996 30220 94036 30260
rect 94078 30220 94118 30260
rect 94160 30220 94200 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 95072 29464 95112 29504
rect 95154 29464 95194 29504
rect 95236 29464 95276 29504
rect 95318 29464 95358 29504
rect 95400 29464 95440 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 93832 28708 93872 28748
rect 93914 28708 93954 28748
rect 93996 28708 94036 28748
rect 94078 28708 94118 28748
rect 94160 28708 94200 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 95072 27952 95112 27992
rect 95154 27952 95194 27992
rect 95236 27952 95276 27992
rect 95318 27952 95358 27992
rect 95400 27952 95440 27992
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 93832 27196 93872 27236
rect 93914 27196 93954 27236
rect 93996 27196 94036 27236
rect 94078 27196 94118 27236
rect 94160 27196 94200 27236
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 95072 26440 95112 26480
rect 95154 26440 95194 26480
rect 95236 26440 95276 26480
rect 95318 26440 95358 26480
rect 95400 26440 95440 26480
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 93832 25684 93872 25724
rect 93914 25684 93954 25724
rect 93996 25684 94036 25724
rect 94078 25684 94118 25724
rect 94160 25684 94200 25724
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 95072 24928 95112 24968
rect 95154 24928 95194 24968
rect 95236 24928 95276 24968
rect 95318 24928 95358 24968
rect 95400 24928 95440 24968
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 63592 24172 63632 24212
rect 63674 24172 63714 24212
rect 63756 24172 63796 24212
rect 63838 24172 63878 24212
rect 63920 24172 63960 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 93832 24172 93872 24212
rect 93914 24172 93954 24212
rect 93996 24172 94036 24212
rect 94078 24172 94118 24212
rect 94160 24172 94200 24212
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 64832 23416 64872 23456
rect 64914 23416 64954 23456
rect 64996 23416 65036 23456
rect 65078 23416 65118 23456
rect 65160 23416 65200 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 95072 23416 95112 23456
rect 95154 23416 95194 23456
rect 95236 23416 95276 23456
rect 95318 23416 95358 23456
rect 95400 23416 95440 23456
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 63592 22660 63632 22700
rect 63674 22660 63714 22700
rect 63756 22660 63796 22700
rect 63838 22660 63878 22700
rect 63920 22660 63960 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 93832 22660 93872 22700
rect 93914 22660 93954 22700
rect 93996 22660 94036 22700
rect 94078 22660 94118 22700
rect 94160 22660 94200 22700
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 64832 21904 64872 21944
rect 64914 21904 64954 21944
rect 64996 21904 65036 21944
rect 65078 21904 65118 21944
rect 65160 21904 65200 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 63592 21148 63632 21188
rect 63674 21148 63714 21188
rect 63756 21148 63796 21188
rect 63838 21148 63878 21188
rect 63920 21148 63960 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 64832 20392 64872 20432
rect 64914 20392 64954 20432
rect 64996 20392 65036 20432
rect 65078 20392 65118 20432
rect 65160 20392 65200 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 63592 19636 63632 19676
rect 63674 19636 63714 19676
rect 63756 19636 63796 19676
rect 63838 19636 63878 19676
rect 63920 19636 63960 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 64832 18880 64872 18920
rect 64914 18880 64954 18920
rect 64996 18880 65036 18920
rect 65078 18880 65118 18920
rect 65160 18880 65200 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 95072 18880 95112 18920
rect 95154 18880 95194 18920
rect 95236 18880 95276 18920
rect 95318 18880 95358 18920
rect 95400 18880 95440 18920
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 63592 18124 63632 18164
rect 63674 18124 63714 18164
rect 63756 18124 63796 18164
rect 63838 18124 63878 18164
rect 63920 18124 63960 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 93832 18124 93872 18164
rect 93914 18124 93954 18164
rect 93996 18124 94036 18164
rect 94078 18124 94118 18164
rect 94160 18124 94200 18164
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 64832 17368 64872 17408
rect 64914 17368 64954 17408
rect 64996 17368 65036 17408
rect 65078 17368 65118 17408
rect 65160 17368 65200 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 95072 17368 95112 17408
rect 95154 17368 95194 17408
rect 95236 17368 95276 17408
rect 95318 17368 95358 17408
rect 95400 17368 95440 17408
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 63592 16612 63632 16652
rect 63674 16612 63714 16652
rect 63756 16612 63796 16652
rect 63838 16612 63878 16652
rect 63920 16612 63960 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 93832 16612 93872 16652
rect 93914 16612 93954 16652
rect 93996 16612 94036 16652
rect 94078 16612 94118 16652
rect 94160 16612 94200 16652
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 64832 15856 64872 15896
rect 64914 15856 64954 15896
rect 64996 15856 65036 15896
rect 65078 15856 65118 15896
rect 65160 15856 65200 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 95072 15856 95112 15896
rect 95154 15856 95194 15896
rect 95236 15856 95276 15896
rect 95318 15856 95358 15896
rect 95400 15856 95440 15896
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 93832 15100 93872 15140
rect 93914 15100 93954 15140
rect 93996 15100 94036 15140
rect 94078 15100 94118 15140
rect 94160 15100 94200 15140
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 95072 14344 95112 14384
rect 95154 14344 95194 14384
rect 95236 14344 95276 14384
rect 95318 14344 95358 14384
rect 95400 14344 95440 14384
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 93832 13588 93872 13628
rect 93914 13588 93954 13628
rect 93996 13588 94036 13628
rect 94078 13588 94118 13628
rect 94160 13588 94200 13628
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 95072 12832 95112 12872
rect 95154 12832 95194 12872
rect 95236 12832 95276 12872
rect 95318 12832 95358 12872
rect 95400 12832 95440 12872
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 93832 12076 93872 12116
rect 93914 12076 93954 12116
rect 93996 12076 94036 12116
rect 94078 12076 94118 12116
rect 94160 12076 94200 12116
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 95072 11320 95112 11360
rect 95154 11320 95194 11360
rect 95236 11320 95276 11360
rect 95318 11320 95358 11360
rect 95400 11320 95440 11360
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 93832 10564 93872 10604
rect 93914 10564 93954 10604
rect 93996 10564 94036 10604
rect 94078 10564 94118 10604
rect 94160 10564 94200 10604
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 95072 9808 95112 9848
rect 95154 9808 95194 9848
rect 95236 9808 95276 9848
rect 95318 9808 95358 9848
rect 95400 9808 95440 9848
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 93832 9052 93872 9092
rect 93914 9052 93954 9092
rect 93996 9052 94036 9092
rect 94078 9052 94118 9092
rect 94160 9052 94200 9092
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 95072 8296 95112 8336
rect 95154 8296 95194 8336
rect 95236 8296 95276 8336
rect 95318 8296 95358 8336
rect 95400 8296 95440 8336
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 93832 7540 93872 7580
rect 93914 7540 93954 7580
rect 93996 7540 94036 7580
rect 94078 7540 94118 7580
rect 94160 7540 94200 7580
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 95072 6784 95112 6824
rect 95154 6784 95194 6824
rect 95236 6784 95276 6824
rect 95318 6784 95358 6824
rect 95400 6784 95440 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 93832 6028 93872 6068
rect 93914 6028 93954 6068
rect 93996 6028 94036 6068
rect 94078 6028 94118 6068
rect 94160 6028 94200 6068
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 95072 5272 95112 5312
rect 95154 5272 95194 5312
rect 95236 5272 95276 5312
rect 95318 5272 95358 5312
rect 95400 5272 95440 5312
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 93832 4516 93872 4556
rect 93914 4516 93954 4556
rect 93996 4516 94036 4556
rect 94078 4516 94118 4556
rect 94160 4516 94200 4556
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 95072 3760 95112 3800
rect 95154 3760 95194 3800
rect 95236 3760 95276 3800
rect 95318 3760 95358 3800
rect 95400 3760 95440 3800
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 93832 3004 93872 3044
rect 93914 3004 93954 3044
rect 93996 3004 94036 3044
rect 94078 3004 94118 3044
rect 94160 3004 94200 3044
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 95072 2248 95112 2288
rect 95154 2248 95194 2288
rect 95236 2248 95276 2288
rect 95318 2248 95358 2288
rect 95400 2248 95440 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 93832 1492 93872 1532
rect 93914 1492 93954 1532
rect 93996 1492 94036 1532
rect 94078 1492 94118 1532
rect 94160 1492 94200 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
rect 95072 736 95112 776
rect 95154 736 95194 776
rect 95236 736 95276 776
rect 95318 736 95358 776
rect 95400 736 95440 776
<< metal4 >>
rect 3112 81668 3480 81677
rect 3152 81628 3194 81668
rect 3234 81628 3276 81668
rect 3316 81628 3358 81668
rect 3398 81628 3440 81668
rect 3112 81619 3480 81628
rect 18232 81668 18600 81677
rect 18272 81628 18314 81668
rect 18354 81628 18396 81668
rect 18436 81628 18478 81668
rect 18518 81628 18560 81668
rect 18232 81619 18600 81628
rect 33352 81668 33720 81677
rect 33392 81628 33434 81668
rect 33474 81628 33516 81668
rect 33556 81628 33598 81668
rect 33638 81628 33680 81668
rect 33352 81619 33720 81628
rect 48472 81668 48840 81677
rect 48512 81628 48554 81668
rect 48594 81628 48636 81668
rect 48676 81628 48718 81668
rect 48758 81628 48800 81668
rect 48472 81619 48840 81628
rect 63592 81668 63960 81677
rect 63632 81628 63674 81668
rect 63714 81628 63756 81668
rect 63796 81628 63838 81668
rect 63878 81628 63920 81668
rect 63592 81619 63960 81628
rect 78712 81668 79080 81677
rect 78752 81628 78794 81668
rect 78834 81628 78876 81668
rect 78916 81628 78958 81668
rect 78998 81628 79040 81668
rect 78712 81619 79080 81628
rect 93832 81668 94200 81677
rect 93872 81628 93914 81668
rect 93954 81628 93996 81668
rect 94036 81628 94078 81668
rect 94118 81628 94160 81668
rect 93832 81619 94200 81628
rect 4352 80912 4720 80921
rect 4392 80872 4434 80912
rect 4474 80872 4516 80912
rect 4556 80872 4598 80912
rect 4638 80872 4680 80912
rect 4352 80863 4720 80872
rect 19472 80912 19840 80921
rect 19512 80872 19554 80912
rect 19594 80872 19636 80912
rect 19676 80872 19718 80912
rect 19758 80872 19800 80912
rect 19472 80863 19840 80872
rect 34592 80912 34960 80921
rect 34632 80872 34674 80912
rect 34714 80872 34756 80912
rect 34796 80872 34838 80912
rect 34878 80872 34920 80912
rect 34592 80863 34960 80872
rect 49712 80912 50080 80921
rect 49752 80872 49794 80912
rect 49834 80872 49876 80912
rect 49916 80872 49958 80912
rect 49998 80872 50040 80912
rect 49712 80863 50080 80872
rect 64832 80912 65200 80921
rect 64872 80872 64914 80912
rect 64954 80872 64996 80912
rect 65036 80872 65078 80912
rect 65118 80872 65160 80912
rect 64832 80863 65200 80872
rect 79952 80912 80320 80921
rect 79992 80872 80034 80912
rect 80074 80872 80116 80912
rect 80156 80872 80198 80912
rect 80238 80872 80280 80912
rect 79952 80863 80320 80872
rect 95072 80912 95440 80921
rect 95112 80872 95154 80912
rect 95194 80872 95236 80912
rect 95276 80872 95318 80912
rect 95358 80872 95400 80912
rect 95072 80863 95440 80872
rect 3112 80156 3480 80165
rect 3152 80116 3194 80156
rect 3234 80116 3276 80156
rect 3316 80116 3358 80156
rect 3398 80116 3440 80156
rect 3112 80107 3480 80116
rect 18232 80156 18600 80165
rect 18272 80116 18314 80156
rect 18354 80116 18396 80156
rect 18436 80116 18478 80156
rect 18518 80116 18560 80156
rect 18232 80107 18600 80116
rect 33352 80156 33720 80165
rect 33392 80116 33434 80156
rect 33474 80116 33516 80156
rect 33556 80116 33598 80156
rect 33638 80116 33680 80156
rect 33352 80107 33720 80116
rect 48472 80156 48840 80165
rect 48512 80116 48554 80156
rect 48594 80116 48636 80156
rect 48676 80116 48718 80156
rect 48758 80116 48800 80156
rect 48472 80107 48840 80116
rect 63592 80156 63960 80165
rect 63632 80116 63674 80156
rect 63714 80116 63756 80156
rect 63796 80116 63838 80156
rect 63878 80116 63920 80156
rect 63592 80107 63960 80116
rect 78712 80156 79080 80165
rect 78752 80116 78794 80156
rect 78834 80116 78876 80156
rect 78916 80116 78958 80156
rect 78998 80116 79040 80156
rect 78712 80107 79080 80116
rect 93832 80156 94200 80165
rect 93872 80116 93914 80156
rect 93954 80116 93996 80156
rect 94036 80116 94078 80156
rect 94118 80116 94160 80156
rect 93832 80107 94200 80116
rect 4352 79400 4720 79409
rect 4392 79360 4434 79400
rect 4474 79360 4516 79400
rect 4556 79360 4598 79400
rect 4638 79360 4680 79400
rect 4352 79351 4720 79360
rect 19472 79400 19840 79409
rect 19512 79360 19554 79400
rect 19594 79360 19636 79400
rect 19676 79360 19718 79400
rect 19758 79360 19800 79400
rect 19472 79351 19840 79360
rect 34592 79400 34960 79409
rect 34632 79360 34674 79400
rect 34714 79360 34756 79400
rect 34796 79360 34838 79400
rect 34878 79360 34920 79400
rect 34592 79351 34960 79360
rect 49712 79400 50080 79409
rect 49752 79360 49794 79400
rect 49834 79360 49876 79400
rect 49916 79360 49958 79400
rect 49998 79360 50040 79400
rect 49712 79351 50080 79360
rect 64832 79400 65200 79409
rect 64872 79360 64914 79400
rect 64954 79360 64996 79400
rect 65036 79360 65078 79400
rect 65118 79360 65160 79400
rect 64832 79351 65200 79360
rect 79952 79400 80320 79409
rect 79992 79360 80034 79400
rect 80074 79360 80116 79400
rect 80156 79360 80198 79400
rect 80238 79360 80280 79400
rect 79952 79351 80320 79360
rect 95072 79400 95440 79409
rect 95112 79360 95154 79400
rect 95194 79360 95236 79400
rect 95276 79360 95318 79400
rect 95358 79360 95400 79400
rect 95072 79351 95440 79360
rect 3112 78644 3480 78653
rect 3152 78604 3194 78644
rect 3234 78604 3276 78644
rect 3316 78604 3358 78644
rect 3398 78604 3440 78644
rect 3112 78595 3480 78604
rect 18232 78644 18600 78653
rect 18272 78604 18314 78644
rect 18354 78604 18396 78644
rect 18436 78604 18478 78644
rect 18518 78604 18560 78644
rect 18232 78595 18600 78604
rect 33352 78644 33720 78653
rect 33392 78604 33434 78644
rect 33474 78604 33516 78644
rect 33556 78604 33598 78644
rect 33638 78604 33680 78644
rect 33352 78595 33720 78604
rect 48472 78644 48840 78653
rect 48512 78604 48554 78644
rect 48594 78604 48636 78644
rect 48676 78604 48718 78644
rect 48758 78604 48800 78644
rect 48472 78595 48840 78604
rect 63592 78644 63960 78653
rect 63632 78604 63674 78644
rect 63714 78604 63756 78644
rect 63796 78604 63838 78644
rect 63878 78604 63920 78644
rect 63592 78595 63960 78604
rect 78712 78644 79080 78653
rect 78752 78604 78794 78644
rect 78834 78604 78876 78644
rect 78916 78604 78958 78644
rect 78998 78604 79040 78644
rect 78712 78595 79080 78604
rect 93832 78644 94200 78653
rect 93872 78604 93914 78644
rect 93954 78604 93996 78644
rect 94036 78604 94078 78644
rect 94118 78604 94160 78644
rect 93832 78595 94200 78604
rect 4352 77888 4720 77897
rect 4392 77848 4434 77888
rect 4474 77848 4516 77888
rect 4556 77848 4598 77888
rect 4638 77848 4680 77888
rect 4352 77839 4720 77848
rect 19472 77888 19840 77897
rect 19512 77848 19554 77888
rect 19594 77848 19636 77888
rect 19676 77848 19718 77888
rect 19758 77848 19800 77888
rect 19472 77839 19840 77848
rect 34592 77888 34960 77897
rect 34632 77848 34674 77888
rect 34714 77848 34756 77888
rect 34796 77848 34838 77888
rect 34878 77848 34920 77888
rect 34592 77839 34960 77848
rect 49712 77888 50080 77897
rect 49752 77848 49794 77888
rect 49834 77848 49876 77888
rect 49916 77848 49958 77888
rect 49998 77848 50040 77888
rect 49712 77839 50080 77848
rect 64832 77888 65200 77897
rect 64872 77848 64914 77888
rect 64954 77848 64996 77888
rect 65036 77848 65078 77888
rect 65118 77848 65160 77888
rect 64832 77839 65200 77848
rect 79952 77888 80320 77897
rect 79992 77848 80034 77888
rect 80074 77848 80116 77888
rect 80156 77848 80198 77888
rect 80238 77848 80280 77888
rect 79952 77839 80320 77848
rect 95072 77888 95440 77897
rect 95112 77848 95154 77888
rect 95194 77848 95236 77888
rect 95276 77848 95318 77888
rect 95358 77848 95400 77888
rect 95072 77839 95440 77848
rect 3112 77132 3480 77141
rect 3152 77092 3194 77132
rect 3234 77092 3276 77132
rect 3316 77092 3358 77132
rect 3398 77092 3440 77132
rect 3112 77083 3480 77092
rect 18232 77132 18600 77141
rect 18272 77092 18314 77132
rect 18354 77092 18396 77132
rect 18436 77092 18478 77132
rect 18518 77092 18560 77132
rect 18232 77083 18600 77092
rect 33352 77132 33720 77141
rect 33392 77092 33434 77132
rect 33474 77092 33516 77132
rect 33556 77092 33598 77132
rect 33638 77092 33680 77132
rect 33352 77083 33720 77092
rect 48472 77132 48840 77141
rect 48512 77092 48554 77132
rect 48594 77092 48636 77132
rect 48676 77092 48718 77132
rect 48758 77092 48800 77132
rect 48472 77083 48840 77092
rect 63592 77132 63960 77141
rect 63632 77092 63674 77132
rect 63714 77092 63756 77132
rect 63796 77092 63838 77132
rect 63878 77092 63920 77132
rect 63592 77083 63960 77092
rect 78712 77132 79080 77141
rect 78752 77092 78794 77132
rect 78834 77092 78876 77132
rect 78916 77092 78958 77132
rect 78998 77092 79040 77132
rect 78712 77083 79080 77092
rect 93832 77132 94200 77141
rect 93872 77092 93914 77132
rect 93954 77092 93996 77132
rect 94036 77092 94078 77132
rect 94118 77092 94160 77132
rect 93832 77083 94200 77092
rect 4352 76376 4720 76385
rect 4392 76336 4434 76376
rect 4474 76336 4516 76376
rect 4556 76336 4598 76376
rect 4638 76336 4680 76376
rect 4352 76327 4720 76336
rect 19472 76376 19840 76385
rect 19512 76336 19554 76376
rect 19594 76336 19636 76376
rect 19676 76336 19718 76376
rect 19758 76336 19800 76376
rect 19472 76327 19840 76336
rect 34592 76376 34960 76385
rect 34632 76336 34674 76376
rect 34714 76336 34756 76376
rect 34796 76336 34838 76376
rect 34878 76336 34920 76376
rect 34592 76327 34960 76336
rect 49712 76376 50080 76385
rect 49752 76336 49794 76376
rect 49834 76336 49876 76376
rect 49916 76336 49958 76376
rect 49998 76336 50040 76376
rect 49712 76327 50080 76336
rect 64832 76376 65200 76385
rect 64872 76336 64914 76376
rect 64954 76336 64996 76376
rect 65036 76336 65078 76376
rect 65118 76336 65160 76376
rect 64832 76327 65200 76336
rect 79952 76376 80320 76385
rect 79992 76336 80034 76376
rect 80074 76336 80116 76376
rect 80156 76336 80198 76376
rect 80238 76336 80280 76376
rect 79952 76327 80320 76336
rect 95072 76376 95440 76385
rect 95112 76336 95154 76376
rect 95194 76336 95236 76376
rect 95276 76336 95318 76376
rect 95358 76336 95400 76376
rect 95072 76327 95440 76336
rect 3112 75620 3480 75629
rect 3152 75580 3194 75620
rect 3234 75580 3276 75620
rect 3316 75580 3358 75620
rect 3398 75580 3440 75620
rect 3112 75571 3480 75580
rect 18232 75620 18600 75629
rect 18272 75580 18314 75620
rect 18354 75580 18396 75620
rect 18436 75580 18478 75620
rect 18518 75580 18560 75620
rect 18232 75571 18600 75580
rect 33352 75620 33720 75629
rect 33392 75580 33434 75620
rect 33474 75580 33516 75620
rect 33556 75580 33598 75620
rect 33638 75580 33680 75620
rect 33352 75571 33720 75580
rect 48472 75620 48840 75629
rect 48512 75580 48554 75620
rect 48594 75580 48636 75620
rect 48676 75580 48718 75620
rect 48758 75580 48800 75620
rect 48472 75571 48840 75580
rect 63592 75620 63960 75629
rect 63632 75580 63674 75620
rect 63714 75580 63756 75620
rect 63796 75580 63838 75620
rect 63878 75580 63920 75620
rect 63592 75571 63960 75580
rect 78712 75620 79080 75629
rect 78752 75580 78794 75620
rect 78834 75580 78876 75620
rect 78916 75580 78958 75620
rect 78998 75580 79040 75620
rect 78712 75571 79080 75580
rect 93832 75620 94200 75629
rect 93872 75580 93914 75620
rect 93954 75580 93996 75620
rect 94036 75580 94078 75620
rect 94118 75580 94160 75620
rect 93832 75571 94200 75580
rect 4352 74864 4720 74873
rect 4392 74824 4434 74864
rect 4474 74824 4516 74864
rect 4556 74824 4598 74864
rect 4638 74824 4680 74864
rect 4352 74815 4720 74824
rect 19472 74864 19840 74873
rect 19512 74824 19554 74864
rect 19594 74824 19636 74864
rect 19676 74824 19718 74864
rect 19758 74824 19800 74864
rect 19472 74815 19840 74824
rect 34592 74864 34960 74873
rect 34632 74824 34674 74864
rect 34714 74824 34756 74864
rect 34796 74824 34838 74864
rect 34878 74824 34920 74864
rect 34592 74815 34960 74824
rect 49712 74864 50080 74873
rect 49752 74824 49794 74864
rect 49834 74824 49876 74864
rect 49916 74824 49958 74864
rect 49998 74824 50040 74864
rect 49712 74815 50080 74824
rect 64832 74864 65200 74873
rect 64872 74824 64914 74864
rect 64954 74824 64996 74864
rect 65036 74824 65078 74864
rect 65118 74824 65160 74864
rect 64832 74815 65200 74824
rect 79952 74864 80320 74873
rect 79992 74824 80034 74864
rect 80074 74824 80116 74864
rect 80156 74824 80198 74864
rect 80238 74824 80280 74864
rect 79952 74815 80320 74824
rect 95072 74864 95440 74873
rect 95112 74824 95154 74864
rect 95194 74824 95236 74864
rect 95276 74824 95318 74864
rect 95358 74824 95400 74864
rect 95072 74815 95440 74824
rect 3112 74108 3480 74117
rect 3152 74068 3194 74108
rect 3234 74068 3276 74108
rect 3316 74068 3358 74108
rect 3398 74068 3440 74108
rect 3112 74059 3480 74068
rect 18232 74108 18600 74117
rect 18272 74068 18314 74108
rect 18354 74068 18396 74108
rect 18436 74068 18478 74108
rect 18518 74068 18560 74108
rect 18232 74059 18600 74068
rect 33352 74108 33720 74117
rect 33392 74068 33434 74108
rect 33474 74068 33516 74108
rect 33556 74068 33598 74108
rect 33638 74068 33680 74108
rect 33352 74059 33720 74068
rect 48472 74108 48840 74117
rect 48512 74068 48554 74108
rect 48594 74068 48636 74108
rect 48676 74068 48718 74108
rect 48758 74068 48800 74108
rect 48472 74059 48840 74068
rect 63592 74108 63960 74117
rect 63632 74068 63674 74108
rect 63714 74068 63756 74108
rect 63796 74068 63838 74108
rect 63878 74068 63920 74108
rect 63592 74059 63960 74068
rect 78712 74108 79080 74117
rect 78752 74068 78794 74108
rect 78834 74068 78876 74108
rect 78916 74068 78958 74108
rect 78998 74068 79040 74108
rect 78712 74059 79080 74068
rect 93832 74108 94200 74117
rect 93872 74068 93914 74108
rect 93954 74068 93996 74108
rect 94036 74068 94078 74108
rect 94118 74068 94160 74108
rect 93832 74059 94200 74068
rect 4352 73352 4720 73361
rect 4392 73312 4434 73352
rect 4474 73312 4516 73352
rect 4556 73312 4598 73352
rect 4638 73312 4680 73352
rect 4352 73303 4720 73312
rect 19472 73352 19840 73361
rect 19512 73312 19554 73352
rect 19594 73312 19636 73352
rect 19676 73312 19718 73352
rect 19758 73312 19800 73352
rect 19472 73303 19840 73312
rect 34592 73352 34960 73361
rect 34632 73312 34674 73352
rect 34714 73312 34756 73352
rect 34796 73312 34838 73352
rect 34878 73312 34920 73352
rect 34592 73303 34960 73312
rect 49712 73352 50080 73361
rect 49752 73312 49794 73352
rect 49834 73312 49876 73352
rect 49916 73312 49958 73352
rect 49998 73312 50040 73352
rect 49712 73303 50080 73312
rect 64832 73352 65200 73361
rect 64872 73312 64914 73352
rect 64954 73312 64996 73352
rect 65036 73312 65078 73352
rect 65118 73312 65160 73352
rect 64832 73303 65200 73312
rect 79952 73352 80320 73361
rect 79992 73312 80034 73352
rect 80074 73312 80116 73352
rect 80156 73312 80198 73352
rect 80238 73312 80280 73352
rect 79952 73303 80320 73312
rect 95072 73352 95440 73361
rect 95112 73312 95154 73352
rect 95194 73312 95236 73352
rect 95276 73312 95318 73352
rect 95358 73312 95400 73352
rect 95072 73303 95440 73312
rect 3112 72596 3480 72605
rect 3152 72556 3194 72596
rect 3234 72556 3276 72596
rect 3316 72556 3358 72596
rect 3398 72556 3440 72596
rect 3112 72547 3480 72556
rect 18232 72596 18600 72605
rect 18272 72556 18314 72596
rect 18354 72556 18396 72596
rect 18436 72556 18478 72596
rect 18518 72556 18560 72596
rect 18232 72547 18600 72556
rect 33352 72596 33720 72605
rect 33392 72556 33434 72596
rect 33474 72556 33516 72596
rect 33556 72556 33598 72596
rect 33638 72556 33680 72596
rect 33352 72547 33720 72556
rect 48472 72596 48840 72605
rect 48512 72556 48554 72596
rect 48594 72556 48636 72596
rect 48676 72556 48718 72596
rect 48758 72556 48800 72596
rect 48472 72547 48840 72556
rect 63592 72596 63960 72605
rect 63632 72556 63674 72596
rect 63714 72556 63756 72596
rect 63796 72556 63838 72596
rect 63878 72556 63920 72596
rect 63592 72547 63960 72556
rect 78712 72596 79080 72605
rect 78752 72556 78794 72596
rect 78834 72556 78876 72596
rect 78916 72556 78958 72596
rect 78998 72556 79040 72596
rect 78712 72547 79080 72556
rect 93832 72596 94200 72605
rect 93872 72556 93914 72596
rect 93954 72556 93996 72596
rect 94036 72556 94078 72596
rect 94118 72556 94160 72596
rect 93832 72547 94200 72556
rect 4352 71840 4720 71849
rect 4392 71800 4434 71840
rect 4474 71800 4516 71840
rect 4556 71800 4598 71840
rect 4638 71800 4680 71840
rect 4352 71791 4720 71800
rect 19472 71840 19840 71849
rect 19512 71800 19554 71840
rect 19594 71800 19636 71840
rect 19676 71800 19718 71840
rect 19758 71800 19800 71840
rect 19472 71791 19840 71800
rect 34592 71840 34960 71849
rect 34632 71800 34674 71840
rect 34714 71800 34756 71840
rect 34796 71800 34838 71840
rect 34878 71800 34920 71840
rect 34592 71791 34960 71800
rect 49712 71840 50080 71849
rect 49752 71800 49794 71840
rect 49834 71800 49876 71840
rect 49916 71800 49958 71840
rect 49998 71800 50040 71840
rect 49712 71791 50080 71800
rect 64832 71840 65200 71849
rect 64872 71800 64914 71840
rect 64954 71800 64996 71840
rect 65036 71800 65078 71840
rect 65118 71800 65160 71840
rect 64832 71791 65200 71800
rect 79952 71840 80320 71849
rect 79992 71800 80034 71840
rect 80074 71800 80116 71840
rect 80156 71800 80198 71840
rect 80238 71800 80280 71840
rect 79952 71791 80320 71800
rect 95072 71840 95440 71849
rect 95112 71800 95154 71840
rect 95194 71800 95236 71840
rect 95276 71800 95318 71840
rect 95358 71800 95400 71840
rect 95072 71791 95440 71800
rect 3112 71084 3480 71093
rect 3152 71044 3194 71084
rect 3234 71044 3276 71084
rect 3316 71044 3358 71084
rect 3398 71044 3440 71084
rect 3112 71035 3480 71044
rect 18232 71084 18600 71093
rect 18272 71044 18314 71084
rect 18354 71044 18396 71084
rect 18436 71044 18478 71084
rect 18518 71044 18560 71084
rect 18232 71035 18600 71044
rect 33352 71084 33720 71093
rect 33392 71044 33434 71084
rect 33474 71044 33516 71084
rect 33556 71044 33598 71084
rect 33638 71044 33680 71084
rect 33352 71035 33720 71044
rect 48472 71084 48840 71093
rect 48512 71044 48554 71084
rect 48594 71044 48636 71084
rect 48676 71044 48718 71084
rect 48758 71044 48800 71084
rect 48472 71035 48840 71044
rect 63592 71084 63960 71093
rect 63632 71044 63674 71084
rect 63714 71044 63756 71084
rect 63796 71044 63838 71084
rect 63878 71044 63920 71084
rect 63592 71035 63960 71044
rect 78712 71084 79080 71093
rect 78752 71044 78794 71084
rect 78834 71044 78876 71084
rect 78916 71044 78958 71084
rect 78998 71044 79040 71084
rect 78712 71035 79080 71044
rect 93832 71084 94200 71093
rect 93872 71044 93914 71084
rect 93954 71044 93996 71084
rect 94036 71044 94078 71084
rect 94118 71044 94160 71084
rect 93832 71035 94200 71044
rect 4352 70328 4720 70337
rect 4392 70288 4434 70328
rect 4474 70288 4516 70328
rect 4556 70288 4598 70328
rect 4638 70288 4680 70328
rect 4352 70279 4720 70288
rect 19472 70328 19840 70337
rect 19512 70288 19554 70328
rect 19594 70288 19636 70328
rect 19676 70288 19718 70328
rect 19758 70288 19800 70328
rect 19472 70279 19840 70288
rect 34592 70328 34960 70337
rect 34632 70288 34674 70328
rect 34714 70288 34756 70328
rect 34796 70288 34838 70328
rect 34878 70288 34920 70328
rect 34592 70279 34960 70288
rect 49712 70328 50080 70337
rect 49752 70288 49794 70328
rect 49834 70288 49876 70328
rect 49916 70288 49958 70328
rect 49998 70288 50040 70328
rect 49712 70279 50080 70288
rect 64832 70328 65200 70337
rect 64872 70288 64914 70328
rect 64954 70288 64996 70328
rect 65036 70288 65078 70328
rect 65118 70288 65160 70328
rect 64832 70279 65200 70288
rect 79952 70328 80320 70337
rect 79992 70288 80034 70328
rect 80074 70288 80116 70328
rect 80156 70288 80198 70328
rect 80238 70288 80280 70328
rect 79952 70279 80320 70288
rect 95072 70328 95440 70337
rect 95112 70288 95154 70328
rect 95194 70288 95236 70328
rect 95276 70288 95318 70328
rect 95358 70288 95400 70328
rect 95072 70279 95440 70288
rect 3112 69572 3480 69581
rect 3152 69532 3194 69572
rect 3234 69532 3276 69572
rect 3316 69532 3358 69572
rect 3398 69532 3440 69572
rect 3112 69523 3480 69532
rect 18232 69572 18600 69581
rect 18272 69532 18314 69572
rect 18354 69532 18396 69572
rect 18436 69532 18478 69572
rect 18518 69532 18560 69572
rect 18232 69523 18600 69532
rect 33352 69572 33720 69581
rect 33392 69532 33434 69572
rect 33474 69532 33516 69572
rect 33556 69532 33598 69572
rect 33638 69532 33680 69572
rect 33352 69523 33720 69532
rect 48472 69572 48840 69581
rect 48512 69532 48554 69572
rect 48594 69532 48636 69572
rect 48676 69532 48718 69572
rect 48758 69532 48800 69572
rect 48472 69523 48840 69532
rect 63592 69572 63960 69581
rect 63632 69532 63674 69572
rect 63714 69532 63756 69572
rect 63796 69532 63838 69572
rect 63878 69532 63920 69572
rect 63592 69523 63960 69532
rect 78712 69572 79080 69581
rect 78752 69532 78794 69572
rect 78834 69532 78876 69572
rect 78916 69532 78958 69572
rect 78998 69532 79040 69572
rect 78712 69523 79080 69532
rect 93832 69572 94200 69581
rect 93872 69532 93914 69572
rect 93954 69532 93996 69572
rect 94036 69532 94078 69572
rect 94118 69532 94160 69572
rect 93832 69523 94200 69532
rect 4352 68816 4720 68825
rect 4392 68776 4434 68816
rect 4474 68776 4516 68816
rect 4556 68776 4598 68816
rect 4638 68776 4680 68816
rect 4352 68767 4720 68776
rect 19472 68816 19840 68825
rect 19512 68776 19554 68816
rect 19594 68776 19636 68816
rect 19676 68776 19718 68816
rect 19758 68776 19800 68816
rect 19472 68767 19840 68776
rect 34592 68816 34960 68825
rect 34632 68776 34674 68816
rect 34714 68776 34756 68816
rect 34796 68776 34838 68816
rect 34878 68776 34920 68816
rect 34592 68767 34960 68776
rect 49712 68816 50080 68825
rect 49752 68776 49794 68816
rect 49834 68776 49876 68816
rect 49916 68776 49958 68816
rect 49998 68776 50040 68816
rect 49712 68767 50080 68776
rect 64832 68816 65200 68825
rect 64872 68776 64914 68816
rect 64954 68776 64996 68816
rect 65036 68776 65078 68816
rect 65118 68776 65160 68816
rect 64832 68767 65200 68776
rect 79952 68816 80320 68825
rect 79992 68776 80034 68816
rect 80074 68776 80116 68816
rect 80156 68776 80198 68816
rect 80238 68776 80280 68816
rect 79952 68767 80320 68776
rect 95072 68816 95440 68825
rect 95112 68776 95154 68816
rect 95194 68776 95236 68816
rect 95276 68776 95318 68816
rect 95358 68776 95400 68816
rect 95072 68767 95440 68776
rect 3112 68060 3480 68069
rect 3152 68020 3194 68060
rect 3234 68020 3276 68060
rect 3316 68020 3358 68060
rect 3398 68020 3440 68060
rect 3112 68011 3480 68020
rect 18232 68060 18600 68069
rect 18272 68020 18314 68060
rect 18354 68020 18396 68060
rect 18436 68020 18478 68060
rect 18518 68020 18560 68060
rect 18232 68011 18600 68020
rect 33352 68060 33720 68069
rect 33392 68020 33434 68060
rect 33474 68020 33516 68060
rect 33556 68020 33598 68060
rect 33638 68020 33680 68060
rect 33352 68011 33720 68020
rect 48472 68060 48840 68069
rect 48512 68020 48554 68060
rect 48594 68020 48636 68060
rect 48676 68020 48718 68060
rect 48758 68020 48800 68060
rect 48472 68011 48840 68020
rect 63592 68060 63960 68069
rect 63632 68020 63674 68060
rect 63714 68020 63756 68060
rect 63796 68020 63838 68060
rect 63878 68020 63920 68060
rect 63592 68011 63960 68020
rect 78712 68060 79080 68069
rect 78752 68020 78794 68060
rect 78834 68020 78876 68060
rect 78916 68020 78958 68060
rect 78998 68020 79040 68060
rect 78712 68011 79080 68020
rect 93832 68060 94200 68069
rect 93872 68020 93914 68060
rect 93954 68020 93996 68060
rect 94036 68020 94078 68060
rect 94118 68020 94160 68060
rect 93832 68011 94200 68020
rect 4352 67304 4720 67313
rect 4392 67264 4434 67304
rect 4474 67264 4516 67304
rect 4556 67264 4598 67304
rect 4638 67264 4680 67304
rect 4352 67255 4720 67264
rect 19472 67304 19840 67313
rect 19512 67264 19554 67304
rect 19594 67264 19636 67304
rect 19676 67264 19718 67304
rect 19758 67264 19800 67304
rect 19472 67255 19840 67264
rect 34592 67304 34960 67313
rect 34632 67264 34674 67304
rect 34714 67264 34756 67304
rect 34796 67264 34838 67304
rect 34878 67264 34920 67304
rect 34592 67255 34960 67264
rect 49712 67304 50080 67313
rect 49752 67264 49794 67304
rect 49834 67264 49876 67304
rect 49916 67264 49958 67304
rect 49998 67264 50040 67304
rect 49712 67255 50080 67264
rect 64832 67304 65200 67313
rect 64872 67264 64914 67304
rect 64954 67264 64996 67304
rect 65036 67264 65078 67304
rect 65118 67264 65160 67304
rect 64832 67255 65200 67264
rect 79952 67304 80320 67313
rect 79992 67264 80034 67304
rect 80074 67264 80116 67304
rect 80156 67264 80198 67304
rect 80238 67264 80280 67304
rect 79952 67255 80320 67264
rect 95072 67304 95440 67313
rect 95112 67264 95154 67304
rect 95194 67264 95236 67304
rect 95276 67264 95318 67304
rect 95358 67264 95400 67304
rect 95072 67255 95440 67264
rect 3112 66548 3480 66557
rect 3152 66508 3194 66548
rect 3234 66508 3276 66548
rect 3316 66508 3358 66548
rect 3398 66508 3440 66548
rect 3112 66499 3480 66508
rect 18232 66548 18600 66557
rect 18272 66508 18314 66548
rect 18354 66508 18396 66548
rect 18436 66508 18478 66548
rect 18518 66508 18560 66548
rect 18232 66499 18600 66508
rect 33352 66548 33720 66557
rect 33392 66508 33434 66548
rect 33474 66508 33516 66548
rect 33556 66508 33598 66548
rect 33638 66508 33680 66548
rect 33352 66499 33720 66508
rect 48472 66548 48840 66557
rect 48512 66508 48554 66548
rect 48594 66508 48636 66548
rect 48676 66508 48718 66548
rect 48758 66508 48800 66548
rect 48472 66499 48840 66508
rect 63592 66548 63960 66557
rect 63632 66508 63674 66548
rect 63714 66508 63756 66548
rect 63796 66508 63838 66548
rect 63878 66508 63920 66548
rect 63592 66499 63960 66508
rect 78712 66548 79080 66557
rect 78752 66508 78794 66548
rect 78834 66508 78876 66548
rect 78916 66508 78958 66548
rect 78998 66508 79040 66548
rect 78712 66499 79080 66508
rect 93832 66548 94200 66557
rect 93872 66508 93914 66548
rect 93954 66508 93996 66548
rect 94036 66508 94078 66548
rect 94118 66508 94160 66548
rect 93832 66499 94200 66508
rect 4352 65792 4720 65801
rect 4392 65752 4434 65792
rect 4474 65752 4516 65792
rect 4556 65752 4598 65792
rect 4638 65752 4680 65792
rect 4352 65743 4720 65752
rect 19472 65792 19840 65801
rect 19512 65752 19554 65792
rect 19594 65752 19636 65792
rect 19676 65752 19718 65792
rect 19758 65752 19800 65792
rect 19472 65743 19840 65752
rect 34592 65792 34960 65801
rect 34632 65752 34674 65792
rect 34714 65752 34756 65792
rect 34796 65752 34838 65792
rect 34878 65752 34920 65792
rect 34592 65743 34960 65752
rect 49712 65792 50080 65801
rect 49752 65752 49794 65792
rect 49834 65752 49876 65792
rect 49916 65752 49958 65792
rect 49998 65752 50040 65792
rect 49712 65743 50080 65752
rect 64832 65792 65200 65801
rect 64872 65752 64914 65792
rect 64954 65752 64996 65792
rect 65036 65752 65078 65792
rect 65118 65752 65160 65792
rect 64832 65743 65200 65752
rect 79952 65792 80320 65801
rect 79992 65752 80034 65792
rect 80074 65752 80116 65792
rect 80156 65752 80198 65792
rect 80238 65752 80280 65792
rect 79952 65743 80320 65752
rect 95072 65792 95440 65801
rect 95112 65752 95154 65792
rect 95194 65752 95236 65792
rect 95276 65752 95318 65792
rect 95358 65752 95400 65792
rect 95072 65743 95440 65752
rect 3112 65036 3480 65045
rect 3152 64996 3194 65036
rect 3234 64996 3276 65036
rect 3316 64996 3358 65036
rect 3398 64996 3440 65036
rect 3112 64987 3480 64996
rect 18232 65036 18600 65045
rect 18272 64996 18314 65036
rect 18354 64996 18396 65036
rect 18436 64996 18478 65036
rect 18518 64996 18560 65036
rect 18232 64987 18600 64996
rect 33352 65036 33720 65045
rect 33392 64996 33434 65036
rect 33474 64996 33516 65036
rect 33556 64996 33598 65036
rect 33638 64996 33680 65036
rect 33352 64987 33720 64996
rect 48472 65036 48840 65045
rect 48512 64996 48554 65036
rect 48594 64996 48636 65036
rect 48676 64996 48718 65036
rect 48758 64996 48800 65036
rect 48472 64987 48840 64996
rect 63592 65036 63960 65045
rect 63632 64996 63674 65036
rect 63714 64996 63756 65036
rect 63796 64996 63838 65036
rect 63878 64996 63920 65036
rect 63592 64987 63960 64996
rect 78712 65036 79080 65045
rect 78752 64996 78794 65036
rect 78834 64996 78876 65036
rect 78916 64996 78958 65036
rect 78998 64996 79040 65036
rect 78712 64987 79080 64996
rect 93832 65036 94200 65045
rect 93872 64996 93914 65036
rect 93954 64996 93996 65036
rect 94036 64996 94078 65036
rect 94118 64996 94160 65036
rect 93832 64987 94200 64996
rect 4352 64280 4720 64289
rect 4392 64240 4434 64280
rect 4474 64240 4516 64280
rect 4556 64240 4598 64280
rect 4638 64240 4680 64280
rect 4352 64231 4720 64240
rect 19472 64280 19840 64289
rect 19512 64240 19554 64280
rect 19594 64240 19636 64280
rect 19676 64240 19718 64280
rect 19758 64240 19800 64280
rect 19472 64231 19840 64240
rect 34592 64280 34960 64289
rect 34632 64240 34674 64280
rect 34714 64240 34756 64280
rect 34796 64240 34838 64280
rect 34878 64240 34920 64280
rect 34592 64231 34960 64240
rect 49712 64280 50080 64289
rect 49752 64240 49794 64280
rect 49834 64240 49876 64280
rect 49916 64240 49958 64280
rect 49998 64240 50040 64280
rect 49712 64231 50080 64240
rect 64832 64280 65200 64289
rect 64872 64240 64914 64280
rect 64954 64240 64996 64280
rect 65036 64240 65078 64280
rect 65118 64240 65160 64280
rect 64832 64231 65200 64240
rect 79952 64280 80320 64289
rect 79992 64240 80034 64280
rect 80074 64240 80116 64280
rect 80156 64240 80198 64280
rect 80238 64240 80280 64280
rect 79952 64231 80320 64240
rect 95072 64280 95440 64289
rect 95112 64240 95154 64280
rect 95194 64240 95236 64280
rect 95276 64240 95318 64280
rect 95358 64240 95400 64280
rect 95072 64231 95440 64240
rect 3112 63524 3480 63533
rect 3152 63484 3194 63524
rect 3234 63484 3276 63524
rect 3316 63484 3358 63524
rect 3398 63484 3440 63524
rect 3112 63475 3480 63484
rect 18232 63524 18600 63533
rect 18272 63484 18314 63524
rect 18354 63484 18396 63524
rect 18436 63484 18478 63524
rect 18518 63484 18560 63524
rect 18232 63475 18600 63484
rect 33352 63524 33720 63533
rect 33392 63484 33434 63524
rect 33474 63484 33516 63524
rect 33556 63484 33598 63524
rect 33638 63484 33680 63524
rect 33352 63475 33720 63484
rect 48472 63524 48840 63533
rect 48512 63484 48554 63524
rect 48594 63484 48636 63524
rect 48676 63484 48718 63524
rect 48758 63484 48800 63524
rect 48472 63475 48840 63484
rect 63592 63524 63960 63533
rect 63632 63484 63674 63524
rect 63714 63484 63756 63524
rect 63796 63484 63838 63524
rect 63878 63484 63920 63524
rect 63592 63475 63960 63484
rect 78712 63524 79080 63533
rect 78752 63484 78794 63524
rect 78834 63484 78876 63524
rect 78916 63484 78958 63524
rect 78998 63484 79040 63524
rect 78712 63475 79080 63484
rect 93832 63524 94200 63533
rect 93872 63484 93914 63524
rect 93954 63484 93996 63524
rect 94036 63484 94078 63524
rect 94118 63484 94160 63524
rect 93832 63475 94200 63484
rect 4352 62768 4720 62777
rect 4392 62728 4434 62768
rect 4474 62728 4516 62768
rect 4556 62728 4598 62768
rect 4638 62728 4680 62768
rect 4352 62719 4720 62728
rect 19472 62768 19840 62777
rect 19512 62728 19554 62768
rect 19594 62728 19636 62768
rect 19676 62728 19718 62768
rect 19758 62728 19800 62768
rect 19472 62719 19840 62728
rect 34592 62768 34960 62777
rect 34632 62728 34674 62768
rect 34714 62728 34756 62768
rect 34796 62728 34838 62768
rect 34878 62728 34920 62768
rect 34592 62719 34960 62728
rect 49712 62768 50080 62777
rect 49752 62728 49794 62768
rect 49834 62728 49876 62768
rect 49916 62728 49958 62768
rect 49998 62728 50040 62768
rect 49712 62719 50080 62728
rect 64832 62768 65200 62777
rect 64872 62728 64914 62768
rect 64954 62728 64996 62768
rect 65036 62728 65078 62768
rect 65118 62728 65160 62768
rect 64832 62719 65200 62728
rect 79952 62768 80320 62777
rect 79992 62728 80034 62768
rect 80074 62728 80116 62768
rect 80156 62728 80198 62768
rect 80238 62728 80280 62768
rect 79952 62719 80320 62728
rect 95072 62768 95440 62777
rect 95112 62728 95154 62768
rect 95194 62728 95236 62768
rect 95276 62728 95318 62768
rect 95358 62728 95400 62768
rect 95072 62719 95440 62728
rect 3112 62012 3480 62021
rect 3152 61972 3194 62012
rect 3234 61972 3276 62012
rect 3316 61972 3358 62012
rect 3398 61972 3440 62012
rect 3112 61963 3480 61972
rect 18232 62012 18600 62021
rect 18272 61972 18314 62012
rect 18354 61972 18396 62012
rect 18436 61972 18478 62012
rect 18518 61972 18560 62012
rect 18232 61963 18600 61972
rect 33352 62012 33720 62021
rect 33392 61972 33434 62012
rect 33474 61972 33516 62012
rect 33556 61972 33598 62012
rect 33638 61972 33680 62012
rect 33352 61963 33720 61972
rect 48472 62012 48840 62021
rect 48512 61972 48554 62012
rect 48594 61972 48636 62012
rect 48676 61972 48718 62012
rect 48758 61972 48800 62012
rect 48472 61963 48840 61972
rect 63592 62012 63960 62021
rect 63632 61972 63674 62012
rect 63714 61972 63756 62012
rect 63796 61972 63838 62012
rect 63878 61972 63920 62012
rect 63592 61963 63960 61972
rect 78712 62012 79080 62021
rect 78752 61972 78794 62012
rect 78834 61972 78876 62012
rect 78916 61972 78958 62012
rect 78998 61972 79040 62012
rect 78712 61963 79080 61972
rect 93832 62012 94200 62021
rect 93872 61972 93914 62012
rect 93954 61972 93996 62012
rect 94036 61972 94078 62012
rect 94118 61972 94160 62012
rect 93832 61963 94200 61972
rect 4352 61256 4720 61265
rect 4392 61216 4434 61256
rect 4474 61216 4516 61256
rect 4556 61216 4598 61256
rect 4638 61216 4680 61256
rect 4352 61207 4720 61216
rect 19472 61256 19840 61265
rect 19512 61216 19554 61256
rect 19594 61216 19636 61256
rect 19676 61216 19718 61256
rect 19758 61216 19800 61256
rect 19472 61207 19840 61216
rect 34592 61256 34960 61265
rect 34632 61216 34674 61256
rect 34714 61216 34756 61256
rect 34796 61216 34838 61256
rect 34878 61216 34920 61256
rect 34592 61207 34960 61216
rect 49712 61256 50080 61265
rect 49752 61216 49794 61256
rect 49834 61216 49876 61256
rect 49916 61216 49958 61256
rect 49998 61216 50040 61256
rect 49712 61207 50080 61216
rect 64832 61256 65200 61265
rect 64872 61216 64914 61256
rect 64954 61216 64996 61256
rect 65036 61216 65078 61256
rect 65118 61216 65160 61256
rect 64832 61207 65200 61216
rect 79952 61256 80320 61265
rect 79992 61216 80034 61256
rect 80074 61216 80116 61256
rect 80156 61216 80198 61256
rect 80238 61216 80280 61256
rect 79952 61207 80320 61216
rect 95072 61256 95440 61265
rect 95112 61216 95154 61256
rect 95194 61216 95236 61256
rect 95276 61216 95318 61256
rect 95358 61216 95400 61256
rect 95072 61207 95440 61216
rect 3112 60500 3480 60509
rect 3152 60460 3194 60500
rect 3234 60460 3276 60500
rect 3316 60460 3358 60500
rect 3398 60460 3440 60500
rect 3112 60451 3480 60460
rect 18232 60500 18600 60509
rect 18272 60460 18314 60500
rect 18354 60460 18396 60500
rect 18436 60460 18478 60500
rect 18518 60460 18560 60500
rect 18232 60451 18600 60460
rect 33352 60500 33720 60509
rect 33392 60460 33434 60500
rect 33474 60460 33516 60500
rect 33556 60460 33598 60500
rect 33638 60460 33680 60500
rect 33352 60451 33720 60460
rect 48472 60500 48840 60509
rect 48512 60460 48554 60500
rect 48594 60460 48636 60500
rect 48676 60460 48718 60500
rect 48758 60460 48800 60500
rect 48472 60451 48840 60460
rect 63592 60500 63960 60509
rect 63632 60460 63674 60500
rect 63714 60460 63756 60500
rect 63796 60460 63838 60500
rect 63878 60460 63920 60500
rect 63592 60451 63960 60460
rect 78712 60500 79080 60509
rect 78752 60460 78794 60500
rect 78834 60460 78876 60500
rect 78916 60460 78958 60500
rect 78998 60460 79040 60500
rect 78712 60451 79080 60460
rect 93832 60500 94200 60509
rect 93872 60460 93914 60500
rect 93954 60460 93996 60500
rect 94036 60460 94078 60500
rect 94118 60460 94160 60500
rect 93832 60451 94200 60460
rect 4352 59744 4720 59753
rect 4392 59704 4434 59744
rect 4474 59704 4516 59744
rect 4556 59704 4598 59744
rect 4638 59704 4680 59744
rect 4352 59695 4720 59704
rect 19472 59744 19840 59753
rect 19512 59704 19554 59744
rect 19594 59704 19636 59744
rect 19676 59704 19718 59744
rect 19758 59704 19800 59744
rect 19472 59695 19840 59704
rect 34592 59744 34960 59753
rect 34632 59704 34674 59744
rect 34714 59704 34756 59744
rect 34796 59704 34838 59744
rect 34878 59704 34920 59744
rect 34592 59695 34960 59704
rect 49712 59744 50080 59753
rect 49752 59704 49794 59744
rect 49834 59704 49876 59744
rect 49916 59704 49958 59744
rect 49998 59704 50040 59744
rect 49712 59695 50080 59704
rect 64832 59744 65200 59753
rect 64872 59704 64914 59744
rect 64954 59704 64996 59744
rect 65036 59704 65078 59744
rect 65118 59704 65160 59744
rect 64832 59695 65200 59704
rect 79952 59744 80320 59753
rect 79992 59704 80034 59744
rect 80074 59704 80116 59744
rect 80156 59704 80198 59744
rect 80238 59704 80280 59744
rect 79952 59695 80320 59704
rect 95072 59744 95440 59753
rect 95112 59704 95154 59744
rect 95194 59704 95236 59744
rect 95276 59704 95318 59744
rect 95358 59704 95400 59744
rect 95072 59695 95440 59704
rect 3112 58988 3480 58997
rect 3152 58948 3194 58988
rect 3234 58948 3276 58988
rect 3316 58948 3358 58988
rect 3398 58948 3440 58988
rect 3112 58939 3480 58948
rect 18232 58988 18600 58997
rect 18272 58948 18314 58988
rect 18354 58948 18396 58988
rect 18436 58948 18478 58988
rect 18518 58948 18560 58988
rect 18232 58939 18600 58948
rect 33352 58988 33720 58997
rect 33392 58948 33434 58988
rect 33474 58948 33516 58988
rect 33556 58948 33598 58988
rect 33638 58948 33680 58988
rect 33352 58939 33720 58948
rect 48472 58988 48840 58997
rect 48512 58948 48554 58988
rect 48594 58948 48636 58988
rect 48676 58948 48718 58988
rect 48758 58948 48800 58988
rect 48472 58939 48840 58948
rect 63592 58988 63960 58997
rect 63632 58948 63674 58988
rect 63714 58948 63756 58988
rect 63796 58948 63838 58988
rect 63878 58948 63920 58988
rect 63592 58939 63960 58948
rect 78712 58988 79080 58997
rect 78752 58948 78794 58988
rect 78834 58948 78876 58988
rect 78916 58948 78958 58988
rect 78998 58948 79040 58988
rect 78712 58939 79080 58948
rect 93832 58988 94200 58997
rect 93872 58948 93914 58988
rect 93954 58948 93996 58988
rect 94036 58948 94078 58988
rect 94118 58948 94160 58988
rect 93832 58939 94200 58948
rect 4352 58232 4720 58241
rect 4392 58192 4434 58232
rect 4474 58192 4516 58232
rect 4556 58192 4598 58232
rect 4638 58192 4680 58232
rect 4352 58183 4720 58192
rect 19472 58232 19840 58241
rect 19512 58192 19554 58232
rect 19594 58192 19636 58232
rect 19676 58192 19718 58232
rect 19758 58192 19800 58232
rect 19472 58183 19840 58192
rect 34592 58232 34960 58241
rect 34632 58192 34674 58232
rect 34714 58192 34756 58232
rect 34796 58192 34838 58232
rect 34878 58192 34920 58232
rect 34592 58183 34960 58192
rect 49712 58232 50080 58241
rect 49752 58192 49794 58232
rect 49834 58192 49876 58232
rect 49916 58192 49958 58232
rect 49998 58192 50040 58232
rect 49712 58183 50080 58192
rect 64832 58232 65200 58241
rect 64872 58192 64914 58232
rect 64954 58192 64996 58232
rect 65036 58192 65078 58232
rect 65118 58192 65160 58232
rect 64832 58183 65200 58192
rect 79952 58232 80320 58241
rect 79992 58192 80034 58232
rect 80074 58192 80116 58232
rect 80156 58192 80198 58232
rect 80238 58192 80280 58232
rect 79952 58183 80320 58192
rect 95072 58232 95440 58241
rect 95112 58192 95154 58232
rect 95194 58192 95236 58232
rect 95276 58192 95318 58232
rect 95358 58192 95400 58232
rect 95072 58183 95440 58192
rect 3112 57476 3480 57485
rect 3152 57436 3194 57476
rect 3234 57436 3276 57476
rect 3316 57436 3358 57476
rect 3398 57436 3440 57476
rect 3112 57427 3480 57436
rect 18232 57476 18600 57485
rect 18272 57436 18314 57476
rect 18354 57436 18396 57476
rect 18436 57436 18478 57476
rect 18518 57436 18560 57476
rect 18232 57427 18600 57436
rect 33352 57476 33720 57485
rect 33392 57436 33434 57476
rect 33474 57436 33516 57476
rect 33556 57436 33598 57476
rect 33638 57436 33680 57476
rect 33352 57427 33720 57436
rect 48472 57476 48840 57485
rect 48512 57436 48554 57476
rect 48594 57436 48636 57476
rect 48676 57436 48718 57476
rect 48758 57436 48800 57476
rect 48472 57427 48840 57436
rect 63592 57476 63960 57485
rect 63632 57436 63674 57476
rect 63714 57436 63756 57476
rect 63796 57436 63838 57476
rect 63878 57436 63920 57476
rect 63592 57427 63960 57436
rect 78712 57476 79080 57485
rect 78752 57436 78794 57476
rect 78834 57436 78876 57476
rect 78916 57436 78958 57476
rect 78998 57436 79040 57476
rect 78712 57427 79080 57436
rect 93832 57476 94200 57485
rect 93872 57436 93914 57476
rect 93954 57436 93996 57476
rect 94036 57436 94078 57476
rect 94118 57436 94160 57476
rect 93832 57427 94200 57436
rect 4352 56720 4720 56729
rect 4392 56680 4434 56720
rect 4474 56680 4516 56720
rect 4556 56680 4598 56720
rect 4638 56680 4680 56720
rect 4352 56671 4720 56680
rect 19472 56720 19840 56729
rect 19512 56680 19554 56720
rect 19594 56680 19636 56720
rect 19676 56680 19718 56720
rect 19758 56680 19800 56720
rect 19472 56671 19840 56680
rect 34592 56720 34960 56729
rect 34632 56680 34674 56720
rect 34714 56680 34756 56720
rect 34796 56680 34838 56720
rect 34878 56680 34920 56720
rect 34592 56671 34960 56680
rect 49712 56720 50080 56729
rect 49752 56680 49794 56720
rect 49834 56680 49876 56720
rect 49916 56680 49958 56720
rect 49998 56680 50040 56720
rect 49712 56671 50080 56680
rect 64832 56720 65200 56729
rect 64872 56680 64914 56720
rect 64954 56680 64996 56720
rect 65036 56680 65078 56720
rect 65118 56680 65160 56720
rect 64832 56671 65200 56680
rect 79952 56720 80320 56729
rect 79992 56680 80034 56720
rect 80074 56680 80116 56720
rect 80156 56680 80198 56720
rect 80238 56680 80280 56720
rect 79952 56671 80320 56680
rect 95072 56720 95440 56729
rect 95112 56680 95154 56720
rect 95194 56680 95236 56720
rect 95276 56680 95318 56720
rect 95358 56680 95400 56720
rect 95072 56671 95440 56680
rect 3112 55964 3480 55973
rect 3152 55924 3194 55964
rect 3234 55924 3276 55964
rect 3316 55924 3358 55964
rect 3398 55924 3440 55964
rect 3112 55915 3480 55924
rect 18232 55964 18600 55973
rect 18272 55924 18314 55964
rect 18354 55924 18396 55964
rect 18436 55924 18478 55964
rect 18518 55924 18560 55964
rect 18232 55915 18600 55924
rect 33352 55964 33720 55973
rect 33392 55924 33434 55964
rect 33474 55924 33516 55964
rect 33556 55924 33598 55964
rect 33638 55924 33680 55964
rect 33352 55915 33720 55924
rect 48472 55964 48840 55973
rect 48512 55924 48554 55964
rect 48594 55924 48636 55964
rect 48676 55924 48718 55964
rect 48758 55924 48800 55964
rect 48472 55915 48840 55924
rect 63592 55964 63960 55973
rect 63632 55924 63674 55964
rect 63714 55924 63756 55964
rect 63796 55924 63838 55964
rect 63878 55924 63920 55964
rect 63592 55915 63960 55924
rect 78712 55964 79080 55973
rect 78752 55924 78794 55964
rect 78834 55924 78876 55964
rect 78916 55924 78958 55964
rect 78998 55924 79040 55964
rect 78712 55915 79080 55924
rect 93832 55964 94200 55973
rect 93872 55924 93914 55964
rect 93954 55924 93996 55964
rect 94036 55924 94078 55964
rect 94118 55924 94160 55964
rect 93832 55915 94200 55924
rect 4352 55208 4720 55217
rect 4392 55168 4434 55208
rect 4474 55168 4516 55208
rect 4556 55168 4598 55208
rect 4638 55168 4680 55208
rect 4352 55159 4720 55168
rect 19472 55208 19840 55217
rect 19512 55168 19554 55208
rect 19594 55168 19636 55208
rect 19676 55168 19718 55208
rect 19758 55168 19800 55208
rect 19472 55159 19840 55168
rect 34592 55208 34960 55217
rect 34632 55168 34674 55208
rect 34714 55168 34756 55208
rect 34796 55168 34838 55208
rect 34878 55168 34920 55208
rect 34592 55159 34960 55168
rect 49712 55208 50080 55217
rect 49752 55168 49794 55208
rect 49834 55168 49876 55208
rect 49916 55168 49958 55208
rect 49998 55168 50040 55208
rect 49712 55159 50080 55168
rect 64832 55208 65200 55217
rect 64872 55168 64914 55208
rect 64954 55168 64996 55208
rect 65036 55168 65078 55208
rect 65118 55168 65160 55208
rect 64832 55159 65200 55168
rect 79952 55208 80320 55217
rect 79992 55168 80034 55208
rect 80074 55168 80116 55208
rect 80156 55168 80198 55208
rect 80238 55168 80280 55208
rect 79952 55159 80320 55168
rect 95072 55208 95440 55217
rect 95112 55168 95154 55208
rect 95194 55168 95236 55208
rect 95276 55168 95318 55208
rect 95358 55168 95400 55208
rect 95072 55159 95440 55168
rect 3112 54452 3480 54461
rect 3152 54412 3194 54452
rect 3234 54412 3276 54452
rect 3316 54412 3358 54452
rect 3398 54412 3440 54452
rect 3112 54403 3480 54412
rect 18232 54452 18600 54461
rect 18272 54412 18314 54452
rect 18354 54412 18396 54452
rect 18436 54412 18478 54452
rect 18518 54412 18560 54452
rect 18232 54403 18600 54412
rect 33352 54452 33720 54461
rect 33392 54412 33434 54452
rect 33474 54412 33516 54452
rect 33556 54412 33598 54452
rect 33638 54412 33680 54452
rect 33352 54403 33720 54412
rect 48472 54452 48840 54461
rect 48512 54412 48554 54452
rect 48594 54412 48636 54452
rect 48676 54412 48718 54452
rect 48758 54412 48800 54452
rect 48472 54403 48840 54412
rect 63592 54452 63960 54461
rect 63632 54412 63674 54452
rect 63714 54412 63756 54452
rect 63796 54412 63838 54452
rect 63878 54412 63920 54452
rect 63592 54403 63960 54412
rect 78712 54452 79080 54461
rect 78752 54412 78794 54452
rect 78834 54412 78876 54452
rect 78916 54412 78958 54452
rect 78998 54412 79040 54452
rect 78712 54403 79080 54412
rect 93832 54452 94200 54461
rect 93872 54412 93914 54452
rect 93954 54412 93996 54452
rect 94036 54412 94078 54452
rect 94118 54412 94160 54452
rect 93832 54403 94200 54412
rect 4352 53696 4720 53705
rect 4392 53656 4434 53696
rect 4474 53656 4516 53696
rect 4556 53656 4598 53696
rect 4638 53656 4680 53696
rect 4352 53647 4720 53656
rect 19472 53696 19840 53705
rect 19512 53656 19554 53696
rect 19594 53656 19636 53696
rect 19676 53656 19718 53696
rect 19758 53656 19800 53696
rect 19472 53647 19840 53656
rect 34592 53696 34960 53705
rect 34632 53656 34674 53696
rect 34714 53656 34756 53696
rect 34796 53656 34838 53696
rect 34878 53656 34920 53696
rect 34592 53647 34960 53656
rect 49712 53696 50080 53705
rect 49752 53656 49794 53696
rect 49834 53656 49876 53696
rect 49916 53656 49958 53696
rect 49998 53656 50040 53696
rect 49712 53647 50080 53656
rect 64832 53696 65200 53705
rect 64872 53656 64914 53696
rect 64954 53656 64996 53696
rect 65036 53656 65078 53696
rect 65118 53656 65160 53696
rect 64832 53647 65200 53656
rect 79952 53696 80320 53705
rect 79992 53656 80034 53696
rect 80074 53656 80116 53696
rect 80156 53656 80198 53696
rect 80238 53656 80280 53696
rect 79952 53647 80320 53656
rect 95072 53696 95440 53705
rect 95112 53656 95154 53696
rect 95194 53656 95236 53696
rect 95276 53656 95318 53696
rect 95358 53656 95400 53696
rect 95072 53647 95440 53656
rect 3112 52940 3480 52949
rect 3152 52900 3194 52940
rect 3234 52900 3276 52940
rect 3316 52900 3358 52940
rect 3398 52900 3440 52940
rect 3112 52891 3480 52900
rect 18232 52940 18600 52949
rect 18272 52900 18314 52940
rect 18354 52900 18396 52940
rect 18436 52900 18478 52940
rect 18518 52900 18560 52940
rect 18232 52891 18600 52900
rect 33352 52940 33720 52949
rect 33392 52900 33434 52940
rect 33474 52900 33516 52940
rect 33556 52900 33598 52940
rect 33638 52900 33680 52940
rect 33352 52891 33720 52900
rect 48472 52940 48840 52949
rect 48512 52900 48554 52940
rect 48594 52900 48636 52940
rect 48676 52900 48718 52940
rect 48758 52900 48800 52940
rect 48472 52891 48840 52900
rect 63592 52940 63960 52949
rect 63632 52900 63674 52940
rect 63714 52900 63756 52940
rect 63796 52900 63838 52940
rect 63878 52900 63920 52940
rect 63592 52891 63960 52900
rect 78712 52940 79080 52949
rect 78752 52900 78794 52940
rect 78834 52900 78876 52940
rect 78916 52900 78958 52940
rect 78998 52900 79040 52940
rect 78712 52891 79080 52900
rect 93832 52940 94200 52949
rect 93872 52900 93914 52940
rect 93954 52900 93996 52940
rect 94036 52900 94078 52940
rect 94118 52900 94160 52940
rect 93832 52891 94200 52900
rect 4352 52184 4720 52193
rect 4392 52144 4434 52184
rect 4474 52144 4516 52184
rect 4556 52144 4598 52184
rect 4638 52144 4680 52184
rect 4352 52135 4720 52144
rect 19472 52184 19840 52193
rect 19512 52144 19554 52184
rect 19594 52144 19636 52184
rect 19676 52144 19718 52184
rect 19758 52144 19800 52184
rect 19472 52135 19840 52144
rect 34592 52184 34960 52193
rect 34632 52144 34674 52184
rect 34714 52144 34756 52184
rect 34796 52144 34838 52184
rect 34878 52144 34920 52184
rect 34592 52135 34960 52144
rect 49712 52184 50080 52193
rect 49752 52144 49794 52184
rect 49834 52144 49876 52184
rect 49916 52144 49958 52184
rect 49998 52144 50040 52184
rect 49712 52135 50080 52144
rect 64832 52184 65200 52193
rect 64872 52144 64914 52184
rect 64954 52144 64996 52184
rect 65036 52144 65078 52184
rect 65118 52144 65160 52184
rect 64832 52135 65200 52144
rect 79952 52184 80320 52193
rect 79992 52144 80034 52184
rect 80074 52144 80116 52184
rect 80156 52144 80198 52184
rect 80238 52144 80280 52184
rect 79952 52135 80320 52144
rect 95072 52184 95440 52193
rect 95112 52144 95154 52184
rect 95194 52144 95236 52184
rect 95276 52144 95318 52184
rect 95358 52144 95400 52184
rect 95072 52135 95440 52144
rect 3112 51428 3480 51437
rect 3152 51388 3194 51428
rect 3234 51388 3276 51428
rect 3316 51388 3358 51428
rect 3398 51388 3440 51428
rect 3112 51379 3480 51388
rect 18232 51428 18600 51437
rect 18272 51388 18314 51428
rect 18354 51388 18396 51428
rect 18436 51388 18478 51428
rect 18518 51388 18560 51428
rect 18232 51379 18600 51388
rect 33352 51428 33720 51437
rect 33392 51388 33434 51428
rect 33474 51388 33516 51428
rect 33556 51388 33598 51428
rect 33638 51388 33680 51428
rect 33352 51379 33720 51388
rect 48472 51428 48840 51437
rect 48512 51388 48554 51428
rect 48594 51388 48636 51428
rect 48676 51388 48718 51428
rect 48758 51388 48800 51428
rect 48472 51379 48840 51388
rect 63592 51428 63960 51437
rect 63632 51388 63674 51428
rect 63714 51388 63756 51428
rect 63796 51388 63838 51428
rect 63878 51388 63920 51428
rect 63592 51379 63960 51388
rect 78712 51428 79080 51437
rect 78752 51388 78794 51428
rect 78834 51388 78876 51428
rect 78916 51388 78958 51428
rect 78998 51388 79040 51428
rect 78712 51379 79080 51388
rect 93832 51428 94200 51437
rect 93872 51388 93914 51428
rect 93954 51388 93996 51428
rect 94036 51388 94078 51428
rect 94118 51388 94160 51428
rect 93832 51379 94200 51388
rect 4352 50672 4720 50681
rect 4392 50632 4434 50672
rect 4474 50632 4516 50672
rect 4556 50632 4598 50672
rect 4638 50632 4680 50672
rect 4352 50623 4720 50632
rect 19472 50672 19840 50681
rect 19512 50632 19554 50672
rect 19594 50632 19636 50672
rect 19676 50632 19718 50672
rect 19758 50632 19800 50672
rect 19472 50623 19840 50632
rect 34592 50672 34960 50681
rect 34632 50632 34674 50672
rect 34714 50632 34756 50672
rect 34796 50632 34838 50672
rect 34878 50632 34920 50672
rect 34592 50623 34960 50632
rect 49712 50672 50080 50681
rect 49752 50632 49794 50672
rect 49834 50632 49876 50672
rect 49916 50632 49958 50672
rect 49998 50632 50040 50672
rect 49712 50623 50080 50632
rect 64832 50672 65200 50681
rect 64872 50632 64914 50672
rect 64954 50632 64996 50672
rect 65036 50632 65078 50672
rect 65118 50632 65160 50672
rect 64832 50623 65200 50632
rect 79952 50672 80320 50681
rect 79992 50632 80034 50672
rect 80074 50632 80116 50672
rect 80156 50632 80198 50672
rect 80238 50632 80280 50672
rect 79952 50623 80320 50632
rect 95072 50672 95440 50681
rect 95112 50632 95154 50672
rect 95194 50632 95236 50672
rect 95276 50632 95318 50672
rect 95358 50632 95400 50672
rect 95072 50623 95440 50632
rect 3112 49916 3480 49925
rect 3152 49876 3194 49916
rect 3234 49876 3276 49916
rect 3316 49876 3358 49916
rect 3398 49876 3440 49916
rect 3112 49867 3480 49876
rect 18232 49916 18600 49925
rect 18272 49876 18314 49916
rect 18354 49876 18396 49916
rect 18436 49876 18478 49916
rect 18518 49876 18560 49916
rect 18232 49867 18600 49876
rect 33352 49916 33720 49925
rect 33392 49876 33434 49916
rect 33474 49876 33516 49916
rect 33556 49876 33598 49916
rect 33638 49876 33680 49916
rect 33352 49867 33720 49876
rect 48472 49916 48840 49925
rect 48512 49876 48554 49916
rect 48594 49876 48636 49916
rect 48676 49876 48718 49916
rect 48758 49876 48800 49916
rect 48472 49867 48840 49876
rect 63592 49916 63960 49925
rect 63632 49876 63674 49916
rect 63714 49876 63756 49916
rect 63796 49876 63838 49916
rect 63878 49876 63920 49916
rect 63592 49867 63960 49876
rect 78712 49916 79080 49925
rect 78752 49876 78794 49916
rect 78834 49876 78876 49916
rect 78916 49876 78958 49916
rect 78998 49876 79040 49916
rect 78712 49867 79080 49876
rect 93832 49916 94200 49925
rect 93872 49876 93914 49916
rect 93954 49876 93996 49916
rect 94036 49876 94078 49916
rect 94118 49876 94160 49916
rect 93832 49867 94200 49876
rect 4352 49160 4720 49169
rect 4392 49120 4434 49160
rect 4474 49120 4516 49160
rect 4556 49120 4598 49160
rect 4638 49120 4680 49160
rect 4352 49111 4720 49120
rect 19472 49160 19840 49169
rect 19512 49120 19554 49160
rect 19594 49120 19636 49160
rect 19676 49120 19718 49160
rect 19758 49120 19800 49160
rect 19472 49111 19840 49120
rect 34592 49160 34960 49169
rect 34632 49120 34674 49160
rect 34714 49120 34756 49160
rect 34796 49120 34838 49160
rect 34878 49120 34920 49160
rect 34592 49111 34960 49120
rect 49712 49160 50080 49169
rect 49752 49120 49794 49160
rect 49834 49120 49876 49160
rect 49916 49120 49958 49160
rect 49998 49120 50040 49160
rect 49712 49111 50080 49120
rect 64832 49160 65200 49169
rect 64872 49120 64914 49160
rect 64954 49120 64996 49160
rect 65036 49120 65078 49160
rect 65118 49120 65160 49160
rect 64832 49111 65200 49120
rect 79952 49160 80320 49169
rect 79992 49120 80034 49160
rect 80074 49120 80116 49160
rect 80156 49120 80198 49160
rect 80238 49120 80280 49160
rect 79952 49111 80320 49120
rect 95072 49160 95440 49169
rect 95112 49120 95154 49160
rect 95194 49120 95236 49160
rect 95276 49120 95318 49160
rect 95358 49120 95400 49160
rect 95072 49111 95440 49120
rect 3112 48404 3480 48413
rect 3152 48364 3194 48404
rect 3234 48364 3276 48404
rect 3316 48364 3358 48404
rect 3398 48364 3440 48404
rect 3112 48355 3480 48364
rect 18232 48404 18600 48413
rect 18272 48364 18314 48404
rect 18354 48364 18396 48404
rect 18436 48364 18478 48404
rect 18518 48364 18560 48404
rect 18232 48355 18600 48364
rect 33352 48404 33720 48413
rect 33392 48364 33434 48404
rect 33474 48364 33516 48404
rect 33556 48364 33598 48404
rect 33638 48364 33680 48404
rect 33352 48355 33720 48364
rect 48472 48404 48840 48413
rect 48512 48364 48554 48404
rect 48594 48364 48636 48404
rect 48676 48364 48718 48404
rect 48758 48364 48800 48404
rect 48472 48355 48840 48364
rect 63592 48404 63960 48413
rect 63632 48364 63674 48404
rect 63714 48364 63756 48404
rect 63796 48364 63838 48404
rect 63878 48364 63920 48404
rect 63592 48355 63960 48364
rect 78712 48404 79080 48413
rect 78752 48364 78794 48404
rect 78834 48364 78876 48404
rect 78916 48364 78958 48404
rect 78998 48364 79040 48404
rect 78712 48355 79080 48364
rect 93832 48404 94200 48413
rect 93872 48364 93914 48404
rect 93954 48364 93996 48404
rect 94036 48364 94078 48404
rect 94118 48364 94160 48404
rect 93832 48355 94200 48364
rect 4352 47648 4720 47657
rect 4392 47608 4434 47648
rect 4474 47608 4516 47648
rect 4556 47608 4598 47648
rect 4638 47608 4680 47648
rect 4352 47599 4720 47608
rect 19472 47648 19840 47657
rect 19512 47608 19554 47648
rect 19594 47608 19636 47648
rect 19676 47608 19718 47648
rect 19758 47608 19800 47648
rect 19472 47599 19840 47608
rect 34592 47648 34960 47657
rect 34632 47608 34674 47648
rect 34714 47608 34756 47648
rect 34796 47608 34838 47648
rect 34878 47608 34920 47648
rect 34592 47599 34960 47608
rect 49712 47648 50080 47657
rect 49752 47608 49794 47648
rect 49834 47608 49876 47648
rect 49916 47608 49958 47648
rect 49998 47608 50040 47648
rect 49712 47599 50080 47608
rect 64832 47648 65200 47657
rect 64872 47608 64914 47648
rect 64954 47608 64996 47648
rect 65036 47608 65078 47648
rect 65118 47608 65160 47648
rect 64832 47599 65200 47608
rect 79952 47648 80320 47657
rect 79992 47608 80034 47648
rect 80074 47608 80116 47648
rect 80156 47608 80198 47648
rect 80238 47608 80280 47648
rect 79952 47599 80320 47608
rect 95072 47648 95440 47657
rect 95112 47608 95154 47648
rect 95194 47608 95236 47648
rect 95276 47608 95318 47648
rect 95358 47608 95400 47648
rect 95072 47599 95440 47608
rect 3112 46892 3480 46901
rect 3152 46852 3194 46892
rect 3234 46852 3276 46892
rect 3316 46852 3358 46892
rect 3398 46852 3440 46892
rect 3112 46843 3480 46852
rect 18232 46892 18600 46901
rect 18272 46852 18314 46892
rect 18354 46852 18396 46892
rect 18436 46852 18478 46892
rect 18518 46852 18560 46892
rect 18232 46843 18600 46852
rect 33352 46892 33720 46901
rect 33392 46852 33434 46892
rect 33474 46852 33516 46892
rect 33556 46852 33598 46892
rect 33638 46852 33680 46892
rect 33352 46843 33720 46852
rect 48472 46892 48840 46901
rect 48512 46852 48554 46892
rect 48594 46852 48636 46892
rect 48676 46852 48718 46892
rect 48758 46852 48800 46892
rect 48472 46843 48840 46852
rect 63592 46892 63960 46901
rect 63632 46852 63674 46892
rect 63714 46852 63756 46892
rect 63796 46852 63838 46892
rect 63878 46852 63920 46892
rect 63592 46843 63960 46852
rect 78712 46892 79080 46901
rect 78752 46852 78794 46892
rect 78834 46852 78876 46892
rect 78916 46852 78958 46892
rect 78998 46852 79040 46892
rect 78712 46843 79080 46852
rect 93832 46892 94200 46901
rect 93872 46852 93914 46892
rect 93954 46852 93996 46892
rect 94036 46852 94078 46892
rect 94118 46852 94160 46892
rect 93832 46843 94200 46852
rect 4352 46136 4720 46145
rect 4392 46096 4434 46136
rect 4474 46096 4516 46136
rect 4556 46096 4598 46136
rect 4638 46096 4680 46136
rect 4352 46087 4720 46096
rect 19472 46136 19840 46145
rect 19512 46096 19554 46136
rect 19594 46096 19636 46136
rect 19676 46096 19718 46136
rect 19758 46096 19800 46136
rect 19472 46087 19840 46096
rect 34592 46136 34960 46145
rect 34632 46096 34674 46136
rect 34714 46096 34756 46136
rect 34796 46096 34838 46136
rect 34878 46096 34920 46136
rect 34592 46087 34960 46096
rect 49712 46136 50080 46145
rect 49752 46096 49794 46136
rect 49834 46096 49876 46136
rect 49916 46096 49958 46136
rect 49998 46096 50040 46136
rect 49712 46087 50080 46096
rect 64832 46136 65200 46145
rect 64872 46096 64914 46136
rect 64954 46096 64996 46136
rect 65036 46096 65078 46136
rect 65118 46096 65160 46136
rect 64832 46087 65200 46096
rect 79952 46136 80320 46145
rect 79992 46096 80034 46136
rect 80074 46096 80116 46136
rect 80156 46096 80198 46136
rect 80238 46096 80280 46136
rect 79952 46087 80320 46096
rect 95072 46136 95440 46145
rect 95112 46096 95154 46136
rect 95194 46096 95236 46136
rect 95276 46096 95318 46136
rect 95358 46096 95400 46136
rect 95072 46087 95440 46096
rect 3112 45380 3480 45389
rect 3152 45340 3194 45380
rect 3234 45340 3276 45380
rect 3316 45340 3358 45380
rect 3398 45340 3440 45380
rect 3112 45331 3480 45340
rect 18232 45380 18600 45389
rect 18272 45340 18314 45380
rect 18354 45340 18396 45380
rect 18436 45340 18478 45380
rect 18518 45340 18560 45380
rect 18232 45331 18600 45340
rect 33352 45380 33720 45389
rect 33392 45340 33434 45380
rect 33474 45340 33516 45380
rect 33556 45340 33598 45380
rect 33638 45340 33680 45380
rect 33352 45331 33720 45340
rect 48472 45380 48840 45389
rect 48512 45340 48554 45380
rect 48594 45340 48636 45380
rect 48676 45340 48718 45380
rect 48758 45340 48800 45380
rect 48472 45331 48840 45340
rect 63592 45380 63960 45389
rect 63632 45340 63674 45380
rect 63714 45340 63756 45380
rect 63796 45340 63838 45380
rect 63878 45340 63920 45380
rect 63592 45331 63960 45340
rect 78712 45380 79080 45389
rect 78752 45340 78794 45380
rect 78834 45340 78876 45380
rect 78916 45340 78958 45380
rect 78998 45340 79040 45380
rect 78712 45331 79080 45340
rect 93832 45380 94200 45389
rect 93872 45340 93914 45380
rect 93954 45340 93996 45380
rect 94036 45340 94078 45380
rect 94118 45340 94160 45380
rect 93832 45331 94200 45340
rect 4352 44624 4720 44633
rect 4392 44584 4434 44624
rect 4474 44584 4516 44624
rect 4556 44584 4598 44624
rect 4638 44584 4680 44624
rect 4352 44575 4720 44584
rect 19472 44624 19840 44633
rect 19512 44584 19554 44624
rect 19594 44584 19636 44624
rect 19676 44584 19718 44624
rect 19758 44584 19800 44624
rect 19472 44575 19840 44584
rect 34592 44624 34960 44633
rect 34632 44584 34674 44624
rect 34714 44584 34756 44624
rect 34796 44584 34838 44624
rect 34878 44584 34920 44624
rect 34592 44575 34960 44584
rect 49712 44624 50080 44633
rect 49752 44584 49794 44624
rect 49834 44584 49876 44624
rect 49916 44584 49958 44624
rect 49998 44584 50040 44624
rect 49712 44575 50080 44584
rect 64832 44624 65200 44633
rect 64872 44584 64914 44624
rect 64954 44584 64996 44624
rect 65036 44584 65078 44624
rect 65118 44584 65160 44624
rect 64832 44575 65200 44584
rect 79952 44624 80320 44633
rect 79992 44584 80034 44624
rect 80074 44584 80116 44624
rect 80156 44584 80198 44624
rect 80238 44584 80280 44624
rect 79952 44575 80320 44584
rect 95072 44624 95440 44633
rect 95112 44584 95154 44624
rect 95194 44584 95236 44624
rect 95276 44584 95318 44624
rect 95358 44584 95400 44624
rect 95072 44575 95440 44584
rect 3112 43868 3480 43877
rect 3152 43828 3194 43868
rect 3234 43828 3276 43868
rect 3316 43828 3358 43868
rect 3398 43828 3440 43868
rect 3112 43819 3480 43828
rect 18232 43868 18600 43877
rect 18272 43828 18314 43868
rect 18354 43828 18396 43868
rect 18436 43828 18478 43868
rect 18518 43828 18560 43868
rect 18232 43819 18600 43828
rect 33352 43868 33720 43877
rect 33392 43828 33434 43868
rect 33474 43828 33516 43868
rect 33556 43828 33598 43868
rect 33638 43828 33680 43868
rect 33352 43819 33720 43828
rect 48472 43868 48840 43877
rect 48512 43828 48554 43868
rect 48594 43828 48636 43868
rect 48676 43828 48718 43868
rect 48758 43828 48800 43868
rect 48472 43819 48840 43828
rect 63592 43868 63960 43877
rect 63632 43828 63674 43868
rect 63714 43828 63756 43868
rect 63796 43828 63838 43868
rect 63878 43828 63920 43868
rect 63592 43819 63960 43828
rect 78712 43868 79080 43877
rect 78752 43828 78794 43868
rect 78834 43828 78876 43868
rect 78916 43828 78958 43868
rect 78998 43828 79040 43868
rect 78712 43819 79080 43828
rect 93832 43868 94200 43877
rect 93872 43828 93914 43868
rect 93954 43828 93996 43868
rect 94036 43828 94078 43868
rect 94118 43828 94160 43868
rect 93832 43819 94200 43828
rect 4352 43112 4720 43121
rect 4392 43072 4434 43112
rect 4474 43072 4516 43112
rect 4556 43072 4598 43112
rect 4638 43072 4680 43112
rect 4352 43063 4720 43072
rect 19472 43112 19840 43121
rect 19512 43072 19554 43112
rect 19594 43072 19636 43112
rect 19676 43072 19718 43112
rect 19758 43072 19800 43112
rect 19472 43063 19840 43072
rect 34592 43112 34960 43121
rect 34632 43072 34674 43112
rect 34714 43072 34756 43112
rect 34796 43072 34838 43112
rect 34878 43072 34920 43112
rect 34592 43063 34960 43072
rect 49712 43112 50080 43121
rect 49752 43072 49794 43112
rect 49834 43072 49876 43112
rect 49916 43072 49958 43112
rect 49998 43072 50040 43112
rect 49712 43063 50080 43072
rect 64832 43112 65200 43121
rect 64872 43072 64914 43112
rect 64954 43072 64996 43112
rect 65036 43072 65078 43112
rect 65118 43072 65160 43112
rect 64832 43063 65200 43072
rect 79952 43112 80320 43121
rect 79992 43072 80034 43112
rect 80074 43072 80116 43112
rect 80156 43072 80198 43112
rect 80238 43072 80280 43112
rect 79952 43063 80320 43072
rect 95072 43112 95440 43121
rect 95112 43072 95154 43112
rect 95194 43072 95236 43112
rect 95276 43072 95318 43112
rect 95358 43072 95400 43112
rect 95072 43063 95440 43072
rect 3112 42356 3480 42365
rect 3152 42316 3194 42356
rect 3234 42316 3276 42356
rect 3316 42316 3358 42356
rect 3398 42316 3440 42356
rect 3112 42307 3480 42316
rect 18232 42356 18600 42365
rect 18272 42316 18314 42356
rect 18354 42316 18396 42356
rect 18436 42316 18478 42356
rect 18518 42316 18560 42356
rect 18232 42307 18600 42316
rect 33352 42356 33720 42365
rect 33392 42316 33434 42356
rect 33474 42316 33516 42356
rect 33556 42316 33598 42356
rect 33638 42316 33680 42356
rect 33352 42307 33720 42316
rect 48472 42356 48840 42365
rect 48512 42316 48554 42356
rect 48594 42316 48636 42356
rect 48676 42316 48718 42356
rect 48758 42316 48800 42356
rect 48472 42307 48840 42316
rect 63592 42356 63960 42365
rect 63632 42316 63674 42356
rect 63714 42316 63756 42356
rect 63796 42316 63838 42356
rect 63878 42316 63920 42356
rect 63592 42307 63960 42316
rect 78712 42356 79080 42365
rect 78752 42316 78794 42356
rect 78834 42316 78876 42356
rect 78916 42316 78958 42356
rect 78998 42316 79040 42356
rect 78712 42307 79080 42316
rect 93832 42356 94200 42365
rect 93872 42316 93914 42356
rect 93954 42316 93996 42356
rect 94036 42316 94078 42356
rect 94118 42316 94160 42356
rect 93832 42307 94200 42316
rect 4352 41600 4720 41609
rect 4392 41560 4434 41600
rect 4474 41560 4516 41600
rect 4556 41560 4598 41600
rect 4638 41560 4680 41600
rect 4352 41551 4720 41560
rect 19472 41600 19840 41609
rect 19512 41560 19554 41600
rect 19594 41560 19636 41600
rect 19676 41560 19718 41600
rect 19758 41560 19800 41600
rect 19472 41551 19840 41560
rect 34592 41600 34960 41609
rect 34632 41560 34674 41600
rect 34714 41560 34756 41600
rect 34796 41560 34838 41600
rect 34878 41560 34920 41600
rect 34592 41551 34960 41560
rect 49712 41600 50080 41609
rect 49752 41560 49794 41600
rect 49834 41560 49876 41600
rect 49916 41560 49958 41600
rect 49998 41560 50040 41600
rect 49712 41551 50080 41560
rect 64832 41600 65200 41609
rect 64872 41560 64914 41600
rect 64954 41560 64996 41600
rect 65036 41560 65078 41600
rect 65118 41560 65160 41600
rect 64832 41551 65200 41560
rect 79952 41600 80320 41609
rect 79992 41560 80034 41600
rect 80074 41560 80116 41600
rect 80156 41560 80198 41600
rect 80238 41560 80280 41600
rect 79952 41551 80320 41560
rect 95072 41600 95440 41609
rect 95112 41560 95154 41600
rect 95194 41560 95236 41600
rect 95276 41560 95318 41600
rect 95358 41560 95400 41600
rect 95072 41551 95440 41560
rect 3112 40844 3480 40853
rect 3152 40804 3194 40844
rect 3234 40804 3276 40844
rect 3316 40804 3358 40844
rect 3398 40804 3440 40844
rect 3112 40795 3480 40804
rect 18232 40844 18600 40853
rect 18272 40804 18314 40844
rect 18354 40804 18396 40844
rect 18436 40804 18478 40844
rect 18518 40804 18560 40844
rect 18232 40795 18600 40804
rect 33352 40844 33720 40853
rect 33392 40804 33434 40844
rect 33474 40804 33516 40844
rect 33556 40804 33598 40844
rect 33638 40804 33680 40844
rect 33352 40795 33720 40804
rect 48472 40844 48840 40853
rect 48512 40804 48554 40844
rect 48594 40804 48636 40844
rect 48676 40804 48718 40844
rect 48758 40804 48800 40844
rect 48472 40795 48840 40804
rect 63592 40844 63960 40853
rect 63632 40804 63674 40844
rect 63714 40804 63756 40844
rect 63796 40804 63838 40844
rect 63878 40804 63920 40844
rect 63592 40795 63960 40804
rect 78712 40844 79080 40853
rect 78752 40804 78794 40844
rect 78834 40804 78876 40844
rect 78916 40804 78958 40844
rect 78998 40804 79040 40844
rect 78712 40795 79080 40804
rect 93832 40844 94200 40853
rect 93872 40804 93914 40844
rect 93954 40804 93996 40844
rect 94036 40804 94078 40844
rect 94118 40804 94160 40844
rect 93832 40795 94200 40804
rect 4352 40088 4720 40097
rect 4392 40048 4434 40088
rect 4474 40048 4516 40088
rect 4556 40048 4598 40088
rect 4638 40048 4680 40088
rect 4352 40039 4720 40048
rect 19472 40088 19840 40097
rect 19512 40048 19554 40088
rect 19594 40048 19636 40088
rect 19676 40048 19718 40088
rect 19758 40048 19800 40088
rect 19472 40039 19840 40048
rect 34592 40088 34960 40097
rect 34632 40048 34674 40088
rect 34714 40048 34756 40088
rect 34796 40048 34838 40088
rect 34878 40048 34920 40088
rect 34592 40039 34960 40048
rect 49712 40088 50080 40097
rect 49752 40048 49794 40088
rect 49834 40048 49876 40088
rect 49916 40048 49958 40088
rect 49998 40048 50040 40088
rect 49712 40039 50080 40048
rect 64832 40088 65200 40097
rect 64872 40048 64914 40088
rect 64954 40048 64996 40088
rect 65036 40048 65078 40088
rect 65118 40048 65160 40088
rect 64832 40039 65200 40048
rect 79952 40088 80320 40097
rect 79992 40048 80034 40088
rect 80074 40048 80116 40088
rect 80156 40048 80198 40088
rect 80238 40048 80280 40088
rect 79952 40039 80320 40048
rect 95072 40088 95440 40097
rect 95112 40048 95154 40088
rect 95194 40048 95236 40088
rect 95276 40048 95318 40088
rect 95358 40048 95400 40088
rect 95072 40039 95440 40048
rect 3112 39332 3480 39341
rect 3152 39292 3194 39332
rect 3234 39292 3276 39332
rect 3316 39292 3358 39332
rect 3398 39292 3440 39332
rect 3112 39283 3480 39292
rect 18232 39332 18600 39341
rect 18272 39292 18314 39332
rect 18354 39292 18396 39332
rect 18436 39292 18478 39332
rect 18518 39292 18560 39332
rect 18232 39283 18600 39292
rect 33352 39332 33720 39341
rect 33392 39292 33434 39332
rect 33474 39292 33516 39332
rect 33556 39292 33598 39332
rect 33638 39292 33680 39332
rect 33352 39283 33720 39292
rect 48472 39332 48840 39341
rect 48512 39292 48554 39332
rect 48594 39292 48636 39332
rect 48676 39292 48718 39332
rect 48758 39292 48800 39332
rect 48472 39283 48840 39292
rect 63592 39332 63960 39341
rect 63632 39292 63674 39332
rect 63714 39292 63756 39332
rect 63796 39292 63838 39332
rect 63878 39292 63920 39332
rect 63592 39283 63960 39292
rect 78712 39332 79080 39341
rect 78752 39292 78794 39332
rect 78834 39292 78876 39332
rect 78916 39292 78958 39332
rect 78998 39292 79040 39332
rect 78712 39283 79080 39292
rect 93832 39332 94200 39341
rect 93872 39292 93914 39332
rect 93954 39292 93996 39332
rect 94036 39292 94078 39332
rect 94118 39292 94160 39332
rect 93832 39283 94200 39292
rect 4352 38576 4720 38585
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4352 38527 4720 38536
rect 19472 38576 19840 38585
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19472 38527 19840 38536
rect 34592 38576 34960 38585
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34592 38527 34960 38536
rect 49712 38576 50080 38585
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 49712 38527 50080 38536
rect 64832 38576 65200 38585
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 64832 38527 65200 38536
rect 79952 38576 80320 38585
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 79952 38527 80320 38536
rect 95072 38576 95440 38585
rect 95112 38536 95154 38576
rect 95194 38536 95236 38576
rect 95276 38536 95318 38576
rect 95358 38536 95400 38576
rect 95072 38527 95440 38536
rect 3112 37820 3480 37829
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3112 37771 3480 37780
rect 18232 37820 18600 37829
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18232 37771 18600 37780
rect 33352 37820 33720 37829
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33352 37771 33720 37780
rect 48472 37820 48840 37829
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48472 37771 48840 37780
rect 63592 37820 63960 37829
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63592 37771 63960 37780
rect 78712 37820 79080 37829
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 78712 37771 79080 37780
rect 93832 37820 94200 37829
rect 93872 37780 93914 37820
rect 93954 37780 93996 37820
rect 94036 37780 94078 37820
rect 94118 37780 94160 37820
rect 93832 37771 94200 37780
rect 4352 37064 4720 37073
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4352 37015 4720 37024
rect 19472 37064 19840 37073
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19472 37015 19840 37024
rect 34592 37064 34960 37073
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34592 37015 34960 37024
rect 49712 37064 50080 37073
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 49712 37015 50080 37024
rect 64832 37064 65200 37073
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 64832 37015 65200 37024
rect 79952 37064 80320 37073
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 79952 37015 80320 37024
rect 95072 37064 95440 37073
rect 95112 37024 95154 37064
rect 95194 37024 95236 37064
rect 95276 37024 95318 37064
rect 95358 37024 95400 37064
rect 95072 37015 95440 37024
rect 3112 36308 3480 36317
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3112 36259 3480 36268
rect 18232 36308 18600 36317
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18232 36259 18600 36268
rect 33352 36308 33720 36317
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33352 36259 33720 36268
rect 48472 36308 48840 36317
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48472 36259 48840 36268
rect 63592 36308 63960 36317
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63592 36259 63960 36268
rect 78712 36308 79080 36317
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 78712 36259 79080 36268
rect 93832 36308 94200 36317
rect 93872 36268 93914 36308
rect 93954 36268 93996 36308
rect 94036 36268 94078 36308
rect 94118 36268 94160 36308
rect 93832 36259 94200 36268
rect 4352 35552 4720 35561
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4352 35503 4720 35512
rect 19472 35552 19840 35561
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19472 35503 19840 35512
rect 34592 35552 34960 35561
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34592 35503 34960 35512
rect 49712 35552 50080 35561
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 49712 35503 50080 35512
rect 64832 35552 65200 35561
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 64832 35503 65200 35512
rect 79952 35552 80320 35561
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 79952 35503 80320 35512
rect 95072 35552 95440 35561
rect 95112 35512 95154 35552
rect 95194 35512 95236 35552
rect 95276 35512 95318 35552
rect 95358 35512 95400 35552
rect 95072 35503 95440 35512
rect 3112 34796 3480 34805
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3112 34747 3480 34756
rect 18232 34796 18600 34805
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18232 34747 18600 34756
rect 33352 34796 33720 34805
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33352 34747 33720 34756
rect 48472 34796 48840 34805
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48472 34747 48840 34756
rect 63592 34796 63960 34805
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63592 34747 63960 34756
rect 78712 34796 79080 34805
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 78712 34747 79080 34756
rect 93832 34796 94200 34805
rect 93872 34756 93914 34796
rect 93954 34756 93996 34796
rect 94036 34756 94078 34796
rect 94118 34756 94160 34796
rect 93832 34747 94200 34756
rect 4352 34040 4720 34049
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4352 33991 4720 34000
rect 19472 34040 19840 34049
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19472 33991 19840 34000
rect 34592 34040 34960 34049
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34592 33991 34960 34000
rect 49712 34040 50080 34049
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 49712 33991 50080 34000
rect 64832 34040 65200 34049
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 64832 33991 65200 34000
rect 79952 34040 80320 34049
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 79952 33991 80320 34000
rect 95072 34040 95440 34049
rect 95112 34000 95154 34040
rect 95194 34000 95236 34040
rect 95276 34000 95318 34040
rect 95358 34000 95400 34040
rect 95072 33991 95440 34000
rect 3112 33284 3480 33293
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3112 33235 3480 33244
rect 18232 33284 18600 33293
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18232 33235 18600 33244
rect 33352 33284 33720 33293
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33352 33235 33720 33244
rect 48472 33284 48840 33293
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48472 33235 48840 33244
rect 63592 33284 63960 33293
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63592 33235 63960 33244
rect 78712 33284 79080 33293
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 78712 33235 79080 33244
rect 93832 33284 94200 33293
rect 93872 33244 93914 33284
rect 93954 33244 93996 33284
rect 94036 33244 94078 33284
rect 94118 33244 94160 33284
rect 93832 33235 94200 33244
rect 4352 32528 4720 32537
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4352 32479 4720 32488
rect 19472 32528 19840 32537
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19472 32479 19840 32488
rect 34592 32528 34960 32537
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34592 32479 34960 32488
rect 49712 32528 50080 32537
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 49712 32479 50080 32488
rect 64832 32528 65200 32537
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 64832 32479 65200 32488
rect 79952 32528 80320 32537
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 79952 32479 80320 32488
rect 95072 32528 95440 32537
rect 95112 32488 95154 32528
rect 95194 32488 95236 32528
rect 95276 32488 95318 32528
rect 95358 32488 95400 32528
rect 95072 32479 95440 32488
rect 3112 31772 3480 31781
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3112 31723 3480 31732
rect 18232 31772 18600 31781
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18232 31723 18600 31732
rect 33352 31772 33720 31781
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33352 31723 33720 31732
rect 48472 31772 48840 31781
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48472 31723 48840 31732
rect 63592 31772 63960 31781
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63592 31723 63960 31732
rect 78712 31772 79080 31781
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 78712 31723 79080 31732
rect 93832 31772 94200 31781
rect 93872 31732 93914 31772
rect 93954 31732 93996 31772
rect 94036 31732 94078 31772
rect 94118 31732 94160 31772
rect 93832 31723 94200 31732
rect 4352 31016 4720 31025
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4352 30967 4720 30976
rect 19472 31016 19840 31025
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19472 30967 19840 30976
rect 34592 31016 34960 31025
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34592 30967 34960 30976
rect 49712 31016 50080 31025
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 49712 30967 50080 30976
rect 64832 31016 65200 31025
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 64832 30967 65200 30976
rect 79952 31016 80320 31025
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 79952 30967 80320 30976
rect 95072 31016 95440 31025
rect 95112 30976 95154 31016
rect 95194 30976 95236 31016
rect 95276 30976 95318 31016
rect 95358 30976 95400 31016
rect 95072 30967 95440 30976
rect 3112 30260 3480 30269
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3112 30211 3480 30220
rect 18232 30260 18600 30269
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18232 30211 18600 30220
rect 33352 30260 33720 30269
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33352 30211 33720 30220
rect 48472 30260 48840 30269
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48472 30211 48840 30220
rect 63592 30260 63960 30269
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63592 30211 63960 30220
rect 78712 30260 79080 30269
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 78712 30211 79080 30220
rect 93832 30260 94200 30269
rect 93872 30220 93914 30260
rect 93954 30220 93996 30260
rect 94036 30220 94078 30260
rect 94118 30220 94160 30260
rect 93832 30211 94200 30220
rect 4352 29504 4720 29513
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4352 29455 4720 29464
rect 19472 29504 19840 29513
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19472 29455 19840 29464
rect 34592 29504 34960 29513
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34592 29455 34960 29464
rect 49712 29504 50080 29513
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 49712 29455 50080 29464
rect 64832 29504 65200 29513
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 64832 29455 65200 29464
rect 79952 29504 80320 29513
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 79952 29455 80320 29464
rect 95072 29504 95440 29513
rect 95112 29464 95154 29504
rect 95194 29464 95236 29504
rect 95276 29464 95318 29504
rect 95358 29464 95400 29504
rect 95072 29455 95440 29464
rect 3112 28748 3480 28757
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3112 28699 3480 28708
rect 18232 28748 18600 28757
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18232 28699 18600 28708
rect 33352 28748 33720 28757
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33352 28699 33720 28708
rect 48472 28748 48840 28757
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48472 28699 48840 28708
rect 63592 28748 63960 28757
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63592 28699 63960 28708
rect 78712 28748 79080 28757
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 78712 28699 79080 28708
rect 93832 28748 94200 28757
rect 93872 28708 93914 28748
rect 93954 28708 93996 28748
rect 94036 28708 94078 28748
rect 94118 28708 94160 28748
rect 93832 28699 94200 28708
rect 4352 27992 4720 28001
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4352 27943 4720 27952
rect 19472 27992 19840 28001
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19472 27943 19840 27952
rect 34592 27992 34960 28001
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34592 27943 34960 27952
rect 49712 27992 50080 28001
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 49712 27943 50080 27952
rect 64832 27992 65200 28001
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 64832 27943 65200 27952
rect 79952 27992 80320 28001
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 79952 27943 80320 27952
rect 95072 27992 95440 28001
rect 95112 27952 95154 27992
rect 95194 27952 95236 27992
rect 95276 27952 95318 27992
rect 95358 27952 95400 27992
rect 95072 27943 95440 27952
rect 3112 27236 3480 27245
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3112 27187 3480 27196
rect 18232 27236 18600 27245
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18232 27187 18600 27196
rect 33352 27236 33720 27245
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33352 27187 33720 27196
rect 48472 27236 48840 27245
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48472 27187 48840 27196
rect 63592 27236 63960 27245
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63592 27187 63960 27196
rect 78712 27236 79080 27245
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 78712 27187 79080 27196
rect 93832 27236 94200 27245
rect 93872 27196 93914 27236
rect 93954 27196 93996 27236
rect 94036 27196 94078 27236
rect 94118 27196 94160 27236
rect 93832 27187 94200 27196
rect 4352 26480 4720 26489
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4352 26431 4720 26440
rect 19472 26480 19840 26489
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19472 26431 19840 26440
rect 34592 26480 34960 26489
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34592 26431 34960 26440
rect 49712 26480 50080 26489
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 49712 26431 50080 26440
rect 64832 26480 65200 26489
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 64832 26431 65200 26440
rect 79952 26480 80320 26489
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 79952 26431 80320 26440
rect 95072 26480 95440 26489
rect 95112 26440 95154 26480
rect 95194 26440 95236 26480
rect 95276 26440 95318 26480
rect 95358 26440 95400 26480
rect 95072 26431 95440 26440
rect 3112 25724 3480 25733
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3112 25675 3480 25684
rect 18232 25724 18600 25733
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18232 25675 18600 25684
rect 33352 25724 33720 25733
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33352 25675 33720 25684
rect 48472 25724 48840 25733
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48472 25675 48840 25684
rect 63592 25724 63960 25733
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63592 25675 63960 25684
rect 78712 25724 79080 25733
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 78712 25675 79080 25684
rect 93832 25724 94200 25733
rect 93872 25684 93914 25724
rect 93954 25684 93996 25724
rect 94036 25684 94078 25724
rect 94118 25684 94160 25724
rect 93832 25675 94200 25684
rect 4352 24968 4720 24977
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4352 24919 4720 24928
rect 19472 24968 19840 24977
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19472 24919 19840 24928
rect 34592 24968 34960 24977
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34592 24919 34960 24928
rect 49712 24968 50080 24977
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 49712 24919 50080 24928
rect 64832 24968 65200 24977
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 64832 24919 65200 24928
rect 79952 24968 80320 24977
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 79952 24919 80320 24928
rect 95072 24968 95440 24977
rect 95112 24928 95154 24968
rect 95194 24928 95236 24968
rect 95276 24928 95318 24968
rect 95358 24928 95400 24968
rect 95072 24919 95440 24928
rect 3112 24212 3480 24221
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3112 24163 3480 24172
rect 18232 24212 18600 24221
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18232 24163 18600 24172
rect 33352 24212 33720 24221
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33352 24163 33720 24172
rect 48472 24212 48840 24221
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48472 24163 48840 24172
rect 63592 24212 63960 24221
rect 63632 24172 63674 24212
rect 63714 24172 63756 24212
rect 63796 24172 63838 24212
rect 63878 24172 63920 24212
rect 63592 24163 63960 24172
rect 78712 24212 79080 24221
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 78712 24163 79080 24172
rect 93832 24212 94200 24221
rect 93872 24172 93914 24212
rect 93954 24172 93996 24212
rect 94036 24172 94078 24212
rect 94118 24172 94160 24212
rect 93832 24163 94200 24172
rect 4352 23456 4720 23465
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4352 23407 4720 23416
rect 19472 23456 19840 23465
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19472 23407 19840 23416
rect 34592 23456 34960 23465
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34592 23407 34960 23416
rect 49712 23456 50080 23465
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 49712 23407 50080 23416
rect 64832 23456 65200 23465
rect 64872 23416 64914 23456
rect 64954 23416 64996 23456
rect 65036 23416 65078 23456
rect 65118 23416 65160 23456
rect 64832 23407 65200 23416
rect 79952 23456 80320 23465
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 79952 23407 80320 23416
rect 95072 23456 95440 23465
rect 95112 23416 95154 23456
rect 95194 23416 95236 23456
rect 95276 23416 95318 23456
rect 95358 23416 95400 23456
rect 95072 23407 95440 23416
rect 3112 22700 3480 22709
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3112 22651 3480 22660
rect 18232 22700 18600 22709
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18232 22651 18600 22660
rect 33352 22700 33720 22709
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33352 22651 33720 22660
rect 48472 22700 48840 22709
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48472 22651 48840 22660
rect 63592 22700 63960 22709
rect 63632 22660 63674 22700
rect 63714 22660 63756 22700
rect 63796 22660 63838 22700
rect 63878 22660 63920 22700
rect 63592 22651 63960 22660
rect 78712 22700 79080 22709
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 78712 22651 79080 22660
rect 93832 22700 94200 22709
rect 93872 22660 93914 22700
rect 93954 22660 93996 22700
rect 94036 22660 94078 22700
rect 94118 22660 94160 22700
rect 93832 22651 94200 22660
rect 4352 21944 4720 21953
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4352 21895 4720 21904
rect 19472 21944 19840 21953
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19472 21895 19840 21904
rect 34592 21944 34960 21953
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34592 21895 34960 21904
rect 49712 21944 50080 21953
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 49712 21895 50080 21904
rect 64832 21944 65200 21953
rect 64872 21904 64914 21944
rect 64954 21904 64996 21944
rect 65036 21904 65078 21944
rect 65118 21904 65160 21944
rect 64832 21895 65200 21904
rect 79952 21944 80320 21953
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 79952 21895 80320 21904
rect 95072 21944 95440 21953
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95072 21895 95440 21904
rect 3112 21188 3480 21197
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3112 21139 3480 21148
rect 18232 21188 18600 21197
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18232 21139 18600 21148
rect 33352 21188 33720 21197
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33352 21139 33720 21148
rect 48472 21188 48840 21197
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48472 21139 48840 21148
rect 63592 21188 63960 21197
rect 63632 21148 63674 21188
rect 63714 21148 63756 21188
rect 63796 21148 63838 21188
rect 63878 21148 63920 21188
rect 63592 21139 63960 21148
rect 78712 21188 79080 21197
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 78712 21139 79080 21148
rect 93832 21188 94200 21197
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 93832 21139 94200 21148
rect 4352 20432 4720 20441
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4352 20383 4720 20392
rect 19472 20432 19840 20441
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19472 20383 19840 20392
rect 34592 20432 34960 20441
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34592 20383 34960 20392
rect 49712 20432 50080 20441
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 49712 20383 50080 20392
rect 64832 20432 65200 20441
rect 64872 20392 64914 20432
rect 64954 20392 64996 20432
rect 65036 20392 65078 20432
rect 65118 20392 65160 20432
rect 64832 20383 65200 20392
rect 79952 20432 80320 20441
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 79952 20383 80320 20392
rect 95072 20432 95440 20441
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95072 20383 95440 20392
rect 3112 19676 3480 19685
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3112 19627 3480 19636
rect 18232 19676 18600 19685
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18232 19627 18600 19636
rect 33352 19676 33720 19685
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33352 19627 33720 19636
rect 48472 19676 48840 19685
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48472 19627 48840 19636
rect 63592 19676 63960 19685
rect 63632 19636 63674 19676
rect 63714 19636 63756 19676
rect 63796 19636 63838 19676
rect 63878 19636 63920 19676
rect 63592 19627 63960 19636
rect 78712 19676 79080 19685
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 78712 19627 79080 19636
rect 93832 19676 94200 19685
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 93832 19627 94200 19636
rect 4352 18920 4720 18929
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4352 18871 4720 18880
rect 19472 18920 19840 18929
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19472 18871 19840 18880
rect 34592 18920 34960 18929
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34592 18871 34960 18880
rect 49712 18920 50080 18929
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 49712 18871 50080 18880
rect 64832 18920 65200 18929
rect 64872 18880 64914 18920
rect 64954 18880 64996 18920
rect 65036 18880 65078 18920
rect 65118 18880 65160 18920
rect 64832 18871 65200 18880
rect 79952 18920 80320 18929
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 79952 18871 80320 18880
rect 95072 18920 95440 18929
rect 95112 18880 95154 18920
rect 95194 18880 95236 18920
rect 95276 18880 95318 18920
rect 95358 18880 95400 18920
rect 95072 18871 95440 18880
rect 3112 18164 3480 18173
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3112 18115 3480 18124
rect 18232 18164 18600 18173
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18232 18115 18600 18124
rect 33352 18164 33720 18173
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33352 18115 33720 18124
rect 48472 18164 48840 18173
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48472 18115 48840 18124
rect 63592 18164 63960 18173
rect 63632 18124 63674 18164
rect 63714 18124 63756 18164
rect 63796 18124 63838 18164
rect 63878 18124 63920 18164
rect 63592 18115 63960 18124
rect 78712 18164 79080 18173
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 78712 18115 79080 18124
rect 93832 18164 94200 18173
rect 93872 18124 93914 18164
rect 93954 18124 93996 18164
rect 94036 18124 94078 18164
rect 94118 18124 94160 18164
rect 93832 18115 94200 18124
rect 4352 17408 4720 17417
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4352 17359 4720 17368
rect 19472 17408 19840 17417
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19472 17359 19840 17368
rect 34592 17408 34960 17417
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34592 17359 34960 17368
rect 49712 17408 50080 17417
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 49712 17359 50080 17368
rect 64832 17408 65200 17417
rect 64872 17368 64914 17408
rect 64954 17368 64996 17408
rect 65036 17368 65078 17408
rect 65118 17368 65160 17408
rect 64832 17359 65200 17368
rect 79952 17408 80320 17417
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 79952 17359 80320 17368
rect 95072 17408 95440 17417
rect 95112 17368 95154 17408
rect 95194 17368 95236 17408
rect 95276 17368 95318 17408
rect 95358 17368 95400 17408
rect 95072 17359 95440 17368
rect 3112 16652 3480 16661
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3112 16603 3480 16612
rect 18232 16652 18600 16661
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18232 16603 18600 16612
rect 33352 16652 33720 16661
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33352 16603 33720 16612
rect 48472 16652 48840 16661
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48472 16603 48840 16612
rect 63592 16652 63960 16661
rect 63632 16612 63674 16652
rect 63714 16612 63756 16652
rect 63796 16612 63838 16652
rect 63878 16612 63920 16652
rect 63592 16603 63960 16612
rect 78712 16652 79080 16661
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 78712 16603 79080 16612
rect 93832 16652 94200 16661
rect 93872 16612 93914 16652
rect 93954 16612 93996 16652
rect 94036 16612 94078 16652
rect 94118 16612 94160 16652
rect 93832 16603 94200 16612
rect 4352 15896 4720 15905
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4352 15847 4720 15856
rect 19472 15896 19840 15905
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19472 15847 19840 15856
rect 34592 15896 34960 15905
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34592 15847 34960 15856
rect 49712 15896 50080 15905
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 49712 15847 50080 15856
rect 64832 15896 65200 15905
rect 64872 15856 64914 15896
rect 64954 15856 64996 15896
rect 65036 15856 65078 15896
rect 65118 15856 65160 15896
rect 64832 15847 65200 15856
rect 79952 15896 80320 15905
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 79952 15847 80320 15856
rect 95072 15896 95440 15905
rect 95112 15856 95154 15896
rect 95194 15856 95236 15896
rect 95276 15856 95318 15896
rect 95358 15856 95400 15896
rect 95072 15847 95440 15856
rect 3112 15140 3480 15149
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3112 15091 3480 15100
rect 18232 15140 18600 15149
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18232 15091 18600 15100
rect 33352 15140 33720 15149
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 33352 15091 33720 15100
rect 48472 15140 48840 15149
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48472 15091 48840 15100
rect 63592 15140 63960 15149
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63592 15091 63960 15100
rect 78712 15140 79080 15149
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 78712 15091 79080 15100
rect 93832 15140 94200 15149
rect 93872 15100 93914 15140
rect 93954 15100 93996 15140
rect 94036 15100 94078 15140
rect 94118 15100 94160 15140
rect 93832 15091 94200 15100
rect 4352 14384 4720 14393
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4352 14335 4720 14344
rect 19472 14384 19840 14393
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19472 14335 19840 14344
rect 34592 14384 34960 14393
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34592 14335 34960 14344
rect 49712 14384 50080 14393
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 49712 14335 50080 14344
rect 64832 14384 65200 14393
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 64832 14335 65200 14344
rect 79952 14384 80320 14393
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 79952 14335 80320 14344
rect 95072 14384 95440 14393
rect 95112 14344 95154 14384
rect 95194 14344 95236 14384
rect 95276 14344 95318 14384
rect 95358 14344 95400 14384
rect 95072 14335 95440 14344
rect 3112 13628 3480 13637
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3112 13579 3480 13588
rect 18232 13628 18600 13637
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18232 13579 18600 13588
rect 33352 13628 33720 13637
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33352 13579 33720 13588
rect 48472 13628 48840 13637
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48472 13579 48840 13588
rect 63592 13628 63960 13637
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63592 13579 63960 13588
rect 78712 13628 79080 13637
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 78712 13579 79080 13588
rect 93832 13628 94200 13637
rect 93872 13588 93914 13628
rect 93954 13588 93996 13628
rect 94036 13588 94078 13628
rect 94118 13588 94160 13628
rect 93832 13579 94200 13588
rect 4352 12872 4720 12881
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4352 12823 4720 12832
rect 19472 12872 19840 12881
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19472 12823 19840 12832
rect 34592 12872 34960 12881
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34592 12823 34960 12832
rect 49712 12872 50080 12881
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 49712 12823 50080 12832
rect 64832 12872 65200 12881
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 64832 12823 65200 12832
rect 79952 12872 80320 12881
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 79952 12823 80320 12832
rect 95072 12872 95440 12881
rect 95112 12832 95154 12872
rect 95194 12832 95236 12872
rect 95276 12832 95318 12872
rect 95358 12832 95400 12872
rect 95072 12823 95440 12832
rect 3112 12116 3480 12125
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3112 12067 3480 12076
rect 18232 12116 18600 12125
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18232 12067 18600 12076
rect 33352 12116 33720 12125
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33352 12067 33720 12076
rect 48472 12116 48840 12125
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48472 12067 48840 12076
rect 63592 12116 63960 12125
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63592 12067 63960 12076
rect 78712 12116 79080 12125
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 78712 12067 79080 12076
rect 93832 12116 94200 12125
rect 93872 12076 93914 12116
rect 93954 12076 93996 12116
rect 94036 12076 94078 12116
rect 94118 12076 94160 12116
rect 93832 12067 94200 12076
rect 4352 11360 4720 11369
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4352 11311 4720 11320
rect 19472 11360 19840 11369
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19472 11311 19840 11320
rect 34592 11360 34960 11369
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34592 11311 34960 11320
rect 49712 11360 50080 11369
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 49712 11311 50080 11320
rect 64832 11360 65200 11369
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 64832 11311 65200 11320
rect 79952 11360 80320 11369
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 79952 11311 80320 11320
rect 95072 11360 95440 11369
rect 95112 11320 95154 11360
rect 95194 11320 95236 11360
rect 95276 11320 95318 11360
rect 95358 11320 95400 11360
rect 95072 11311 95440 11320
rect 3112 10604 3480 10613
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3112 10555 3480 10564
rect 18232 10604 18600 10613
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18232 10555 18600 10564
rect 33352 10604 33720 10613
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33352 10555 33720 10564
rect 48472 10604 48840 10613
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48472 10555 48840 10564
rect 63592 10604 63960 10613
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63592 10555 63960 10564
rect 78712 10604 79080 10613
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 78712 10555 79080 10564
rect 93832 10604 94200 10613
rect 93872 10564 93914 10604
rect 93954 10564 93996 10604
rect 94036 10564 94078 10604
rect 94118 10564 94160 10604
rect 93832 10555 94200 10564
rect 4352 9848 4720 9857
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4352 9799 4720 9808
rect 19472 9848 19840 9857
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19472 9799 19840 9808
rect 34592 9848 34960 9857
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34592 9799 34960 9808
rect 49712 9848 50080 9857
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 49712 9799 50080 9808
rect 64832 9848 65200 9857
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 64832 9799 65200 9808
rect 79952 9848 80320 9857
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 79952 9799 80320 9808
rect 95072 9848 95440 9857
rect 95112 9808 95154 9848
rect 95194 9808 95236 9848
rect 95276 9808 95318 9848
rect 95358 9808 95400 9848
rect 95072 9799 95440 9808
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 18232 9092 18600 9101
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18232 9043 18600 9052
rect 33352 9092 33720 9101
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33352 9043 33720 9052
rect 48472 9092 48840 9101
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48472 9043 48840 9052
rect 63592 9092 63960 9101
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63592 9043 63960 9052
rect 78712 9092 79080 9101
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 78712 9043 79080 9052
rect 93832 9092 94200 9101
rect 93872 9052 93914 9092
rect 93954 9052 93996 9092
rect 94036 9052 94078 9092
rect 94118 9052 94160 9092
rect 93832 9043 94200 9052
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 19472 8336 19840 8345
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19472 8287 19840 8296
rect 34592 8336 34960 8345
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34592 8287 34960 8296
rect 49712 8336 50080 8345
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 49712 8287 50080 8296
rect 64832 8336 65200 8345
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 64832 8287 65200 8296
rect 79952 8336 80320 8345
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 79952 8287 80320 8296
rect 95072 8336 95440 8345
rect 95112 8296 95154 8336
rect 95194 8296 95236 8336
rect 95276 8296 95318 8336
rect 95358 8296 95400 8336
rect 95072 8287 95440 8296
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 18232 7580 18600 7589
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18232 7531 18600 7540
rect 33352 7580 33720 7589
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33352 7531 33720 7540
rect 48472 7580 48840 7589
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48472 7531 48840 7540
rect 63592 7580 63960 7589
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63592 7531 63960 7540
rect 78712 7580 79080 7589
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 78712 7531 79080 7540
rect 93832 7580 94200 7589
rect 93872 7540 93914 7580
rect 93954 7540 93996 7580
rect 94036 7540 94078 7580
rect 94118 7540 94160 7580
rect 93832 7531 94200 7540
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 19472 6824 19840 6833
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19472 6775 19840 6784
rect 34592 6824 34960 6833
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34592 6775 34960 6784
rect 49712 6824 50080 6833
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 49712 6775 50080 6784
rect 64832 6824 65200 6833
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 64832 6775 65200 6784
rect 79952 6824 80320 6833
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 79952 6775 80320 6784
rect 95072 6824 95440 6833
rect 95112 6784 95154 6824
rect 95194 6784 95236 6824
rect 95276 6784 95318 6824
rect 95358 6784 95400 6824
rect 95072 6775 95440 6784
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 18232 6068 18600 6077
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18232 6019 18600 6028
rect 33352 6068 33720 6077
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33352 6019 33720 6028
rect 48472 6068 48840 6077
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48472 6019 48840 6028
rect 63592 6068 63960 6077
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63592 6019 63960 6028
rect 78712 6068 79080 6077
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 78712 6019 79080 6028
rect 93832 6068 94200 6077
rect 93872 6028 93914 6068
rect 93954 6028 93996 6068
rect 94036 6028 94078 6068
rect 94118 6028 94160 6068
rect 93832 6019 94200 6028
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 19472 5312 19840 5321
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19472 5263 19840 5272
rect 34592 5312 34960 5321
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34592 5263 34960 5272
rect 49712 5312 50080 5321
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 49712 5263 50080 5272
rect 64832 5312 65200 5321
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 64832 5263 65200 5272
rect 79952 5312 80320 5321
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 79952 5263 80320 5272
rect 95072 5312 95440 5321
rect 95112 5272 95154 5312
rect 95194 5272 95236 5312
rect 95276 5272 95318 5312
rect 95358 5272 95400 5312
rect 95072 5263 95440 5272
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 18232 4556 18600 4565
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18232 4507 18600 4516
rect 33352 4556 33720 4565
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33352 4507 33720 4516
rect 48472 4556 48840 4565
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48472 4507 48840 4516
rect 63592 4556 63960 4565
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63592 4507 63960 4516
rect 78712 4556 79080 4565
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 78712 4507 79080 4516
rect 93832 4556 94200 4565
rect 93872 4516 93914 4556
rect 93954 4516 93996 4556
rect 94036 4516 94078 4556
rect 94118 4516 94160 4556
rect 93832 4507 94200 4516
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 19472 3800 19840 3809
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19472 3751 19840 3760
rect 34592 3800 34960 3809
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34592 3751 34960 3760
rect 49712 3800 50080 3809
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 49712 3751 50080 3760
rect 64832 3800 65200 3809
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 64832 3751 65200 3760
rect 79952 3800 80320 3809
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 79952 3751 80320 3760
rect 95072 3800 95440 3809
rect 95112 3760 95154 3800
rect 95194 3760 95236 3800
rect 95276 3760 95318 3800
rect 95358 3760 95400 3800
rect 95072 3751 95440 3760
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 18232 3044 18600 3053
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18232 2995 18600 3004
rect 33352 3044 33720 3053
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33352 2995 33720 3004
rect 48472 3044 48840 3053
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48472 2995 48840 3004
rect 63592 3044 63960 3053
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63592 2995 63960 3004
rect 78712 3044 79080 3053
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 78712 2995 79080 3004
rect 93832 3044 94200 3053
rect 93872 3004 93914 3044
rect 93954 3004 93996 3044
rect 94036 3004 94078 3044
rect 94118 3004 94160 3044
rect 93832 2995 94200 3004
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 19472 2288 19840 2297
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19472 2239 19840 2248
rect 34592 2288 34960 2297
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34592 2239 34960 2248
rect 49712 2288 50080 2297
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 49712 2239 50080 2248
rect 64832 2288 65200 2297
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 64832 2239 65200 2248
rect 79952 2288 80320 2297
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 79952 2239 80320 2248
rect 95072 2288 95440 2297
rect 95112 2248 95154 2288
rect 95194 2248 95236 2288
rect 95276 2248 95318 2288
rect 95358 2248 95400 2288
rect 95072 2239 95440 2248
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 18232 1532 18600 1541
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18232 1483 18600 1492
rect 33352 1532 33720 1541
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33352 1483 33720 1492
rect 48472 1532 48840 1541
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48472 1483 48840 1492
rect 63592 1532 63960 1541
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63592 1483 63960 1492
rect 78712 1532 79080 1541
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 78712 1483 79080 1492
rect 93832 1532 94200 1541
rect 93872 1492 93914 1532
rect 93954 1492 93996 1532
rect 94036 1492 94078 1532
rect 94118 1492 94160 1532
rect 93832 1483 94200 1492
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
rect 19472 776 19840 785
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19472 727 19840 736
rect 34592 776 34960 785
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34592 727 34960 736
rect 49712 776 50080 785
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 49712 727 50080 736
rect 64832 776 65200 785
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 64832 727 65200 736
rect 79952 776 80320 785
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 79952 727 80320 736
rect 95072 776 95440 785
rect 95112 736 95154 776
rect 95194 736 95236 776
rect 95276 736 95318 776
rect 95358 736 95400 776
rect 95072 727 95440 736
<< via4 >>
rect 3112 81628 3152 81668
rect 3194 81628 3234 81668
rect 3276 81628 3316 81668
rect 3358 81628 3398 81668
rect 3440 81628 3480 81668
rect 18232 81628 18272 81668
rect 18314 81628 18354 81668
rect 18396 81628 18436 81668
rect 18478 81628 18518 81668
rect 18560 81628 18600 81668
rect 33352 81628 33392 81668
rect 33434 81628 33474 81668
rect 33516 81628 33556 81668
rect 33598 81628 33638 81668
rect 33680 81628 33720 81668
rect 48472 81628 48512 81668
rect 48554 81628 48594 81668
rect 48636 81628 48676 81668
rect 48718 81628 48758 81668
rect 48800 81628 48840 81668
rect 63592 81628 63632 81668
rect 63674 81628 63714 81668
rect 63756 81628 63796 81668
rect 63838 81628 63878 81668
rect 63920 81628 63960 81668
rect 78712 81628 78752 81668
rect 78794 81628 78834 81668
rect 78876 81628 78916 81668
rect 78958 81628 78998 81668
rect 79040 81628 79080 81668
rect 93832 81628 93872 81668
rect 93914 81628 93954 81668
rect 93996 81628 94036 81668
rect 94078 81628 94118 81668
rect 94160 81628 94200 81668
rect 4352 80872 4392 80912
rect 4434 80872 4474 80912
rect 4516 80872 4556 80912
rect 4598 80872 4638 80912
rect 4680 80872 4720 80912
rect 19472 80872 19512 80912
rect 19554 80872 19594 80912
rect 19636 80872 19676 80912
rect 19718 80872 19758 80912
rect 19800 80872 19840 80912
rect 34592 80872 34632 80912
rect 34674 80872 34714 80912
rect 34756 80872 34796 80912
rect 34838 80872 34878 80912
rect 34920 80872 34960 80912
rect 49712 80872 49752 80912
rect 49794 80872 49834 80912
rect 49876 80872 49916 80912
rect 49958 80872 49998 80912
rect 50040 80872 50080 80912
rect 64832 80872 64872 80912
rect 64914 80872 64954 80912
rect 64996 80872 65036 80912
rect 65078 80872 65118 80912
rect 65160 80872 65200 80912
rect 79952 80872 79992 80912
rect 80034 80872 80074 80912
rect 80116 80872 80156 80912
rect 80198 80872 80238 80912
rect 80280 80872 80320 80912
rect 95072 80872 95112 80912
rect 95154 80872 95194 80912
rect 95236 80872 95276 80912
rect 95318 80872 95358 80912
rect 95400 80872 95440 80912
rect 3112 80116 3152 80156
rect 3194 80116 3234 80156
rect 3276 80116 3316 80156
rect 3358 80116 3398 80156
rect 3440 80116 3480 80156
rect 18232 80116 18272 80156
rect 18314 80116 18354 80156
rect 18396 80116 18436 80156
rect 18478 80116 18518 80156
rect 18560 80116 18600 80156
rect 33352 80116 33392 80156
rect 33434 80116 33474 80156
rect 33516 80116 33556 80156
rect 33598 80116 33638 80156
rect 33680 80116 33720 80156
rect 48472 80116 48512 80156
rect 48554 80116 48594 80156
rect 48636 80116 48676 80156
rect 48718 80116 48758 80156
rect 48800 80116 48840 80156
rect 63592 80116 63632 80156
rect 63674 80116 63714 80156
rect 63756 80116 63796 80156
rect 63838 80116 63878 80156
rect 63920 80116 63960 80156
rect 78712 80116 78752 80156
rect 78794 80116 78834 80156
rect 78876 80116 78916 80156
rect 78958 80116 78998 80156
rect 79040 80116 79080 80156
rect 93832 80116 93872 80156
rect 93914 80116 93954 80156
rect 93996 80116 94036 80156
rect 94078 80116 94118 80156
rect 94160 80116 94200 80156
rect 4352 79360 4392 79400
rect 4434 79360 4474 79400
rect 4516 79360 4556 79400
rect 4598 79360 4638 79400
rect 4680 79360 4720 79400
rect 19472 79360 19512 79400
rect 19554 79360 19594 79400
rect 19636 79360 19676 79400
rect 19718 79360 19758 79400
rect 19800 79360 19840 79400
rect 34592 79360 34632 79400
rect 34674 79360 34714 79400
rect 34756 79360 34796 79400
rect 34838 79360 34878 79400
rect 34920 79360 34960 79400
rect 49712 79360 49752 79400
rect 49794 79360 49834 79400
rect 49876 79360 49916 79400
rect 49958 79360 49998 79400
rect 50040 79360 50080 79400
rect 64832 79360 64872 79400
rect 64914 79360 64954 79400
rect 64996 79360 65036 79400
rect 65078 79360 65118 79400
rect 65160 79360 65200 79400
rect 79952 79360 79992 79400
rect 80034 79360 80074 79400
rect 80116 79360 80156 79400
rect 80198 79360 80238 79400
rect 80280 79360 80320 79400
rect 95072 79360 95112 79400
rect 95154 79360 95194 79400
rect 95236 79360 95276 79400
rect 95318 79360 95358 79400
rect 95400 79360 95440 79400
rect 3112 78604 3152 78644
rect 3194 78604 3234 78644
rect 3276 78604 3316 78644
rect 3358 78604 3398 78644
rect 3440 78604 3480 78644
rect 18232 78604 18272 78644
rect 18314 78604 18354 78644
rect 18396 78604 18436 78644
rect 18478 78604 18518 78644
rect 18560 78604 18600 78644
rect 33352 78604 33392 78644
rect 33434 78604 33474 78644
rect 33516 78604 33556 78644
rect 33598 78604 33638 78644
rect 33680 78604 33720 78644
rect 48472 78604 48512 78644
rect 48554 78604 48594 78644
rect 48636 78604 48676 78644
rect 48718 78604 48758 78644
rect 48800 78604 48840 78644
rect 63592 78604 63632 78644
rect 63674 78604 63714 78644
rect 63756 78604 63796 78644
rect 63838 78604 63878 78644
rect 63920 78604 63960 78644
rect 78712 78604 78752 78644
rect 78794 78604 78834 78644
rect 78876 78604 78916 78644
rect 78958 78604 78998 78644
rect 79040 78604 79080 78644
rect 93832 78604 93872 78644
rect 93914 78604 93954 78644
rect 93996 78604 94036 78644
rect 94078 78604 94118 78644
rect 94160 78604 94200 78644
rect 4352 77848 4392 77888
rect 4434 77848 4474 77888
rect 4516 77848 4556 77888
rect 4598 77848 4638 77888
rect 4680 77848 4720 77888
rect 19472 77848 19512 77888
rect 19554 77848 19594 77888
rect 19636 77848 19676 77888
rect 19718 77848 19758 77888
rect 19800 77848 19840 77888
rect 34592 77848 34632 77888
rect 34674 77848 34714 77888
rect 34756 77848 34796 77888
rect 34838 77848 34878 77888
rect 34920 77848 34960 77888
rect 49712 77848 49752 77888
rect 49794 77848 49834 77888
rect 49876 77848 49916 77888
rect 49958 77848 49998 77888
rect 50040 77848 50080 77888
rect 64832 77848 64872 77888
rect 64914 77848 64954 77888
rect 64996 77848 65036 77888
rect 65078 77848 65118 77888
rect 65160 77848 65200 77888
rect 79952 77848 79992 77888
rect 80034 77848 80074 77888
rect 80116 77848 80156 77888
rect 80198 77848 80238 77888
rect 80280 77848 80320 77888
rect 95072 77848 95112 77888
rect 95154 77848 95194 77888
rect 95236 77848 95276 77888
rect 95318 77848 95358 77888
rect 95400 77848 95440 77888
rect 3112 77092 3152 77132
rect 3194 77092 3234 77132
rect 3276 77092 3316 77132
rect 3358 77092 3398 77132
rect 3440 77092 3480 77132
rect 18232 77092 18272 77132
rect 18314 77092 18354 77132
rect 18396 77092 18436 77132
rect 18478 77092 18518 77132
rect 18560 77092 18600 77132
rect 33352 77092 33392 77132
rect 33434 77092 33474 77132
rect 33516 77092 33556 77132
rect 33598 77092 33638 77132
rect 33680 77092 33720 77132
rect 48472 77092 48512 77132
rect 48554 77092 48594 77132
rect 48636 77092 48676 77132
rect 48718 77092 48758 77132
rect 48800 77092 48840 77132
rect 63592 77092 63632 77132
rect 63674 77092 63714 77132
rect 63756 77092 63796 77132
rect 63838 77092 63878 77132
rect 63920 77092 63960 77132
rect 78712 77092 78752 77132
rect 78794 77092 78834 77132
rect 78876 77092 78916 77132
rect 78958 77092 78998 77132
rect 79040 77092 79080 77132
rect 93832 77092 93872 77132
rect 93914 77092 93954 77132
rect 93996 77092 94036 77132
rect 94078 77092 94118 77132
rect 94160 77092 94200 77132
rect 4352 76336 4392 76376
rect 4434 76336 4474 76376
rect 4516 76336 4556 76376
rect 4598 76336 4638 76376
rect 4680 76336 4720 76376
rect 19472 76336 19512 76376
rect 19554 76336 19594 76376
rect 19636 76336 19676 76376
rect 19718 76336 19758 76376
rect 19800 76336 19840 76376
rect 34592 76336 34632 76376
rect 34674 76336 34714 76376
rect 34756 76336 34796 76376
rect 34838 76336 34878 76376
rect 34920 76336 34960 76376
rect 49712 76336 49752 76376
rect 49794 76336 49834 76376
rect 49876 76336 49916 76376
rect 49958 76336 49998 76376
rect 50040 76336 50080 76376
rect 64832 76336 64872 76376
rect 64914 76336 64954 76376
rect 64996 76336 65036 76376
rect 65078 76336 65118 76376
rect 65160 76336 65200 76376
rect 79952 76336 79992 76376
rect 80034 76336 80074 76376
rect 80116 76336 80156 76376
rect 80198 76336 80238 76376
rect 80280 76336 80320 76376
rect 95072 76336 95112 76376
rect 95154 76336 95194 76376
rect 95236 76336 95276 76376
rect 95318 76336 95358 76376
rect 95400 76336 95440 76376
rect 3112 75580 3152 75620
rect 3194 75580 3234 75620
rect 3276 75580 3316 75620
rect 3358 75580 3398 75620
rect 3440 75580 3480 75620
rect 18232 75580 18272 75620
rect 18314 75580 18354 75620
rect 18396 75580 18436 75620
rect 18478 75580 18518 75620
rect 18560 75580 18600 75620
rect 33352 75580 33392 75620
rect 33434 75580 33474 75620
rect 33516 75580 33556 75620
rect 33598 75580 33638 75620
rect 33680 75580 33720 75620
rect 48472 75580 48512 75620
rect 48554 75580 48594 75620
rect 48636 75580 48676 75620
rect 48718 75580 48758 75620
rect 48800 75580 48840 75620
rect 63592 75580 63632 75620
rect 63674 75580 63714 75620
rect 63756 75580 63796 75620
rect 63838 75580 63878 75620
rect 63920 75580 63960 75620
rect 78712 75580 78752 75620
rect 78794 75580 78834 75620
rect 78876 75580 78916 75620
rect 78958 75580 78998 75620
rect 79040 75580 79080 75620
rect 93832 75580 93872 75620
rect 93914 75580 93954 75620
rect 93996 75580 94036 75620
rect 94078 75580 94118 75620
rect 94160 75580 94200 75620
rect 4352 74824 4392 74864
rect 4434 74824 4474 74864
rect 4516 74824 4556 74864
rect 4598 74824 4638 74864
rect 4680 74824 4720 74864
rect 19472 74824 19512 74864
rect 19554 74824 19594 74864
rect 19636 74824 19676 74864
rect 19718 74824 19758 74864
rect 19800 74824 19840 74864
rect 34592 74824 34632 74864
rect 34674 74824 34714 74864
rect 34756 74824 34796 74864
rect 34838 74824 34878 74864
rect 34920 74824 34960 74864
rect 49712 74824 49752 74864
rect 49794 74824 49834 74864
rect 49876 74824 49916 74864
rect 49958 74824 49998 74864
rect 50040 74824 50080 74864
rect 64832 74824 64872 74864
rect 64914 74824 64954 74864
rect 64996 74824 65036 74864
rect 65078 74824 65118 74864
rect 65160 74824 65200 74864
rect 79952 74824 79992 74864
rect 80034 74824 80074 74864
rect 80116 74824 80156 74864
rect 80198 74824 80238 74864
rect 80280 74824 80320 74864
rect 95072 74824 95112 74864
rect 95154 74824 95194 74864
rect 95236 74824 95276 74864
rect 95318 74824 95358 74864
rect 95400 74824 95440 74864
rect 3112 74068 3152 74108
rect 3194 74068 3234 74108
rect 3276 74068 3316 74108
rect 3358 74068 3398 74108
rect 3440 74068 3480 74108
rect 18232 74068 18272 74108
rect 18314 74068 18354 74108
rect 18396 74068 18436 74108
rect 18478 74068 18518 74108
rect 18560 74068 18600 74108
rect 33352 74068 33392 74108
rect 33434 74068 33474 74108
rect 33516 74068 33556 74108
rect 33598 74068 33638 74108
rect 33680 74068 33720 74108
rect 48472 74068 48512 74108
rect 48554 74068 48594 74108
rect 48636 74068 48676 74108
rect 48718 74068 48758 74108
rect 48800 74068 48840 74108
rect 63592 74068 63632 74108
rect 63674 74068 63714 74108
rect 63756 74068 63796 74108
rect 63838 74068 63878 74108
rect 63920 74068 63960 74108
rect 78712 74068 78752 74108
rect 78794 74068 78834 74108
rect 78876 74068 78916 74108
rect 78958 74068 78998 74108
rect 79040 74068 79080 74108
rect 93832 74068 93872 74108
rect 93914 74068 93954 74108
rect 93996 74068 94036 74108
rect 94078 74068 94118 74108
rect 94160 74068 94200 74108
rect 4352 73312 4392 73352
rect 4434 73312 4474 73352
rect 4516 73312 4556 73352
rect 4598 73312 4638 73352
rect 4680 73312 4720 73352
rect 19472 73312 19512 73352
rect 19554 73312 19594 73352
rect 19636 73312 19676 73352
rect 19718 73312 19758 73352
rect 19800 73312 19840 73352
rect 34592 73312 34632 73352
rect 34674 73312 34714 73352
rect 34756 73312 34796 73352
rect 34838 73312 34878 73352
rect 34920 73312 34960 73352
rect 49712 73312 49752 73352
rect 49794 73312 49834 73352
rect 49876 73312 49916 73352
rect 49958 73312 49998 73352
rect 50040 73312 50080 73352
rect 64832 73312 64872 73352
rect 64914 73312 64954 73352
rect 64996 73312 65036 73352
rect 65078 73312 65118 73352
rect 65160 73312 65200 73352
rect 79952 73312 79992 73352
rect 80034 73312 80074 73352
rect 80116 73312 80156 73352
rect 80198 73312 80238 73352
rect 80280 73312 80320 73352
rect 95072 73312 95112 73352
rect 95154 73312 95194 73352
rect 95236 73312 95276 73352
rect 95318 73312 95358 73352
rect 95400 73312 95440 73352
rect 3112 72556 3152 72596
rect 3194 72556 3234 72596
rect 3276 72556 3316 72596
rect 3358 72556 3398 72596
rect 3440 72556 3480 72596
rect 18232 72556 18272 72596
rect 18314 72556 18354 72596
rect 18396 72556 18436 72596
rect 18478 72556 18518 72596
rect 18560 72556 18600 72596
rect 33352 72556 33392 72596
rect 33434 72556 33474 72596
rect 33516 72556 33556 72596
rect 33598 72556 33638 72596
rect 33680 72556 33720 72596
rect 48472 72556 48512 72596
rect 48554 72556 48594 72596
rect 48636 72556 48676 72596
rect 48718 72556 48758 72596
rect 48800 72556 48840 72596
rect 63592 72556 63632 72596
rect 63674 72556 63714 72596
rect 63756 72556 63796 72596
rect 63838 72556 63878 72596
rect 63920 72556 63960 72596
rect 78712 72556 78752 72596
rect 78794 72556 78834 72596
rect 78876 72556 78916 72596
rect 78958 72556 78998 72596
rect 79040 72556 79080 72596
rect 93832 72556 93872 72596
rect 93914 72556 93954 72596
rect 93996 72556 94036 72596
rect 94078 72556 94118 72596
rect 94160 72556 94200 72596
rect 4352 71800 4392 71840
rect 4434 71800 4474 71840
rect 4516 71800 4556 71840
rect 4598 71800 4638 71840
rect 4680 71800 4720 71840
rect 19472 71800 19512 71840
rect 19554 71800 19594 71840
rect 19636 71800 19676 71840
rect 19718 71800 19758 71840
rect 19800 71800 19840 71840
rect 34592 71800 34632 71840
rect 34674 71800 34714 71840
rect 34756 71800 34796 71840
rect 34838 71800 34878 71840
rect 34920 71800 34960 71840
rect 49712 71800 49752 71840
rect 49794 71800 49834 71840
rect 49876 71800 49916 71840
rect 49958 71800 49998 71840
rect 50040 71800 50080 71840
rect 64832 71800 64872 71840
rect 64914 71800 64954 71840
rect 64996 71800 65036 71840
rect 65078 71800 65118 71840
rect 65160 71800 65200 71840
rect 79952 71800 79992 71840
rect 80034 71800 80074 71840
rect 80116 71800 80156 71840
rect 80198 71800 80238 71840
rect 80280 71800 80320 71840
rect 95072 71800 95112 71840
rect 95154 71800 95194 71840
rect 95236 71800 95276 71840
rect 95318 71800 95358 71840
rect 95400 71800 95440 71840
rect 3112 71044 3152 71084
rect 3194 71044 3234 71084
rect 3276 71044 3316 71084
rect 3358 71044 3398 71084
rect 3440 71044 3480 71084
rect 18232 71044 18272 71084
rect 18314 71044 18354 71084
rect 18396 71044 18436 71084
rect 18478 71044 18518 71084
rect 18560 71044 18600 71084
rect 33352 71044 33392 71084
rect 33434 71044 33474 71084
rect 33516 71044 33556 71084
rect 33598 71044 33638 71084
rect 33680 71044 33720 71084
rect 48472 71044 48512 71084
rect 48554 71044 48594 71084
rect 48636 71044 48676 71084
rect 48718 71044 48758 71084
rect 48800 71044 48840 71084
rect 63592 71044 63632 71084
rect 63674 71044 63714 71084
rect 63756 71044 63796 71084
rect 63838 71044 63878 71084
rect 63920 71044 63960 71084
rect 78712 71044 78752 71084
rect 78794 71044 78834 71084
rect 78876 71044 78916 71084
rect 78958 71044 78998 71084
rect 79040 71044 79080 71084
rect 93832 71044 93872 71084
rect 93914 71044 93954 71084
rect 93996 71044 94036 71084
rect 94078 71044 94118 71084
rect 94160 71044 94200 71084
rect 4352 70288 4392 70328
rect 4434 70288 4474 70328
rect 4516 70288 4556 70328
rect 4598 70288 4638 70328
rect 4680 70288 4720 70328
rect 19472 70288 19512 70328
rect 19554 70288 19594 70328
rect 19636 70288 19676 70328
rect 19718 70288 19758 70328
rect 19800 70288 19840 70328
rect 34592 70288 34632 70328
rect 34674 70288 34714 70328
rect 34756 70288 34796 70328
rect 34838 70288 34878 70328
rect 34920 70288 34960 70328
rect 49712 70288 49752 70328
rect 49794 70288 49834 70328
rect 49876 70288 49916 70328
rect 49958 70288 49998 70328
rect 50040 70288 50080 70328
rect 64832 70288 64872 70328
rect 64914 70288 64954 70328
rect 64996 70288 65036 70328
rect 65078 70288 65118 70328
rect 65160 70288 65200 70328
rect 79952 70288 79992 70328
rect 80034 70288 80074 70328
rect 80116 70288 80156 70328
rect 80198 70288 80238 70328
rect 80280 70288 80320 70328
rect 95072 70288 95112 70328
rect 95154 70288 95194 70328
rect 95236 70288 95276 70328
rect 95318 70288 95358 70328
rect 95400 70288 95440 70328
rect 3112 69532 3152 69572
rect 3194 69532 3234 69572
rect 3276 69532 3316 69572
rect 3358 69532 3398 69572
rect 3440 69532 3480 69572
rect 18232 69532 18272 69572
rect 18314 69532 18354 69572
rect 18396 69532 18436 69572
rect 18478 69532 18518 69572
rect 18560 69532 18600 69572
rect 33352 69532 33392 69572
rect 33434 69532 33474 69572
rect 33516 69532 33556 69572
rect 33598 69532 33638 69572
rect 33680 69532 33720 69572
rect 48472 69532 48512 69572
rect 48554 69532 48594 69572
rect 48636 69532 48676 69572
rect 48718 69532 48758 69572
rect 48800 69532 48840 69572
rect 63592 69532 63632 69572
rect 63674 69532 63714 69572
rect 63756 69532 63796 69572
rect 63838 69532 63878 69572
rect 63920 69532 63960 69572
rect 78712 69532 78752 69572
rect 78794 69532 78834 69572
rect 78876 69532 78916 69572
rect 78958 69532 78998 69572
rect 79040 69532 79080 69572
rect 93832 69532 93872 69572
rect 93914 69532 93954 69572
rect 93996 69532 94036 69572
rect 94078 69532 94118 69572
rect 94160 69532 94200 69572
rect 4352 68776 4392 68816
rect 4434 68776 4474 68816
rect 4516 68776 4556 68816
rect 4598 68776 4638 68816
rect 4680 68776 4720 68816
rect 19472 68776 19512 68816
rect 19554 68776 19594 68816
rect 19636 68776 19676 68816
rect 19718 68776 19758 68816
rect 19800 68776 19840 68816
rect 34592 68776 34632 68816
rect 34674 68776 34714 68816
rect 34756 68776 34796 68816
rect 34838 68776 34878 68816
rect 34920 68776 34960 68816
rect 49712 68776 49752 68816
rect 49794 68776 49834 68816
rect 49876 68776 49916 68816
rect 49958 68776 49998 68816
rect 50040 68776 50080 68816
rect 64832 68776 64872 68816
rect 64914 68776 64954 68816
rect 64996 68776 65036 68816
rect 65078 68776 65118 68816
rect 65160 68776 65200 68816
rect 79952 68776 79992 68816
rect 80034 68776 80074 68816
rect 80116 68776 80156 68816
rect 80198 68776 80238 68816
rect 80280 68776 80320 68816
rect 95072 68776 95112 68816
rect 95154 68776 95194 68816
rect 95236 68776 95276 68816
rect 95318 68776 95358 68816
rect 95400 68776 95440 68816
rect 3112 68020 3152 68060
rect 3194 68020 3234 68060
rect 3276 68020 3316 68060
rect 3358 68020 3398 68060
rect 3440 68020 3480 68060
rect 18232 68020 18272 68060
rect 18314 68020 18354 68060
rect 18396 68020 18436 68060
rect 18478 68020 18518 68060
rect 18560 68020 18600 68060
rect 33352 68020 33392 68060
rect 33434 68020 33474 68060
rect 33516 68020 33556 68060
rect 33598 68020 33638 68060
rect 33680 68020 33720 68060
rect 48472 68020 48512 68060
rect 48554 68020 48594 68060
rect 48636 68020 48676 68060
rect 48718 68020 48758 68060
rect 48800 68020 48840 68060
rect 63592 68020 63632 68060
rect 63674 68020 63714 68060
rect 63756 68020 63796 68060
rect 63838 68020 63878 68060
rect 63920 68020 63960 68060
rect 78712 68020 78752 68060
rect 78794 68020 78834 68060
rect 78876 68020 78916 68060
rect 78958 68020 78998 68060
rect 79040 68020 79080 68060
rect 93832 68020 93872 68060
rect 93914 68020 93954 68060
rect 93996 68020 94036 68060
rect 94078 68020 94118 68060
rect 94160 68020 94200 68060
rect 4352 67264 4392 67304
rect 4434 67264 4474 67304
rect 4516 67264 4556 67304
rect 4598 67264 4638 67304
rect 4680 67264 4720 67304
rect 19472 67264 19512 67304
rect 19554 67264 19594 67304
rect 19636 67264 19676 67304
rect 19718 67264 19758 67304
rect 19800 67264 19840 67304
rect 34592 67264 34632 67304
rect 34674 67264 34714 67304
rect 34756 67264 34796 67304
rect 34838 67264 34878 67304
rect 34920 67264 34960 67304
rect 49712 67264 49752 67304
rect 49794 67264 49834 67304
rect 49876 67264 49916 67304
rect 49958 67264 49998 67304
rect 50040 67264 50080 67304
rect 64832 67264 64872 67304
rect 64914 67264 64954 67304
rect 64996 67264 65036 67304
rect 65078 67264 65118 67304
rect 65160 67264 65200 67304
rect 79952 67264 79992 67304
rect 80034 67264 80074 67304
rect 80116 67264 80156 67304
rect 80198 67264 80238 67304
rect 80280 67264 80320 67304
rect 95072 67264 95112 67304
rect 95154 67264 95194 67304
rect 95236 67264 95276 67304
rect 95318 67264 95358 67304
rect 95400 67264 95440 67304
rect 3112 66508 3152 66548
rect 3194 66508 3234 66548
rect 3276 66508 3316 66548
rect 3358 66508 3398 66548
rect 3440 66508 3480 66548
rect 18232 66508 18272 66548
rect 18314 66508 18354 66548
rect 18396 66508 18436 66548
rect 18478 66508 18518 66548
rect 18560 66508 18600 66548
rect 33352 66508 33392 66548
rect 33434 66508 33474 66548
rect 33516 66508 33556 66548
rect 33598 66508 33638 66548
rect 33680 66508 33720 66548
rect 48472 66508 48512 66548
rect 48554 66508 48594 66548
rect 48636 66508 48676 66548
rect 48718 66508 48758 66548
rect 48800 66508 48840 66548
rect 63592 66508 63632 66548
rect 63674 66508 63714 66548
rect 63756 66508 63796 66548
rect 63838 66508 63878 66548
rect 63920 66508 63960 66548
rect 78712 66508 78752 66548
rect 78794 66508 78834 66548
rect 78876 66508 78916 66548
rect 78958 66508 78998 66548
rect 79040 66508 79080 66548
rect 93832 66508 93872 66548
rect 93914 66508 93954 66548
rect 93996 66508 94036 66548
rect 94078 66508 94118 66548
rect 94160 66508 94200 66548
rect 4352 65752 4392 65792
rect 4434 65752 4474 65792
rect 4516 65752 4556 65792
rect 4598 65752 4638 65792
rect 4680 65752 4720 65792
rect 19472 65752 19512 65792
rect 19554 65752 19594 65792
rect 19636 65752 19676 65792
rect 19718 65752 19758 65792
rect 19800 65752 19840 65792
rect 34592 65752 34632 65792
rect 34674 65752 34714 65792
rect 34756 65752 34796 65792
rect 34838 65752 34878 65792
rect 34920 65752 34960 65792
rect 49712 65752 49752 65792
rect 49794 65752 49834 65792
rect 49876 65752 49916 65792
rect 49958 65752 49998 65792
rect 50040 65752 50080 65792
rect 64832 65752 64872 65792
rect 64914 65752 64954 65792
rect 64996 65752 65036 65792
rect 65078 65752 65118 65792
rect 65160 65752 65200 65792
rect 79952 65752 79992 65792
rect 80034 65752 80074 65792
rect 80116 65752 80156 65792
rect 80198 65752 80238 65792
rect 80280 65752 80320 65792
rect 95072 65752 95112 65792
rect 95154 65752 95194 65792
rect 95236 65752 95276 65792
rect 95318 65752 95358 65792
rect 95400 65752 95440 65792
rect 3112 64996 3152 65036
rect 3194 64996 3234 65036
rect 3276 64996 3316 65036
rect 3358 64996 3398 65036
rect 3440 64996 3480 65036
rect 18232 64996 18272 65036
rect 18314 64996 18354 65036
rect 18396 64996 18436 65036
rect 18478 64996 18518 65036
rect 18560 64996 18600 65036
rect 33352 64996 33392 65036
rect 33434 64996 33474 65036
rect 33516 64996 33556 65036
rect 33598 64996 33638 65036
rect 33680 64996 33720 65036
rect 48472 64996 48512 65036
rect 48554 64996 48594 65036
rect 48636 64996 48676 65036
rect 48718 64996 48758 65036
rect 48800 64996 48840 65036
rect 63592 64996 63632 65036
rect 63674 64996 63714 65036
rect 63756 64996 63796 65036
rect 63838 64996 63878 65036
rect 63920 64996 63960 65036
rect 78712 64996 78752 65036
rect 78794 64996 78834 65036
rect 78876 64996 78916 65036
rect 78958 64996 78998 65036
rect 79040 64996 79080 65036
rect 93832 64996 93872 65036
rect 93914 64996 93954 65036
rect 93996 64996 94036 65036
rect 94078 64996 94118 65036
rect 94160 64996 94200 65036
rect 4352 64240 4392 64280
rect 4434 64240 4474 64280
rect 4516 64240 4556 64280
rect 4598 64240 4638 64280
rect 4680 64240 4720 64280
rect 19472 64240 19512 64280
rect 19554 64240 19594 64280
rect 19636 64240 19676 64280
rect 19718 64240 19758 64280
rect 19800 64240 19840 64280
rect 34592 64240 34632 64280
rect 34674 64240 34714 64280
rect 34756 64240 34796 64280
rect 34838 64240 34878 64280
rect 34920 64240 34960 64280
rect 49712 64240 49752 64280
rect 49794 64240 49834 64280
rect 49876 64240 49916 64280
rect 49958 64240 49998 64280
rect 50040 64240 50080 64280
rect 64832 64240 64872 64280
rect 64914 64240 64954 64280
rect 64996 64240 65036 64280
rect 65078 64240 65118 64280
rect 65160 64240 65200 64280
rect 79952 64240 79992 64280
rect 80034 64240 80074 64280
rect 80116 64240 80156 64280
rect 80198 64240 80238 64280
rect 80280 64240 80320 64280
rect 95072 64240 95112 64280
rect 95154 64240 95194 64280
rect 95236 64240 95276 64280
rect 95318 64240 95358 64280
rect 95400 64240 95440 64280
rect 3112 63484 3152 63524
rect 3194 63484 3234 63524
rect 3276 63484 3316 63524
rect 3358 63484 3398 63524
rect 3440 63484 3480 63524
rect 18232 63484 18272 63524
rect 18314 63484 18354 63524
rect 18396 63484 18436 63524
rect 18478 63484 18518 63524
rect 18560 63484 18600 63524
rect 33352 63484 33392 63524
rect 33434 63484 33474 63524
rect 33516 63484 33556 63524
rect 33598 63484 33638 63524
rect 33680 63484 33720 63524
rect 48472 63484 48512 63524
rect 48554 63484 48594 63524
rect 48636 63484 48676 63524
rect 48718 63484 48758 63524
rect 48800 63484 48840 63524
rect 63592 63484 63632 63524
rect 63674 63484 63714 63524
rect 63756 63484 63796 63524
rect 63838 63484 63878 63524
rect 63920 63484 63960 63524
rect 78712 63484 78752 63524
rect 78794 63484 78834 63524
rect 78876 63484 78916 63524
rect 78958 63484 78998 63524
rect 79040 63484 79080 63524
rect 93832 63484 93872 63524
rect 93914 63484 93954 63524
rect 93996 63484 94036 63524
rect 94078 63484 94118 63524
rect 94160 63484 94200 63524
rect 4352 62728 4392 62768
rect 4434 62728 4474 62768
rect 4516 62728 4556 62768
rect 4598 62728 4638 62768
rect 4680 62728 4720 62768
rect 19472 62728 19512 62768
rect 19554 62728 19594 62768
rect 19636 62728 19676 62768
rect 19718 62728 19758 62768
rect 19800 62728 19840 62768
rect 34592 62728 34632 62768
rect 34674 62728 34714 62768
rect 34756 62728 34796 62768
rect 34838 62728 34878 62768
rect 34920 62728 34960 62768
rect 49712 62728 49752 62768
rect 49794 62728 49834 62768
rect 49876 62728 49916 62768
rect 49958 62728 49998 62768
rect 50040 62728 50080 62768
rect 64832 62728 64872 62768
rect 64914 62728 64954 62768
rect 64996 62728 65036 62768
rect 65078 62728 65118 62768
rect 65160 62728 65200 62768
rect 79952 62728 79992 62768
rect 80034 62728 80074 62768
rect 80116 62728 80156 62768
rect 80198 62728 80238 62768
rect 80280 62728 80320 62768
rect 95072 62728 95112 62768
rect 95154 62728 95194 62768
rect 95236 62728 95276 62768
rect 95318 62728 95358 62768
rect 95400 62728 95440 62768
rect 3112 61972 3152 62012
rect 3194 61972 3234 62012
rect 3276 61972 3316 62012
rect 3358 61972 3398 62012
rect 3440 61972 3480 62012
rect 18232 61972 18272 62012
rect 18314 61972 18354 62012
rect 18396 61972 18436 62012
rect 18478 61972 18518 62012
rect 18560 61972 18600 62012
rect 33352 61972 33392 62012
rect 33434 61972 33474 62012
rect 33516 61972 33556 62012
rect 33598 61972 33638 62012
rect 33680 61972 33720 62012
rect 48472 61972 48512 62012
rect 48554 61972 48594 62012
rect 48636 61972 48676 62012
rect 48718 61972 48758 62012
rect 48800 61972 48840 62012
rect 63592 61972 63632 62012
rect 63674 61972 63714 62012
rect 63756 61972 63796 62012
rect 63838 61972 63878 62012
rect 63920 61972 63960 62012
rect 78712 61972 78752 62012
rect 78794 61972 78834 62012
rect 78876 61972 78916 62012
rect 78958 61972 78998 62012
rect 79040 61972 79080 62012
rect 93832 61972 93872 62012
rect 93914 61972 93954 62012
rect 93996 61972 94036 62012
rect 94078 61972 94118 62012
rect 94160 61972 94200 62012
rect 4352 61216 4392 61256
rect 4434 61216 4474 61256
rect 4516 61216 4556 61256
rect 4598 61216 4638 61256
rect 4680 61216 4720 61256
rect 19472 61216 19512 61256
rect 19554 61216 19594 61256
rect 19636 61216 19676 61256
rect 19718 61216 19758 61256
rect 19800 61216 19840 61256
rect 34592 61216 34632 61256
rect 34674 61216 34714 61256
rect 34756 61216 34796 61256
rect 34838 61216 34878 61256
rect 34920 61216 34960 61256
rect 49712 61216 49752 61256
rect 49794 61216 49834 61256
rect 49876 61216 49916 61256
rect 49958 61216 49998 61256
rect 50040 61216 50080 61256
rect 64832 61216 64872 61256
rect 64914 61216 64954 61256
rect 64996 61216 65036 61256
rect 65078 61216 65118 61256
rect 65160 61216 65200 61256
rect 79952 61216 79992 61256
rect 80034 61216 80074 61256
rect 80116 61216 80156 61256
rect 80198 61216 80238 61256
rect 80280 61216 80320 61256
rect 95072 61216 95112 61256
rect 95154 61216 95194 61256
rect 95236 61216 95276 61256
rect 95318 61216 95358 61256
rect 95400 61216 95440 61256
rect 3112 60460 3152 60500
rect 3194 60460 3234 60500
rect 3276 60460 3316 60500
rect 3358 60460 3398 60500
rect 3440 60460 3480 60500
rect 18232 60460 18272 60500
rect 18314 60460 18354 60500
rect 18396 60460 18436 60500
rect 18478 60460 18518 60500
rect 18560 60460 18600 60500
rect 33352 60460 33392 60500
rect 33434 60460 33474 60500
rect 33516 60460 33556 60500
rect 33598 60460 33638 60500
rect 33680 60460 33720 60500
rect 48472 60460 48512 60500
rect 48554 60460 48594 60500
rect 48636 60460 48676 60500
rect 48718 60460 48758 60500
rect 48800 60460 48840 60500
rect 63592 60460 63632 60500
rect 63674 60460 63714 60500
rect 63756 60460 63796 60500
rect 63838 60460 63878 60500
rect 63920 60460 63960 60500
rect 78712 60460 78752 60500
rect 78794 60460 78834 60500
rect 78876 60460 78916 60500
rect 78958 60460 78998 60500
rect 79040 60460 79080 60500
rect 93832 60460 93872 60500
rect 93914 60460 93954 60500
rect 93996 60460 94036 60500
rect 94078 60460 94118 60500
rect 94160 60460 94200 60500
rect 4352 59704 4392 59744
rect 4434 59704 4474 59744
rect 4516 59704 4556 59744
rect 4598 59704 4638 59744
rect 4680 59704 4720 59744
rect 19472 59704 19512 59744
rect 19554 59704 19594 59744
rect 19636 59704 19676 59744
rect 19718 59704 19758 59744
rect 19800 59704 19840 59744
rect 34592 59704 34632 59744
rect 34674 59704 34714 59744
rect 34756 59704 34796 59744
rect 34838 59704 34878 59744
rect 34920 59704 34960 59744
rect 49712 59704 49752 59744
rect 49794 59704 49834 59744
rect 49876 59704 49916 59744
rect 49958 59704 49998 59744
rect 50040 59704 50080 59744
rect 64832 59704 64872 59744
rect 64914 59704 64954 59744
rect 64996 59704 65036 59744
rect 65078 59704 65118 59744
rect 65160 59704 65200 59744
rect 79952 59704 79992 59744
rect 80034 59704 80074 59744
rect 80116 59704 80156 59744
rect 80198 59704 80238 59744
rect 80280 59704 80320 59744
rect 95072 59704 95112 59744
rect 95154 59704 95194 59744
rect 95236 59704 95276 59744
rect 95318 59704 95358 59744
rect 95400 59704 95440 59744
rect 3112 58948 3152 58988
rect 3194 58948 3234 58988
rect 3276 58948 3316 58988
rect 3358 58948 3398 58988
rect 3440 58948 3480 58988
rect 18232 58948 18272 58988
rect 18314 58948 18354 58988
rect 18396 58948 18436 58988
rect 18478 58948 18518 58988
rect 18560 58948 18600 58988
rect 33352 58948 33392 58988
rect 33434 58948 33474 58988
rect 33516 58948 33556 58988
rect 33598 58948 33638 58988
rect 33680 58948 33720 58988
rect 48472 58948 48512 58988
rect 48554 58948 48594 58988
rect 48636 58948 48676 58988
rect 48718 58948 48758 58988
rect 48800 58948 48840 58988
rect 63592 58948 63632 58988
rect 63674 58948 63714 58988
rect 63756 58948 63796 58988
rect 63838 58948 63878 58988
rect 63920 58948 63960 58988
rect 78712 58948 78752 58988
rect 78794 58948 78834 58988
rect 78876 58948 78916 58988
rect 78958 58948 78998 58988
rect 79040 58948 79080 58988
rect 93832 58948 93872 58988
rect 93914 58948 93954 58988
rect 93996 58948 94036 58988
rect 94078 58948 94118 58988
rect 94160 58948 94200 58988
rect 4352 58192 4392 58232
rect 4434 58192 4474 58232
rect 4516 58192 4556 58232
rect 4598 58192 4638 58232
rect 4680 58192 4720 58232
rect 19472 58192 19512 58232
rect 19554 58192 19594 58232
rect 19636 58192 19676 58232
rect 19718 58192 19758 58232
rect 19800 58192 19840 58232
rect 34592 58192 34632 58232
rect 34674 58192 34714 58232
rect 34756 58192 34796 58232
rect 34838 58192 34878 58232
rect 34920 58192 34960 58232
rect 49712 58192 49752 58232
rect 49794 58192 49834 58232
rect 49876 58192 49916 58232
rect 49958 58192 49998 58232
rect 50040 58192 50080 58232
rect 64832 58192 64872 58232
rect 64914 58192 64954 58232
rect 64996 58192 65036 58232
rect 65078 58192 65118 58232
rect 65160 58192 65200 58232
rect 79952 58192 79992 58232
rect 80034 58192 80074 58232
rect 80116 58192 80156 58232
rect 80198 58192 80238 58232
rect 80280 58192 80320 58232
rect 95072 58192 95112 58232
rect 95154 58192 95194 58232
rect 95236 58192 95276 58232
rect 95318 58192 95358 58232
rect 95400 58192 95440 58232
rect 3112 57436 3152 57476
rect 3194 57436 3234 57476
rect 3276 57436 3316 57476
rect 3358 57436 3398 57476
rect 3440 57436 3480 57476
rect 18232 57436 18272 57476
rect 18314 57436 18354 57476
rect 18396 57436 18436 57476
rect 18478 57436 18518 57476
rect 18560 57436 18600 57476
rect 33352 57436 33392 57476
rect 33434 57436 33474 57476
rect 33516 57436 33556 57476
rect 33598 57436 33638 57476
rect 33680 57436 33720 57476
rect 48472 57436 48512 57476
rect 48554 57436 48594 57476
rect 48636 57436 48676 57476
rect 48718 57436 48758 57476
rect 48800 57436 48840 57476
rect 63592 57436 63632 57476
rect 63674 57436 63714 57476
rect 63756 57436 63796 57476
rect 63838 57436 63878 57476
rect 63920 57436 63960 57476
rect 78712 57436 78752 57476
rect 78794 57436 78834 57476
rect 78876 57436 78916 57476
rect 78958 57436 78998 57476
rect 79040 57436 79080 57476
rect 93832 57436 93872 57476
rect 93914 57436 93954 57476
rect 93996 57436 94036 57476
rect 94078 57436 94118 57476
rect 94160 57436 94200 57476
rect 4352 56680 4392 56720
rect 4434 56680 4474 56720
rect 4516 56680 4556 56720
rect 4598 56680 4638 56720
rect 4680 56680 4720 56720
rect 19472 56680 19512 56720
rect 19554 56680 19594 56720
rect 19636 56680 19676 56720
rect 19718 56680 19758 56720
rect 19800 56680 19840 56720
rect 34592 56680 34632 56720
rect 34674 56680 34714 56720
rect 34756 56680 34796 56720
rect 34838 56680 34878 56720
rect 34920 56680 34960 56720
rect 49712 56680 49752 56720
rect 49794 56680 49834 56720
rect 49876 56680 49916 56720
rect 49958 56680 49998 56720
rect 50040 56680 50080 56720
rect 64832 56680 64872 56720
rect 64914 56680 64954 56720
rect 64996 56680 65036 56720
rect 65078 56680 65118 56720
rect 65160 56680 65200 56720
rect 79952 56680 79992 56720
rect 80034 56680 80074 56720
rect 80116 56680 80156 56720
rect 80198 56680 80238 56720
rect 80280 56680 80320 56720
rect 95072 56680 95112 56720
rect 95154 56680 95194 56720
rect 95236 56680 95276 56720
rect 95318 56680 95358 56720
rect 95400 56680 95440 56720
rect 3112 55924 3152 55964
rect 3194 55924 3234 55964
rect 3276 55924 3316 55964
rect 3358 55924 3398 55964
rect 3440 55924 3480 55964
rect 18232 55924 18272 55964
rect 18314 55924 18354 55964
rect 18396 55924 18436 55964
rect 18478 55924 18518 55964
rect 18560 55924 18600 55964
rect 33352 55924 33392 55964
rect 33434 55924 33474 55964
rect 33516 55924 33556 55964
rect 33598 55924 33638 55964
rect 33680 55924 33720 55964
rect 48472 55924 48512 55964
rect 48554 55924 48594 55964
rect 48636 55924 48676 55964
rect 48718 55924 48758 55964
rect 48800 55924 48840 55964
rect 63592 55924 63632 55964
rect 63674 55924 63714 55964
rect 63756 55924 63796 55964
rect 63838 55924 63878 55964
rect 63920 55924 63960 55964
rect 78712 55924 78752 55964
rect 78794 55924 78834 55964
rect 78876 55924 78916 55964
rect 78958 55924 78998 55964
rect 79040 55924 79080 55964
rect 93832 55924 93872 55964
rect 93914 55924 93954 55964
rect 93996 55924 94036 55964
rect 94078 55924 94118 55964
rect 94160 55924 94200 55964
rect 4352 55168 4392 55208
rect 4434 55168 4474 55208
rect 4516 55168 4556 55208
rect 4598 55168 4638 55208
rect 4680 55168 4720 55208
rect 19472 55168 19512 55208
rect 19554 55168 19594 55208
rect 19636 55168 19676 55208
rect 19718 55168 19758 55208
rect 19800 55168 19840 55208
rect 34592 55168 34632 55208
rect 34674 55168 34714 55208
rect 34756 55168 34796 55208
rect 34838 55168 34878 55208
rect 34920 55168 34960 55208
rect 49712 55168 49752 55208
rect 49794 55168 49834 55208
rect 49876 55168 49916 55208
rect 49958 55168 49998 55208
rect 50040 55168 50080 55208
rect 64832 55168 64872 55208
rect 64914 55168 64954 55208
rect 64996 55168 65036 55208
rect 65078 55168 65118 55208
rect 65160 55168 65200 55208
rect 79952 55168 79992 55208
rect 80034 55168 80074 55208
rect 80116 55168 80156 55208
rect 80198 55168 80238 55208
rect 80280 55168 80320 55208
rect 95072 55168 95112 55208
rect 95154 55168 95194 55208
rect 95236 55168 95276 55208
rect 95318 55168 95358 55208
rect 95400 55168 95440 55208
rect 3112 54412 3152 54452
rect 3194 54412 3234 54452
rect 3276 54412 3316 54452
rect 3358 54412 3398 54452
rect 3440 54412 3480 54452
rect 18232 54412 18272 54452
rect 18314 54412 18354 54452
rect 18396 54412 18436 54452
rect 18478 54412 18518 54452
rect 18560 54412 18600 54452
rect 33352 54412 33392 54452
rect 33434 54412 33474 54452
rect 33516 54412 33556 54452
rect 33598 54412 33638 54452
rect 33680 54412 33720 54452
rect 48472 54412 48512 54452
rect 48554 54412 48594 54452
rect 48636 54412 48676 54452
rect 48718 54412 48758 54452
rect 48800 54412 48840 54452
rect 63592 54412 63632 54452
rect 63674 54412 63714 54452
rect 63756 54412 63796 54452
rect 63838 54412 63878 54452
rect 63920 54412 63960 54452
rect 78712 54412 78752 54452
rect 78794 54412 78834 54452
rect 78876 54412 78916 54452
rect 78958 54412 78998 54452
rect 79040 54412 79080 54452
rect 93832 54412 93872 54452
rect 93914 54412 93954 54452
rect 93996 54412 94036 54452
rect 94078 54412 94118 54452
rect 94160 54412 94200 54452
rect 4352 53656 4392 53696
rect 4434 53656 4474 53696
rect 4516 53656 4556 53696
rect 4598 53656 4638 53696
rect 4680 53656 4720 53696
rect 19472 53656 19512 53696
rect 19554 53656 19594 53696
rect 19636 53656 19676 53696
rect 19718 53656 19758 53696
rect 19800 53656 19840 53696
rect 34592 53656 34632 53696
rect 34674 53656 34714 53696
rect 34756 53656 34796 53696
rect 34838 53656 34878 53696
rect 34920 53656 34960 53696
rect 49712 53656 49752 53696
rect 49794 53656 49834 53696
rect 49876 53656 49916 53696
rect 49958 53656 49998 53696
rect 50040 53656 50080 53696
rect 64832 53656 64872 53696
rect 64914 53656 64954 53696
rect 64996 53656 65036 53696
rect 65078 53656 65118 53696
rect 65160 53656 65200 53696
rect 79952 53656 79992 53696
rect 80034 53656 80074 53696
rect 80116 53656 80156 53696
rect 80198 53656 80238 53696
rect 80280 53656 80320 53696
rect 95072 53656 95112 53696
rect 95154 53656 95194 53696
rect 95236 53656 95276 53696
rect 95318 53656 95358 53696
rect 95400 53656 95440 53696
rect 3112 52900 3152 52940
rect 3194 52900 3234 52940
rect 3276 52900 3316 52940
rect 3358 52900 3398 52940
rect 3440 52900 3480 52940
rect 18232 52900 18272 52940
rect 18314 52900 18354 52940
rect 18396 52900 18436 52940
rect 18478 52900 18518 52940
rect 18560 52900 18600 52940
rect 33352 52900 33392 52940
rect 33434 52900 33474 52940
rect 33516 52900 33556 52940
rect 33598 52900 33638 52940
rect 33680 52900 33720 52940
rect 48472 52900 48512 52940
rect 48554 52900 48594 52940
rect 48636 52900 48676 52940
rect 48718 52900 48758 52940
rect 48800 52900 48840 52940
rect 63592 52900 63632 52940
rect 63674 52900 63714 52940
rect 63756 52900 63796 52940
rect 63838 52900 63878 52940
rect 63920 52900 63960 52940
rect 78712 52900 78752 52940
rect 78794 52900 78834 52940
rect 78876 52900 78916 52940
rect 78958 52900 78998 52940
rect 79040 52900 79080 52940
rect 93832 52900 93872 52940
rect 93914 52900 93954 52940
rect 93996 52900 94036 52940
rect 94078 52900 94118 52940
rect 94160 52900 94200 52940
rect 4352 52144 4392 52184
rect 4434 52144 4474 52184
rect 4516 52144 4556 52184
rect 4598 52144 4638 52184
rect 4680 52144 4720 52184
rect 19472 52144 19512 52184
rect 19554 52144 19594 52184
rect 19636 52144 19676 52184
rect 19718 52144 19758 52184
rect 19800 52144 19840 52184
rect 34592 52144 34632 52184
rect 34674 52144 34714 52184
rect 34756 52144 34796 52184
rect 34838 52144 34878 52184
rect 34920 52144 34960 52184
rect 49712 52144 49752 52184
rect 49794 52144 49834 52184
rect 49876 52144 49916 52184
rect 49958 52144 49998 52184
rect 50040 52144 50080 52184
rect 64832 52144 64872 52184
rect 64914 52144 64954 52184
rect 64996 52144 65036 52184
rect 65078 52144 65118 52184
rect 65160 52144 65200 52184
rect 79952 52144 79992 52184
rect 80034 52144 80074 52184
rect 80116 52144 80156 52184
rect 80198 52144 80238 52184
rect 80280 52144 80320 52184
rect 95072 52144 95112 52184
rect 95154 52144 95194 52184
rect 95236 52144 95276 52184
rect 95318 52144 95358 52184
rect 95400 52144 95440 52184
rect 3112 51388 3152 51428
rect 3194 51388 3234 51428
rect 3276 51388 3316 51428
rect 3358 51388 3398 51428
rect 3440 51388 3480 51428
rect 18232 51388 18272 51428
rect 18314 51388 18354 51428
rect 18396 51388 18436 51428
rect 18478 51388 18518 51428
rect 18560 51388 18600 51428
rect 33352 51388 33392 51428
rect 33434 51388 33474 51428
rect 33516 51388 33556 51428
rect 33598 51388 33638 51428
rect 33680 51388 33720 51428
rect 48472 51388 48512 51428
rect 48554 51388 48594 51428
rect 48636 51388 48676 51428
rect 48718 51388 48758 51428
rect 48800 51388 48840 51428
rect 63592 51388 63632 51428
rect 63674 51388 63714 51428
rect 63756 51388 63796 51428
rect 63838 51388 63878 51428
rect 63920 51388 63960 51428
rect 78712 51388 78752 51428
rect 78794 51388 78834 51428
rect 78876 51388 78916 51428
rect 78958 51388 78998 51428
rect 79040 51388 79080 51428
rect 93832 51388 93872 51428
rect 93914 51388 93954 51428
rect 93996 51388 94036 51428
rect 94078 51388 94118 51428
rect 94160 51388 94200 51428
rect 4352 50632 4392 50672
rect 4434 50632 4474 50672
rect 4516 50632 4556 50672
rect 4598 50632 4638 50672
rect 4680 50632 4720 50672
rect 19472 50632 19512 50672
rect 19554 50632 19594 50672
rect 19636 50632 19676 50672
rect 19718 50632 19758 50672
rect 19800 50632 19840 50672
rect 34592 50632 34632 50672
rect 34674 50632 34714 50672
rect 34756 50632 34796 50672
rect 34838 50632 34878 50672
rect 34920 50632 34960 50672
rect 49712 50632 49752 50672
rect 49794 50632 49834 50672
rect 49876 50632 49916 50672
rect 49958 50632 49998 50672
rect 50040 50632 50080 50672
rect 64832 50632 64872 50672
rect 64914 50632 64954 50672
rect 64996 50632 65036 50672
rect 65078 50632 65118 50672
rect 65160 50632 65200 50672
rect 79952 50632 79992 50672
rect 80034 50632 80074 50672
rect 80116 50632 80156 50672
rect 80198 50632 80238 50672
rect 80280 50632 80320 50672
rect 95072 50632 95112 50672
rect 95154 50632 95194 50672
rect 95236 50632 95276 50672
rect 95318 50632 95358 50672
rect 95400 50632 95440 50672
rect 3112 49876 3152 49916
rect 3194 49876 3234 49916
rect 3276 49876 3316 49916
rect 3358 49876 3398 49916
rect 3440 49876 3480 49916
rect 18232 49876 18272 49916
rect 18314 49876 18354 49916
rect 18396 49876 18436 49916
rect 18478 49876 18518 49916
rect 18560 49876 18600 49916
rect 33352 49876 33392 49916
rect 33434 49876 33474 49916
rect 33516 49876 33556 49916
rect 33598 49876 33638 49916
rect 33680 49876 33720 49916
rect 48472 49876 48512 49916
rect 48554 49876 48594 49916
rect 48636 49876 48676 49916
rect 48718 49876 48758 49916
rect 48800 49876 48840 49916
rect 63592 49876 63632 49916
rect 63674 49876 63714 49916
rect 63756 49876 63796 49916
rect 63838 49876 63878 49916
rect 63920 49876 63960 49916
rect 78712 49876 78752 49916
rect 78794 49876 78834 49916
rect 78876 49876 78916 49916
rect 78958 49876 78998 49916
rect 79040 49876 79080 49916
rect 93832 49876 93872 49916
rect 93914 49876 93954 49916
rect 93996 49876 94036 49916
rect 94078 49876 94118 49916
rect 94160 49876 94200 49916
rect 4352 49120 4392 49160
rect 4434 49120 4474 49160
rect 4516 49120 4556 49160
rect 4598 49120 4638 49160
rect 4680 49120 4720 49160
rect 19472 49120 19512 49160
rect 19554 49120 19594 49160
rect 19636 49120 19676 49160
rect 19718 49120 19758 49160
rect 19800 49120 19840 49160
rect 34592 49120 34632 49160
rect 34674 49120 34714 49160
rect 34756 49120 34796 49160
rect 34838 49120 34878 49160
rect 34920 49120 34960 49160
rect 49712 49120 49752 49160
rect 49794 49120 49834 49160
rect 49876 49120 49916 49160
rect 49958 49120 49998 49160
rect 50040 49120 50080 49160
rect 64832 49120 64872 49160
rect 64914 49120 64954 49160
rect 64996 49120 65036 49160
rect 65078 49120 65118 49160
rect 65160 49120 65200 49160
rect 79952 49120 79992 49160
rect 80034 49120 80074 49160
rect 80116 49120 80156 49160
rect 80198 49120 80238 49160
rect 80280 49120 80320 49160
rect 95072 49120 95112 49160
rect 95154 49120 95194 49160
rect 95236 49120 95276 49160
rect 95318 49120 95358 49160
rect 95400 49120 95440 49160
rect 3112 48364 3152 48404
rect 3194 48364 3234 48404
rect 3276 48364 3316 48404
rect 3358 48364 3398 48404
rect 3440 48364 3480 48404
rect 18232 48364 18272 48404
rect 18314 48364 18354 48404
rect 18396 48364 18436 48404
rect 18478 48364 18518 48404
rect 18560 48364 18600 48404
rect 33352 48364 33392 48404
rect 33434 48364 33474 48404
rect 33516 48364 33556 48404
rect 33598 48364 33638 48404
rect 33680 48364 33720 48404
rect 48472 48364 48512 48404
rect 48554 48364 48594 48404
rect 48636 48364 48676 48404
rect 48718 48364 48758 48404
rect 48800 48364 48840 48404
rect 63592 48364 63632 48404
rect 63674 48364 63714 48404
rect 63756 48364 63796 48404
rect 63838 48364 63878 48404
rect 63920 48364 63960 48404
rect 78712 48364 78752 48404
rect 78794 48364 78834 48404
rect 78876 48364 78916 48404
rect 78958 48364 78998 48404
rect 79040 48364 79080 48404
rect 93832 48364 93872 48404
rect 93914 48364 93954 48404
rect 93996 48364 94036 48404
rect 94078 48364 94118 48404
rect 94160 48364 94200 48404
rect 4352 47608 4392 47648
rect 4434 47608 4474 47648
rect 4516 47608 4556 47648
rect 4598 47608 4638 47648
rect 4680 47608 4720 47648
rect 19472 47608 19512 47648
rect 19554 47608 19594 47648
rect 19636 47608 19676 47648
rect 19718 47608 19758 47648
rect 19800 47608 19840 47648
rect 34592 47608 34632 47648
rect 34674 47608 34714 47648
rect 34756 47608 34796 47648
rect 34838 47608 34878 47648
rect 34920 47608 34960 47648
rect 49712 47608 49752 47648
rect 49794 47608 49834 47648
rect 49876 47608 49916 47648
rect 49958 47608 49998 47648
rect 50040 47608 50080 47648
rect 64832 47608 64872 47648
rect 64914 47608 64954 47648
rect 64996 47608 65036 47648
rect 65078 47608 65118 47648
rect 65160 47608 65200 47648
rect 79952 47608 79992 47648
rect 80034 47608 80074 47648
rect 80116 47608 80156 47648
rect 80198 47608 80238 47648
rect 80280 47608 80320 47648
rect 95072 47608 95112 47648
rect 95154 47608 95194 47648
rect 95236 47608 95276 47648
rect 95318 47608 95358 47648
rect 95400 47608 95440 47648
rect 3112 46852 3152 46892
rect 3194 46852 3234 46892
rect 3276 46852 3316 46892
rect 3358 46852 3398 46892
rect 3440 46852 3480 46892
rect 18232 46852 18272 46892
rect 18314 46852 18354 46892
rect 18396 46852 18436 46892
rect 18478 46852 18518 46892
rect 18560 46852 18600 46892
rect 33352 46852 33392 46892
rect 33434 46852 33474 46892
rect 33516 46852 33556 46892
rect 33598 46852 33638 46892
rect 33680 46852 33720 46892
rect 48472 46852 48512 46892
rect 48554 46852 48594 46892
rect 48636 46852 48676 46892
rect 48718 46852 48758 46892
rect 48800 46852 48840 46892
rect 63592 46852 63632 46892
rect 63674 46852 63714 46892
rect 63756 46852 63796 46892
rect 63838 46852 63878 46892
rect 63920 46852 63960 46892
rect 78712 46852 78752 46892
rect 78794 46852 78834 46892
rect 78876 46852 78916 46892
rect 78958 46852 78998 46892
rect 79040 46852 79080 46892
rect 93832 46852 93872 46892
rect 93914 46852 93954 46892
rect 93996 46852 94036 46892
rect 94078 46852 94118 46892
rect 94160 46852 94200 46892
rect 4352 46096 4392 46136
rect 4434 46096 4474 46136
rect 4516 46096 4556 46136
rect 4598 46096 4638 46136
rect 4680 46096 4720 46136
rect 19472 46096 19512 46136
rect 19554 46096 19594 46136
rect 19636 46096 19676 46136
rect 19718 46096 19758 46136
rect 19800 46096 19840 46136
rect 34592 46096 34632 46136
rect 34674 46096 34714 46136
rect 34756 46096 34796 46136
rect 34838 46096 34878 46136
rect 34920 46096 34960 46136
rect 49712 46096 49752 46136
rect 49794 46096 49834 46136
rect 49876 46096 49916 46136
rect 49958 46096 49998 46136
rect 50040 46096 50080 46136
rect 64832 46096 64872 46136
rect 64914 46096 64954 46136
rect 64996 46096 65036 46136
rect 65078 46096 65118 46136
rect 65160 46096 65200 46136
rect 79952 46096 79992 46136
rect 80034 46096 80074 46136
rect 80116 46096 80156 46136
rect 80198 46096 80238 46136
rect 80280 46096 80320 46136
rect 95072 46096 95112 46136
rect 95154 46096 95194 46136
rect 95236 46096 95276 46136
rect 95318 46096 95358 46136
rect 95400 46096 95440 46136
rect 3112 45340 3152 45380
rect 3194 45340 3234 45380
rect 3276 45340 3316 45380
rect 3358 45340 3398 45380
rect 3440 45340 3480 45380
rect 18232 45340 18272 45380
rect 18314 45340 18354 45380
rect 18396 45340 18436 45380
rect 18478 45340 18518 45380
rect 18560 45340 18600 45380
rect 33352 45340 33392 45380
rect 33434 45340 33474 45380
rect 33516 45340 33556 45380
rect 33598 45340 33638 45380
rect 33680 45340 33720 45380
rect 48472 45340 48512 45380
rect 48554 45340 48594 45380
rect 48636 45340 48676 45380
rect 48718 45340 48758 45380
rect 48800 45340 48840 45380
rect 63592 45340 63632 45380
rect 63674 45340 63714 45380
rect 63756 45340 63796 45380
rect 63838 45340 63878 45380
rect 63920 45340 63960 45380
rect 78712 45340 78752 45380
rect 78794 45340 78834 45380
rect 78876 45340 78916 45380
rect 78958 45340 78998 45380
rect 79040 45340 79080 45380
rect 93832 45340 93872 45380
rect 93914 45340 93954 45380
rect 93996 45340 94036 45380
rect 94078 45340 94118 45380
rect 94160 45340 94200 45380
rect 4352 44584 4392 44624
rect 4434 44584 4474 44624
rect 4516 44584 4556 44624
rect 4598 44584 4638 44624
rect 4680 44584 4720 44624
rect 19472 44584 19512 44624
rect 19554 44584 19594 44624
rect 19636 44584 19676 44624
rect 19718 44584 19758 44624
rect 19800 44584 19840 44624
rect 34592 44584 34632 44624
rect 34674 44584 34714 44624
rect 34756 44584 34796 44624
rect 34838 44584 34878 44624
rect 34920 44584 34960 44624
rect 49712 44584 49752 44624
rect 49794 44584 49834 44624
rect 49876 44584 49916 44624
rect 49958 44584 49998 44624
rect 50040 44584 50080 44624
rect 64832 44584 64872 44624
rect 64914 44584 64954 44624
rect 64996 44584 65036 44624
rect 65078 44584 65118 44624
rect 65160 44584 65200 44624
rect 79952 44584 79992 44624
rect 80034 44584 80074 44624
rect 80116 44584 80156 44624
rect 80198 44584 80238 44624
rect 80280 44584 80320 44624
rect 95072 44584 95112 44624
rect 95154 44584 95194 44624
rect 95236 44584 95276 44624
rect 95318 44584 95358 44624
rect 95400 44584 95440 44624
rect 3112 43828 3152 43868
rect 3194 43828 3234 43868
rect 3276 43828 3316 43868
rect 3358 43828 3398 43868
rect 3440 43828 3480 43868
rect 18232 43828 18272 43868
rect 18314 43828 18354 43868
rect 18396 43828 18436 43868
rect 18478 43828 18518 43868
rect 18560 43828 18600 43868
rect 33352 43828 33392 43868
rect 33434 43828 33474 43868
rect 33516 43828 33556 43868
rect 33598 43828 33638 43868
rect 33680 43828 33720 43868
rect 48472 43828 48512 43868
rect 48554 43828 48594 43868
rect 48636 43828 48676 43868
rect 48718 43828 48758 43868
rect 48800 43828 48840 43868
rect 63592 43828 63632 43868
rect 63674 43828 63714 43868
rect 63756 43828 63796 43868
rect 63838 43828 63878 43868
rect 63920 43828 63960 43868
rect 78712 43828 78752 43868
rect 78794 43828 78834 43868
rect 78876 43828 78916 43868
rect 78958 43828 78998 43868
rect 79040 43828 79080 43868
rect 93832 43828 93872 43868
rect 93914 43828 93954 43868
rect 93996 43828 94036 43868
rect 94078 43828 94118 43868
rect 94160 43828 94200 43868
rect 4352 43072 4392 43112
rect 4434 43072 4474 43112
rect 4516 43072 4556 43112
rect 4598 43072 4638 43112
rect 4680 43072 4720 43112
rect 19472 43072 19512 43112
rect 19554 43072 19594 43112
rect 19636 43072 19676 43112
rect 19718 43072 19758 43112
rect 19800 43072 19840 43112
rect 34592 43072 34632 43112
rect 34674 43072 34714 43112
rect 34756 43072 34796 43112
rect 34838 43072 34878 43112
rect 34920 43072 34960 43112
rect 49712 43072 49752 43112
rect 49794 43072 49834 43112
rect 49876 43072 49916 43112
rect 49958 43072 49998 43112
rect 50040 43072 50080 43112
rect 64832 43072 64872 43112
rect 64914 43072 64954 43112
rect 64996 43072 65036 43112
rect 65078 43072 65118 43112
rect 65160 43072 65200 43112
rect 79952 43072 79992 43112
rect 80034 43072 80074 43112
rect 80116 43072 80156 43112
rect 80198 43072 80238 43112
rect 80280 43072 80320 43112
rect 95072 43072 95112 43112
rect 95154 43072 95194 43112
rect 95236 43072 95276 43112
rect 95318 43072 95358 43112
rect 95400 43072 95440 43112
rect 3112 42316 3152 42356
rect 3194 42316 3234 42356
rect 3276 42316 3316 42356
rect 3358 42316 3398 42356
rect 3440 42316 3480 42356
rect 18232 42316 18272 42356
rect 18314 42316 18354 42356
rect 18396 42316 18436 42356
rect 18478 42316 18518 42356
rect 18560 42316 18600 42356
rect 33352 42316 33392 42356
rect 33434 42316 33474 42356
rect 33516 42316 33556 42356
rect 33598 42316 33638 42356
rect 33680 42316 33720 42356
rect 48472 42316 48512 42356
rect 48554 42316 48594 42356
rect 48636 42316 48676 42356
rect 48718 42316 48758 42356
rect 48800 42316 48840 42356
rect 63592 42316 63632 42356
rect 63674 42316 63714 42356
rect 63756 42316 63796 42356
rect 63838 42316 63878 42356
rect 63920 42316 63960 42356
rect 78712 42316 78752 42356
rect 78794 42316 78834 42356
rect 78876 42316 78916 42356
rect 78958 42316 78998 42356
rect 79040 42316 79080 42356
rect 93832 42316 93872 42356
rect 93914 42316 93954 42356
rect 93996 42316 94036 42356
rect 94078 42316 94118 42356
rect 94160 42316 94200 42356
rect 4352 41560 4392 41600
rect 4434 41560 4474 41600
rect 4516 41560 4556 41600
rect 4598 41560 4638 41600
rect 4680 41560 4720 41600
rect 19472 41560 19512 41600
rect 19554 41560 19594 41600
rect 19636 41560 19676 41600
rect 19718 41560 19758 41600
rect 19800 41560 19840 41600
rect 34592 41560 34632 41600
rect 34674 41560 34714 41600
rect 34756 41560 34796 41600
rect 34838 41560 34878 41600
rect 34920 41560 34960 41600
rect 49712 41560 49752 41600
rect 49794 41560 49834 41600
rect 49876 41560 49916 41600
rect 49958 41560 49998 41600
rect 50040 41560 50080 41600
rect 64832 41560 64872 41600
rect 64914 41560 64954 41600
rect 64996 41560 65036 41600
rect 65078 41560 65118 41600
rect 65160 41560 65200 41600
rect 79952 41560 79992 41600
rect 80034 41560 80074 41600
rect 80116 41560 80156 41600
rect 80198 41560 80238 41600
rect 80280 41560 80320 41600
rect 95072 41560 95112 41600
rect 95154 41560 95194 41600
rect 95236 41560 95276 41600
rect 95318 41560 95358 41600
rect 95400 41560 95440 41600
rect 3112 40804 3152 40844
rect 3194 40804 3234 40844
rect 3276 40804 3316 40844
rect 3358 40804 3398 40844
rect 3440 40804 3480 40844
rect 18232 40804 18272 40844
rect 18314 40804 18354 40844
rect 18396 40804 18436 40844
rect 18478 40804 18518 40844
rect 18560 40804 18600 40844
rect 33352 40804 33392 40844
rect 33434 40804 33474 40844
rect 33516 40804 33556 40844
rect 33598 40804 33638 40844
rect 33680 40804 33720 40844
rect 48472 40804 48512 40844
rect 48554 40804 48594 40844
rect 48636 40804 48676 40844
rect 48718 40804 48758 40844
rect 48800 40804 48840 40844
rect 63592 40804 63632 40844
rect 63674 40804 63714 40844
rect 63756 40804 63796 40844
rect 63838 40804 63878 40844
rect 63920 40804 63960 40844
rect 78712 40804 78752 40844
rect 78794 40804 78834 40844
rect 78876 40804 78916 40844
rect 78958 40804 78998 40844
rect 79040 40804 79080 40844
rect 93832 40804 93872 40844
rect 93914 40804 93954 40844
rect 93996 40804 94036 40844
rect 94078 40804 94118 40844
rect 94160 40804 94200 40844
rect 4352 40048 4392 40088
rect 4434 40048 4474 40088
rect 4516 40048 4556 40088
rect 4598 40048 4638 40088
rect 4680 40048 4720 40088
rect 19472 40048 19512 40088
rect 19554 40048 19594 40088
rect 19636 40048 19676 40088
rect 19718 40048 19758 40088
rect 19800 40048 19840 40088
rect 34592 40048 34632 40088
rect 34674 40048 34714 40088
rect 34756 40048 34796 40088
rect 34838 40048 34878 40088
rect 34920 40048 34960 40088
rect 49712 40048 49752 40088
rect 49794 40048 49834 40088
rect 49876 40048 49916 40088
rect 49958 40048 49998 40088
rect 50040 40048 50080 40088
rect 64832 40048 64872 40088
rect 64914 40048 64954 40088
rect 64996 40048 65036 40088
rect 65078 40048 65118 40088
rect 65160 40048 65200 40088
rect 79952 40048 79992 40088
rect 80034 40048 80074 40088
rect 80116 40048 80156 40088
rect 80198 40048 80238 40088
rect 80280 40048 80320 40088
rect 95072 40048 95112 40088
rect 95154 40048 95194 40088
rect 95236 40048 95276 40088
rect 95318 40048 95358 40088
rect 95400 40048 95440 40088
rect 3112 39292 3152 39332
rect 3194 39292 3234 39332
rect 3276 39292 3316 39332
rect 3358 39292 3398 39332
rect 3440 39292 3480 39332
rect 18232 39292 18272 39332
rect 18314 39292 18354 39332
rect 18396 39292 18436 39332
rect 18478 39292 18518 39332
rect 18560 39292 18600 39332
rect 33352 39292 33392 39332
rect 33434 39292 33474 39332
rect 33516 39292 33556 39332
rect 33598 39292 33638 39332
rect 33680 39292 33720 39332
rect 48472 39292 48512 39332
rect 48554 39292 48594 39332
rect 48636 39292 48676 39332
rect 48718 39292 48758 39332
rect 48800 39292 48840 39332
rect 63592 39292 63632 39332
rect 63674 39292 63714 39332
rect 63756 39292 63796 39332
rect 63838 39292 63878 39332
rect 63920 39292 63960 39332
rect 78712 39292 78752 39332
rect 78794 39292 78834 39332
rect 78876 39292 78916 39332
rect 78958 39292 78998 39332
rect 79040 39292 79080 39332
rect 93832 39292 93872 39332
rect 93914 39292 93954 39332
rect 93996 39292 94036 39332
rect 94078 39292 94118 39332
rect 94160 39292 94200 39332
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 95072 38536 95112 38576
rect 95154 38536 95194 38576
rect 95236 38536 95276 38576
rect 95318 38536 95358 38576
rect 95400 38536 95440 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 93832 37780 93872 37820
rect 93914 37780 93954 37820
rect 93996 37780 94036 37820
rect 94078 37780 94118 37820
rect 94160 37780 94200 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 95072 37024 95112 37064
rect 95154 37024 95194 37064
rect 95236 37024 95276 37064
rect 95318 37024 95358 37064
rect 95400 37024 95440 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 93832 36268 93872 36308
rect 93914 36268 93954 36308
rect 93996 36268 94036 36308
rect 94078 36268 94118 36308
rect 94160 36268 94200 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 95072 35512 95112 35552
rect 95154 35512 95194 35552
rect 95236 35512 95276 35552
rect 95318 35512 95358 35552
rect 95400 35512 95440 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 93832 34756 93872 34796
rect 93914 34756 93954 34796
rect 93996 34756 94036 34796
rect 94078 34756 94118 34796
rect 94160 34756 94200 34796
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 95072 34000 95112 34040
rect 95154 34000 95194 34040
rect 95236 34000 95276 34040
rect 95318 34000 95358 34040
rect 95400 34000 95440 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 93832 33244 93872 33284
rect 93914 33244 93954 33284
rect 93996 33244 94036 33284
rect 94078 33244 94118 33284
rect 94160 33244 94200 33284
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 95072 32488 95112 32528
rect 95154 32488 95194 32528
rect 95236 32488 95276 32528
rect 95318 32488 95358 32528
rect 95400 32488 95440 32528
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 93832 31732 93872 31772
rect 93914 31732 93954 31772
rect 93996 31732 94036 31772
rect 94078 31732 94118 31772
rect 94160 31732 94200 31772
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 95072 30976 95112 31016
rect 95154 30976 95194 31016
rect 95236 30976 95276 31016
rect 95318 30976 95358 31016
rect 95400 30976 95440 31016
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 93832 30220 93872 30260
rect 93914 30220 93954 30260
rect 93996 30220 94036 30260
rect 94078 30220 94118 30260
rect 94160 30220 94200 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 95072 29464 95112 29504
rect 95154 29464 95194 29504
rect 95236 29464 95276 29504
rect 95318 29464 95358 29504
rect 95400 29464 95440 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 93832 28708 93872 28748
rect 93914 28708 93954 28748
rect 93996 28708 94036 28748
rect 94078 28708 94118 28748
rect 94160 28708 94200 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 95072 27952 95112 27992
rect 95154 27952 95194 27992
rect 95236 27952 95276 27992
rect 95318 27952 95358 27992
rect 95400 27952 95440 27992
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 93832 27196 93872 27236
rect 93914 27196 93954 27236
rect 93996 27196 94036 27236
rect 94078 27196 94118 27236
rect 94160 27196 94200 27236
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 95072 26440 95112 26480
rect 95154 26440 95194 26480
rect 95236 26440 95276 26480
rect 95318 26440 95358 26480
rect 95400 26440 95440 26480
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 93832 25684 93872 25724
rect 93914 25684 93954 25724
rect 93996 25684 94036 25724
rect 94078 25684 94118 25724
rect 94160 25684 94200 25724
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 95072 24928 95112 24968
rect 95154 24928 95194 24968
rect 95236 24928 95276 24968
rect 95318 24928 95358 24968
rect 95400 24928 95440 24968
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 63592 24172 63632 24212
rect 63674 24172 63714 24212
rect 63756 24172 63796 24212
rect 63838 24172 63878 24212
rect 63920 24172 63960 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 93832 24172 93872 24212
rect 93914 24172 93954 24212
rect 93996 24172 94036 24212
rect 94078 24172 94118 24212
rect 94160 24172 94200 24212
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 64832 23416 64872 23456
rect 64914 23416 64954 23456
rect 64996 23416 65036 23456
rect 65078 23416 65118 23456
rect 65160 23416 65200 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 95072 23416 95112 23456
rect 95154 23416 95194 23456
rect 95236 23416 95276 23456
rect 95318 23416 95358 23456
rect 95400 23416 95440 23456
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 63592 22660 63632 22700
rect 63674 22660 63714 22700
rect 63756 22660 63796 22700
rect 63838 22660 63878 22700
rect 63920 22660 63960 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 93832 22660 93872 22700
rect 93914 22660 93954 22700
rect 93996 22660 94036 22700
rect 94078 22660 94118 22700
rect 94160 22660 94200 22700
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 64832 21904 64872 21944
rect 64914 21904 64954 21944
rect 64996 21904 65036 21944
rect 65078 21904 65118 21944
rect 65160 21904 65200 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 63592 21148 63632 21188
rect 63674 21148 63714 21188
rect 63756 21148 63796 21188
rect 63838 21148 63878 21188
rect 63920 21148 63960 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 64832 20392 64872 20432
rect 64914 20392 64954 20432
rect 64996 20392 65036 20432
rect 65078 20392 65118 20432
rect 65160 20392 65200 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 63592 19636 63632 19676
rect 63674 19636 63714 19676
rect 63756 19636 63796 19676
rect 63838 19636 63878 19676
rect 63920 19636 63960 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 64832 18880 64872 18920
rect 64914 18880 64954 18920
rect 64996 18880 65036 18920
rect 65078 18880 65118 18920
rect 65160 18880 65200 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 95072 18880 95112 18920
rect 95154 18880 95194 18920
rect 95236 18880 95276 18920
rect 95318 18880 95358 18920
rect 95400 18880 95440 18920
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 63592 18124 63632 18164
rect 63674 18124 63714 18164
rect 63756 18124 63796 18164
rect 63838 18124 63878 18164
rect 63920 18124 63960 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 93832 18124 93872 18164
rect 93914 18124 93954 18164
rect 93996 18124 94036 18164
rect 94078 18124 94118 18164
rect 94160 18124 94200 18164
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 64832 17368 64872 17408
rect 64914 17368 64954 17408
rect 64996 17368 65036 17408
rect 65078 17368 65118 17408
rect 65160 17368 65200 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 95072 17368 95112 17408
rect 95154 17368 95194 17408
rect 95236 17368 95276 17408
rect 95318 17368 95358 17408
rect 95400 17368 95440 17408
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 63592 16612 63632 16652
rect 63674 16612 63714 16652
rect 63756 16612 63796 16652
rect 63838 16612 63878 16652
rect 63920 16612 63960 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 93832 16612 93872 16652
rect 93914 16612 93954 16652
rect 93996 16612 94036 16652
rect 94078 16612 94118 16652
rect 94160 16612 94200 16652
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 64832 15856 64872 15896
rect 64914 15856 64954 15896
rect 64996 15856 65036 15896
rect 65078 15856 65118 15896
rect 65160 15856 65200 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 95072 15856 95112 15896
rect 95154 15856 95194 15896
rect 95236 15856 95276 15896
rect 95318 15856 95358 15896
rect 95400 15856 95440 15896
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 93832 15100 93872 15140
rect 93914 15100 93954 15140
rect 93996 15100 94036 15140
rect 94078 15100 94118 15140
rect 94160 15100 94200 15140
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 95072 14344 95112 14384
rect 95154 14344 95194 14384
rect 95236 14344 95276 14384
rect 95318 14344 95358 14384
rect 95400 14344 95440 14384
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 93832 13588 93872 13628
rect 93914 13588 93954 13628
rect 93996 13588 94036 13628
rect 94078 13588 94118 13628
rect 94160 13588 94200 13628
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 95072 12832 95112 12872
rect 95154 12832 95194 12872
rect 95236 12832 95276 12872
rect 95318 12832 95358 12872
rect 95400 12832 95440 12872
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 93832 12076 93872 12116
rect 93914 12076 93954 12116
rect 93996 12076 94036 12116
rect 94078 12076 94118 12116
rect 94160 12076 94200 12116
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 95072 11320 95112 11360
rect 95154 11320 95194 11360
rect 95236 11320 95276 11360
rect 95318 11320 95358 11360
rect 95400 11320 95440 11360
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 93832 10564 93872 10604
rect 93914 10564 93954 10604
rect 93996 10564 94036 10604
rect 94078 10564 94118 10604
rect 94160 10564 94200 10604
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 95072 9808 95112 9848
rect 95154 9808 95194 9848
rect 95236 9808 95276 9848
rect 95318 9808 95358 9848
rect 95400 9808 95440 9848
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 93832 9052 93872 9092
rect 93914 9052 93954 9092
rect 93996 9052 94036 9092
rect 94078 9052 94118 9092
rect 94160 9052 94200 9092
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 95072 8296 95112 8336
rect 95154 8296 95194 8336
rect 95236 8296 95276 8336
rect 95318 8296 95358 8336
rect 95400 8296 95440 8336
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 93832 7540 93872 7580
rect 93914 7540 93954 7580
rect 93996 7540 94036 7580
rect 94078 7540 94118 7580
rect 94160 7540 94200 7580
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 95072 6784 95112 6824
rect 95154 6784 95194 6824
rect 95236 6784 95276 6824
rect 95318 6784 95358 6824
rect 95400 6784 95440 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 93832 6028 93872 6068
rect 93914 6028 93954 6068
rect 93996 6028 94036 6068
rect 94078 6028 94118 6068
rect 94160 6028 94200 6068
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 95072 5272 95112 5312
rect 95154 5272 95194 5312
rect 95236 5272 95276 5312
rect 95318 5272 95358 5312
rect 95400 5272 95440 5312
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 93832 4516 93872 4556
rect 93914 4516 93954 4556
rect 93996 4516 94036 4556
rect 94078 4516 94118 4556
rect 94160 4516 94200 4556
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 95072 3760 95112 3800
rect 95154 3760 95194 3800
rect 95236 3760 95276 3800
rect 95318 3760 95358 3800
rect 95400 3760 95440 3800
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 93832 3004 93872 3044
rect 93914 3004 93954 3044
rect 93996 3004 94036 3044
rect 94078 3004 94118 3044
rect 94160 3004 94200 3044
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 95072 2248 95112 2288
rect 95154 2248 95194 2288
rect 95236 2248 95276 2288
rect 95318 2248 95358 2288
rect 95400 2248 95440 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 93832 1492 93872 1532
rect 93914 1492 93954 1532
rect 93996 1492 94036 1532
rect 94078 1492 94118 1532
rect 94160 1492 94200 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
rect 95072 736 95112 776
rect 95154 736 95194 776
rect 95236 736 95276 776
rect 95318 736 95358 776
rect 95400 736 95440 776
<< metal5 >>
rect 3103 81691 3489 81710
rect 3103 81668 3169 81691
rect 3255 81668 3337 81691
rect 3423 81668 3489 81691
rect 3103 81628 3112 81668
rect 3152 81628 3169 81668
rect 3255 81628 3276 81668
rect 3316 81628 3337 81668
rect 3423 81628 3440 81668
rect 3480 81628 3489 81668
rect 3103 81605 3169 81628
rect 3255 81605 3337 81628
rect 3423 81605 3489 81628
rect 3103 81586 3489 81605
rect 18223 81691 18609 81710
rect 18223 81668 18289 81691
rect 18375 81668 18457 81691
rect 18543 81668 18609 81691
rect 18223 81628 18232 81668
rect 18272 81628 18289 81668
rect 18375 81628 18396 81668
rect 18436 81628 18457 81668
rect 18543 81628 18560 81668
rect 18600 81628 18609 81668
rect 18223 81605 18289 81628
rect 18375 81605 18457 81628
rect 18543 81605 18609 81628
rect 18223 81586 18609 81605
rect 33343 81691 33729 81710
rect 33343 81668 33409 81691
rect 33495 81668 33577 81691
rect 33663 81668 33729 81691
rect 33343 81628 33352 81668
rect 33392 81628 33409 81668
rect 33495 81628 33516 81668
rect 33556 81628 33577 81668
rect 33663 81628 33680 81668
rect 33720 81628 33729 81668
rect 33343 81605 33409 81628
rect 33495 81605 33577 81628
rect 33663 81605 33729 81628
rect 33343 81586 33729 81605
rect 48463 81691 48849 81710
rect 48463 81668 48529 81691
rect 48615 81668 48697 81691
rect 48783 81668 48849 81691
rect 48463 81628 48472 81668
rect 48512 81628 48529 81668
rect 48615 81628 48636 81668
rect 48676 81628 48697 81668
rect 48783 81628 48800 81668
rect 48840 81628 48849 81668
rect 48463 81605 48529 81628
rect 48615 81605 48697 81628
rect 48783 81605 48849 81628
rect 48463 81586 48849 81605
rect 63583 81691 63969 81710
rect 63583 81668 63649 81691
rect 63735 81668 63817 81691
rect 63903 81668 63969 81691
rect 63583 81628 63592 81668
rect 63632 81628 63649 81668
rect 63735 81628 63756 81668
rect 63796 81628 63817 81668
rect 63903 81628 63920 81668
rect 63960 81628 63969 81668
rect 63583 81605 63649 81628
rect 63735 81605 63817 81628
rect 63903 81605 63969 81628
rect 63583 81586 63969 81605
rect 78703 81691 79089 81710
rect 78703 81668 78769 81691
rect 78855 81668 78937 81691
rect 79023 81668 79089 81691
rect 78703 81628 78712 81668
rect 78752 81628 78769 81668
rect 78855 81628 78876 81668
rect 78916 81628 78937 81668
rect 79023 81628 79040 81668
rect 79080 81628 79089 81668
rect 78703 81605 78769 81628
rect 78855 81605 78937 81628
rect 79023 81605 79089 81628
rect 78703 81586 79089 81605
rect 93823 81691 94209 81710
rect 93823 81668 93889 81691
rect 93975 81668 94057 81691
rect 94143 81668 94209 81691
rect 93823 81628 93832 81668
rect 93872 81628 93889 81668
rect 93975 81628 93996 81668
rect 94036 81628 94057 81668
rect 94143 81628 94160 81668
rect 94200 81628 94209 81668
rect 93823 81605 93889 81628
rect 93975 81605 94057 81628
rect 94143 81605 94209 81628
rect 93823 81586 94209 81605
rect 4343 80935 4729 80954
rect 4343 80912 4409 80935
rect 4495 80912 4577 80935
rect 4663 80912 4729 80935
rect 4343 80872 4352 80912
rect 4392 80872 4409 80912
rect 4495 80872 4516 80912
rect 4556 80872 4577 80912
rect 4663 80872 4680 80912
rect 4720 80872 4729 80912
rect 4343 80849 4409 80872
rect 4495 80849 4577 80872
rect 4663 80849 4729 80872
rect 4343 80830 4729 80849
rect 19463 80935 19849 80954
rect 19463 80912 19529 80935
rect 19615 80912 19697 80935
rect 19783 80912 19849 80935
rect 19463 80872 19472 80912
rect 19512 80872 19529 80912
rect 19615 80872 19636 80912
rect 19676 80872 19697 80912
rect 19783 80872 19800 80912
rect 19840 80872 19849 80912
rect 19463 80849 19529 80872
rect 19615 80849 19697 80872
rect 19783 80849 19849 80872
rect 19463 80830 19849 80849
rect 34583 80935 34969 80954
rect 34583 80912 34649 80935
rect 34735 80912 34817 80935
rect 34903 80912 34969 80935
rect 34583 80872 34592 80912
rect 34632 80872 34649 80912
rect 34735 80872 34756 80912
rect 34796 80872 34817 80912
rect 34903 80872 34920 80912
rect 34960 80872 34969 80912
rect 34583 80849 34649 80872
rect 34735 80849 34817 80872
rect 34903 80849 34969 80872
rect 34583 80830 34969 80849
rect 49703 80935 50089 80954
rect 49703 80912 49769 80935
rect 49855 80912 49937 80935
rect 50023 80912 50089 80935
rect 49703 80872 49712 80912
rect 49752 80872 49769 80912
rect 49855 80872 49876 80912
rect 49916 80872 49937 80912
rect 50023 80872 50040 80912
rect 50080 80872 50089 80912
rect 49703 80849 49769 80872
rect 49855 80849 49937 80872
rect 50023 80849 50089 80872
rect 49703 80830 50089 80849
rect 64823 80935 65209 80954
rect 64823 80912 64889 80935
rect 64975 80912 65057 80935
rect 65143 80912 65209 80935
rect 64823 80872 64832 80912
rect 64872 80872 64889 80912
rect 64975 80872 64996 80912
rect 65036 80872 65057 80912
rect 65143 80872 65160 80912
rect 65200 80872 65209 80912
rect 64823 80849 64889 80872
rect 64975 80849 65057 80872
rect 65143 80849 65209 80872
rect 64823 80830 65209 80849
rect 79943 80935 80329 80954
rect 79943 80912 80009 80935
rect 80095 80912 80177 80935
rect 80263 80912 80329 80935
rect 79943 80872 79952 80912
rect 79992 80872 80009 80912
rect 80095 80872 80116 80912
rect 80156 80872 80177 80912
rect 80263 80872 80280 80912
rect 80320 80872 80329 80912
rect 79943 80849 80009 80872
rect 80095 80849 80177 80872
rect 80263 80849 80329 80872
rect 79943 80830 80329 80849
rect 95063 80935 95449 80954
rect 95063 80912 95129 80935
rect 95215 80912 95297 80935
rect 95383 80912 95449 80935
rect 95063 80872 95072 80912
rect 95112 80872 95129 80912
rect 95215 80872 95236 80912
rect 95276 80872 95297 80912
rect 95383 80872 95400 80912
rect 95440 80872 95449 80912
rect 95063 80849 95129 80872
rect 95215 80849 95297 80872
rect 95383 80849 95449 80872
rect 95063 80830 95449 80849
rect 3103 80179 3489 80198
rect 3103 80156 3169 80179
rect 3255 80156 3337 80179
rect 3423 80156 3489 80179
rect 3103 80116 3112 80156
rect 3152 80116 3169 80156
rect 3255 80116 3276 80156
rect 3316 80116 3337 80156
rect 3423 80116 3440 80156
rect 3480 80116 3489 80156
rect 3103 80093 3169 80116
rect 3255 80093 3337 80116
rect 3423 80093 3489 80116
rect 3103 80074 3489 80093
rect 18223 80179 18609 80198
rect 18223 80156 18289 80179
rect 18375 80156 18457 80179
rect 18543 80156 18609 80179
rect 18223 80116 18232 80156
rect 18272 80116 18289 80156
rect 18375 80116 18396 80156
rect 18436 80116 18457 80156
rect 18543 80116 18560 80156
rect 18600 80116 18609 80156
rect 18223 80093 18289 80116
rect 18375 80093 18457 80116
rect 18543 80093 18609 80116
rect 18223 80074 18609 80093
rect 33343 80179 33729 80198
rect 33343 80156 33409 80179
rect 33495 80156 33577 80179
rect 33663 80156 33729 80179
rect 33343 80116 33352 80156
rect 33392 80116 33409 80156
rect 33495 80116 33516 80156
rect 33556 80116 33577 80156
rect 33663 80116 33680 80156
rect 33720 80116 33729 80156
rect 33343 80093 33409 80116
rect 33495 80093 33577 80116
rect 33663 80093 33729 80116
rect 33343 80074 33729 80093
rect 48463 80179 48849 80198
rect 48463 80156 48529 80179
rect 48615 80156 48697 80179
rect 48783 80156 48849 80179
rect 48463 80116 48472 80156
rect 48512 80116 48529 80156
rect 48615 80116 48636 80156
rect 48676 80116 48697 80156
rect 48783 80116 48800 80156
rect 48840 80116 48849 80156
rect 48463 80093 48529 80116
rect 48615 80093 48697 80116
rect 48783 80093 48849 80116
rect 48463 80074 48849 80093
rect 63583 80179 63969 80198
rect 63583 80156 63649 80179
rect 63735 80156 63817 80179
rect 63903 80156 63969 80179
rect 63583 80116 63592 80156
rect 63632 80116 63649 80156
rect 63735 80116 63756 80156
rect 63796 80116 63817 80156
rect 63903 80116 63920 80156
rect 63960 80116 63969 80156
rect 63583 80093 63649 80116
rect 63735 80093 63817 80116
rect 63903 80093 63969 80116
rect 63583 80074 63969 80093
rect 78703 80179 79089 80198
rect 78703 80156 78769 80179
rect 78855 80156 78937 80179
rect 79023 80156 79089 80179
rect 78703 80116 78712 80156
rect 78752 80116 78769 80156
rect 78855 80116 78876 80156
rect 78916 80116 78937 80156
rect 79023 80116 79040 80156
rect 79080 80116 79089 80156
rect 78703 80093 78769 80116
rect 78855 80093 78937 80116
rect 79023 80093 79089 80116
rect 78703 80074 79089 80093
rect 93823 80179 94209 80198
rect 93823 80156 93889 80179
rect 93975 80156 94057 80179
rect 94143 80156 94209 80179
rect 93823 80116 93832 80156
rect 93872 80116 93889 80156
rect 93975 80116 93996 80156
rect 94036 80116 94057 80156
rect 94143 80116 94160 80156
rect 94200 80116 94209 80156
rect 93823 80093 93889 80116
rect 93975 80093 94057 80116
rect 94143 80093 94209 80116
rect 93823 80074 94209 80093
rect 4343 79423 4729 79442
rect 4343 79400 4409 79423
rect 4495 79400 4577 79423
rect 4663 79400 4729 79423
rect 4343 79360 4352 79400
rect 4392 79360 4409 79400
rect 4495 79360 4516 79400
rect 4556 79360 4577 79400
rect 4663 79360 4680 79400
rect 4720 79360 4729 79400
rect 4343 79337 4409 79360
rect 4495 79337 4577 79360
rect 4663 79337 4729 79360
rect 4343 79318 4729 79337
rect 19463 79423 19849 79442
rect 19463 79400 19529 79423
rect 19615 79400 19697 79423
rect 19783 79400 19849 79423
rect 19463 79360 19472 79400
rect 19512 79360 19529 79400
rect 19615 79360 19636 79400
rect 19676 79360 19697 79400
rect 19783 79360 19800 79400
rect 19840 79360 19849 79400
rect 19463 79337 19529 79360
rect 19615 79337 19697 79360
rect 19783 79337 19849 79360
rect 19463 79318 19849 79337
rect 34583 79423 34969 79442
rect 34583 79400 34649 79423
rect 34735 79400 34817 79423
rect 34903 79400 34969 79423
rect 34583 79360 34592 79400
rect 34632 79360 34649 79400
rect 34735 79360 34756 79400
rect 34796 79360 34817 79400
rect 34903 79360 34920 79400
rect 34960 79360 34969 79400
rect 34583 79337 34649 79360
rect 34735 79337 34817 79360
rect 34903 79337 34969 79360
rect 34583 79318 34969 79337
rect 49703 79423 50089 79442
rect 49703 79400 49769 79423
rect 49855 79400 49937 79423
rect 50023 79400 50089 79423
rect 49703 79360 49712 79400
rect 49752 79360 49769 79400
rect 49855 79360 49876 79400
rect 49916 79360 49937 79400
rect 50023 79360 50040 79400
rect 50080 79360 50089 79400
rect 49703 79337 49769 79360
rect 49855 79337 49937 79360
rect 50023 79337 50089 79360
rect 49703 79318 50089 79337
rect 64823 79423 65209 79442
rect 64823 79400 64889 79423
rect 64975 79400 65057 79423
rect 65143 79400 65209 79423
rect 64823 79360 64832 79400
rect 64872 79360 64889 79400
rect 64975 79360 64996 79400
rect 65036 79360 65057 79400
rect 65143 79360 65160 79400
rect 65200 79360 65209 79400
rect 64823 79337 64889 79360
rect 64975 79337 65057 79360
rect 65143 79337 65209 79360
rect 64823 79318 65209 79337
rect 79943 79423 80329 79442
rect 79943 79400 80009 79423
rect 80095 79400 80177 79423
rect 80263 79400 80329 79423
rect 79943 79360 79952 79400
rect 79992 79360 80009 79400
rect 80095 79360 80116 79400
rect 80156 79360 80177 79400
rect 80263 79360 80280 79400
rect 80320 79360 80329 79400
rect 79943 79337 80009 79360
rect 80095 79337 80177 79360
rect 80263 79337 80329 79360
rect 79943 79318 80329 79337
rect 95063 79423 95449 79442
rect 95063 79400 95129 79423
rect 95215 79400 95297 79423
rect 95383 79400 95449 79423
rect 95063 79360 95072 79400
rect 95112 79360 95129 79400
rect 95215 79360 95236 79400
rect 95276 79360 95297 79400
rect 95383 79360 95400 79400
rect 95440 79360 95449 79400
rect 95063 79337 95129 79360
rect 95215 79337 95297 79360
rect 95383 79337 95449 79360
rect 95063 79318 95449 79337
rect 3103 78667 3489 78686
rect 3103 78644 3169 78667
rect 3255 78644 3337 78667
rect 3423 78644 3489 78667
rect 3103 78604 3112 78644
rect 3152 78604 3169 78644
rect 3255 78604 3276 78644
rect 3316 78604 3337 78644
rect 3423 78604 3440 78644
rect 3480 78604 3489 78644
rect 3103 78581 3169 78604
rect 3255 78581 3337 78604
rect 3423 78581 3489 78604
rect 3103 78562 3489 78581
rect 18223 78667 18609 78686
rect 18223 78644 18289 78667
rect 18375 78644 18457 78667
rect 18543 78644 18609 78667
rect 18223 78604 18232 78644
rect 18272 78604 18289 78644
rect 18375 78604 18396 78644
rect 18436 78604 18457 78644
rect 18543 78604 18560 78644
rect 18600 78604 18609 78644
rect 18223 78581 18289 78604
rect 18375 78581 18457 78604
rect 18543 78581 18609 78604
rect 18223 78562 18609 78581
rect 33343 78667 33729 78686
rect 33343 78644 33409 78667
rect 33495 78644 33577 78667
rect 33663 78644 33729 78667
rect 33343 78604 33352 78644
rect 33392 78604 33409 78644
rect 33495 78604 33516 78644
rect 33556 78604 33577 78644
rect 33663 78604 33680 78644
rect 33720 78604 33729 78644
rect 33343 78581 33409 78604
rect 33495 78581 33577 78604
rect 33663 78581 33729 78604
rect 33343 78562 33729 78581
rect 48463 78667 48849 78686
rect 48463 78644 48529 78667
rect 48615 78644 48697 78667
rect 48783 78644 48849 78667
rect 48463 78604 48472 78644
rect 48512 78604 48529 78644
rect 48615 78604 48636 78644
rect 48676 78604 48697 78644
rect 48783 78604 48800 78644
rect 48840 78604 48849 78644
rect 48463 78581 48529 78604
rect 48615 78581 48697 78604
rect 48783 78581 48849 78604
rect 48463 78562 48849 78581
rect 63583 78667 63969 78686
rect 63583 78644 63649 78667
rect 63735 78644 63817 78667
rect 63903 78644 63969 78667
rect 63583 78604 63592 78644
rect 63632 78604 63649 78644
rect 63735 78604 63756 78644
rect 63796 78604 63817 78644
rect 63903 78604 63920 78644
rect 63960 78604 63969 78644
rect 63583 78581 63649 78604
rect 63735 78581 63817 78604
rect 63903 78581 63969 78604
rect 63583 78562 63969 78581
rect 78703 78667 79089 78686
rect 78703 78644 78769 78667
rect 78855 78644 78937 78667
rect 79023 78644 79089 78667
rect 78703 78604 78712 78644
rect 78752 78604 78769 78644
rect 78855 78604 78876 78644
rect 78916 78604 78937 78644
rect 79023 78604 79040 78644
rect 79080 78604 79089 78644
rect 78703 78581 78769 78604
rect 78855 78581 78937 78604
rect 79023 78581 79089 78604
rect 78703 78562 79089 78581
rect 93823 78667 94209 78686
rect 93823 78644 93889 78667
rect 93975 78644 94057 78667
rect 94143 78644 94209 78667
rect 93823 78604 93832 78644
rect 93872 78604 93889 78644
rect 93975 78604 93996 78644
rect 94036 78604 94057 78644
rect 94143 78604 94160 78644
rect 94200 78604 94209 78644
rect 93823 78581 93889 78604
rect 93975 78581 94057 78604
rect 94143 78581 94209 78604
rect 93823 78562 94209 78581
rect 4343 77911 4729 77930
rect 4343 77888 4409 77911
rect 4495 77888 4577 77911
rect 4663 77888 4729 77911
rect 4343 77848 4352 77888
rect 4392 77848 4409 77888
rect 4495 77848 4516 77888
rect 4556 77848 4577 77888
rect 4663 77848 4680 77888
rect 4720 77848 4729 77888
rect 4343 77825 4409 77848
rect 4495 77825 4577 77848
rect 4663 77825 4729 77848
rect 4343 77806 4729 77825
rect 19463 77911 19849 77930
rect 19463 77888 19529 77911
rect 19615 77888 19697 77911
rect 19783 77888 19849 77911
rect 19463 77848 19472 77888
rect 19512 77848 19529 77888
rect 19615 77848 19636 77888
rect 19676 77848 19697 77888
rect 19783 77848 19800 77888
rect 19840 77848 19849 77888
rect 19463 77825 19529 77848
rect 19615 77825 19697 77848
rect 19783 77825 19849 77848
rect 19463 77806 19849 77825
rect 34583 77911 34969 77930
rect 34583 77888 34649 77911
rect 34735 77888 34817 77911
rect 34903 77888 34969 77911
rect 34583 77848 34592 77888
rect 34632 77848 34649 77888
rect 34735 77848 34756 77888
rect 34796 77848 34817 77888
rect 34903 77848 34920 77888
rect 34960 77848 34969 77888
rect 34583 77825 34649 77848
rect 34735 77825 34817 77848
rect 34903 77825 34969 77848
rect 34583 77806 34969 77825
rect 49703 77911 50089 77930
rect 49703 77888 49769 77911
rect 49855 77888 49937 77911
rect 50023 77888 50089 77911
rect 49703 77848 49712 77888
rect 49752 77848 49769 77888
rect 49855 77848 49876 77888
rect 49916 77848 49937 77888
rect 50023 77848 50040 77888
rect 50080 77848 50089 77888
rect 49703 77825 49769 77848
rect 49855 77825 49937 77848
rect 50023 77825 50089 77848
rect 49703 77806 50089 77825
rect 64823 77911 65209 77930
rect 64823 77888 64889 77911
rect 64975 77888 65057 77911
rect 65143 77888 65209 77911
rect 64823 77848 64832 77888
rect 64872 77848 64889 77888
rect 64975 77848 64996 77888
rect 65036 77848 65057 77888
rect 65143 77848 65160 77888
rect 65200 77848 65209 77888
rect 64823 77825 64889 77848
rect 64975 77825 65057 77848
rect 65143 77825 65209 77848
rect 64823 77806 65209 77825
rect 79943 77911 80329 77930
rect 79943 77888 80009 77911
rect 80095 77888 80177 77911
rect 80263 77888 80329 77911
rect 79943 77848 79952 77888
rect 79992 77848 80009 77888
rect 80095 77848 80116 77888
rect 80156 77848 80177 77888
rect 80263 77848 80280 77888
rect 80320 77848 80329 77888
rect 79943 77825 80009 77848
rect 80095 77825 80177 77848
rect 80263 77825 80329 77848
rect 79943 77806 80329 77825
rect 95063 77911 95449 77930
rect 95063 77888 95129 77911
rect 95215 77888 95297 77911
rect 95383 77888 95449 77911
rect 95063 77848 95072 77888
rect 95112 77848 95129 77888
rect 95215 77848 95236 77888
rect 95276 77848 95297 77888
rect 95383 77848 95400 77888
rect 95440 77848 95449 77888
rect 95063 77825 95129 77848
rect 95215 77825 95297 77848
rect 95383 77825 95449 77848
rect 95063 77806 95449 77825
rect 3103 77155 3489 77174
rect 3103 77132 3169 77155
rect 3255 77132 3337 77155
rect 3423 77132 3489 77155
rect 3103 77092 3112 77132
rect 3152 77092 3169 77132
rect 3255 77092 3276 77132
rect 3316 77092 3337 77132
rect 3423 77092 3440 77132
rect 3480 77092 3489 77132
rect 3103 77069 3169 77092
rect 3255 77069 3337 77092
rect 3423 77069 3489 77092
rect 3103 77050 3489 77069
rect 18223 77155 18609 77174
rect 18223 77132 18289 77155
rect 18375 77132 18457 77155
rect 18543 77132 18609 77155
rect 18223 77092 18232 77132
rect 18272 77092 18289 77132
rect 18375 77092 18396 77132
rect 18436 77092 18457 77132
rect 18543 77092 18560 77132
rect 18600 77092 18609 77132
rect 18223 77069 18289 77092
rect 18375 77069 18457 77092
rect 18543 77069 18609 77092
rect 18223 77050 18609 77069
rect 33343 77155 33729 77174
rect 33343 77132 33409 77155
rect 33495 77132 33577 77155
rect 33663 77132 33729 77155
rect 33343 77092 33352 77132
rect 33392 77092 33409 77132
rect 33495 77092 33516 77132
rect 33556 77092 33577 77132
rect 33663 77092 33680 77132
rect 33720 77092 33729 77132
rect 33343 77069 33409 77092
rect 33495 77069 33577 77092
rect 33663 77069 33729 77092
rect 33343 77050 33729 77069
rect 48463 77155 48849 77174
rect 48463 77132 48529 77155
rect 48615 77132 48697 77155
rect 48783 77132 48849 77155
rect 48463 77092 48472 77132
rect 48512 77092 48529 77132
rect 48615 77092 48636 77132
rect 48676 77092 48697 77132
rect 48783 77092 48800 77132
rect 48840 77092 48849 77132
rect 48463 77069 48529 77092
rect 48615 77069 48697 77092
rect 48783 77069 48849 77092
rect 48463 77050 48849 77069
rect 63583 77155 63969 77174
rect 63583 77132 63649 77155
rect 63735 77132 63817 77155
rect 63903 77132 63969 77155
rect 63583 77092 63592 77132
rect 63632 77092 63649 77132
rect 63735 77092 63756 77132
rect 63796 77092 63817 77132
rect 63903 77092 63920 77132
rect 63960 77092 63969 77132
rect 63583 77069 63649 77092
rect 63735 77069 63817 77092
rect 63903 77069 63969 77092
rect 63583 77050 63969 77069
rect 78703 77155 79089 77174
rect 78703 77132 78769 77155
rect 78855 77132 78937 77155
rect 79023 77132 79089 77155
rect 78703 77092 78712 77132
rect 78752 77092 78769 77132
rect 78855 77092 78876 77132
rect 78916 77092 78937 77132
rect 79023 77092 79040 77132
rect 79080 77092 79089 77132
rect 78703 77069 78769 77092
rect 78855 77069 78937 77092
rect 79023 77069 79089 77092
rect 78703 77050 79089 77069
rect 93823 77155 94209 77174
rect 93823 77132 93889 77155
rect 93975 77132 94057 77155
rect 94143 77132 94209 77155
rect 93823 77092 93832 77132
rect 93872 77092 93889 77132
rect 93975 77092 93996 77132
rect 94036 77092 94057 77132
rect 94143 77092 94160 77132
rect 94200 77092 94209 77132
rect 93823 77069 93889 77092
rect 93975 77069 94057 77092
rect 94143 77069 94209 77092
rect 93823 77050 94209 77069
rect 4343 76399 4729 76418
rect 4343 76376 4409 76399
rect 4495 76376 4577 76399
rect 4663 76376 4729 76399
rect 4343 76336 4352 76376
rect 4392 76336 4409 76376
rect 4495 76336 4516 76376
rect 4556 76336 4577 76376
rect 4663 76336 4680 76376
rect 4720 76336 4729 76376
rect 4343 76313 4409 76336
rect 4495 76313 4577 76336
rect 4663 76313 4729 76336
rect 4343 76294 4729 76313
rect 19463 76399 19849 76418
rect 19463 76376 19529 76399
rect 19615 76376 19697 76399
rect 19783 76376 19849 76399
rect 19463 76336 19472 76376
rect 19512 76336 19529 76376
rect 19615 76336 19636 76376
rect 19676 76336 19697 76376
rect 19783 76336 19800 76376
rect 19840 76336 19849 76376
rect 19463 76313 19529 76336
rect 19615 76313 19697 76336
rect 19783 76313 19849 76336
rect 19463 76294 19849 76313
rect 34583 76399 34969 76418
rect 34583 76376 34649 76399
rect 34735 76376 34817 76399
rect 34903 76376 34969 76399
rect 34583 76336 34592 76376
rect 34632 76336 34649 76376
rect 34735 76336 34756 76376
rect 34796 76336 34817 76376
rect 34903 76336 34920 76376
rect 34960 76336 34969 76376
rect 34583 76313 34649 76336
rect 34735 76313 34817 76336
rect 34903 76313 34969 76336
rect 34583 76294 34969 76313
rect 49703 76399 50089 76418
rect 49703 76376 49769 76399
rect 49855 76376 49937 76399
rect 50023 76376 50089 76399
rect 49703 76336 49712 76376
rect 49752 76336 49769 76376
rect 49855 76336 49876 76376
rect 49916 76336 49937 76376
rect 50023 76336 50040 76376
rect 50080 76336 50089 76376
rect 49703 76313 49769 76336
rect 49855 76313 49937 76336
rect 50023 76313 50089 76336
rect 49703 76294 50089 76313
rect 64823 76399 65209 76418
rect 64823 76376 64889 76399
rect 64975 76376 65057 76399
rect 65143 76376 65209 76399
rect 64823 76336 64832 76376
rect 64872 76336 64889 76376
rect 64975 76336 64996 76376
rect 65036 76336 65057 76376
rect 65143 76336 65160 76376
rect 65200 76336 65209 76376
rect 64823 76313 64889 76336
rect 64975 76313 65057 76336
rect 65143 76313 65209 76336
rect 64823 76294 65209 76313
rect 79943 76399 80329 76418
rect 79943 76376 80009 76399
rect 80095 76376 80177 76399
rect 80263 76376 80329 76399
rect 79943 76336 79952 76376
rect 79992 76336 80009 76376
rect 80095 76336 80116 76376
rect 80156 76336 80177 76376
rect 80263 76336 80280 76376
rect 80320 76336 80329 76376
rect 79943 76313 80009 76336
rect 80095 76313 80177 76336
rect 80263 76313 80329 76336
rect 79943 76294 80329 76313
rect 95063 76399 95449 76418
rect 95063 76376 95129 76399
rect 95215 76376 95297 76399
rect 95383 76376 95449 76399
rect 95063 76336 95072 76376
rect 95112 76336 95129 76376
rect 95215 76336 95236 76376
rect 95276 76336 95297 76376
rect 95383 76336 95400 76376
rect 95440 76336 95449 76376
rect 95063 76313 95129 76336
rect 95215 76313 95297 76336
rect 95383 76313 95449 76336
rect 95063 76294 95449 76313
rect 3103 75643 3489 75662
rect 3103 75620 3169 75643
rect 3255 75620 3337 75643
rect 3423 75620 3489 75643
rect 3103 75580 3112 75620
rect 3152 75580 3169 75620
rect 3255 75580 3276 75620
rect 3316 75580 3337 75620
rect 3423 75580 3440 75620
rect 3480 75580 3489 75620
rect 3103 75557 3169 75580
rect 3255 75557 3337 75580
rect 3423 75557 3489 75580
rect 3103 75538 3489 75557
rect 18223 75643 18609 75662
rect 18223 75620 18289 75643
rect 18375 75620 18457 75643
rect 18543 75620 18609 75643
rect 18223 75580 18232 75620
rect 18272 75580 18289 75620
rect 18375 75580 18396 75620
rect 18436 75580 18457 75620
rect 18543 75580 18560 75620
rect 18600 75580 18609 75620
rect 18223 75557 18289 75580
rect 18375 75557 18457 75580
rect 18543 75557 18609 75580
rect 18223 75538 18609 75557
rect 33343 75643 33729 75662
rect 33343 75620 33409 75643
rect 33495 75620 33577 75643
rect 33663 75620 33729 75643
rect 33343 75580 33352 75620
rect 33392 75580 33409 75620
rect 33495 75580 33516 75620
rect 33556 75580 33577 75620
rect 33663 75580 33680 75620
rect 33720 75580 33729 75620
rect 33343 75557 33409 75580
rect 33495 75557 33577 75580
rect 33663 75557 33729 75580
rect 33343 75538 33729 75557
rect 48463 75643 48849 75662
rect 48463 75620 48529 75643
rect 48615 75620 48697 75643
rect 48783 75620 48849 75643
rect 48463 75580 48472 75620
rect 48512 75580 48529 75620
rect 48615 75580 48636 75620
rect 48676 75580 48697 75620
rect 48783 75580 48800 75620
rect 48840 75580 48849 75620
rect 48463 75557 48529 75580
rect 48615 75557 48697 75580
rect 48783 75557 48849 75580
rect 48463 75538 48849 75557
rect 63583 75643 63969 75662
rect 63583 75620 63649 75643
rect 63735 75620 63817 75643
rect 63903 75620 63969 75643
rect 63583 75580 63592 75620
rect 63632 75580 63649 75620
rect 63735 75580 63756 75620
rect 63796 75580 63817 75620
rect 63903 75580 63920 75620
rect 63960 75580 63969 75620
rect 63583 75557 63649 75580
rect 63735 75557 63817 75580
rect 63903 75557 63969 75580
rect 63583 75538 63969 75557
rect 78703 75643 79089 75662
rect 78703 75620 78769 75643
rect 78855 75620 78937 75643
rect 79023 75620 79089 75643
rect 78703 75580 78712 75620
rect 78752 75580 78769 75620
rect 78855 75580 78876 75620
rect 78916 75580 78937 75620
rect 79023 75580 79040 75620
rect 79080 75580 79089 75620
rect 78703 75557 78769 75580
rect 78855 75557 78937 75580
rect 79023 75557 79089 75580
rect 78703 75538 79089 75557
rect 93823 75643 94209 75662
rect 93823 75620 93889 75643
rect 93975 75620 94057 75643
rect 94143 75620 94209 75643
rect 93823 75580 93832 75620
rect 93872 75580 93889 75620
rect 93975 75580 93996 75620
rect 94036 75580 94057 75620
rect 94143 75580 94160 75620
rect 94200 75580 94209 75620
rect 93823 75557 93889 75580
rect 93975 75557 94057 75580
rect 94143 75557 94209 75580
rect 93823 75538 94209 75557
rect 4343 74887 4729 74906
rect 4343 74864 4409 74887
rect 4495 74864 4577 74887
rect 4663 74864 4729 74887
rect 4343 74824 4352 74864
rect 4392 74824 4409 74864
rect 4495 74824 4516 74864
rect 4556 74824 4577 74864
rect 4663 74824 4680 74864
rect 4720 74824 4729 74864
rect 4343 74801 4409 74824
rect 4495 74801 4577 74824
rect 4663 74801 4729 74824
rect 4343 74782 4729 74801
rect 19463 74887 19849 74906
rect 19463 74864 19529 74887
rect 19615 74864 19697 74887
rect 19783 74864 19849 74887
rect 19463 74824 19472 74864
rect 19512 74824 19529 74864
rect 19615 74824 19636 74864
rect 19676 74824 19697 74864
rect 19783 74824 19800 74864
rect 19840 74824 19849 74864
rect 19463 74801 19529 74824
rect 19615 74801 19697 74824
rect 19783 74801 19849 74824
rect 19463 74782 19849 74801
rect 34583 74887 34969 74906
rect 34583 74864 34649 74887
rect 34735 74864 34817 74887
rect 34903 74864 34969 74887
rect 34583 74824 34592 74864
rect 34632 74824 34649 74864
rect 34735 74824 34756 74864
rect 34796 74824 34817 74864
rect 34903 74824 34920 74864
rect 34960 74824 34969 74864
rect 34583 74801 34649 74824
rect 34735 74801 34817 74824
rect 34903 74801 34969 74824
rect 34583 74782 34969 74801
rect 49703 74887 50089 74906
rect 49703 74864 49769 74887
rect 49855 74864 49937 74887
rect 50023 74864 50089 74887
rect 49703 74824 49712 74864
rect 49752 74824 49769 74864
rect 49855 74824 49876 74864
rect 49916 74824 49937 74864
rect 50023 74824 50040 74864
rect 50080 74824 50089 74864
rect 49703 74801 49769 74824
rect 49855 74801 49937 74824
rect 50023 74801 50089 74824
rect 49703 74782 50089 74801
rect 64823 74887 65209 74906
rect 64823 74864 64889 74887
rect 64975 74864 65057 74887
rect 65143 74864 65209 74887
rect 64823 74824 64832 74864
rect 64872 74824 64889 74864
rect 64975 74824 64996 74864
rect 65036 74824 65057 74864
rect 65143 74824 65160 74864
rect 65200 74824 65209 74864
rect 64823 74801 64889 74824
rect 64975 74801 65057 74824
rect 65143 74801 65209 74824
rect 64823 74782 65209 74801
rect 79943 74887 80329 74906
rect 79943 74864 80009 74887
rect 80095 74864 80177 74887
rect 80263 74864 80329 74887
rect 79943 74824 79952 74864
rect 79992 74824 80009 74864
rect 80095 74824 80116 74864
rect 80156 74824 80177 74864
rect 80263 74824 80280 74864
rect 80320 74824 80329 74864
rect 79943 74801 80009 74824
rect 80095 74801 80177 74824
rect 80263 74801 80329 74824
rect 79943 74782 80329 74801
rect 95063 74887 95449 74906
rect 95063 74864 95129 74887
rect 95215 74864 95297 74887
rect 95383 74864 95449 74887
rect 95063 74824 95072 74864
rect 95112 74824 95129 74864
rect 95215 74824 95236 74864
rect 95276 74824 95297 74864
rect 95383 74824 95400 74864
rect 95440 74824 95449 74864
rect 95063 74801 95129 74824
rect 95215 74801 95297 74824
rect 95383 74801 95449 74824
rect 95063 74782 95449 74801
rect 3103 74131 3489 74150
rect 3103 74108 3169 74131
rect 3255 74108 3337 74131
rect 3423 74108 3489 74131
rect 3103 74068 3112 74108
rect 3152 74068 3169 74108
rect 3255 74068 3276 74108
rect 3316 74068 3337 74108
rect 3423 74068 3440 74108
rect 3480 74068 3489 74108
rect 3103 74045 3169 74068
rect 3255 74045 3337 74068
rect 3423 74045 3489 74068
rect 3103 74026 3489 74045
rect 18223 74131 18609 74150
rect 18223 74108 18289 74131
rect 18375 74108 18457 74131
rect 18543 74108 18609 74131
rect 18223 74068 18232 74108
rect 18272 74068 18289 74108
rect 18375 74068 18396 74108
rect 18436 74068 18457 74108
rect 18543 74068 18560 74108
rect 18600 74068 18609 74108
rect 18223 74045 18289 74068
rect 18375 74045 18457 74068
rect 18543 74045 18609 74068
rect 18223 74026 18609 74045
rect 33343 74131 33729 74150
rect 33343 74108 33409 74131
rect 33495 74108 33577 74131
rect 33663 74108 33729 74131
rect 33343 74068 33352 74108
rect 33392 74068 33409 74108
rect 33495 74068 33516 74108
rect 33556 74068 33577 74108
rect 33663 74068 33680 74108
rect 33720 74068 33729 74108
rect 33343 74045 33409 74068
rect 33495 74045 33577 74068
rect 33663 74045 33729 74068
rect 33343 74026 33729 74045
rect 48463 74131 48849 74150
rect 48463 74108 48529 74131
rect 48615 74108 48697 74131
rect 48783 74108 48849 74131
rect 48463 74068 48472 74108
rect 48512 74068 48529 74108
rect 48615 74068 48636 74108
rect 48676 74068 48697 74108
rect 48783 74068 48800 74108
rect 48840 74068 48849 74108
rect 48463 74045 48529 74068
rect 48615 74045 48697 74068
rect 48783 74045 48849 74068
rect 48463 74026 48849 74045
rect 63583 74131 63969 74150
rect 63583 74108 63649 74131
rect 63735 74108 63817 74131
rect 63903 74108 63969 74131
rect 63583 74068 63592 74108
rect 63632 74068 63649 74108
rect 63735 74068 63756 74108
rect 63796 74068 63817 74108
rect 63903 74068 63920 74108
rect 63960 74068 63969 74108
rect 63583 74045 63649 74068
rect 63735 74045 63817 74068
rect 63903 74045 63969 74068
rect 63583 74026 63969 74045
rect 78703 74131 79089 74150
rect 78703 74108 78769 74131
rect 78855 74108 78937 74131
rect 79023 74108 79089 74131
rect 78703 74068 78712 74108
rect 78752 74068 78769 74108
rect 78855 74068 78876 74108
rect 78916 74068 78937 74108
rect 79023 74068 79040 74108
rect 79080 74068 79089 74108
rect 78703 74045 78769 74068
rect 78855 74045 78937 74068
rect 79023 74045 79089 74068
rect 78703 74026 79089 74045
rect 93823 74131 94209 74150
rect 93823 74108 93889 74131
rect 93975 74108 94057 74131
rect 94143 74108 94209 74131
rect 93823 74068 93832 74108
rect 93872 74068 93889 74108
rect 93975 74068 93996 74108
rect 94036 74068 94057 74108
rect 94143 74068 94160 74108
rect 94200 74068 94209 74108
rect 93823 74045 93889 74068
rect 93975 74045 94057 74068
rect 94143 74045 94209 74068
rect 93823 74026 94209 74045
rect 4343 73375 4729 73394
rect 4343 73352 4409 73375
rect 4495 73352 4577 73375
rect 4663 73352 4729 73375
rect 4343 73312 4352 73352
rect 4392 73312 4409 73352
rect 4495 73312 4516 73352
rect 4556 73312 4577 73352
rect 4663 73312 4680 73352
rect 4720 73312 4729 73352
rect 4343 73289 4409 73312
rect 4495 73289 4577 73312
rect 4663 73289 4729 73312
rect 4343 73270 4729 73289
rect 19463 73375 19849 73394
rect 19463 73352 19529 73375
rect 19615 73352 19697 73375
rect 19783 73352 19849 73375
rect 19463 73312 19472 73352
rect 19512 73312 19529 73352
rect 19615 73312 19636 73352
rect 19676 73312 19697 73352
rect 19783 73312 19800 73352
rect 19840 73312 19849 73352
rect 19463 73289 19529 73312
rect 19615 73289 19697 73312
rect 19783 73289 19849 73312
rect 19463 73270 19849 73289
rect 34583 73375 34969 73394
rect 34583 73352 34649 73375
rect 34735 73352 34817 73375
rect 34903 73352 34969 73375
rect 34583 73312 34592 73352
rect 34632 73312 34649 73352
rect 34735 73312 34756 73352
rect 34796 73312 34817 73352
rect 34903 73312 34920 73352
rect 34960 73312 34969 73352
rect 34583 73289 34649 73312
rect 34735 73289 34817 73312
rect 34903 73289 34969 73312
rect 34583 73270 34969 73289
rect 49703 73375 50089 73394
rect 49703 73352 49769 73375
rect 49855 73352 49937 73375
rect 50023 73352 50089 73375
rect 49703 73312 49712 73352
rect 49752 73312 49769 73352
rect 49855 73312 49876 73352
rect 49916 73312 49937 73352
rect 50023 73312 50040 73352
rect 50080 73312 50089 73352
rect 49703 73289 49769 73312
rect 49855 73289 49937 73312
rect 50023 73289 50089 73312
rect 49703 73270 50089 73289
rect 64823 73375 65209 73394
rect 64823 73352 64889 73375
rect 64975 73352 65057 73375
rect 65143 73352 65209 73375
rect 64823 73312 64832 73352
rect 64872 73312 64889 73352
rect 64975 73312 64996 73352
rect 65036 73312 65057 73352
rect 65143 73312 65160 73352
rect 65200 73312 65209 73352
rect 64823 73289 64889 73312
rect 64975 73289 65057 73312
rect 65143 73289 65209 73312
rect 64823 73270 65209 73289
rect 79943 73375 80329 73394
rect 79943 73352 80009 73375
rect 80095 73352 80177 73375
rect 80263 73352 80329 73375
rect 79943 73312 79952 73352
rect 79992 73312 80009 73352
rect 80095 73312 80116 73352
rect 80156 73312 80177 73352
rect 80263 73312 80280 73352
rect 80320 73312 80329 73352
rect 79943 73289 80009 73312
rect 80095 73289 80177 73312
rect 80263 73289 80329 73312
rect 79943 73270 80329 73289
rect 95063 73375 95449 73394
rect 95063 73352 95129 73375
rect 95215 73352 95297 73375
rect 95383 73352 95449 73375
rect 95063 73312 95072 73352
rect 95112 73312 95129 73352
rect 95215 73312 95236 73352
rect 95276 73312 95297 73352
rect 95383 73312 95400 73352
rect 95440 73312 95449 73352
rect 95063 73289 95129 73312
rect 95215 73289 95297 73312
rect 95383 73289 95449 73312
rect 95063 73270 95449 73289
rect 3103 72619 3489 72638
rect 3103 72596 3169 72619
rect 3255 72596 3337 72619
rect 3423 72596 3489 72619
rect 3103 72556 3112 72596
rect 3152 72556 3169 72596
rect 3255 72556 3276 72596
rect 3316 72556 3337 72596
rect 3423 72556 3440 72596
rect 3480 72556 3489 72596
rect 3103 72533 3169 72556
rect 3255 72533 3337 72556
rect 3423 72533 3489 72556
rect 3103 72514 3489 72533
rect 18223 72619 18609 72638
rect 18223 72596 18289 72619
rect 18375 72596 18457 72619
rect 18543 72596 18609 72619
rect 18223 72556 18232 72596
rect 18272 72556 18289 72596
rect 18375 72556 18396 72596
rect 18436 72556 18457 72596
rect 18543 72556 18560 72596
rect 18600 72556 18609 72596
rect 18223 72533 18289 72556
rect 18375 72533 18457 72556
rect 18543 72533 18609 72556
rect 18223 72514 18609 72533
rect 33343 72619 33729 72638
rect 33343 72596 33409 72619
rect 33495 72596 33577 72619
rect 33663 72596 33729 72619
rect 33343 72556 33352 72596
rect 33392 72556 33409 72596
rect 33495 72556 33516 72596
rect 33556 72556 33577 72596
rect 33663 72556 33680 72596
rect 33720 72556 33729 72596
rect 33343 72533 33409 72556
rect 33495 72533 33577 72556
rect 33663 72533 33729 72556
rect 33343 72514 33729 72533
rect 48463 72619 48849 72638
rect 48463 72596 48529 72619
rect 48615 72596 48697 72619
rect 48783 72596 48849 72619
rect 48463 72556 48472 72596
rect 48512 72556 48529 72596
rect 48615 72556 48636 72596
rect 48676 72556 48697 72596
rect 48783 72556 48800 72596
rect 48840 72556 48849 72596
rect 48463 72533 48529 72556
rect 48615 72533 48697 72556
rect 48783 72533 48849 72556
rect 48463 72514 48849 72533
rect 63583 72619 63969 72638
rect 63583 72596 63649 72619
rect 63735 72596 63817 72619
rect 63903 72596 63969 72619
rect 63583 72556 63592 72596
rect 63632 72556 63649 72596
rect 63735 72556 63756 72596
rect 63796 72556 63817 72596
rect 63903 72556 63920 72596
rect 63960 72556 63969 72596
rect 63583 72533 63649 72556
rect 63735 72533 63817 72556
rect 63903 72533 63969 72556
rect 63583 72514 63969 72533
rect 78703 72619 79089 72638
rect 78703 72596 78769 72619
rect 78855 72596 78937 72619
rect 79023 72596 79089 72619
rect 78703 72556 78712 72596
rect 78752 72556 78769 72596
rect 78855 72556 78876 72596
rect 78916 72556 78937 72596
rect 79023 72556 79040 72596
rect 79080 72556 79089 72596
rect 78703 72533 78769 72556
rect 78855 72533 78937 72556
rect 79023 72533 79089 72556
rect 78703 72514 79089 72533
rect 93823 72619 94209 72638
rect 93823 72596 93889 72619
rect 93975 72596 94057 72619
rect 94143 72596 94209 72619
rect 93823 72556 93832 72596
rect 93872 72556 93889 72596
rect 93975 72556 93996 72596
rect 94036 72556 94057 72596
rect 94143 72556 94160 72596
rect 94200 72556 94209 72596
rect 93823 72533 93889 72556
rect 93975 72533 94057 72556
rect 94143 72533 94209 72556
rect 93823 72514 94209 72533
rect 4343 71863 4729 71882
rect 4343 71840 4409 71863
rect 4495 71840 4577 71863
rect 4663 71840 4729 71863
rect 4343 71800 4352 71840
rect 4392 71800 4409 71840
rect 4495 71800 4516 71840
rect 4556 71800 4577 71840
rect 4663 71800 4680 71840
rect 4720 71800 4729 71840
rect 4343 71777 4409 71800
rect 4495 71777 4577 71800
rect 4663 71777 4729 71800
rect 4343 71758 4729 71777
rect 19463 71863 19849 71882
rect 19463 71840 19529 71863
rect 19615 71840 19697 71863
rect 19783 71840 19849 71863
rect 19463 71800 19472 71840
rect 19512 71800 19529 71840
rect 19615 71800 19636 71840
rect 19676 71800 19697 71840
rect 19783 71800 19800 71840
rect 19840 71800 19849 71840
rect 19463 71777 19529 71800
rect 19615 71777 19697 71800
rect 19783 71777 19849 71800
rect 19463 71758 19849 71777
rect 34583 71863 34969 71882
rect 34583 71840 34649 71863
rect 34735 71840 34817 71863
rect 34903 71840 34969 71863
rect 34583 71800 34592 71840
rect 34632 71800 34649 71840
rect 34735 71800 34756 71840
rect 34796 71800 34817 71840
rect 34903 71800 34920 71840
rect 34960 71800 34969 71840
rect 34583 71777 34649 71800
rect 34735 71777 34817 71800
rect 34903 71777 34969 71800
rect 34583 71758 34969 71777
rect 49703 71863 50089 71882
rect 49703 71840 49769 71863
rect 49855 71840 49937 71863
rect 50023 71840 50089 71863
rect 49703 71800 49712 71840
rect 49752 71800 49769 71840
rect 49855 71800 49876 71840
rect 49916 71800 49937 71840
rect 50023 71800 50040 71840
rect 50080 71800 50089 71840
rect 49703 71777 49769 71800
rect 49855 71777 49937 71800
rect 50023 71777 50089 71800
rect 49703 71758 50089 71777
rect 64823 71863 65209 71882
rect 64823 71840 64889 71863
rect 64975 71840 65057 71863
rect 65143 71840 65209 71863
rect 64823 71800 64832 71840
rect 64872 71800 64889 71840
rect 64975 71800 64996 71840
rect 65036 71800 65057 71840
rect 65143 71800 65160 71840
rect 65200 71800 65209 71840
rect 64823 71777 64889 71800
rect 64975 71777 65057 71800
rect 65143 71777 65209 71800
rect 64823 71758 65209 71777
rect 79943 71863 80329 71882
rect 79943 71840 80009 71863
rect 80095 71840 80177 71863
rect 80263 71840 80329 71863
rect 79943 71800 79952 71840
rect 79992 71800 80009 71840
rect 80095 71800 80116 71840
rect 80156 71800 80177 71840
rect 80263 71800 80280 71840
rect 80320 71800 80329 71840
rect 79943 71777 80009 71800
rect 80095 71777 80177 71800
rect 80263 71777 80329 71800
rect 79943 71758 80329 71777
rect 95063 71863 95449 71882
rect 95063 71840 95129 71863
rect 95215 71840 95297 71863
rect 95383 71840 95449 71863
rect 95063 71800 95072 71840
rect 95112 71800 95129 71840
rect 95215 71800 95236 71840
rect 95276 71800 95297 71840
rect 95383 71800 95400 71840
rect 95440 71800 95449 71840
rect 95063 71777 95129 71800
rect 95215 71777 95297 71800
rect 95383 71777 95449 71800
rect 95063 71758 95449 71777
rect 3103 71107 3489 71126
rect 3103 71084 3169 71107
rect 3255 71084 3337 71107
rect 3423 71084 3489 71107
rect 3103 71044 3112 71084
rect 3152 71044 3169 71084
rect 3255 71044 3276 71084
rect 3316 71044 3337 71084
rect 3423 71044 3440 71084
rect 3480 71044 3489 71084
rect 3103 71021 3169 71044
rect 3255 71021 3337 71044
rect 3423 71021 3489 71044
rect 3103 71002 3489 71021
rect 18223 71107 18609 71126
rect 18223 71084 18289 71107
rect 18375 71084 18457 71107
rect 18543 71084 18609 71107
rect 18223 71044 18232 71084
rect 18272 71044 18289 71084
rect 18375 71044 18396 71084
rect 18436 71044 18457 71084
rect 18543 71044 18560 71084
rect 18600 71044 18609 71084
rect 18223 71021 18289 71044
rect 18375 71021 18457 71044
rect 18543 71021 18609 71044
rect 18223 71002 18609 71021
rect 33343 71107 33729 71126
rect 33343 71084 33409 71107
rect 33495 71084 33577 71107
rect 33663 71084 33729 71107
rect 33343 71044 33352 71084
rect 33392 71044 33409 71084
rect 33495 71044 33516 71084
rect 33556 71044 33577 71084
rect 33663 71044 33680 71084
rect 33720 71044 33729 71084
rect 33343 71021 33409 71044
rect 33495 71021 33577 71044
rect 33663 71021 33729 71044
rect 33343 71002 33729 71021
rect 48463 71107 48849 71126
rect 48463 71084 48529 71107
rect 48615 71084 48697 71107
rect 48783 71084 48849 71107
rect 48463 71044 48472 71084
rect 48512 71044 48529 71084
rect 48615 71044 48636 71084
rect 48676 71044 48697 71084
rect 48783 71044 48800 71084
rect 48840 71044 48849 71084
rect 48463 71021 48529 71044
rect 48615 71021 48697 71044
rect 48783 71021 48849 71044
rect 48463 71002 48849 71021
rect 63583 71107 63969 71126
rect 63583 71084 63649 71107
rect 63735 71084 63817 71107
rect 63903 71084 63969 71107
rect 63583 71044 63592 71084
rect 63632 71044 63649 71084
rect 63735 71044 63756 71084
rect 63796 71044 63817 71084
rect 63903 71044 63920 71084
rect 63960 71044 63969 71084
rect 63583 71021 63649 71044
rect 63735 71021 63817 71044
rect 63903 71021 63969 71044
rect 63583 71002 63969 71021
rect 78703 71107 79089 71126
rect 78703 71084 78769 71107
rect 78855 71084 78937 71107
rect 79023 71084 79089 71107
rect 78703 71044 78712 71084
rect 78752 71044 78769 71084
rect 78855 71044 78876 71084
rect 78916 71044 78937 71084
rect 79023 71044 79040 71084
rect 79080 71044 79089 71084
rect 78703 71021 78769 71044
rect 78855 71021 78937 71044
rect 79023 71021 79089 71044
rect 78703 71002 79089 71021
rect 93823 71107 94209 71126
rect 93823 71084 93889 71107
rect 93975 71084 94057 71107
rect 94143 71084 94209 71107
rect 93823 71044 93832 71084
rect 93872 71044 93889 71084
rect 93975 71044 93996 71084
rect 94036 71044 94057 71084
rect 94143 71044 94160 71084
rect 94200 71044 94209 71084
rect 93823 71021 93889 71044
rect 93975 71021 94057 71044
rect 94143 71021 94209 71044
rect 93823 71002 94209 71021
rect 4343 70351 4729 70370
rect 4343 70328 4409 70351
rect 4495 70328 4577 70351
rect 4663 70328 4729 70351
rect 4343 70288 4352 70328
rect 4392 70288 4409 70328
rect 4495 70288 4516 70328
rect 4556 70288 4577 70328
rect 4663 70288 4680 70328
rect 4720 70288 4729 70328
rect 4343 70265 4409 70288
rect 4495 70265 4577 70288
rect 4663 70265 4729 70288
rect 4343 70246 4729 70265
rect 19463 70351 19849 70370
rect 19463 70328 19529 70351
rect 19615 70328 19697 70351
rect 19783 70328 19849 70351
rect 19463 70288 19472 70328
rect 19512 70288 19529 70328
rect 19615 70288 19636 70328
rect 19676 70288 19697 70328
rect 19783 70288 19800 70328
rect 19840 70288 19849 70328
rect 19463 70265 19529 70288
rect 19615 70265 19697 70288
rect 19783 70265 19849 70288
rect 19463 70246 19849 70265
rect 34583 70351 34969 70370
rect 34583 70328 34649 70351
rect 34735 70328 34817 70351
rect 34903 70328 34969 70351
rect 34583 70288 34592 70328
rect 34632 70288 34649 70328
rect 34735 70288 34756 70328
rect 34796 70288 34817 70328
rect 34903 70288 34920 70328
rect 34960 70288 34969 70328
rect 34583 70265 34649 70288
rect 34735 70265 34817 70288
rect 34903 70265 34969 70288
rect 34583 70246 34969 70265
rect 49703 70351 50089 70370
rect 49703 70328 49769 70351
rect 49855 70328 49937 70351
rect 50023 70328 50089 70351
rect 49703 70288 49712 70328
rect 49752 70288 49769 70328
rect 49855 70288 49876 70328
rect 49916 70288 49937 70328
rect 50023 70288 50040 70328
rect 50080 70288 50089 70328
rect 49703 70265 49769 70288
rect 49855 70265 49937 70288
rect 50023 70265 50089 70288
rect 49703 70246 50089 70265
rect 64823 70351 65209 70370
rect 64823 70328 64889 70351
rect 64975 70328 65057 70351
rect 65143 70328 65209 70351
rect 64823 70288 64832 70328
rect 64872 70288 64889 70328
rect 64975 70288 64996 70328
rect 65036 70288 65057 70328
rect 65143 70288 65160 70328
rect 65200 70288 65209 70328
rect 64823 70265 64889 70288
rect 64975 70265 65057 70288
rect 65143 70265 65209 70288
rect 64823 70246 65209 70265
rect 79943 70351 80329 70370
rect 79943 70328 80009 70351
rect 80095 70328 80177 70351
rect 80263 70328 80329 70351
rect 79943 70288 79952 70328
rect 79992 70288 80009 70328
rect 80095 70288 80116 70328
rect 80156 70288 80177 70328
rect 80263 70288 80280 70328
rect 80320 70288 80329 70328
rect 79943 70265 80009 70288
rect 80095 70265 80177 70288
rect 80263 70265 80329 70288
rect 79943 70246 80329 70265
rect 95063 70351 95449 70370
rect 95063 70328 95129 70351
rect 95215 70328 95297 70351
rect 95383 70328 95449 70351
rect 95063 70288 95072 70328
rect 95112 70288 95129 70328
rect 95215 70288 95236 70328
rect 95276 70288 95297 70328
rect 95383 70288 95400 70328
rect 95440 70288 95449 70328
rect 95063 70265 95129 70288
rect 95215 70265 95297 70288
rect 95383 70265 95449 70288
rect 95063 70246 95449 70265
rect 3103 69595 3489 69614
rect 3103 69572 3169 69595
rect 3255 69572 3337 69595
rect 3423 69572 3489 69595
rect 3103 69532 3112 69572
rect 3152 69532 3169 69572
rect 3255 69532 3276 69572
rect 3316 69532 3337 69572
rect 3423 69532 3440 69572
rect 3480 69532 3489 69572
rect 3103 69509 3169 69532
rect 3255 69509 3337 69532
rect 3423 69509 3489 69532
rect 3103 69490 3489 69509
rect 18223 69595 18609 69614
rect 18223 69572 18289 69595
rect 18375 69572 18457 69595
rect 18543 69572 18609 69595
rect 18223 69532 18232 69572
rect 18272 69532 18289 69572
rect 18375 69532 18396 69572
rect 18436 69532 18457 69572
rect 18543 69532 18560 69572
rect 18600 69532 18609 69572
rect 18223 69509 18289 69532
rect 18375 69509 18457 69532
rect 18543 69509 18609 69532
rect 18223 69490 18609 69509
rect 33343 69595 33729 69614
rect 33343 69572 33409 69595
rect 33495 69572 33577 69595
rect 33663 69572 33729 69595
rect 33343 69532 33352 69572
rect 33392 69532 33409 69572
rect 33495 69532 33516 69572
rect 33556 69532 33577 69572
rect 33663 69532 33680 69572
rect 33720 69532 33729 69572
rect 33343 69509 33409 69532
rect 33495 69509 33577 69532
rect 33663 69509 33729 69532
rect 33343 69490 33729 69509
rect 48463 69595 48849 69614
rect 48463 69572 48529 69595
rect 48615 69572 48697 69595
rect 48783 69572 48849 69595
rect 48463 69532 48472 69572
rect 48512 69532 48529 69572
rect 48615 69532 48636 69572
rect 48676 69532 48697 69572
rect 48783 69532 48800 69572
rect 48840 69532 48849 69572
rect 48463 69509 48529 69532
rect 48615 69509 48697 69532
rect 48783 69509 48849 69532
rect 48463 69490 48849 69509
rect 63583 69595 63969 69614
rect 63583 69572 63649 69595
rect 63735 69572 63817 69595
rect 63903 69572 63969 69595
rect 63583 69532 63592 69572
rect 63632 69532 63649 69572
rect 63735 69532 63756 69572
rect 63796 69532 63817 69572
rect 63903 69532 63920 69572
rect 63960 69532 63969 69572
rect 63583 69509 63649 69532
rect 63735 69509 63817 69532
rect 63903 69509 63969 69532
rect 63583 69490 63969 69509
rect 78703 69595 79089 69614
rect 78703 69572 78769 69595
rect 78855 69572 78937 69595
rect 79023 69572 79089 69595
rect 78703 69532 78712 69572
rect 78752 69532 78769 69572
rect 78855 69532 78876 69572
rect 78916 69532 78937 69572
rect 79023 69532 79040 69572
rect 79080 69532 79089 69572
rect 78703 69509 78769 69532
rect 78855 69509 78937 69532
rect 79023 69509 79089 69532
rect 78703 69490 79089 69509
rect 93823 69595 94209 69614
rect 93823 69572 93889 69595
rect 93975 69572 94057 69595
rect 94143 69572 94209 69595
rect 93823 69532 93832 69572
rect 93872 69532 93889 69572
rect 93975 69532 93996 69572
rect 94036 69532 94057 69572
rect 94143 69532 94160 69572
rect 94200 69532 94209 69572
rect 93823 69509 93889 69532
rect 93975 69509 94057 69532
rect 94143 69509 94209 69532
rect 93823 69490 94209 69509
rect 4343 68839 4729 68858
rect 4343 68816 4409 68839
rect 4495 68816 4577 68839
rect 4663 68816 4729 68839
rect 4343 68776 4352 68816
rect 4392 68776 4409 68816
rect 4495 68776 4516 68816
rect 4556 68776 4577 68816
rect 4663 68776 4680 68816
rect 4720 68776 4729 68816
rect 4343 68753 4409 68776
rect 4495 68753 4577 68776
rect 4663 68753 4729 68776
rect 4343 68734 4729 68753
rect 19463 68839 19849 68858
rect 19463 68816 19529 68839
rect 19615 68816 19697 68839
rect 19783 68816 19849 68839
rect 19463 68776 19472 68816
rect 19512 68776 19529 68816
rect 19615 68776 19636 68816
rect 19676 68776 19697 68816
rect 19783 68776 19800 68816
rect 19840 68776 19849 68816
rect 19463 68753 19529 68776
rect 19615 68753 19697 68776
rect 19783 68753 19849 68776
rect 19463 68734 19849 68753
rect 34583 68839 34969 68858
rect 34583 68816 34649 68839
rect 34735 68816 34817 68839
rect 34903 68816 34969 68839
rect 34583 68776 34592 68816
rect 34632 68776 34649 68816
rect 34735 68776 34756 68816
rect 34796 68776 34817 68816
rect 34903 68776 34920 68816
rect 34960 68776 34969 68816
rect 34583 68753 34649 68776
rect 34735 68753 34817 68776
rect 34903 68753 34969 68776
rect 34583 68734 34969 68753
rect 49703 68839 50089 68858
rect 49703 68816 49769 68839
rect 49855 68816 49937 68839
rect 50023 68816 50089 68839
rect 49703 68776 49712 68816
rect 49752 68776 49769 68816
rect 49855 68776 49876 68816
rect 49916 68776 49937 68816
rect 50023 68776 50040 68816
rect 50080 68776 50089 68816
rect 49703 68753 49769 68776
rect 49855 68753 49937 68776
rect 50023 68753 50089 68776
rect 49703 68734 50089 68753
rect 64823 68839 65209 68858
rect 64823 68816 64889 68839
rect 64975 68816 65057 68839
rect 65143 68816 65209 68839
rect 64823 68776 64832 68816
rect 64872 68776 64889 68816
rect 64975 68776 64996 68816
rect 65036 68776 65057 68816
rect 65143 68776 65160 68816
rect 65200 68776 65209 68816
rect 64823 68753 64889 68776
rect 64975 68753 65057 68776
rect 65143 68753 65209 68776
rect 64823 68734 65209 68753
rect 79943 68839 80329 68858
rect 79943 68816 80009 68839
rect 80095 68816 80177 68839
rect 80263 68816 80329 68839
rect 79943 68776 79952 68816
rect 79992 68776 80009 68816
rect 80095 68776 80116 68816
rect 80156 68776 80177 68816
rect 80263 68776 80280 68816
rect 80320 68776 80329 68816
rect 79943 68753 80009 68776
rect 80095 68753 80177 68776
rect 80263 68753 80329 68776
rect 79943 68734 80329 68753
rect 95063 68839 95449 68858
rect 95063 68816 95129 68839
rect 95215 68816 95297 68839
rect 95383 68816 95449 68839
rect 95063 68776 95072 68816
rect 95112 68776 95129 68816
rect 95215 68776 95236 68816
rect 95276 68776 95297 68816
rect 95383 68776 95400 68816
rect 95440 68776 95449 68816
rect 95063 68753 95129 68776
rect 95215 68753 95297 68776
rect 95383 68753 95449 68776
rect 95063 68734 95449 68753
rect 3103 68083 3489 68102
rect 3103 68060 3169 68083
rect 3255 68060 3337 68083
rect 3423 68060 3489 68083
rect 3103 68020 3112 68060
rect 3152 68020 3169 68060
rect 3255 68020 3276 68060
rect 3316 68020 3337 68060
rect 3423 68020 3440 68060
rect 3480 68020 3489 68060
rect 3103 67997 3169 68020
rect 3255 67997 3337 68020
rect 3423 67997 3489 68020
rect 3103 67978 3489 67997
rect 18223 68083 18609 68102
rect 18223 68060 18289 68083
rect 18375 68060 18457 68083
rect 18543 68060 18609 68083
rect 18223 68020 18232 68060
rect 18272 68020 18289 68060
rect 18375 68020 18396 68060
rect 18436 68020 18457 68060
rect 18543 68020 18560 68060
rect 18600 68020 18609 68060
rect 18223 67997 18289 68020
rect 18375 67997 18457 68020
rect 18543 67997 18609 68020
rect 18223 67978 18609 67997
rect 33343 68083 33729 68102
rect 33343 68060 33409 68083
rect 33495 68060 33577 68083
rect 33663 68060 33729 68083
rect 33343 68020 33352 68060
rect 33392 68020 33409 68060
rect 33495 68020 33516 68060
rect 33556 68020 33577 68060
rect 33663 68020 33680 68060
rect 33720 68020 33729 68060
rect 33343 67997 33409 68020
rect 33495 67997 33577 68020
rect 33663 67997 33729 68020
rect 33343 67978 33729 67997
rect 48463 68083 48849 68102
rect 48463 68060 48529 68083
rect 48615 68060 48697 68083
rect 48783 68060 48849 68083
rect 48463 68020 48472 68060
rect 48512 68020 48529 68060
rect 48615 68020 48636 68060
rect 48676 68020 48697 68060
rect 48783 68020 48800 68060
rect 48840 68020 48849 68060
rect 48463 67997 48529 68020
rect 48615 67997 48697 68020
rect 48783 67997 48849 68020
rect 48463 67978 48849 67997
rect 63583 68083 63969 68102
rect 63583 68060 63649 68083
rect 63735 68060 63817 68083
rect 63903 68060 63969 68083
rect 63583 68020 63592 68060
rect 63632 68020 63649 68060
rect 63735 68020 63756 68060
rect 63796 68020 63817 68060
rect 63903 68020 63920 68060
rect 63960 68020 63969 68060
rect 63583 67997 63649 68020
rect 63735 67997 63817 68020
rect 63903 67997 63969 68020
rect 63583 67978 63969 67997
rect 78703 68083 79089 68102
rect 78703 68060 78769 68083
rect 78855 68060 78937 68083
rect 79023 68060 79089 68083
rect 78703 68020 78712 68060
rect 78752 68020 78769 68060
rect 78855 68020 78876 68060
rect 78916 68020 78937 68060
rect 79023 68020 79040 68060
rect 79080 68020 79089 68060
rect 78703 67997 78769 68020
rect 78855 67997 78937 68020
rect 79023 67997 79089 68020
rect 78703 67978 79089 67997
rect 93823 68083 94209 68102
rect 93823 68060 93889 68083
rect 93975 68060 94057 68083
rect 94143 68060 94209 68083
rect 93823 68020 93832 68060
rect 93872 68020 93889 68060
rect 93975 68020 93996 68060
rect 94036 68020 94057 68060
rect 94143 68020 94160 68060
rect 94200 68020 94209 68060
rect 93823 67997 93889 68020
rect 93975 67997 94057 68020
rect 94143 67997 94209 68020
rect 93823 67978 94209 67997
rect 4343 67327 4729 67346
rect 4343 67304 4409 67327
rect 4495 67304 4577 67327
rect 4663 67304 4729 67327
rect 4343 67264 4352 67304
rect 4392 67264 4409 67304
rect 4495 67264 4516 67304
rect 4556 67264 4577 67304
rect 4663 67264 4680 67304
rect 4720 67264 4729 67304
rect 4343 67241 4409 67264
rect 4495 67241 4577 67264
rect 4663 67241 4729 67264
rect 4343 67222 4729 67241
rect 19463 67327 19849 67346
rect 19463 67304 19529 67327
rect 19615 67304 19697 67327
rect 19783 67304 19849 67327
rect 19463 67264 19472 67304
rect 19512 67264 19529 67304
rect 19615 67264 19636 67304
rect 19676 67264 19697 67304
rect 19783 67264 19800 67304
rect 19840 67264 19849 67304
rect 19463 67241 19529 67264
rect 19615 67241 19697 67264
rect 19783 67241 19849 67264
rect 19463 67222 19849 67241
rect 34583 67327 34969 67346
rect 34583 67304 34649 67327
rect 34735 67304 34817 67327
rect 34903 67304 34969 67327
rect 34583 67264 34592 67304
rect 34632 67264 34649 67304
rect 34735 67264 34756 67304
rect 34796 67264 34817 67304
rect 34903 67264 34920 67304
rect 34960 67264 34969 67304
rect 34583 67241 34649 67264
rect 34735 67241 34817 67264
rect 34903 67241 34969 67264
rect 34583 67222 34969 67241
rect 49703 67327 50089 67346
rect 49703 67304 49769 67327
rect 49855 67304 49937 67327
rect 50023 67304 50089 67327
rect 49703 67264 49712 67304
rect 49752 67264 49769 67304
rect 49855 67264 49876 67304
rect 49916 67264 49937 67304
rect 50023 67264 50040 67304
rect 50080 67264 50089 67304
rect 49703 67241 49769 67264
rect 49855 67241 49937 67264
rect 50023 67241 50089 67264
rect 49703 67222 50089 67241
rect 64823 67327 65209 67346
rect 64823 67304 64889 67327
rect 64975 67304 65057 67327
rect 65143 67304 65209 67327
rect 64823 67264 64832 67304
rect 64872 67264 64889 67304
rect 64975 67264 64996 67304
rect 65036 67264 65057 67304
rect 65143 67264 65160 67304
rect 65200 67264 65209 67304
rect 64823 67241 64889 67264
rect 64975 67241 65057 67264
rect 65143 67241 65209 67264
rect 64823 67222 65209 67241
rect 79943 67327 80329 67346
rect 79943 67304 80009 67327
rect 80095 67304 80177 67327
rect 80263 67304 80329 67327
rect 79943 67264 79952 67304
rect 79992 67264 80009 67304
rect 80095 67264 80116 67304
rect 80156 67264 80177 67304
rect 80263 67264 80280 67304
rect 80320 67264 80329 67304
rect 79943 67241 80009 67264
rect 80095 67241 80177 67264
rect 80263 67241 80329 67264
rect 79943 67222 80329 67241
rect 95063 67327 95449 67346
rect 95063 67304 95129 67327
rect 95215 67304 95297 67327
rect 95383 67304 95449 67327
rect 95063 67264 95072 67304
rect 95112 67264 95129 67304
rect 95215 67264 95236 67304
rect 95276 67264 95297 67304
rect 95383 67264 95400 67304
rect 95440 67264 95449 67304
rect 95063 67241 95129 67264
rect 95215 67241 95297 67264
rect 95383 67241 95449 67264
rect 95063 67222 95449 67241
rect 3103 66571 3489 66590
rect 3103 66548 3169 66571
rect 3255 66548 3337 66571
rect 3423 66548 3489 66571
rect 3103 66508 3112 66548
rect 3152 66508 3169 66548
rect 3255 66508 3276 66548
rect 3316 66508 3337 66548
rect 3423 66508 3440 66548
rect 3480 66508 3489 66548
rect 3103 66485 3169 66508
rect 3255 66485 3337 66508
rect 3423 66485 3489 66508
rect 3103 66466 3489 66485
rect 18223 66571 18609 66590
rect 18223 66548 18289 66571
rect 18375 66548 18457 66571
rect 18543 66548 18609 66571
rect 18223 66508 18232 66548
rect 18272 66508 18289 66548
rect 18375 66508 18396 66548
rect 18436 66508 18457 66548
rect 18543 66508 18560 66548
rect 18600 66508 18609 66548
rect 18223 66485 18289 66508
rect 18375 66485 18457 66508
rect 18543 66485 18609 66508
rect 18223 66466 18609 66485
rect 33343 66571 33729 66590
rect 33343 66548 33409 66571
rect 33495 66548 33577 66571
rect 33663 66548 33729 66571
rect 33343 66508 33352 66548
rect 33392 66508 33409 66548
rect 33495 66508 33516 66548
rect 33556 66508 33577 66548
rect 33663 66508 33680 66548
rect 33720 66508 33729 66548
rect 33343 66485 33409 66508
rect 33495 66485 33577 66508
rect 33663 66485 33729 66508
rect 33343 66466 33729 66485
rect 48463 66571 48849 66590
rect 48463 66548 48529 66571
rect 48615 66548 48697 66571
rect 48783 66548 48849 66571
rect 48463 66508 48472 66548
rect 48512 66508 48529 66548
rect 48615 66508 48636 66548
rect 48676 66508 48697 66548
rect 48783 66508 48800 66548
rect 48840 66508 48849 66548
rect 48463 66485 48529 66508
rect 48615 66485 48697 66508
rect 48783 66485 48849 66508
rect 48463 66466 48849 66485
rect 63583 66571 63969 66590
rect 63583 66548 63649 66571
rect 63735 66548 63817 66571
rect 63903 66548 63969 66571
rect 63583 66508 63592 66548
rect 63632 66508 63649 66548
rect 63735 66508 63756 66548
rect 63796 66508 63817 66548
rect 63903 66508 63920 66548
rect 63960 66508 63969 66548
rect 63583 66485 63649 66508
rect 63735 66485 63817 66508
rect 63903 66485 63969 66508
rect 63583 66466 63969 66485
rect 78703 66571 79089 66590
rect 78703 66548 78769 66571
rect 78855 66548 78937 66571
rect 79023 66548 79089 66571
rect 78703 66508 78712 66548
rect 78752 66508 78769 66548
rect 78855 66508 78876 66548
rect 78916 66508 78937 66548
rect 79023 66508 79040 66548
rect 79080 66508 79089 66548
rect 78703 66485 78769 66508
rect 78855 66485 78937 66508
rect 79023 66485 79089 66508
rect 78703 66466 79089 66485
rect 93823 66571 94209 66590
rect 93823 66548 93889 66571
rect 93975 66548 94057 66571
rect 94143 66548 94209 66571
rect 93823 66508 93832 66548
rect 93872 66508 93889 66548
rect 93975 66508 93996 66548
rect 94036 66508 94057 66548
rect 94143 66508 94160 66548
rect 94200 66508 94209 66548
rect 93823 66485 93889 66508
rect 93975 66485 94057 66508
rect 94143 66485 94209 66508
rect 93823 66466 94209 66485
rect 4343 65815 4729 65834
rect 4343 65792 4409 65815
rect 4495 65792 4577 65815
rect 4663 65792 4729 65815
rect 4343 65752 4352 65792
rect 4392 65752 4409 65792
rect 4495 65752 4516 65792
rect 4556 65752 4577 65792
rect 4663 65752 4680 65792
rect 4720 65752 4729 65792
rect 4343 65729 4409 65752
rect 4495 65729 4577 65752
rect 4663 65729 4729 65752
rect 4343 65710 4729 65729
rect 19463 65815 19849 65834
rect 19463 65792 19529 65815
rect 19615 65792 19697 65815
rect 19783 65792 19849 65815
rect 19463 65752 19472 65792
rect 19512 65752 19529 65792
rect 19615 65752 19636 65792
rect 19676 65752 19697 65792
rect 19783 65752 19800 65792
rect 19840 65752 19849 65792
rect 19463 65729 19529 65752
rect 19615 65729 19697 65752
rect 19783 65729 19849 65752
rect 19463 65710 19849 65729
rect 34583 65815 34969 65834
rect 34583 65792 34649 65815
rect 34735 65792 34817 65815
rect 34903 65792 34969 65815
rect 34583 65752 34592 65792
rect 34632 65752 34649 65792
rect 34735 65752 34756 65792
rect 34796 65752 34817 65792
rect 34903 65752 34920 65792
rect 34960 65752 34969 65792
rect 34583 65729 34649 65752
rect 34735 65729 34817 65752
rect 34903 65729 34969 65752
rect 34583 65710 34969 65729
rect 49703 65815 50089 65834
rect 49703 65792 49769 65815
rect 49855 65792 49937 65815
rect 50023 65792 50089 65815
rect 49703 65752 49712 65792
rect 49752 65752 49769 65792
rect 49855 65752 49876 65792
rect 49916 65752 49937 65792
rect 50023 65752 50040 65792
rect 50080 65752 50089 65792
rect 49703 65729 49769 65752
rect 49855 65729 49937 65752
rect 50023 65729 50089 65752
rect 49703 65710 50089 65729
rect 64823 65815 65209 65834
rect 64823 65792 64889 65815
rect 64975 65792 65057 65815
rect 65143 65792 65209 65815
rect 64823 65752 64832 65792
rect 64872 65752 64889 65792
rect 64975 65752 64996 65792
rect 65036 65752 65057 65792
rect 65143 65752 65160 65792
rect 65200 65752 65209 65792
rect 64823 65729 64889 65752
rect 64975 65729 65057 65752
rect 65143 65729 65209 65752
rect 64823 65710 65209 65729
rect 79943 65815 80329 65834
rect 79943 65792 80009 65815
rect 80095 65792 80177 65815
rect 80263 65792 80329 65815
rect 79943 65752 79952 65792
rect 79992 65752 80009 65792
rect 80095 65752 80116 65792
rect 80156 65752 80177 65792
rect 80263 65752 80280 65792
rect 80320 65752 80329 65792
rect 79943 65729 80009 65752
rect 80095 65729 80177 65752
rect 80263 65729 80329 65752
rect 79943 65710 80329 65729
rect 95063 65815 95449 65834
rect 95063 65792 95129 65815
rect 95215 65792 95297 65815
rect 95383 65792 95449 65815
rect 95063 65752 95072 65792
rect 95112 65752 95129 65792
rect 95215 65752 95236 65792
rect 95276 65752 95297 65792
rect 95383 65752 95400 65792
rect 95440 65752 95449 65792
rect 95063 65729 95129 65752
rect 95215 65729 95297 65752
rect 95383 65729 95449 65752
rect 95063 65710 95449 65729
rect 3103 65059 3489 65078
rect 3103 65036 3169 65059
rect 3255 65036 3337 65059
rect 3423 65036 3489 65059
rect 3103 64996 3112 65036
rect 3152 64996 3169 65036
rect 3255 64996 3276 65036
rect 3316 64996 3337 65036
rect 3423 64996 3440 65036
rect 3480 64996 3489 65036
rect 3103 64973 3169 64996
rect 3255 64973 3337 64996
rect 3423 64973 3489 64996
rect 3103 64954 3489 64973
rect 18223 65059 18609 65078
rect 18223 65036 18289 65059
rect 18375 65036 18457 65059
rect 18543 65036 18609 65059
rect 18223 64996 18232 65036
rect 18272 64996 18289 65036
rect 18375 64996 18396 65036
rect 18436 64996 18457 65036
rect 18543 64996 18560 65036
rect 18600 64996 18609 65036
rect 18223 64973 18289 64996
rect 18375 64973 18457 64996
rect 18543 64973 18609 64996
rect 18223 64954 18609 64973
rect 33343 65059 33729 65078
rect 33343 65036 33409 65059
rect 33495 65036 33577 65059
rect 33663 65036 33729 65059
rect 33343 64996 33352 65036
rect 33392 64996 33409 65036
rect 33495 64996 33516 65036
rect 33556 64996 33577 65036
rect 33663 64996 33680 65036
rect 33720 64996 33729 65036
rect 33343 64973 33409 64996
rect 33495 64973 33577 64996
rect 33663 64973 33729 64996
rect 33343 64954 33729 64973
rect 48463 65059 48849 65078
rect 48463 65036 48529 65059
rect 48615 65036 48697 65059
rect 48783 65036 48849 65059
rect 48463 64996 48472 65036
rect 48512 64996 48529 65036
rect 48615 64996 48636 65036
rect 48676 64996 48697 65036
rect 48783 64996 48800 65036
rect 48840 64996 48849 65036
rect 48463 64973 48529 64996
rect 48615 64973 48697 64996
rect 48783 64973 48849 64996
rect 48463 64954 48849 64973
rect 63583 65059 63969 65078
rect 63583 65036 63649 65059
rect 63735 65036 63817 65059
rect 63903 65036 63969 65059
rect 63583 64996 63592 65036
rect 63632 64996 63649 65036
rect 63735 64996 63756 65036
rect 63796 64996 63817 65036
rect 63903 64996 63920 65036
rect 63960 64996 63969 65036
rect 63583 64973 63649 64996
rect 63735 64973 63817 64996
rect 63903 64973 63969 64996
rect 63583 64954 63969 64973
rect 78703 65059 79089 65078
rect 78703 65036 78769 65059
rect 78855 65036 78937 65059
rect 79023 65036 79089 65059
rect 78703 64996 78712 65036
rect 78752 64996 78769 65036
rect 78855 64996 78876 65036
rect 78916 64996 78937 65036
rect 79023 64996 79040 65036
rect 79080 64996 79089 65036
rect 78703 64973 78769 64996
rect 78855 64973 78937 64996
rect 79023 64973 79089 64996
rect 78703 64954 79089 64973
rect 93823 65059 94209 65078
rect 93823 65036 93889 65059
rect 93975 65036 94057 65059
rect 94143 65036 94209 65059
rect 93823 64996 93832 65036
rect 93872 64996 93889 65036
rect 93975 64996 93996 65036
rect 94036 64996 94057 65036
rect 94143 64996 94160 65036
rect 94200 64996 94209 65036
rect 93823 64973 93889 64996
rect 93975 64973 94057 64996
rect 94143 64973 94209 64996
rect 93823 64954 94209 64973
rect 4343 64303 4729 64322
rect 4343 64280 4409 64303
rect 4495 64280 4577 64303
rect 4663 64280 4729 64303
rect 4343 64240 4352 64280
rect 4392 64240 4409 64280
rect 4495 64240 4516 64280
rect 4556 64240 4577 64280
rect 4663 64240 4680 64280
rect 4720 64240 4729 64280
rect 4343 64217 4409 64240
rect 4495 64217 4577 64240
rect 4663 64217 4729 64240
rect 4343 64198 4729 64217
rect 19463 64303 19849 64322
rect 19463 64280 19529 64303
rect 19615 64280 19697 64303
rect 19783 64280 19849 64303
rect 19463 64240 19472 64280
rect 19512 64240 19529 64280
rect 19615 64240 19636 64280
rect 19676 64240 19697 64280
rect 19783 64240 19800 64280
rect 19840 64240 19849 64280
rect 19463 64217 19529 64240
rect 19615 64217 19697 64240
rect 19783 64217 19849 64240
rect 19463 64198 19849 64217
rect 34583 64303 34969 64322
rect 34583 64280 34649 64303
rect 34735 64280 34817 64303
rect 34903 64280 34969 64303
rect 34583 64240 34592 64280
rect 34632 64240 34649 64280
rect 34735 64240 34756 64280
rect 34796 64240 34817 64280
rect 34903 64240 34920 64280
rect 34960 64240 34969 64280
rect 34583 64217 34649 64240
rect 34735 64217 34817 64240
rect 34903 64217 34969 64240
rect 34583 64198 34969 64217
rect 49703 64303 50089 64322
rect 49703 64280 49769 64303
rect 49855 64280 49937 64303
rect 50023 64280 50089 64303
rect 49703 64240 49712 64280
rect 49752 64240 49769 64280
rect 49855 64240 49876 64280
rect 49916 64240 49937 64280
rect 50023 64240 50040 64280
rect 50080 64240 50089 64280
rect 49703 64217 49769 64240
rect 49855 64217 49937 64240
rect 50023 64217 50089 64240
rect 49703 64198 50089 64217
rect 64823 64303 65209 64322
rect 64823 64280 64889 64303
rect 64975 64280 65057 64303
rect 65143 64280 65209 64303
rect 64823 64240 64832 64280
rect 64872 64240 64889 64280
rect 64975 64240 64996 64280
rect 65036 64240 65057 64280
rect 65143 64240 65160 64280
rect 65200 64240 65209 64280
rect 64823 64217 64889 64240
rect 64975 64217 65057 64240
rect 65143 64217 65209 64240
rect 64823 64198 65209 64217
rect 79943 64303 80329 64322
rect 79943 64280 80009 64303
rect 80095 64280 80177 64303
rect 80263 64280 80329 64303
rect 79943 64240 79952 64280
rect 79992 64240 80009 64280
rect 80095 64240 80116 64280
rect 80156 64240 80177 64280
rect 80263 64240 80280 64280
rect 80320 64240 80329 64280
rect 79943 64217 80009 64240
rect 80095 64217 80177 64240
rect 80263 64217 80329 64240
rect 79943 64198 80329 64217
rect 95063 64303 95449 64322
rect 95063 64280 95129 64303
rect 95215 64280 95297 64303
rect 95383 64280 95449 64303
rect 95063 64240 95072 64280
rect 95112 64240 95129 64280
rect 95215 64240 95236 64280
rect 95276 64240 95297 64280
rect 95383 64240 95400 64280
rect 95440 64240 95449 64280
rect 95063 64217 95129 64240
rect 95215 64217 95297 64240
rect 95383 64217 95449 64240
rect 95063 64198 95449 64217
rect 3103 63547 3489 63566
rect 3103 63524 3169 63547
rect 3255 63524 3337 63547
rect 3423 63524 3489 63547
rect 3103 63484 3112 63524
rect 3152 63484 3169 63524
rect 3255 63484 3276 63524
rect 3316 63484 3337 63524
rect 3423 63484 3440 63524
rect 3480 63484 3489 63524
rect 3103 63461 3169 63484
rect 3255 63461 3337 63484
rect 3423 63461 3489 63484
rect 3103 63442 3489 63461
rect 18223 63547 18609 63566
rect 18223 63524 18289 63547
rect 18375 63524 18457 63547
rect 18543 63524 18609 63547
rect 18223 63484 18232 63524
rect 18272 63484 18289 63524
rect 18375 63484 18396 63524
rect 18436 63484 18457 63524
rect 18543 63484 18560 63524
rect 18600 63484 18609 63524
rect 18223 63461 18289 63484
rect 18375 63461 18457 63484
rect 18543 63461 18609 63484
rect 18223 63442 18609 63461
rect 33343 63547 33729 63566
rect 33343 63524 33409 63547
rect 33495 63524 33577 63547
rect 33663 63524 33729 63547
rect 33343 63484 33352 63524
rect 33392 63484 33409 63524
rect 33495 63484 33516 63524
rect 33556 63484 33577 63524
rect 33663 63484 33680 63524
rect 33720 63484 33729 63524
rect 33343 63461 33409 63484
rect 33495 63461 33577 63484
rect 33663 63461 33729 63484
rect 33343 63442 33729 63461
rect 48463 63547 48849 63566
rect 48463 63524 48529 63547
rect 48615 63524 48697 63547
rect 48783 63524 48849 63547
rect 48463 63484 48472 63524
rect 48512 63484 48529 63524
rect 48615 63484 48636 63524
rect 48676 63484 48697 63524
rect 48783 63484 48800 63524
rect 48840 63484 48849 63524
rect 48463 63461 48529 63484
rect 48615 63461 48697 63484
rect 48783 63461 48849 63484
rect 48463 63442 48849 63461
rect 63583 63547 63969 63566
rect 63583 63524 63649 63547
rect 63735 63524 63817 63547
rect 63903 63524 63969 63547
rect 63583 63484 63592 63524
rect 63632 63484 63649 63524
rect 63735 63484 63756 63524
rect 63796 63484 63817 63524
rect 63903 63484 63920 63524
rect 63960 63484 63969 63524
rect 63583 63461 63649 63484
rect 63735 63461 63817 63484
rect 63903 63461 63969 63484
rect 63583 63442 63969 63461
rect 78703 63547 79089 63566
rect 78703 63524 78769 63547
rect 78855 63524 78937 63547
rect 79023 63524 79089 63547
rect 78703 63484 78712 63524
rect 78752 63484 78769 63524
rect 78855 63484 78876 63524
rect 78916 63484 78937 63524
rect 79023 63484 79040 63524
rect 79080 63484 79089 63524
rect 78703 63461 78769 63484
rect 78855 63461 78937 63484
rect 79023 63461 79089 63484
rect 78703 63442 79089 63461
rect 93823 63547 94209 63566
rect 93823 63524 93889 63547
rect 93975 63524 94057 63547
rect 94143 63524 94209 63547
rect 93823 63484 93832 63524
rect 93872 63484 93889 63524
rect 93975 63484 93996 63524
rect 94036 63484 94057 63524
rect 94143 63484 94160 63524
rect 94200 63484 94209 63524
rect 93823 63461 93889 63484
rect 93975 63461 94057 63484
rect 94143 63461 94209 63484
rect 93823 63442 94209 63461
rect 4343 62791 4729 62810
rect 4343 62768 4409 62791
rect 4495 62768 4577 62791
rect 4663 62768 4729 62791
rect 4343 62728 4352 62768
rect 4392 62728 4409 62768
rect 4495 62728 4516 62768
rect 4556 62728 4577 62768
rect 4663 62728 4680 62768
rect 4720 62728 4729 62768
rect 4343 62705 4409 62728
rect 4495 62705 4577 62728
rect 4663 62705 4729 62728
rect 4343 62686 4729 62705
rect 19463 62791 19849 62810
rect 19463 62768 19529 62791
rect 19615 62768 19697 62791
rect 19783 62768 19849 62791
rect 19463 62728 19472 62768
rect 19512 62728 19529 62768
rect 19615 62728 19636 62768
rect 19676 62728 19697 62768
rect 19783 62728 19800 62768
rect 19840 62728 19849 62768
rect 19463 62705 19529 62728
rect 19615 62705 19697 62728
rect 19783 62705 19849 62728
rect 19463 62686 19849 62705
rect 34583 62791 34969 62810
rect 34583 62768 34649 62791
rect 34735 62768 34817 62791
rect 34903 62768 34969 62791
rect 34583 62728 34592 62768
rect 34632 62728 34649 62768
rect 34735 62728 34756 62768
rect 34796 62728 34817 62768
rect 34903 62728 34920 62768
rect 34960 62728 34969 62768
rect 34583 62705 34649 62728
rect 34735 62705 34817 62728
rect 34903 62705 34969 62728
rect 34583 62686 34969 62705
rect 49703 62791 50089 62810
rect 49703 62768 49769 62791
rect 49855 62768 49937 62791
rect 50023 62768 50089 62791
rect 49703 62728 49712 62768
rect 49752 62728 49769 62768
rect 49855 62728 49876 62768
rect 49916 62728 49937 62768
rect 50023 62728 50040 62768
rect 50080 62728 50089 62768
rect 49703 62705 49769 62728
rect 49855 62705 49937 62728
rect 50023 62705 50089 62728
rect 49703 62686 50089 62705
rect 64823 62791 65209 62810
rect 64823 62768 64889 62791
rect 64975 62768 65057 62791
rect 65143 62768 65209 62791
rect 64823 62728 64832 62768
rect 64872 62728 64889 62768
rect 64975 62728 64996 62768
rect 65036 62728 65057 62768
rect 65143 62728 65160 62768
rect 65200 62728 65209 62768
rect 64823 62705 64889 62728
rect 64975 62705 65057 62728
rect 65143 62705 65209 62728
rect 64823 62686 65209 62705
rect 79943 62791 80329 62810
rect 79943 62768 80009 62791
rect 80095 62768 80177 62791
rect 80263 62768 80329 62791
rect 79943 62728 79952 62768
rect 79992 62728 80009 62768
rect 80095 62728 80116 62768
rect 80156 62728 80177 62768
rect 80263 62728 80280 62768
rect 80320 62728 80329 62768
rect 79943 62705 80009 62728
rect 80095 62705 80177 62728
rect 80263 62705 80329 62728
rect 79943 62686 80329 62705
rect 95063 62791 95449 62810
rect 95063 62768 95129 62791
rect 95215 62768 95297 62791
rect 95383 62768 95449 62791
rect 95063 62728 95072 62768
rect 95112 62728 95129 62768
rect 95215 62728 95236 62768
rect 95276 62728 95297 62768
rect 95383 62728 95400 62768
rect 95440 62728 95449 62768
rect 95063 62705 95129 62728
rect 95215 62705 95297 62728
rect 95383 62705 95449 62728
rect 95063 62686 95449 62705
rect 3103 62035 3489 62054
rect 3103 62012 3169 62035
rect 3255 62012 3337 62035
rect 3423 62012 3489 62035
rect 3103 61972 3112 62012
rect 3152 61972 3169 62012
rect 3255 61972 3276 62012
rect 3316 61972 3337 62012
rect 3423 61972 3440 62012
rect 3480 61972 3489 62012
rect 3103 61949 3169 61972
rect 3255 61949 3337 61972
rect 3423 61949 3489 61972
rect 3103 61930 3489 61949
rect 18223 62035 18609 62054
rect 18223 62012 18289 62035
rect 18375 62012 18457 62035
rect 18543 62012 18609 62035
rect 18223 61972 18232 62012
rect 18272 61972 18289 62012
rect 18375 61972 18396 62012
rect 18436 61972 18457 62012
rect 18543 61972 18560 62012
rect 18600 61972 18609 62012
rect 18223 61949 18289 61972
rect 18375 61949 18457 61972
rect 18543 61949 18609 61972
rect 18223 61930 18609 61949
rect 33343 62035 33729 62054
rect 33343 62012 33409 62035
rect 33495 62012 33577 62035
rect 33663 62012 33729 62035
rect 33343 61972 33352 62012
rect 33392 61972 33409 62012
rect 33495 61972 33516 62012
rect 33556 61972 33577 62012
rect 33663 61972 33680 62012
rect 33720 61972 33729 62012
rect 33343 61949 33409 61972
rect 33495 61949 33577 61972
rect 33663 61949 33729 61972
rect 33343 61930 33729 61949
rect 48463 62035 48849 62054
rect 48463 62012 48529 62035
rect 48615 62012 48697 62035
rect 48783 62012 48849 62035
rect 48463 61972 48472 62012
rect 48512 61972 48529 62012
rect 48615 61972 48636 62012
rect 48676 61972 48697 62012
rect 48783 61972 48800 62012
rect 48840 61972 48849 62012
rect 48463 61949 48529 61972
rect 48615 61949 48697 61972
rect 48783 61949 48849 61972
rect 48463 61930 48849 61949
rect 63583 62035 63969 62054
rect 63583 62012 63649 62035
rect 63735 62012 63817 62035
rect 63903 62012 63969 62035
rect 63583 61972 63592 62012
rect 63632 61972 63649 62012
rect 63735 61972 63756 62012
rect 63796 61972 63817 62012
rect 63903 61972 63920 62012
rect 63960 61972 63969 62012
rect 63583 61949 63649 61972
rect 63735 61949 63817 61972
rect 63903 61949 63969 61972
rect 63583 61930 63969 61949
rect 78703 62035 79089 62054
rect 78703 62012 78769 62035
rect 78855 62012 78937 62035
rect 79023 62012 79089 62035
rect 78703 61972 78712 62012
rect 78752 61972 78769 62012
rect 78855 61972 78876 62012
rect 78916 61972 78937 62012
rect 79023 61972 79040 62012
rect 79080 61972 79089 62012
rect 78703 61949 78769 61972
rect 78855 61949 78937 61972
rect 79023 61949 79089 61972
rect 78703 61930 79089 61949
rect 93823 62035 94209 62054
rect 93823 62012 93889 62035
rect 93975 62012 94057 62035
rect 94143 62012 94209 62035
rect 93823 61972 93832 62012
rect 93872 61972 93889 62012
rect 93975 61972 93996 62012
rect 94036 61972 94057 62012
rect 94143 61972 94160 62012
rect 94200 61972 94209 62012
rect 93823 61949 93889 61972
rect 93975 61949 94057 61972
rect 94143 61949 94209 61972
rect 93823 61930 94209 61949
rect 4343 61279 4729 61298
rect 4343 61256 4409 61279
rect 4495 61256 4577 61279
rect 4663 61256 4729 61279
rect 4343 61216 4352 61256
rect 4392 61216 4409 61256
rect 4495 61216 4516 61256
rect 4556 61216 4577 61256
rect 4663 61216 4680 61256
rect 4720 61216 4729 61256
rect 4343 61193 4409 61216
rect 4495 61193 4577 61216
rect 4663 61193 4729 61216
rect 4343 61174 4729 61193
rect 19463 61279 19849 61298
rect 19463 61256 19529 61279
rect 19615 61256 19697 61279
rect 19783 61256 19849 61279
rect 19463 61216 19472 61256
rect 19512 61216 19529 61256
rect 19615 61216 19636 61256
rect 19676 61216 19697 61256
rect 19783 61216 19800 61256
rect 19840 61216 19849 61256
rect 19463 61193 19529 61216
rect 19615 61193 19697 61216
rect 19783 61193 19849 61216
rect 19463 61174 19849 61193
rect 34583 61279 34969 61298
rect 34583 61256 34649 61279
rect 34735 61256 34817 61279
rect 34903 61256 34969 61279
rect 34583 61216 34592 61256
rect 34632 61216 34649 61256
rect 34735 61216 34756 61256
rect 34796 61216 34817 61256
rect 34903 61216 34920 61256
rect 34960 61216 34969 61256
rect 34583 61193 34649 61216
rect 34735 61193 34817 61216
rect 34903 61193 34969 61216
rect 34583 61174 34969 61193
rect 49703 61279 50089 61298
rect 49703 61256 49769 61279
rect 49855 61256 49937 61279
rect 50023 61256 50089 61279
rect 49703 61216 49712 61256
rect 49752 61216 49769 61256
rect 49855 61216 49876 61256
rect 49916 61216 49937 61256
rect 50023 61216 50040 61256
rect 50080 61216 50089 61256
rect 49703 61193 49769 61216
rect 49855 61193 49937 61216
rect 50023 61193 50089 61216
rect 49703 61174 50089 61193
rect 64823 61279 65209 61298
rect 64823 61256 64889 61279
rect 64975 61256 65057 61279
rect 65143 61256 65209 61279
rect 64823 61216 64832 61256
rect 64872 61216 64889 61256
rect 64975 61216 64996 61256
rect 65036 61216 65057 61256
rect 65143 61216 65160 61256
rect 65200 61216 65209 61256
rect 64823 61193 64889 61216
rect 64975 61193 65057 61216
rect 65143 61193 65209 61216
rect 64823 61174 65209 61193
rect 79943 61279 80329 61298
rect 79943 61256 80009 61279
rect 80095 61256 80177 61279
rect 80263 61256 80329 61279
rect 79943 61216 79952 61256
rect 79992 61216 80009 61256
rect 80095 61216 80116 61256
rect 80156 61216 80177 61256
rect 80263 61216 80280 61256
rect 80320 61216 80329 61256
rect 79943 61193 80009 61216
rect 80095 61193 80177 61216
rect 80263 61193 80329 61216
rect 79943 61174 80329 61193
rect 95063 61279 95449 61298
rect 95063 61256 95129 61279
rect 95215 61256 95297 61279
rect 95383 61256 95449 61279
rect 95063 61216 95072 61256
rect 95112 61216 95129 61256
rect 95215 61216 95236 61256
rect 95276 61216 95297 61256
rect 95383 61216 95400 61256
rect 95440 61216 95449 61256
rect 95063 61193 95129 61216
rect 95215 61193 95297 61216
rect 95383 61193 95449 61216
rect 95063 61174 95449 61193
rect 3103 60523 3489 60542
rect 3103 60500 3169 60523
rect 3255 60500 3337 60523
rect 3423 60500 3489 60523
rect 3103 60460 3112 60500
rect 3152 60460 3169 60500
rect 3255 60460 3276 60500
rect 3316 60460 3337 60500
rect 3423 60460 3440 60500
rect 3480 60460 3489 60500
rect 3103 60437 3169 60460
rect 3255 60437 3337 60460
rect 3423 60437 3489 60460
rect 3103 60418 3489 60437
rect 18223 60523 18609 60542
rect 18223 60500 18289 60523
rect 18375 60500 18457 60523
rect 18543 60500 18609 60523
rect 18223 60460 18232 60500
rect 18272 60460 18289 60500
rect 18375 60460 18396 60500
rect 18436 60460 18457 60500
rect 18543 60460 18560 60500
rect 18600 60460 18609 60500
rect 18223 60437 18289 60460
rect 18375 60437 18457 60460
rect 18543 60437 18609 60460
rect 18223 60418 18609 60437
rect 33343 60523 33729 60542
rect 33343 60500 33409 60523
rect 33495 60500 33577 60523
rect 33663 60500 33729 60523
rect 33343 60460 33352 60500
rect 33392 60460 33409 60500
rect 33495 60460 33516 60500
rect 33556 60460 33577 60500
rect 33663 60460 33680 60500
rect 33720 60460 33729 60500
rect 33343 60437 33409 60460
rect 33495 60437 33577 60460
rect 33663 60437 33729 60460
rect 33343 60418 33729 60437
rect 48463 60523 48849 60542
rect 48463 60500 48529 60523
rect 48615 60500 48697 60523
rect 48783 60500 48849 60523
rect 48463 60460 48472 60500
rect 48512 60460 48529 60500
rect 48615 60460 48636 60500
rect 48676 60460 48697 60500
rect 48783 60460 48800 60500
rect 48840 60460 48849 60500
rect 48463 60437 48529 60460
rect 48615 60437 48697 60460
rect 48783 60437 48849 60460
rect 48463 60418 48849 60437
rect 63583 60523 63969 60542
rect 63583 60500 63649 60523
rect 63735 60500 63817 60523
rect 63903 60500 63969 60523
rect 63583 60460 63592 60500
rect 63632 60460 63649 60500
rect 63735 60460 63756 60500
rect 63796 60460 63817 60500
rect 63903 60460 63920 60500
rect 63960 60460 63969 60500
rect 63583 60437 63649 60460
rect 63735 60437 63817 60460
rect 63903 60437 63969 60460
rect 63583 60418 63969 60437
rect 78703 60523 79089 60542
rect 78703 60500 78769 60523
rect 78855 60500 78937 60523
rect 79023 60500 79089 60523
rect 78703 60460 78712 60500
rect 78752 60460 78769 60500
rect 78855 60460 78876 60500
rect 78916 60460 78937 60500
rect 79023 60460 79040 60500
rect 79080 60460 79089 60500
rect 78703 60437 78769 60460
rect 78855 60437 78937 60460
rect 79023 60437 79089 60460
rect 78703 60418 79089 60437
rect 93823 60523 94209 60542
rect 93823 60500 93889 60523
rect 93975 60500 94057 60523
rect 94143 60500 94209 60523
rect 93823 60460 93832 60500
rect 93872 60460 93889 60500
rect 93975 60460 93996 60500
rect 94036 60460 94057 60500
rect 94143 60460 94160 60500
rect 94200 60460 94209 60500
rect 93823 60437 93889 60460
rect 93975 60437 94057 60460
rect 94143 60437 94209 60460
rect 93823 60418 94209 60437
rect 4343 59767 4729 59786
rect 4343 59744 4409 59767
rect 4495 59744 4577 59767
rect 4663 59744 4729 59767
rect 4343 59704 4352 59744
rect 4392 59704 4409 59744
rect 4495 59704 4516 59744
rect 4556 59704 4577 59744
rect 4663 59704 4680 59744
rect 4720 59704 4729 59744
rect 4343 59681 4409 59704
rect 4495 59681 4577 59704
rect 4663 59681 4729 59704
rect 4343 59662 4729 59681
rect 19463 59767 19849 59786
rect 19463 59744 19529 59767
rect 19615 59744 19697 59767
rect 19783 59744 19849 59767
rect 19463 59704 19472 59744
rect 19512 59704 19529 59744
rect 19615 59704 19636 59744
rect 19676 59704 19697 59744
rect 19783 59704 19800 59744
rect 19840 59704 19849 59744
rect 19463 59681 19529 59704
rect 19615 59681 19697 59704
rect 19783 59681 19849 59704
rect 19463 59662 19849 59681
rect 34583 59767 34969 59786
rect 34583 59744 34649 59767
rect 34735 59744 34817 59767
rect 34903 59744 34969 59767
rect 34583 59704 34592 59744
rect 34632 59704 34649 59744
rect 34735 59704 34756 59744
rect 34796 59704 34817 59744
rect 34903 59704 34920 59744
rect 34960 59704 34969 59744
rect 34583 59681 34649 59704
rect 34735 59681 34817 59704
rect 34903 59681 34969 59704
rect 34583 59662 34969 59681
rect 49703 59767 50089 59786
rect 49703 59744 49769 59767
rect 49855 59744 49937 59767
rect 50023 59744 50089 59767
rect 49703 59704 49712 59744
rect 49752 59704 49769 59744
rect 49855 59704 49876 59744
rect 49916 59704 49937 59744
rect 50023 59704 50040 59744
rect 50080 59704 50089 59744
rect 49703 59681 49769 59704
rect 49855 59681 49937 59704
rect 50023 59681 50089 59704
rect 49703 59662 50089 59681
rect 64823 59767 65209 59786
rect 64823 59744 64889 59767
rect 64975 59744 65057 59767
rect 65143 59744 65209 59767
rect 64823 59704 64832 59744
rect 64872 59704 64889 59744
rect 64975 59704 64996 59744
rect 65036 59704 65057 59744
rect 65143 59704 65160 59744
rect 65200 59704 65209 59744
rect 64823 59681 64889 59704
rect 64975 59681 65057 59704
rect 65143 59681 65209 59704
rect 64823 59662 65209 59681
rect 79943 59767 80329 59786
rect 79943 59744 80009 59767
rect 80095 59744 80177 59767
rect 80263 59744 80329 59767
rect 79943 59704 79952 59744
rect 79992 59704 80009 59744
rect 80095 59704 80116 59744
rect 80156 59704 80177 59744
rect 80263 59704 80280 59744
rect 80320 59704 80329 59744
rect 79943 59681 80009 59704
rect 80095 59681 80177 59704
rect 80263 59681 80329 59704
rect 79943 59662 80329 59681
rect 95063 59767 95449 59786
rect 95063 59744 95129 59767
rect 95215 59744 95297 59767
rect 95383 59744 95449 59767
rect 95063 59704 95072 59744
rect 95112 59704 95129 59744
rect 95215 59704 95236 59744
rect 95276 59704 95297 59744
rect 95383 59704 95400 59744
rect 95440 59704 95449 59744
rect 95063 59681 95129 59704
rect 95215 59681 95297 59704
rect 95383 59681 95449 59704
rect 95063 59662 95449 59681
rect 3103 59011 3489 59030
rect 3103 58988 3169 59011
rect 3255 58988 3337 59011
rect 3423 58988 3489 59011
rect 3103 58948 3112 58988
rect 3152 58948 3169 58988
rect 3255 58948 3276 58988
rect 3316 58948 3337 58988
rect 3423 58948 3440 58988
rect 3480 58948 3489 58988
rect 3103 58925 3169 58948
rect 3255 58925 3337 58948
rect 3423 58925 3489 58948
rect 3103 58906 3489 58925
rect 18223 59011 18609 59030
rect 18223 58988 18289 59011
rect 18375 58988 18457 59011
rect 18543 58988 18609 59011
rect 18223 58948 18232 58988
rect 18272 58948 18289 58988
rect 18375 58948 18396 58988
rect 18436 58948 18457 58988
rect 18543 58948 18560 58988
rect 18600 58948 18609 58988
rect 18223 58925 18289 58948
rect 18375 58925 18457 58948
rect 18543 58925 18609 58948
rect 18223 58906 18609 58925
rect 33343 59011 33729 59030
rect 33343 58988 33409 59011
rect 33495 58988 33577 59011
rect 33663 58988 33729 59011
rect 33343 58948 33352 58988
rect 33392 58948 33409 58988
rect 33495 58948 33516 58988
rect 33556 58948 33577 58988
rect 33663 58948 33680 58988
rect 33720 58948 33729 58988
rect 33343 58925 33409 58948
rect 33495 58925 33577 58948
rect 33663 58925 33729 58948
rect 33343 58906 33729 58925
rect 48463 59011 48849 59030
rect 48463 58988 48529 59011
rect 48615 58988 48697 59011
rect 48783 58988 48849 59011
rect 48463 58948 48472 58988
rect 48512 58948 48529 58988
rect 48615 58948 48636 58988
rect 48676 58948 48697 58988
rect 48783 58948 48800 58988
rect 48840 58948 48849 58988
rect 48463 58925 48529 58948
rect 48615 58925 48697 58948
rect 48783 58925 48849 58948
rect 48463 58906 48849 58925
rect 63583 59011 63969 59030
rect 63583 58988 63649 59011
rect 63735 58988 63817 59011
rect 63903 58988 63969 59011
rect 63583 58948 63592 58988
rect 63632 58948 63649 58988
rect 63735 58948 63756 58988
rect 63796 58948 63817 58988
rect 63903 58948 63920 58988
rect 63960 58948 63969 58988
rect 63583 58925 63649 58948
rect 63735 58925 63817 58948
rect 63903 58925 63969 58948
rect 63583 58906 63969 58925
rect 78703 59011 79089 59030
rect 78703 58988 78769 59011
rect 78855 58988 78937 59011
rect 79023 58988 79089 59011
rect 78703 58948 78712 58988
rect 78752 58948 78769 58988
rect 78855 58948 78876 58988
rect 78916 58948 78937 58988
rect 79023 58948 79040 58988
rect 79080 58948 79089 58988
rect 78703 58925 78769 58948
rect 78855 58925 78937 58948
rect 79023 58925 79089 58948
rect 78703 58906 79089 58925
rect 93823 59011 94209 59030
rect 93823 58988 93889 59011
rect 93975 58988 94057 59011
rect 94143 58988 94209 59011
rect 93823 58948 93832 58988
rect 93872 58948 93889 58988
rect 93975 58948 93996 58988
rect 94036 58948 94057 58988
rect 94143 58948 94160 58988
rect 94200 58948 94209 58988
rect 93823 58925 93889 58948
rect 93975 58925 94057 58948
rect 94143 58925 94209 58948
rect 93823 58906 94209 58925
rect 4343 58255 4729 58274
rect 4343 58232 4409 58255
rect 4495 58232 4577 58255
rect 4663 58232 4729 58255
rect 4343 58192 4352 58232
rect 4392 58192 4409 58232
rect 4495 58192 4516 58232
rect 4556 58192 4577 58232
rect 4663 58192 4680 58232
rect 4720 58192 4729 58232
rect 4343 58169 4409 58192
rect 4495 58169 4577 58192
rect 4663 58169 4729 58192
rect 4343 58150 4729 58169
rect 19463 58255 19849 58274
rect 19463 58232 19529 58255
rect 19615 58232 19697 58255
rect 19783 58232 19849 58255
rect 19463 58192 19472 58232
rect 19512 58192 19529 58232
rect 19615 58192 19636 58232
rect 19676 58192 19697 58232
rect 19783 58192 19800 58232
rect 19840 58192 19849 58232
rect 19463 58169 19529 58192
rect 19615 58169 19697 58192
rect 19783 58169 19849 58192
rect 19463 58150 19849 58169
rect 34583 58255 34969 58274
rect 34583 58232 34649 58255
rect 34735 58232 34817 58255
rect 34903 58232 34969 58255
rect 34583 58192 34592 58232
rect 34632 58192 34649 58232
rect 34735 58192 34756 58232
rect 34796 58192 34817 58232
rect 34903 58192 34920 58232
rect 34960 58192 34969 58232
rect 34583 58169 34649 58192
rect 34735 58169 34817 58192
rect 34903 58169 34969 58192
rect 34583 58150 34969 58169
rect 49703 58255 50089 58274
rect 49703 58232 49769 58255
rect 49855 58232 49937 58255
rect 50023 58232 50089 58255
rect 49703 58192 49712 58232
rect 49752 58192 49769 58232
rect 49855 58192 49876 58232
rect 49916 58192 49937 58232
rect 50023 58192 50040 58232
rect 50080 58192 50089 58232
rect 49703 58169 49769 58192
rect 49855 58169 49937 58192
rect 50023 58169 50089 58192
rect 49703 58150 50089 58169
rect 64823 58255 65209 58274
rect 64823 58232 64889 58255
rect 64975 58232 65057 58255
rect 65143 58232 65209 58255
rect 64823 58192 64832 58232
rect 64872 58192 64889 58232
rect 64975 58192 64996 58232
rect 65036 58192 65057 58232
rect 65143 58192 65160 58232
rect 65200 58192 65209 58232
rect 64823 58169 64889 58192
rect 64975 58169 65057 58192
rect 65143 58169 65209 58192
rect 64823 58150 65209 58169
rect 79943 58255 80329 58274
rect 79943 58232 80009 58255
rect 80095 58232 80177 58255
rect 80263 58232 80329 58255
rect 79943 58192 79952 58232
rect 79992 58192 80009 58232
rect 80095 58192 80116 58232
rect 80156 58192 80177 58232
rect 80263 58192 80280 58232
rect 80320 58192 80329 58232
rect 79943 58169 80009 58192
rect 80095 58169 80177 58192
rect 80263 58169 80329 58192
rect 79943 58150 80329 58169
rect 95063 58255 95449 58274
rect 95063 58232 95129 58255
rect 95215 58232 95297 58255
rect 95383 58232 95449 58255
rect 95063 58192 95072 58232
rect 95112 58192 95129 58232
rect 95215 58192 95236 58232
rect 95276 58192 95297 58232
rect 95383 58192 95400 58232
rect 95440 58192 95449 58232
rect 95063 58169 95129 58192
rect 95215 58169 95297 58192
rect 95383 58169 95449 58192
rect 95063 58150 95449 58169
rect 3103 57499 3489 57518
rect 3103 57476 3169 57499
rect 3255 57476 3337 57499
rect 3423 57476 3489 57499
rect 3103 57436 3112 57476
rect 3152 57436 3169 57476
rect 3255 57436 3276 57476
rect 3316 57436 3337 57476
rect 3423 57436 3440 57476
rect 3480 57436 3489 57476
rect 3103 57413 3169 57436
rect 3255 57413 3337 57436
rect 3423 57413 3489 57436
rect 3103 57394 3489 57413
rect 18223 57499 18609 57518
rect 18223 57476 18289 57499
rect 18375 57476 18457 57499
rect 18543 57476 18609 57499
rect 18223 57436 18232 57476
rect 18272 57436 18289 57476
rect 18375 57436 18396 57476
rect 18436 57436 18457 57476
rect 18543 57436 18560 57476
rect 18600 57436 18609 57476
rect 18223 57413 18289 57436
rect 18375 57413 18457 57436
rect 18543 57413 18609 57436
rect 18223 57394 18609 57413
rect 33343 57499 33729 57518
rect 33343 57476 33409 57499
rect 33495 57476 33577 57499
rect 33663 57476 33729 57499
rect 33343 57436 33352 57476
rect 33392 57436 33409 57476
rect 33495 57436 33516 57476
rect 33556 57436 33577 57476
rect 33663 57436 33680 57476
rect 33720 57436 33729 57476
rect 33343 57413 33409 57436
rect 33495 57413 33577 57436
rect 33663 57413 33729 57436
rect 33343 57394 33729 57413
rect 48463 57499 48849 57518
rect 48463 57476 48529 57499
rect 48615 57476 48697 57499
rect 48783 57476 48849 57499
rect 48463 57436 48472 57476
rect 48512 57436 48529 57476
rect 48615 57436 48636 57476
rect 48676 57436 48697 57476
rect 48783 57436 48800 57476
rect 48840 57436 48849 57476
rect 48463 57413 48529 57436
rect 48615 57413 48697 57436
rect 48783 57413 48849 57436
rect 48463 57394 48849 57413
rect 63583 57499 63969 57518
rect 63583 57476 63649 57499
rect 63735 57476 63817 57499
rect 63903 57476 63969 57499
rect 63583 57436 63592 57476
rect 63632 57436 63649 57476
rect 63735 57436 63756 57476
rect 63796 57436 63817 57476
rect 63903 57436 63920 57476
rect 63960 57436 63969 57476
rect 63583 57413 63649 57436
rect 63735 57413 63817 57436
rect 63903 57413 63969 57436
rect 63583 57394 63969 57413
rect 78703 57499 79089 57518
rect 78703 57476 78769 57499
rect 78855 57476 78937 57499
rect 79023 57476 79089 57499
rect 78703 57436 78712 57476
rect 78752 57436 78769 57476
rect 78855 57436 78876 57476
rect 78916 57436 78937 57476
rect 79023 57436 79040 57476
rect 79080 57436 79089 57476
rect 78703 57413 78769 57436
rect 78855 57413 78937 57436
rect 79023 57413 79089 57436
rect 78703 57394 79089 57413
rect 93823 57499 94209 57518
rect 93823 57476 93889 57499
rect 93975 57476 94057 57499
rect 94143 57476 94209 57499
rect 93823 57436 93832 57476
rect 93872 57436 93889 57476
rect 93975 57436 93996 57476
rect 94036 57436 94057 57476
rect 94143 57436 94160 57476
rect 94200 57436 94209 57476
rect 93823 57413 93889 57436
rect 93975 57413 94057 57436
rect 94143 57413 94209 57436
rect 93823 57394 94209 57413
rect 4343 56743 4729 56762
rect 4343 56720 4409 56743
rect 4495 56720 4577 56743
rect 4663 56720 4729 56743
rect 4343 56680 4352 56720
rect 4392 56680 4409 56720
rect 4495 56680 4516 56720
rect 4556 56680 4577 56720
rect 4663 56680 4680 56720
rect 4720 56680 4729 56720
rect 4343 56657 4409 56680
rect 4495 56657 4577 56680
rect 4663 56657 4729 56680
rect 4343 56638 4729 56657
rect 19463 56743 19849 56762
rect 19463 56720 19529 56743
rect 19615 56720 19697 56743
rect 19783 56720 19849 56743
rect 19463 56680 19472 56720
rect 19512 56680 19529 56720
rect 19615 56680 19636 56720
rect 19676 56680 19697 56720
rect 19783 56680 19800 56720
rect 19840 56680 19849 56720
rect 19463 56657 19529 56680
rect 19615 56657 19697 56680
rect 19783 56657 19849 56680
rect 19463 56638 19849 56657
rect 34583 56743 34969 56762
rect 34583 56720 34649 56743
rect 34735 56720 34817 56743
rect 34903 56720 34969 56743
rect 34583 56680 34592 56720
rect 34632 56680 34649 56720
rect 34735 56680 34756 56720
rect 34796 56680 34817 56720
rect 34903 56680 34920 56720
rect 34960 56680 34969 56720
rect 34583 56657 34649 56680
rect 34735 56657 34817 56680
rect 34903 56657 34969 56680
rect 34583 56638 34969 56657
rect 49703 56743 50089 56762
rect 49703 56720 49769 56743
rect 49855 56720 49937 56743
rect 50023 56720 50089 56743
rect 49703 56680 49712 56720
rect 49752 56680 49769 56720
rect 49855 56680 49876 56720
rect 49916 56680 49937 56720
rect 50023 56680 50040 56720
rect 50080 56680 50089 56720
rect 49703 56657 49769 56680
rect 49855 56657 49937 56680
rect 50023 56657 50089 56680
rect 49703 56638 50089 56657
rect 64823 56743 65209 56762
rect 64823 56720 64889 56743
rect 64975 56720 65057 56743
rect 65143 56720 65209 56743
rect 64823 56680 64832 56720
rect 64872 56680 64889 56720
rect 64975 56680 64996 56720
rect 65036 56680 65057 56720
rect 65143 56680 65160 56720
rect 65200 56680 65209 56720
rect 64823 56657 64889 56680
rect 64975 56657 65057 56680
rect 65143 56657 65209 56680
rect 64823 56638 65209 56657
rect 79943 56743 80329 56762
rect 79943 56720 80009 56743
rect 80095 56720 80177 56743
rect 80263 56720 80329 56743
rect 79943 56680 79952 56720
rect 79992 56680 80009 56720
rect 80095 56680 80116 56720
rect 80156 56680 80177 56720
rect 80263 56680 80280 56720
rect 80320 56680 80329 56720
rect 79943 56657 80009 56680
rect 80095 56657 80177 56680
rect 80263 56657 80329 56680
rect 79943 56638 80329 56657
rect 95063 56743 95449 56762
rect 95063 56720 95129 56743
rect 95215 56720 95297 56743
rect 95383 56720 95449 56743
rect 95063 56680 95072 56720
rect 95112 56680 95129 56720
rect 95215 56680 95236 56720
rect 95276 56680 95297 56720
rect 95383 56680 95400 56720
rect 95440 56680 95449 56720
rect 95063 56657 95129 56680
rect 95215 56657 95297 56680
rect 95383 56657 95449 56680
rect 95063 56638 95449 56657
rect 3103 55987 3489 56006
rect 3103 55964 3169 55987
rect 3255 55964 3337 55987
rect 3423 55964 3489 55987
rect 3103 55924 3112 55964
rect 3152 55924 3169 55964
rect 3255 55924 3276 55964
rect 3316 55924 3337 55964
rect 3423 55924 3440 55964
rect 3480 55924 3489 55964
rect 3103 55901 3169 55924
rect 3255 55901 3337 55924
rect 3423 55901 3489 55924
rect 3103 55882 3489 55901
rect 18223 55987 18609 56006
rect 18223 55964 18289 55987
rect 18375 55964 18457 55987
rect 18543 55964 18609 55987
rect 18223 55924 18232 55964
rect 18272 55924 18289 55964
rect 18375 55924 18396 55964
rect 18436 55924 18457 55964
rect 18543 55924 18560 55964
rect 18600 55924 18609 55964
rect 18223 55901 18289 55924
rect 18375 55901 18457 55924
rect 18543 55901 18609 55924
rect 18223 55882 18609 55901
rect 33343 55987 33729 56006
rect 33343 55964 33409 55987
rect 33495 55964 33577 55987
rect 33663 55964 33729 55987
rect 33343 55924 33352 55964
rect 33392 55924 33409 55964
rect 33495 55924 33516 55964
rect 33556 55924 33577 55964
rect 33663 55924 33680 55964
rect 33720 55924 33729 55964
rect 33343 55901 33409 55924
rect 33495 55901 33577 55924
rect 33663 55901 33729 55924
rect 33343 55882 33729 55901
rect 48463 55987 48849 56006
rect 48463 55964 48529 55987
rect 48615 55964 48697 55987
rect 48783 55964 48849 55987
rect 48463 55924 48472 55964
rect 48512 55924 48529 55964
rect 48615 55924 48636 55964
rect 48676 55924 48697 55964
rect 48783 55924 48800 55964
rect 48840 55924 48849 55964
rect 48463 55901 48529 55924
rect 48615 55901 48697 55924
rect 48783 55901 48849 55924
rect 48463 55882 48849 55901
rect 63583 55987 63969 56006
rect 63583 55964 63649 55987
rect 63735 55964 63817 55987
rect 63903 55964 63969 55987
rect 63583 55924 63592 55964
rect 63632 55924 63649 55964
rect 63735 55924 63756 55964
rect 63796 55924 63817 55964
rect 63903 55924 63920 55964
rect 63960 55924 63969 55964
rect 63583 55901 63649 55924
rect 63735 55901 63817 55924
rect 63903 55901 63969 55924
rect 63583 55882 63969 55901
rect 78703 55987 79089 56006
rect 78703 55964 78769 55987
rect 78855 55964 78937 55987
rect 79023 55964 79089 55987
rect 78703 55924 78712 55964
rect 78752 55924 78769 55964
rect 78855 55924 78876 55964
rect 78916 55924 78937 55964
rect 79023 55924 79040 55964
rect 79080 55924 79089 55964
rect 78703 55901 78769 55924
rect 78855 55901 78937 55924
rect 79023 55901 79089 55924
rect 78703 55882 79089 55901
rect 93823 55987 94209 56006
rect 93823 55964 93889 55987
rect 93975 55964 94057 55987
rect 94143 55964 94209 55987
rect 93823 55924 93832 55964
rect 93872 55924 93889 55964
rect 93975 55924 93996 55964
rect 94036 55924 94057 55964
rect 94143 55924 94160 55964
rect 94200 55924 94209 55964
rect 93823 55901 93889 55924
rect 93975 55901 94057 55924
rect 94143 55901 94209 55924
rect 93823 55882 94209 55901
rect 4343 55231 4729 55250
rect 4343 55208 4409 55231
rect 4495 55208 4577 55231
rect 4663 55208 4729 55231
rect 4343 55168 4352 55208
rect 4392 55168 4409 55208
rect 4495 55168 4516 55208
rect 4556 55168 4577 55208
rect 4663 55168 4680 55208
rect 4720 55168 4729 55208
rect 4343 55145 4409 55168
rect 4495 55145 4577 55168
rect 4663 55145 4729 55168
rect 4343 55126 4729 55145
rect 19463 55231 19849 55250
rect 19463 55208 19529 55231
rect 19615 55208 19697 55231
rect 19783 55208 19849 55231
rect 19463 55168 19472 55208
rect 19512 55168 19529 55208
rect 19615 55168 19636 55208
rect 19676 55168 19697 55208
rect 19783 55168 19800 55208
rect 19840 55168 19849 55208
rect 19463 55145 19529 55168
rect 19615 55145 19697 55168
rect 19783 55145 19849 55168
rect 19463 55126 19849 55145
rect 34583 55231 34969 55250
rect 34583 55208 34649 55231
rect 34735 55208 34817 55231
rect 34903 55208 34969 55231
rect 34583 55168 34592 55208
rect 34632 55168 34649 55208
rect 34735 55168 34756 55208
rect 34796 55168 34817 55208
rect 34903 55168 34920 55208
rect 34960 55168 34969 55208
rect 34583 55145 34649 55168
rect 34735 55145 34817 55168
rect 34903 55145 34969 55168
rect 34583 55126 34969 55145
rect 49703 55231 50089 55250
rect 49703 55208 49769 55231
rect 49855 55208 49937 55231
rect 50023 55208 50089 55231
rect 49703 55168 49712 55208
rect 49752 55168 49769 55208
rect 49855 55168 49876 55208
rect 49916 55168 49937 55208
rect 50023 55168 50040 55208
rect 50080 55168 50089 55208
rect 49703 55145 49769 55168
rect 49855 55145 49937 55168
rect 50023 55145 50089 55168
rect 49703 55126 50089 55145
rect 64823 55231 65209 55250
rect 64823 55208 64889 55231
rect 64975 55208 65057 55231
rect 65143 55208 65209 55231
rect 64823 55168 64832 55208
rect 64872 55168 64889 55208
rect 64975 55168 64996 55208
rect 65036 55168 65057 55208
rect 65143 55168 65160 55208
rect 65200 55168 65209 55208
rect 64823 55145 64889 55168
rect 64975 55145 65057 55168
rect 65143 55145 65209 55168
rect 64823 55126 65209 55145
rect 79943 55231 80329 55250
rect 79943 55208 80009 55231
rect 80095 55208 80177 55231
rect 80263 55208 80329 55231
rect 79943 55168 79952 55208
rect 79992 55168 80009 55208
rect 80095 55168 80116 55208
rect 80156 55168 80177 55208
rect 80263 55168 80280 55208
rect 80320 55168 80329 55208
rect 79943 55145 80009 55168
rect 80095 55145 80177 55168
rect 80263 55145 80329 55168
rect 79943 55126 80329 55145
rect 95063 55231 95449 55250
rect 95063 55208 95129 55231
rect 95215 55208 95297 55231
rect 95383 55208 95449 55231
rect 95063 55168 95072 55208
rect 95112 55168 95129 55208
rect 95215 55168 95236 55208
rect 95276 55168 95297 55208
rect 95383 55168 95400 55208
rect 95440 55168 95449 55208
rect 95063 55145 95129 55168
rect 95215 55145 95297 55168
rect 95383 55145 95449 55168
rect 95063 55126 95449 55145
rect 3103 54475 3489 54494
rect 3103 54452 3169 54475
rect 3255 54452 3337 54475
rect 3423 54452 3489 54475
rect 3103 54412 3112 54452
rect 3152 54412 3169 54452
rect 3255 54412 3276 54452
rect 3316 54412 3337 54452
rect 3423 54412 3440 54452
rect 3480 54412 3489 54452
rect 3103 54389 3169 54412
rect 3255 54389 3337 54412
rect 3423 54389 3489 54412
rect 3103 54370 3489 54389
rect 18223 54475 18609 54494
rect 18223 54452 18289 54475
rect 18375 54452 18457 54475
rect 18543 54452 18609 54475
rect 18223 54412 18232 54452
rect 18272 54412 18289 54452
rect 18375 54412 18396 54452
rect 18436 54412 18457 54452
rect 18543 54412 18560 54452
rect 18600 54412 18609 54452
rect 18223 54389 18289 54412
rect 18375 54389 18457 54412
rect 18543 54389 18609 54412
rect 18223 54370 18609 54389
rect 33343 54475 33729 54494
rect 33343 54452 33409 54475
rect 33495 54452 33577 54475
rect 33663 54452 33729 54475
rect 33343 54412 33352 54452
rect 33392 54412 33409 54452
rect 33495 54412 33516 54452
rect 33556 54412 33577 54452
rect 33663 54412 33680 54452
rect 33720 54412 33729 54452
rect 33343 54389 33409 54412
rect 33495 54389 33577 54412
rect 33663 54389 33729 54412
rect 33343 54370 33729 54389
rect 48463 54475 48849 54494
rect 48463 54452 48529 54475
rect 48615 54452 48697 54475
rect 48783 54452 48849 54475
rect 48463 54412 48472 54452
rect 48512 54412 48529 54452
rect 48615 54412 48636 54452
rect 48676 54412 48697 54452
rect 48783 54412 48800 54452
rect 48840 54412 48849 54452
rect 48463 54389 48529 54412
rect 48615 54389 48697 54412
rect 48783 54389 48849 54412
rect 48463 54370 48849 54389
rect 63583 54475 63969 54494
rect 63583 54452 63649 54475
rect 63735 54452 63817 54475
rect 63903 54452 63969 54475
rect 63583 54412 63592 54452
rect 63632 54412 63649 54452
rect 63735 54412 63756 54452
rect 63796 54412 63817 54452
rect 63903 54412 63920 54452
rect 63960 54412 63969 54452
rect 63583 54389 63649 54412
rect 63735 54389 63817 54412
rect 63903 54389 63969 54412
rect 63583 54370 63969 54389
rect 78703 54475 79089 54494
rect 78703 54452 78769 54475
rect 78855 54452 78937 54475
rect 79023 54452 79089 54475
rect 78703 54412 78712 54452
rect 78752 54412 78769 54452
rect 78855 54412 78876 54452
rect 78916 54412 78937 54452
rect 79023 54412 79040 54452
rect 79080 54412 79089 54452
rect 78703 54389 78769 54412
rect 78855 54389 78937 54412
rect 79023 54389 79089 54412
rect 78703 54370 79089 54389
rect 93823 54475 94209 54494
rect 93823 54452 93889 54475
rect 93975 54452 94057 54475
rect 94143 54452 94209 54475
rect 93823 54412 93832 54452
rect 93872 54412 93889 54452
rect 93975 54412 93996 54452
rect 94036 54412 94057 54452
rect 94143 54412 94160 54452
rect 94200 54412 94209 54452
rect 93823 54389 93889 54412
rect 93975 54389 94057 54412
rect 94143 54389 94209 54412
rect 93823 54370 94209 54389
rect 4343 53719 4729 53738
rect 4343 53696 4409 53719
rect 4495 53696 4577 53719
rect 4663 53696 4729 53719
rect 4343 53656 4352 53696
rect 4392 53656 4409 53696
rect 4495 53656 4516 53696
rect 4556 53656 4577 53696
rect 4663 53656 4680 53696
rect 4720 53656 4729 53696
rect 4343 53633 4409 53656
rect 4495 53633 4577 53656
rect 4663 53633 4729 53656
rect 4343 53614 4729 53633
rect 19463 53719 19849 53738
rect 19463 53696 19529 53719
rect 19615 53696 19697 53719
rect 19783 53696 19849 53719
rect 19463 53656 19472 53696
rect 19512 53656 19529 53696
rect 19615 53656 19636 53696
rect 19676 53656 19697 53696
rect 19783 53656 19800 53696
rect 19840 53656 19849 53696
rect 19463 53633 19529 53656
rect 19615 53633 19697 53656
rect 19783 53633 19849 53656
rect 19463 53614 19849 53633
rect 34583 53719 34969 53738
rect 34583 53696 34649 53719
rect 34735 53696 34817 53719
rect 34903 53696 34969 53719
rect 34583 53656 34592 53696
rect 34632 53656 34649 53696
rect 34735 53656 34756 53696
rect 34796 53656 34817 53696
rect 34903 53656 34920 53696
rect 34960 53656 34969 53696
rect 34583 53633 34649 53656
rect 34735 53633 34817 53656
rect 34903 53633 34969 53656
rect 34583 53614 34969 53633
rect 49703 53719 50089 53738
rect 49703 53696 49769 53719
rect 49855 53696 49937 53719
rect 50023 53696 50089 53719
rect 49703 53656 49712 53696
rect 49752 53656 49769 53696
rect 49855 53656 49876 53696
rect 49916 53656 49937 53696
rect 50023 53656 50040 53696
rect 50080 53656 50089 53696
rect 49703 53633 49769 53656
rect 49855 53633 49937 53656
rect 50023 53633 50089 53656
rect 49703 53614 50089 53633
rect 64823 53719 65209 53738
rect 64823 53696 64889 53719
rect 64975 53696 65057 53719
rect 65143 53696 65209 53719
rect 64823 53656 64832 53696
rect 64872 53656 64889 53696
rect 64975 53656 64996 53696
rect 65036 53656 65057 53696
rect 65143 53656 65160 53696
rect 65200 53656 65209 53696
rect 64823 53633 64889 53656
rect 64975 53633 65057 53656
rect 65143 53633 65209 53656
rect 64823 53614 65209 53633
rect 79943 53719 80329 53738
rect 79943 53696 80009 53719
rect 80095 53696 80177 53719
rect 80263 53696 80329 53719
rect 79943 53656 79952 53696
rect 79992 53656 80009 53696
rect 80095 53656 80116 53696
rect 80156 53656 80177 53696
rect 80263 53656 80280 53696
rect 80320 53656 80329 53696
rect 79943 53633 80009 53656
rect 80095 53633 80177 53656
rect 80263 53633 80329 53656
rect 79943 53614 80329 53633
rect 95063 53719 95449 53738
rect 95063 53696 95129 53719
rect 95215 53696 95297 53719
rect 95383 53696 95449 53719
rect 95063 53656 95072 53696
rect 95112 53656 95129 53696
rect 95215 53656 95236 53696
rect 95276 53656 95297 53696
rect 95383 53656 95400 53696
rect 95440 53656 95449 53696
rect 95063 53633 95129 53656
rect 95215 53633 95297 53656
rect 95383 53633 95449 53656
rect 95063 53614 95449 53633
rect 3103 52963 3489 52982
rect 3103 52940 3169 52963
rect 3255 52940 3337 52963
rect 3423 52940 3489 52963
rect 3103 52900 3112 52940
rect 3152 52900 3169 52940
rect 3255 52900 3276 52940
rect 3316 52900 3337 52940
rect 3423 52900 3440 52940
rect 3480 52900 3489 52940
rect 3103 52877 3169 52900
rect 3255 52877 3337 52900
rect 3423 52877 3489 52900
rect 3103 52858 3489 52877
rect 18223 52963 18609 52982
rect 18223 52940 18289 52963
rect 18375 52940 18457 52963
rect 18543 52940 18609 52963
rect 18223 52900 18232 52940
rect 18272 52900 18289 52940
rect 18375 52900 18396 52940
rect 18436 52900 18457 52940
rect 18543 52900 18560 52940
rect 18600 52900 18609 52940
rect 18223 52877 18289 52900
rect 18375 52877 18457 52900
rect 18543 52877 18609 52900
rect 18223 52858 18609 52877
rect 33343 52963 33729 52982
rect 33343 52940 33409 52963
rect 33495 52940 33577 52963
rect 33663 52940 33729 52963
rect 33343 52900 33352 52940
rect 33392 52900 33409 52940
rect 33495 52900 33516 52940
rect 33556 52900 33577 52940
rect 33663 52900 33680 52940
rect 33720 52900 33729 52940
rect 33343 52877 33409 52900
rect 33495 52877 33577 52900
rect 33663 52877 33729 52900
rect 33343 52858 33729 52877
rect 48463 52963 48849 52982
rect 48463 52940 48529 52963
rect 48615 52940 48697 52963
rect 48783 52940 48849 52963
rect 48463 52900 48472 52940
rect 48512 52900 48529 52940
rect 48615 52900 48636 52940
rect 48676 52900 48697 52940
rect 48783 52900 48800 52940
rect 48840 52900 48849 52940
rect 48463 52877 48529 52900
rect 48615 52877 48697 52900
rect 48783 52877 48849 52900
rect 48463 52858 48849 52877
rect 63583 52963 63969 52982
rect 63583 52940 63649 52963
rect 63735 52940 63817 52963
rect 63903 52940 63969 52963
rect 63583 52900 63592 52940
rect 63632 52900 63649 52940
rect 63735 52900 63756 52940
rect 63796 52900 63817 52940
rect 63903 52900 63920 52940
rect 63960 52900 63969 52940
rect 63583 52877 63649 52900
rect 63735 52877 63817 52900
rect 63903 52877 63969 52900
rect 63583 52858 63969 52877
rect 78703 52963 79089 52982
rect 78703 52940 78769 52963
rect 78855 52940 78937 52963
rect 79023 52940 79089 52963
rect 78703 52900 78712 52940
rect 78752 52900 78769 52940
rect 78855 52900 78876 52940
rect 78916 52900 78937 52940
rect 79023 52900 79040 52940
rect 79080 52900 79089 52940
rect 78703 52877 78769 52900
rect 78855 52877 78937 52900
rect 79023 52877 79089 52900
rect 78703 52858 79089 52877
rect 93823 52963 94209 52982
rect 93823 52940 93889 52963
rect 93975 52940 94057 52963
rect 94143 52940 94209 52963
rect 93823 52900 93832 52940
rect 93872 52900 93889 52940
rect 93975 52900 93996 52940
rect 94036 52900 94057 52940
rect 94143 52900 94160 52940
rect 94200 52900 94209 52940
rect 93823 52877 93889 52900
rect 93975 52877 94057 52900
rect 94143 52877 94209 52900
rect 93823 52858 94209 52877
rect 4343 52207 4729 52226
rect 4343 52184 4409 52207
rect 4495 52184 4577 52207
rect 4663 52184 4729 52207
rect 4343 52144 4352 52184
rect 4392 52144 4409 52184
rect 4495 52144 4516 52184
rect 4556 52144 4577 52184
rect 4663 52144 4680 52184
rect 4720 52144 4729 52184
rect 4343 52121 4409 52144
rect 4495 52121 4577 52144
rect 4663 52121 4729 52144
rect 4343 52102 4729 52121
rect 19463 52207 19849 52226
rect 19463 52184 19529 52207
rect 19615 52184 19697 52207
rect 19783 52184 19849 52207
rect 19463 52144 19472 52184
rect 19512 52144 19529 52184
rect 19615 52144 19636 52184
rect 19676 52144 19697 52184
rect 19783 52144 19800 52184
rect 19840 52144 19849 52184
rect 19463 52121 19529 52144
rect 19615 52121 19697 52144
rect 19783 52121 19849 52144
rect 19463 52102 19849 52121
rect 34583 52207 34969 52226
rect 34583 52184 34649 52207
rect 34735 52184 34817 52207
rect 34903 52184 34969 52207
rect 34583 52144 34592 52184
rect 34632 52144 34649 52184
rect 34735 52144 34756 52184
rect 34796 52144 34817 52184
rect 34903 52144 34920 52184
rect 34960 52144 34969 52184
rect 34583 52121 34649 52144
rect 34735 52121 34817 52144
rect 34903 52121 34969 52144
rect 34583 52102 34969 52121
rect 49703 52207 50089 52226
rect 49703 52184 49769 52207
rect 49855 52184 49937 52207
rect 50023 52184 50089 52207
rect 49703 52144 49712 52184
rect 49752 52144 49769 52184
rect 49855 52144 49876 52184
rect 49916 52144 49937 52184
rect 50023 52144 50040 52184
rect 50080 52144 50089 52184
rect 49703 52121 49769 52144
rect 49855 52121 49937 52144
rect 50023 52121 50089 52144
rect 49703 52102 50089 52121
rect 64823 52207 65209 52226
rect 64823 52184 64889 52207
rect 64975 52184 65057 52207
rect 65143 52184 65209 52207
rect 64823 52144 64832 52184
rect 64872 52144 64889 52184
rect 64975 52144 64996 52184
rect 65036 52144 65057 52184
rect 65143 52144 65160 52184
rect 65200 52144 65209 52184
rect 64823 52121 64889 52144
rect 64975 52121 65057 52144
rect 65143 52121 65209 52144
rect 64823 52102 65209 52121
rect 79943 52207 80329 52226
rect 79943 52184 80009 52207
rect 80095 52184 80177 52207
rect 80263 52184 80329 52207
rect 79943 52144 79952 52184
rect 79992 52144 80009 52184
rect 80095 52144 80116 52184
rect 80156 52144 80177 52184
rect 80263 52144 80280 52184
rect 80320 52144 80329 52184
rect 79943 52121 80009 52144
rect 80095 52121 80177 52144
rect 80263 52121 80329 52144
rect 79943 52102 80329 52121
rect 95063 52207 95449 52226
rect 95063 52184 95129 52207
rect 95215 52184 95297 52207
rect 95383 52184 95449 52207
rect 95063 52144 95072 52184
rect 95112 52144 95129 52184
rect 95215 52144 95236 52184
rect 95276 52144 95297 52184
rect 95383 52144 95400 52184
rect 95440 52144 95449 52184
rect 95063 52121 95129 52144
rect 95215 52121 95297 52144
rect 95383 52121 95449 52144
rect 95063 52102 95449 52121
rect 3103 51451 3489 51470
rect 3103 51428 3169 51451
rect 3255 51428 3337 51451
rect 3423 51428 3489 51451
rect 3103 51388 3112 51428
rect 3152 51388 3169 51428
rect 3255 51388 3276 51428
rect 3316 51388 3337 51428
rect 3423 51388 3440 51428
rect 3480 51388 3489 51428
rect 3103 51365 3169 51388
rect 3255 51365 3337 51388
rect 3423 51365 3489 51388
rect 3103 51346 3489 51365
rect 18223 51451 18609 51470
rect 18223 51428 18289 51451
rect 18375 51428 18457 51451
rect 18543 51428 18609 51451
rect 18223 51388 18232 51428
rect 18272 51388 18289 51428
rect 18375 51388 18396 51428
rect 18436 51388 18457 51428
rect 18543 51388 18560 51428
rect 18600 51388 18609 51428
rect 18223 51365 18289 51388
rect 18375 51365 18457 51388
rect 18543 51365 18609 51388
rect 18223 51346 18609 51365
rect 33343 51451 33729 51470
rect 33343 51428 33409 51451
rect 33495 51428 33577 51451
rect 33663 51428 33729 51451
rect 33343 51388 33352 51428
rect 33392 51388 33409 51428
rect 33495 51388 33516 51428
rect 33556 51388 33577 51428
rect 33663 51388 33680 51428
rect 33720 51388 33729 51428
rect 33343 51365 33409 51388
rect 33495 51365 33577 51388
rect 33663 51365 33729 51388
rect 33343 51346 33729 51365
rect 48463 51451 48849 51470
rect 48463 51428 48529 51451
rect 48615 51428 48697 51451
rect 48783 51428 48849 51451
rect 48463 51388 48472 51428
rect 48512 51388 48529 51428
rect 48615 51388 48636 51428
rect 48676 51388 48697 51428
rect 48783 51388 48800 51428
rect 48840 51388 48849 51428
rect 48463 51365 48529 51388
rect 48615 51365 48697 51388
rect 48783 51365 48849 51388
rect 48463 51346 48849 51365
rect 63583 51451 63969 51470
rect 63583 51428 63649 51451
rect 63735 51428 63817 51451
rect 63903 51428 63969 51451
rect 63583 51388 63592 51428
rect 63632 51388 63649 51428
rect 63735 51388 63756 51428
rect 63796 51388 63817 51428
rect 63903 51388 63920 51428
rect 63960 51388 63969 51428
rect 63583 51365 63649 51388
rect 63735 51365 63817 51388
rect 63903 51365 63969 51388
rect 63583 51346 63969 51365
rect 78703 51451 79089 51470
rect 78703 51428 78769 51451
rect 78855 51428 78937 51451
rect 79023 51428 79089 51451
rect 78703 51388 78712 51428
rect 78752 51388 78769 51428
rect 78855 51388 78876 51428
rect 78916 51388 78937 51428
rect 79023 51388 79040 51428
rect 79080 51388 79089 51428
rect 78703 51365 78769 51388
rect 78855 51365 78937 51388
rect 79023 51365 79089 51388
rect 78703 51346 79089 51365
rect 93823 51451 94209 51470
rect 93823 51428 93889 51451
rect 93975 51428 94057 51451
rect 94143 51428 94209 51451
rect 93823 51388 93832 51428
rect 93872 51388 93889 51428
rect 93975 51388 93996 51428
rect 94036 51388 94057 51428
rect 94143 51388 94160 51428
rect 94200 51388 94209 51428
rect 93823 51365 93889 51388
rect 93975 51365 94057 51388
rect 94143 51365 94209 51388
rect 93823 51346 94209 51365
rect 4343 50695 4729 50714
rect 4343 50672 4409 50695
rect 4495 50672 4577 50695
rect 4663 50672 4729 50695
rect 4343 50632 4352 50672
rect 4392 50632 4409 50672
rect 4495 50632 4516 50672
rect 4556 50632 4577 50672
rect 4663 50632 4680 50672
rect 4720 50632 4729 50672
rect 4343 50609 4409 50632
rect 4495 50609 4577 50632
rect 4663 50609 4729 50632
rect 4343 50590 4729 50609
rect 19463 50695 19849 50714
rect 19463 50672 19529 50695
rect 19615 50672 19697 50695
rect 19783 50672 19849 50695
rect 19463 50632 19472 50672
rect 19512 50632 19529 50672
rect 19615 50632 19636 50672
rect 19676 50632 19697 50672
rect 19783 50632 19800 50672
rect 19840 50632 19849 50672
rect 19463 50609 19529 50632
rect 19615 50609 19697 50632
rect 19783 50609 19849 50632
rect 19463 50590 19849 50609
rect 34583 50695 34969 50714
rect 34583 50672 34649 50695
rect 34735 50672 34817 50695
rect 34903 50672 34969 50695
rect 34583 50632 34592 50672
rect 34632 50632 34649 50672
rect 34735 50632 34756 50672
rect 34796 50632 34817 50672
rect 34903 50632 34920 50672
rect 34960 50632 34969 50672
rect 34583 50609 34649 50632
rect 34735 50609 34817 50632
rect 34903 50609 34969 50632
rect 34583 50590 34969 50609
rect 49703 50695 50089 50714
rect 49703 50672 49769 50695
rect 49855 50672 49937 50695
rect 50023 50672 50089 50695
rect 49703 50632 49712 50672
rect 49752 50632 49769 50672
rect 49855 50632 49876 50672
rect 49916 50632 49937 50672
rect 50023 50632 50040 50672
rect 50080 50632 50089 50672
rect 49703 50609 49769 50632
rect 49855 50609 49937 50632
rect 50023 50609 50089 50632
rect 49703 50590 50089 50609
rect 64823 50695 65209 50714
rect 64823 50672 64889 50695
rect 64975 50672 65057 50695
rect 65143 50672 65209 50695
rect 64823 50632 64832 50672
rect 64872 50632 64889 50672
rect 64975 50632 64996 50672
rect 65036 50632 65057 50672
rect 65143 50632 65160 50672
rect 65200 50632 65209 50672
rect 64823 50609 64889 50632
rect 64975 50609 65057 50632
rect 65143 50609 65209 50632
rect 64823 50590 65209 50609
rect 79943 50695 80329 50714
rect 79943 50672 80009 50695
rect 80095 50672 80177 50695
rect 80263 50672 80329 50695
rect 79943 50632 79952 50672
rect 79992 50632 80009 50672
rect 80095 50632 80116 50672
rect 80156 50632 80177 50672
rect 80263 50632 80280 50672
rect 80320 50632 80329 50672
rect 79943 50609 80009 50632
rect 80095 50609 80177 50632
rect 80263 50609 80329 50632
rect 79943 50590 80329 50609
rect 95063 50695 95449 50714
rect 95063 50672 95129 50695
rect 95215 50672 95297 50695
rect 95383 50672 95449 50695
rect 95063 50632 95072 50672
rect 95112 50632 95129 50672
rect 95215 50632 95236 50672
rect 95276 50632 95297 50672
rect 95383 50632 95400 50672
rect 95440 50632 95449 50672
rect 95063 50609 95129 50632
rect 95215 50609 95297 50632
rect 95383 50609 95449 50632
rect 95063 50590 95449 50609
rect 3103 49939 3489 49958
rect 3103 49916 3169 49939
rect 3255 49916 3337 49939
rect 3423 49916 3489 49939
rect 3103 49876 3112 49916
rect 3152 49876 3169 49916
rect 3255 49876 3276 49916
rect 3316 49876 3337 49916
rect 3423 49876 3440 49916
rect 3480 49876 3489 49916
rect 3103 49853 3169 49876
rect 3255 49853 3337 49876
rect 3423 49853 3489 49876
rect 3103 49834 3489 49853
rect 18223 49939 18609 49958
rect 18223 49916 18289 49939
rect 18375 49916 18457 49939
rect 18543 49916 18609 49939
rect 18223 49876 18232 49916
rect 18272 49876 18289 49916
rect 18375 49876 18396 49916
rect 18436 49876 18457 49916
rect 18543 49876 18560 49916
rect 18600 49876 18609 49916
rect 18223 49853 18289 49876
rect 18375 49853 18457 49876
rect 18543 49853 18609 49876
rect 18223 49834 18609 49853
rect 33343 49939 33729 49958
rect 33343 49916 33409 49939
rect 33495 49916 33577 49939
rect 33663 49916 33729 49939
rect 33343 49876 33352 49916
rect 33392 49876 33409 49916
rect 33495 49876 33516 49916
rect 33556 49876 33577 49916
rect 33663 49876 33680 49916
rect 33720 49876 33729 49916
rect 33343 49853 33409 49876
rect 33495 49853 33577 49876
rect 33663 49853 33729 49876
rect 33343 49834 33729 49853
rect 48463 49939 48849 49958
rect 48463 49916 48529 49939
rect 48615 49916 48697 49939
rect 48783 49916 48849 49939
rect 48463 49876 48472 49916
rect 48512 49876 48529 49916
rect 48615 49876 48636 49916
rect 48676 49876 48697 49916
rect 48783 49876 48800 49916
rect 48840 49876 48849 49916
rect 48463 49853 48529 49876
rect 48615 49853 48697 49876
rect 48783 49853 48849 49876
rect 48463 49834 48849 49853
rect 63583 49939 63969 49958
rect 63583 49916 63649 49939
rect 63735 49916 63817 49939
rect 63903 49916 63969 49939
rect 63583 49876 63592 49916
rect 63632 49876 63649 49916
rect 63735 49876 63756 49916
rect 63796 49876 63817 49916
rect 63903 49876 63920 49916
rect 63960 49876 63969 49916
rect 63583 49853 63649 49876
rect 63735 49853 63817 49876
rect 63903 49853 63969 49876
rect 63583 49834 63969 49853
rect 78703 49939 79089 49958
rect 78703 49916 78769 49939
rect 78855 49916 78937 49939
rect 79023 49916 79089 49939
rect 78703 49876 78712 49916
rect 78752 49876 78769 49916
rect 78855 49876 78876 49916
rect 78916 49876 78937 49916
rect 79023 49876 79040 49916
rect 79080 49876 79089 49916
rect 78703 49853 78769 49876
rect 78855 49853 78937 49876
rect 79023 49853 79089 49876
rect 78703 49834 79089 49853
rect 93823 49939 94209 49958
rect 93823 49916 93889 49939
rect 93975 49916 94057 49939
rect 94143 49916 94209 49939
rect 93823 49876 93832 49916
rect 93872 49876 93889 49916
rect 93975 49876 93996 49916
rect 94036 49876 94057 49916
rect 94143 49876 94160 49916
rect 94200 49876 94209 49916
rect 93823 49853 93889 49876
rect 93975 49853 94057 49876
rect 94143 49853 94209 49876
rect 93823 49834 94209 49853
rect 4343 49183 4729 49202
rect 4343 49160 4409 49183
rect 4495 49160 4577 49183
rect 4663 49160 4729 49183
rect 4343 49120 4352 49160
rect 4392 49120 4409 49160
rect 4495 49120 4516 49160
rect 4556 49120 4577 49160
rect 4663 49120 4680 49160
rect 4720 49120 4729 49160
rect 4343 49097 4409 49120
rect 4495 49097 4577 49120
rect 4663 49097 4729 49120
rect 4343 49078 4729 49097
rect 19463 49183 19849 49202
rect 19463 49160 19529 49183
rect 19615 49160 19697 49183
rect 19783 49160 19849 49183
rect 19463 49120 19472 49160
rect 19512 49120 19529 49160
rect 19615 49120 19636 49160
rect 19676 49120 19697 49160
rect 19783 49120 19800 49160
rect 19840 49120 19849 49160
rect 19463 49097 19529 49120
rect 19615 49097 19697 49120
rect 19783 49097 19849 49120
rect 19463 49078 19849 49097
rect 34583 49183 34969 49202
rect 34583 49160 34649 49183
rect 34735 49160 34817 49183
rect 34903 49160 34969 49183
rect 34583 49120 34592 49160
rect 34632 49120 34649 49160
rect 34735 49120 34756 49160
rect 34796 49120 34817 49160
rect 34903 49120 34920 49160
rect 34960 49120 34969 49160
rect 34583 49097 34649 49120
rect 34735 49097 34817 49120
rect 34903 49097 34969 49120
rect 34583 49078 34969 49097
rect 49703 49183 50089 49202
rect 49703 49160 49769 49183
rect 49855 49160 49937 49183
rect 50023 49160 50089 49183
rect 49703 49120 49712 49160
rect 49752 49120 49769 49160
rect 49855 49120 49876 49160
rect 49916 49120 49937 49160
rect 50023 49120 50040 49160
rect 50080 49120 50089 49160
rect 49703 49097 49769 49120
rect 49855 49097 49937 49120
rect 50023 49097 50089 49120
rect 49703 49078 50089 49097
rect 64823 49183 65209 49202
rect 64823 49160 64889 49183
rect 64975 49160 65057 49183
rect 65143 49160 65209 49183
rect 64823 49120 64832 49160
rect 64872 49120 64889 49160
rect 64975 49120 64996 49160
rect 65036 49120 65057 49160
rect 65143 49120 65160 49160
rect 65200 49120 65209 49160
rect 64823 49097 64889 49120
rect 64975 49097 65057 49120
rect 65143 49097 65209 49120
rect 64823 49078 65209 49097
rect 79943 49183 80329 49202
rect 79943 49160 80009 49183
rect 80095 49160 80177 49183
rect 80263 49160 80329 49183
rect 79943 49120 79952 49160
rect 79992 49120 80009 49160
rect 80095 49120 80116 49160
rect 80156 49120 80177 49160
rect 80263 49120 80280 49160
rect 80320 49120 80329 49160
rect 79943 49097 80009 49120
rect 80095 49097 80177 49120
rect 80263 49097 80329 49120
rect 79943 49078 80329 49097
rect 95063 49183 95449 49202
rect 95063 49160 95129 49183
rect 95215 49160 95297 49183
rect 95383 49160 95449 49183
rect 95063 49120 95072 49160
rect 95112 49120 95129 49160
rect 95215 49120 95236 49160
rect 95276 49120 95297 49160
rect 95383 49120 95400 49160
rect 95440 49120 95449 49160
rect 95063 49097 95129 49120
rect 95215 49097 95297 49120
rect 95383 49097 95449 49120
rect 95063 49078 95449 49097
rect 3103 48427 3489 48446
rect 3103 48404 3169 48427
rect 3255 48404 3337 48427
rect 3423 48404 3489 48427
rect 3103 48364 3112 48404
rect 3152 48364 3169 48404
rect 3255 48364 3276 48404
rect 3316 48364 3337 48404
rect 3423 48364 3440 48404
rect 3480 48364 3489 48404
rect 3103 48341 3169 48364
rect 3255 48341 3337 48364
rect 3423 48341 3489 48364
rect 3103 48322 3489 48341
rect 18223 48427 18609 48446
rect 18223 48404 18289 48427
rect 18375 48404 18457 48427
rect 18543 48404 18609 48427
rect 18223 48364 18232 48404
rect 18272 48364 18289 48404
rect 18375 48364 18396 48404
rect 18436 48364 18457 48404
rect 18543 48364 18560 48404
rect 18600 48364 18609 48404
rect 18223 48341 18289 48364
rect 18375 48341 18457 48364
rect 18543 48341 18609 48364
rect 18223 48322 18609 48341
rect 33343 48427 33729 48446
rect 33343 48404 33409 48427
rect 33495 48404 33577 48427
rect 33663 48404 33729 48427
rect 33343 48364 33352 48404
rect 33392 48364 33409 48404
rect 33495 48364 33516 48404
rect 33556 48364 33577 48404
rect 33663 48364 33680 48404
rect 33720 48364 33729 48404
rect 33343 48341 33409 48364
rect 33495 48341 33577 48364
rect 33663 48341 33729 48364
rect 33343 48322 33729 48341
rect 48463 48427 48849 48446
rect 48463 48404 48529 48427
rect 48615 48404 48697 48427
rect 48783 48404 48849 48427
rect 48463 48364 48472 48404
rect 48512 48364 48529 48404
rect 48615 48364 48636 48404
rect 48676 48364 48697 48404
rect 48783 48364 48800 48404
rect 48840 48364 48849 48404
rect 48463 48341 48529 48364
rect 48615 48341 48697 48364
rect 48783 48341 48849 48364
rect 48463 48322 48849 48341
rect 63583 48427 63969 48446
rect 63583 48404 63649 48427
rect 63735 48404 63817 48427
rect 63903 48404 63969 48427
rect 63583 48364 63592 48404
rect 63632 48364 63649 48404
rect 63735 48364 63756 48404
rect 63796 48364 63817 48404
rect 63903 48364 63920 48404
rect 63960 48364 63969 48404
rect 63583 48341 63649 48364
rect 63735 48341 63817 48364
rect 63903 48341 63969 48364
rect 63583 48322 63969 48341
rect 78703 48427 79089 48446
rect 78703 48404 78769 48427
rect 78855 48404 78937 48427
rect 79023 48404 79089 48427
rect 78703 48364 78712 48404
rect 78752 48364 78769 48404
rect 78855 48364 78876 48404
rect 78916 48364 78937 48404
rect 79023 48364 79040 48404
rect 79080 48364 79089 48404
rect 78703 48341 78769 48364
rect 78855 48341 78937 48364
rect 79023 48341 79089 48364
rect 78703 48322 79089 48341
rect 93823 48427 94209 48446
rect 93823 48404 93889 48427
rect 93975 48404 94057 48427
rect 94143 48404 94209 48427
rect 93823 48364 93832 48404
rect 93872 48364 93889 48404
rect 93975 48364 93996 48404
rect 94036 48364 94057 48404
rect 94143 48364 94160 48404
rect 94200 48364 94209 48404
rect 93823 48341 93889 48364
rect 93975 48341 94057 48364
rect 94143 48341 94209 48364
rect 93823 48322 94209 48341
rect 4343 47671 4729 47690
rect 4343 47648 4409 47671
rect 4495 47648 4577 47671
rect 4663 47648 4729 47671
rect 4343 47608 4352 47648
rect 4392 47608 4409 47648
rect 4495 47608 4516 47648
rect 4556 47608 4577 47648
rect 4663 47608 4680 47648
rect 4720 47608 4729 47648
rect 4343 47585 4409 47608
rect 4495 47585 4577 47608
rect 4663 47585 4729 47608
rect 4343 47566 4729 47585
rect 19463 47671 19849 47690
rect 19463 47648 19529 47671
rect 19615 47648 19697 47671
rect 19783 47648 19849 47671
rect 19463 47608 19472 47648
rect 19512 47608 19529 47648
rect 19615 47608 19636 47648
rect 19676 47608 19697 47648
rect 19783 47608 19800 47648
rect 19840 47608 19849 47648
rect 19463 47585 19529 47608
rect 19615 47585 19697 47608
rect 19783 47585 19849 47608
rect 19463 47566 19849 47585
rect 34583 47671 34969 47690
rect 34583 47648 34649 47671
rect 34735 47648 34817 47671
rect 34903 47648 34969 47671
rect 34583 47608 34592 47648
rect 34632 47608 34649 47648
rect 34735 47608 34756 47648
rect 34796 47608 34817 47648
rect 34903 47608 34920 47648
rect 34960 47608 34969 47648
rect 34583 47585 34649 47608
rect 34735 47585 34817 47608
rect 34903 47585 34969 47608
rect 34583 47566 34969 47585
rect 49703 47671 50089 47690
rect 49703 47648 49769 47671
rect 49855 47648 49937 47671
rect 50023 47648 50089 47671
rect 49703 47608 49712 47648
rect 49752 47608 49769 47648
rect 49855 47608 49876 47648
rect 49916 47608 49937 47648
rect 50023 47608 50040 47648
rect 50080 47608 50089 47648
rect 49703 47585 49769 47608
rect 49855 47585 49937 47608
rect 50023 47585 50089 47608
rect 49703 47566 50089 47585
rect 64823 47671 65209 47690
rect 64823 47648 64889 47671
rect 64975 47648 65057 47671
rect 65143 47648 65209 47671
rect 64823 47608 64832 47648
rect 64872 47608 64889 47648
rect 64975 47608 64996 47648
rect 65036 47608 65057 47648
rect 65143 47608 65160 47648
rect 65200 47608 65209 47648
rect 64823 47585 64889 47608
rect 64975 47585 65057 47608
rect 65143 47585 65209 47608
rect 64823 47566 65209 47585
rect 79943 47671 80329 47690
rect 79943 47648 80009 47671
rect 80095 47648 80177 47671
rect 80263 47648 80329 47671
rect 79943 47608 79952 47648
rect 79992 47608 80009 47648
rect 80095 47608 80116 47648
rect 80156 47608 80177 47648
rect 80263 47608 80280 47648
rect 80320 47608 80329 47648
rect 79943 47585 80009 47608
rect 80095 47585 80177 47608
rect 80263 47585 80329 47608
rect 79943 47566 80329 47585
rect 95063 47671 95449 47690
rect 95063 47648 95129 47671
rect 95215 47648 95297 47671
rect 95383 47648 95449 47671
rect 95063 47608 95072 47648
rect 95112 47608 95129 47648
rect 95215 47608 95236 47648
rect 95276 47608 95297 47648
rect 95383 47608 95400 47648
rect 95440 47608 95449 47648
rect 95063 47585 95129 47608
rect 95215 47585 95297 47608
rect 95383 47585 95449 47608
rect 95063 47566 95449 47585
rect 3103 46915 3489 46934
rect 3103 46892 3169 46915
rect 3255 46892 3337 46915
rect 3423 46892 3489 46915
rect 3103 46852 3112 46892
rect 3152 46852 3169 46892
rect 3255 46852 3276 46892
rect 3316 46852 3337 46892
rect 3423 46852 3440 46892
rect 3480 46852 3489 46892
rect 3103 46829 3169 46852
rect 3255 46829 3337 46852
rect 3423 46829 3489 46852
rect 3103 46810 3489 46829
rect 18223 46915 18609 46934
rect 18223 46892 18289 46915
rect 18375 46892 18457 46915
rect 18543 46892 18609 46915
rect 18223 46852 18232 46892
rect 18272 46852 18289 46892
rect 18375 46852 18396 46892
rect 18436 46852 18457 46892
rect 18543 46852 18560 46892
rect 18600 46852 18609 46892
rect 18223 46829 18289 46852
rect 18375 46829 18457 46852
rect 18543 46829 18609 46852
rect 18223 46810 18609 46829
rect 33343 46915 33729 46934
rect 33343 46892 33409 46915
rect 33495 46892 33577 46915
rect 33663 46892 33729 46915
rect 33343 46852 33352 46892
rect 33392 46852 33409 46892
rect 33495 46852 33516 46892
rect 33556 46852 33577 46892
rect 33663 46852 33680 46892
rect 33720 46852 33729 46892
rect 33343 46829 33409 46852
rect 33495 46829 33577 46852
rect 33663 46829 33729 46852
rect 33343 46810 33729 46829
rect 48463 46915 48849 46934
rect 48463 46892 48529 46915
rect 48615 46892 48697 46915
rect 48783 46892 48849 46915
rect 48463 46852 48472 46892
rect 48512 46852 48529 46892
rect 48615 46852 48636 46892
rect 48676 46852 48697 46892
rect 48783 46852 48800 46892
rect 48840 46852 48849 46892
rect 48463 46829 48529 46852
rect 48615 46829 48697 46852
rect 48783 46829 48849 46852
rect 48463 46810 48849 46829
rect 63583 46915 63969 46934
rect 63583 46892 63649 46915
rect 63735 46892 63817 46915
rect 63903 46892 63969 46915
rect 63583 46852 63592 46892
rect 63632 46852 63649 46892
rect 63735 46852 63756 46892
rect 63796 46852 63817 46892
rect 63903 46852 63920 46892
rect 63960 46852 63969 46892
rect 63583 46829 63649 46852
rect 63735 46829 63817 46852
rect 63903 46829 63969 46852
rect 63583 46810 63969 46829
rect 78703 46915 79089 46934
rect 78703 46892 78769 46915
rect 78855 46892 78937 46915
rect 79023 46892 79089 46915
rect 78703 46852 78712 46892
rect 78752 46852 78769 46892
rect 78855 46852 78876 46892
rect 78916 46852 78937 46892
rect 79023 46852 79040 46892
rect 79080 46852 79089 46892
rect 78703 46829 78769 46852
rect 78855 46829 78937 46852
rect 79023 46829 79089 46852
rect 78703 46810 79089 46829
rect 93823 46915 94209 46934
rect 93823 46892 93889 46915
rect 93975 46892 94057 46915
rect 94143 46892 94209 46915
rect 93823 46852 93832 46892
rect 93872 46852 93889 46892
rect 93975 46852 93996 46892
rect 94036 46852 94057 46892
rect 94143 46852 94160 46892
rect 94200 46852 94209 46892
rect 93823 46829 93889 46852
rect 93975 46829 94057 46852
rect 94143 46829 94209 46852
rect 93823 46810 94209 46829
rect 4343 46159 4729 46178
rect 4343 46136 4409 46159
rect 4495 46136 4577 46159
rect 4663 46136 4729 46159
rect 4343 46096 4352 46136
rect 4392 46096 4409 46136
rect 4495 46096 4516 46136
rect 4556 46096 4577 46136
rect 4663 46096 4680 46136
rect 4720 46096 4729 46136
rect 4343 46073 4409 46096
rect 4495 46073 4577 46096
rect 4663 46073 4729 46096
rect 4343 46054 4729 46073
rect 19463 46159 19849 46178
rect 19463 46136 19529 46159
rect 19615 46136 19697 46159
rect 19783 46136 19849 46159
rect 19463 46096 19472 46136
rect 19512 46096 19529 46136
rect 19615 46096 19636 46136
rect 19676 46096 19697 46136
rect 19783 46096 19800 46136
rect 19840 46096 19849 46136
rect 19463 46073 19529 46096
rect 19615 46073 19697 46096
rect 19783 46073 19849 46096
rect 19463 46054 19849 46073
rect 34583 46159 34969 46178
rect 34583 46136 34649 46159
rect 34735 46136 34817 46159
rect 34903 46136 34969 46159
rect 34583 46096 34592 46136
rect 34632 46096 34649 46136
rect 34735 46096 34756 46136
rect 34796 46096 34817 46136
rect 34903 46096 34920 46136
rect 34960 46096 34969 46136
rect 34583 46073 34649 46096
rect 34735 46073 34817 46096
rect 34903 46073 34969 46096
rect 34583 46054 34969 46073
rect 49703 46159 50089 46178
rect 49703 46136 49769 46159
rect 49855 46136 49937 46159
rect 50023 46136 50089 46159
rect 49703 46096 49712 46136
rect 49752 46096 49769 46136
rect 49855 46096 49876 46136
rect 49916 46096 49937 46136
rect 50023 46096 50040 46136
rect 50080 46096 50089 46136
rect 49703 46073 49769 46096
rect 49855 46073 49937 46096
rect 50023 46073 50089 46096
rect 49703 46054 50089 46073
rect 64823 46159 65209 46178
rect 64823 46136 64889 46159
rect 64975 46136 65057 46159
rect 65143 46136 65209 46159
rect 64823 46096 64832 46136
rect 64872 46096 64889 46136
rect 64975 46096 64996 46136
rect 65036 46096 65057 46136
rect 65143 46096 65160 46136
rect 65200 46096 65209 46136
rect 64823 46073 64889 46096
rect 64975 46073 65057 46096
rect 65143 46073 65209 46096
rect 64823 46054 65209 46073
rect 79943 46159 80329 46178
rect 79943 46136 80009 46159
rect 80095 46136 80177 46159
rect 80263 46136 80329 46159
rect 79943 46096 79952 46136
rect 79992 46096 80009 46136
rect 80095 46096 80116 46136
rect 80156 46096 80177 46136
rect 80263 46096 80280 46136
rect 80320 46096 80329 46136
rect 79943 46073 80009 46096
rect 80095 46073 80177 46096
rect 80263 46073 80329 46096
rect 79943 46054 80329 46073
rect 95063 46159 95449 46178
rect 95063 46136 95129 46159
rect 95215 46136 95297 46159
rect 95383 46136 95449 46159
rect 95063 46096 95072 46136
rect 95112 46096 95129 46136
rect 95215 46096 95236 46136
rect 95276 46096 95297 46136
rect 95383 46096 95400 46136
rect 95440 46096 95449 46136
rect 95063 46073 95129 46096
rect 95215 46073 95297 46096
rect 95383 46073 95449 46096
rect 95063 46054 95449 46073
rect 3103 45403 3489 45422
rect 3103 45380 3169 45403
rect 3255 45380 3337 45403
rect 3423 45380 3489 45403
rect 3103 45340 3112 45380
rect 3152 45340 3169 45380
rect 3255 45340 3276 45380
rect 3316 45340 3337 45380
rect 3423 45340 3440 45380
rect 3480 45340 3489 45380
rect 3103 45317 3169 45340
rect 3255 45317 3337 45340
rect 3423 45317 3489 45340
rect 3103 45298 3489 45317
rect 18223 45403 18609 45422
rect 18223 45380 18289 45403
rect 18375 45380 18457 45403
rect 18543 45380 18609 45403
rect 18223 45340 18232 45380
rect 18272 45340 18289 45380
rect 18375 45340 18396 45380
rect 18436 45340 18457 45380
rect 18543 45340 18560 45380
rect 18600 45340 18609 45380
rect 18223 45317 18289 45340
rect 18375 45317 18457 45340
rect 18543 45317 18609 45340
rect 18223 45298 18609 45317
rect 33343 45403 33729 45422
rect 33343 45380 33409 45403
rect 33495 45380 33577 45403
rect 33663 45380 33729 45403
rect 33343 45340 33352 45380
rect 33392 45340 33409 45380
rect 33495 45340 33516 45380
rect 33556 45340 33577 45380
rect 33663 45340 33680 45380
rect 33720 45340 33729 45380
rect 33343 45317 33409 45340
rect 33495 45317 33577 45340
rect 33663 45317 33729 45340
rect 33343 45298 33729 45317
rect 48463 45403 48849 45422
rect 48463 45380 48529 45403
rect 48615 45380 48697 45403
rect 48783 45380 48849 45403
rect 48463 45340 48472 45380
rect 48512 45340 48529 45380
rect 48615 45340 48636 45380
rect 48676 45340 48697 45380
rect 48783 45340 48800 45380
rect 48840 45340 48849 45380
rect 48463 45317 48529 45340
rect 48615 45317 48697 45340
rect 48783 45317 48849 45340
rect 48463 45298 48849 45317
rect 63583 45403 63969 45422
rect 63583 45380 63649 45403
rect 63735 45380 63817 45403
rect 63903 45380 63969 45403
rect 63583 45340 63592 45380
rect 63632 45340 63649 45380
rect 63735 45340 63756 45380
rect 63796 45340 63817 45380
rect 63903 45340 63920 45380
rect 63960 45340 63969 45380
rect 63583 45317 63649 45340
rect 63735 45317 63817 45340
rect 63903 45317 63969 45340
rect 63583 45298 63969 45317
rect 78703 45403 79089 45422
rect 78703 45380 78769 45403
rect 78855 45380 78937 45403
rect 79023 45380 79089 45403
rect 78703 45340 78712 45380
rect 78752 45340 78769 45380
rect 78855 45340 78876 45380
rect 78916 45340 78937 45380
rect 79023 45340 79040 45380
rect 79080 45340 79089 45380
rect 78703 45317 78769 45340
rect 78855 45317 78937 45340
rect 79023 45317 79089 45340
rect 78703 45298 79089 45317
rect 93823 45403 94209 45422
rect 93823 45380 93889 45403
rect 93975 45380 94057 45403
rect 94143 45380 94209 45403
rect 93823 45340 93832 45380
rect 93872 45340 93889 45380
rect 93975 45340 93996 45380
rect 94036 45340 94057 45380
rect 94143 45340 94160 45380
rect 94200 45340 94209 45380
rect 93823 45317 93889 45340
rect 93975 45317 94057 45340
rect 94143 45317 94209 45340
rect 93823 45298 94209 45317
rect 4343 44647 4729 44666
rect 4343 44624 4409 44647
rect 4495 44624 4577 44647
rect 4663 44624 4729 44647
rect 4343 44584 4352 44624
rect 4392 44584 4409 44624
rect 4495 44584 4516 44624
rect 4556 44584 4577 44624
rect 4663 44584 4680 44624
rect 4720 44584 4729 44624
rect 4343 44561 4409 44584
rect 4495 44561 4577 44584
rect 4663 44561 4729 44584
rect 4343 44542 4729 44561
rect 19463 44647 19849 44666
rect 19463 44624 19529 44647
rect 19615 44624 19697 44647
rect 19783 44624 19849 44647
rect 19463 44584 19472 44624
rect 19512 44584 19529 44624
rect 19615 44584 19636 44624
rect 19676 44584 19697 44624
rect 19783 44584 19800 44624
rect 19840 44584 19849 44624
rect 19463 44561 19529 44584
rect 19615 44561 19697 44584
rect 19783 44561 19849 44584
rect 19463 44542 19849 44561
rect 34583 44647 34969 44666
rect 34583 44624 34649 44647
rect 34735 44624 34817 44647
rect 34903 44624 34969 44647
rect 34583 44584 34592 44624
rect 34632 44584 34649 44624
rect 34735 44584 34756 44624
rect 34796 44584 34817 44624
rect 34903 44584 34920 44624
rect 34960 44584 34969 44624
rect 34583 44561 34649 44584
rect 34735 44561 34817 44584
rect 34903 44561 34969 44584
rect 34583 44542 34969 44561
rect 49703 44647 50089 44666
rect 49703 44624 49769 44647
rect 49855 44624 49937 44647
rect 50023 44624 50089 44647
rect 49703 44584 49712 44624
rect 49752 44584 49769 44624
rect 49855 44584 49876 44624
rect 49916 44584 49937 44624
rect 50023 44584 50040 44624
rect 50080 44584 50089 44624
rect 49703 44561 49769 44584
rect 49855 44561 49937 44584
rect 50023 44561 50089 44584
rect 49703 44542 50089 44561
rect 64823 44647 65209 44666
rect 64823 44624 64889 44647
rect 64975 44624 65057 44647
rect 65143 44624 65209 44647
rect 64823 44584 64832 44624
rect 64872 44584 64889 44624
rect 64975 44584 64996 44624
rect 65036 44584 65057 44624
rect 65143 44584 65160 44624
rect 65200 44584 65209 44624
rect 64823 44561 64889 44584
rect 64975 44561 65057 44584
rect 65143 44561 65209 44584
rect 64823 44542 65209 44561
rect 79943 44647 80329 44666
rect 79943 44624 80009 44647
rect 80095 44624 80177 44647
rect 80263 44624 80329 44647
rect 79943 44584 79952 44624
rect 79992 44584 80009 44624
rect 80095 44584 80116 44624
rect 80156 44584 80177 44624
rect 80263 44584 80280 44624
rect 80320 44584 80329 44624
rect 79943 44561 80009 44584
rect 80095 44561 80177 44584
rect 80263 44561 80329 44584
rect 79943 44542 80329 44561
rect 95063 44647 95449 44666
rect 95063 44624 95129 44647
rect 95215 44624 95297 44647
rect 95383 44624 95449 44647
rect 95063 44584 95072 44624
rect 95112 44584 95129 44624
rect 95215 44584 95236 44624
rect 95276 44584 95297 44624
rect 95383 44584 95400 44624
rect 95440 44584 95449 44624
rect 95063 44561 95129 44584
rect 95215 44561 95297 44584
rect 95383 44561 95449 44584
rect 95063 44542 95449 44561
rect 3103 43891 3489 43910
rect 3103 43868 3169 43891
rect 3255 43868 3337 43891
rect 3423 43868 3489 43891
rect 3103 43828 3112 43868
rect 3152 43828 3169 43868
rect 3255 43828 3276 43868
rect 3316 43828 3337 43868
rect 3423 43828 3440 43868
rect 3480 43828 3489 43868
rect 3103 43805 3169 43828
rect 3255 43805 3337 43828
rect 3423 43805 3489 43828
rect 3103 43786 3489 43805
rect 18223 43891 18609 43910
rect 18223 43868 18289 43891
rect 18375 43868 18457 43891
rect 18543 43868 18609 43891
rect 18223 43828 18232 43868
rect 18272 43828 18289 43868
rect 18375 43828 18396 43868
rect 18436 43828 18457 43868
rect 18543 43828 18560 43868
rect 18600 43828 18609 43868
rect 18223 43805 18289 43828
rect 18375 43805 18457 43828
rect 18543 43805 18609 43828
rect 18223 43786 18609 43805
rect 33343 43891 33729 43910
rect 33343 43868 33409 43891
rect 33495 43868 33577 43891
rect 33663 43868 33729 43891
rect 33343 43828 33352 43868
rect 33392 43828 33409 43868
rect 33495 43828 33516 43868
rect 33556 43828 33577 43868
rect 33663 43828 33680 43868
rect 33720 43828 33729 43868
rect 33343 43805 33409 43828
rect 33495 43805 33577 43828
rect 33663 43805 33729 43828
rect 33343 43786 33729 43805
rect 48463 43891 48849 43910
rect 48463 43868 48529 43891
rect 48615 43868 48697 43891
rect 48783 43868 48849 43891
rect 48463 43828 48472 43868
rect 48512 43828 48529 43868
rect 48615 43828 48636 43868
rect 48676 43828 48697 43868
rect 48783 43828 48800 43868
rect 48840 43828 48849 43868
rect 48463 43805 48529 43828
rect 48615 43805 48697 43828
rect 48783 43805 48849 43828
rect 48463 43786 48849 43805
rect 63583 43891 63969 43910
rect 63583 43868 63649 43891
rect 63735 43868 63817 43891
rect 63903 43868 63969 43891
rect 63583 43828 63592 43868
rect 63632 43828 63649 43868
rect 63735 43828 63756 43868
rect 63796 43828 63817 43868
rect 63903 43828 63920 43868
rect 63960 43828 63969 43868
rect 63583 43805 63649 43828
rect 63735 43805 63817 43828
rect 63903 43805 63969 43828
rect 63583 43786 63969 43805
rect 78703 43891 79089 43910
rect 78703 43868 78769 43891
rect 78855 43868 78937 43891
rect 79023 43868 79089 43891
rect 78703 43828 78712 43868
rect 78752 43828 78769 43868
rect 78855 43828 78876 43868
rect 78916 43828 78937 43868
rect 79023 43828 79040 43868
rect 79080 43828 79089 43868
rect 78703 43805 78769 43828
rect 78855 43805 78937 43828
rect 79023 43805 79089 43828
rect 78703 43786 79089 43805
rect 93823 43891 94209 43910
rect 93823 43868 93889 43891
rect 93975 43868 94057 43891
rect 94143 43868 94209 43891
rect 93823 43828 93832 43868
rect 93872 43828 93889 43868
rect 93975 43828 93996 43868
rect 94036 43828 94057 43868
rect 94143 43828 94160 43868
rect 94200 43828 94209 43868
rect 93823 43805 93889 43828
rect 93975 43805 94057 43828
rect 94143 43805 94209 43828
rect 93823 43786 94209 43805
rect 4343 43135 4729 43154
rect 4343 43112 4409 43135
rect 4495 43112 4577 43135
rect 4663 43112 4729 43135
rect 4343 43072 4352 43112
rect 4392 43072 4409 43112
rect 4495 43072 4516 43112
rect 4556 43072 4577 43112
rect 4663 43072 4680 43112
rect 4720 43072 4729 43112
rect 4343 43049 4409 43072
rect 4495 43049 4577 43072
rect 4663 43049 4729 43072
rect 4343 43030 4729 43049
rect 19463 43135 19849 43154
rect 19463 43112 19529 43135
rect 19615 43112 19697 43135
rect 19783 43112 19849 43135
rect 19463 43072 19472 43112
rect 19512 43072 19529 43112
rect 19615 43072 19636 43112
rect 19676 43072 19697 43112
rect 19783 43072 19800 43112
rect 19840 43072 19849 43112
rect 19463 43049 19529 43072
rect 19615 43049 19697 43072
rect 19783 43049 19849 43072
rect 19463 43030 19849 43049
rect 34583 43135 34969 43154
rect 34583 43112 34649 43135
rect 34735 43112 34817 43135
rect 34903 43112 34969 43135
rect 34583 43072 34592 43112
rect 34632 43072 34649 43112
rect 34735 43072 34756 43112
rect 34796 43072 34817 43112
rect 34903 43072 34920 43112
rect 34960 43072 34969 43112
rect 34583 43049 34649 43072
rect 34735 43049 34817 43072
rect 34903 43049 34969 43072
rect 34583 43030 34969 43049
rect 49703 43135 50089 43154
rect 49703 43112 49769 43135
rect 49855 43112 49937 43135
rect 50023 43112 50089 43135
rect 49703 43072 49712 43112
rect 49752 43072 49769 43112
rect 49855 43072 49876 43112
rect 49916 43072 49937 43112
rect 50023 43072 50040 43112
rect 50080 43072 50089 43112
rect 49703 43049 49769 43072
rect 49855 43049 49937 43072
rect 50023 43049 50089 43072
rect 49703 43030 50089 43049
rect 64823 43135 65209 43154
rect 64823 43112 64889 43135
rect 64975 43112 65057 43135
rect 65143 43112 65209 43135
rect 64823 43072 64832 43112
rect 64872 43072 64889 43112
rect 64975 43072 64996 43112
rect 65036 43072 65057 43112
rect 65143 43072 65160 43112
rect 65200 43072 65209 43112
rect 64823 43049 64889 43072
rect 64975 43049 65057 43072
rect 65143 43049 65209 43072
rect 64823 43030 65209 43049
rect 79943 43135 80329 43154
rect 79943 43112 80009 43135
rect 80095 43112 80177 43135
rect 80263 43112 80329 43135
rect 79943 43072 79952 43112
rect 79992 43072 80009 43112
rect 80095 43072 80116 43112
rect 80156 43072 80177 43112
rect 80263 43072 80280 43112
rect 80320 43072 80329 43112
rect 79943 43049 80009 43072
rect 80095 43049 80177 43072
rect 80263 43049 80329 43072
rect 79943 43030 80329 43049
rect 95063 43135 95449 43154
rect 95063 43112 95129 43135
rect 95215 43112 95297 43135
rect 95383 43112 95449 43135
rect 95063 43072 95072 43112
rect 95112 43072 95129 43112
rect 95215 43072 95236 43112
rect 95276 43072 95297 43112
rect 95383 43072 95400 43112
rect 95440 43072 95449 43112
rect 95063 43049 95129 43072
rect 95215 43049 95297 43072
rect 95383 43049 95449 43072
rect 95063 43030 95449 43049
rect 3103 42379 3489 42398
rect 3103 42356 3169 42379
rect 3255 42356 3337 42379
rect 3423 42356 3489 42379
rect 3103 42316 3112 42356
rect 3152 42316 3169 42356
rect 3255 42316 3276 42356
rect 3316 42316 3337 42356
rect 3423 42316 3440 42356
rect 3480 42316 3489 42356
rect 3103 42293 3169 42316
rect 3255 42293 3337 42316
rect 3423 42293 3489 42316
rect 3103 42274 3489 42293
rect 18223 42379 18609 42398
rect 18223 42356 18289 42379
rect 18375 42356 18457 42379
rect 18543 42356 18609 42379
rect 18223 42316 18232 42356
rect 18272 42316 18289 42356
rect 18375 42316 18396 42356
rect 18436 42316 18457 42356
rect 18543 42316 18560 42356
rect 18600 42316 18609 42356
rect 18223 42293 18289 42316
rect 18375 42293 18457 42316
rect 18543 42293 18609 42316
rect 18223 42274 18609 42293
rect 33343 42379 33729 42398
rect 33343 42356 33409 42379
rect 33495 42356 33577 42379
rect 33663 42356 33729 42379
rect 33343 42316 33352 42356
rect 33392 42316 33409 42356
rect 33495 42316 33516 42356
rect 33556 42316 33577 42356
rect 33663 42316 33680 42356
rect 33720 42316 33729 42356
rect 33343 42293 33409 42316
rect 33495 42293 33577 42316
rect 33663 42293 33729 42316
rect 33343 42274 33729 42293
rect 48463 42379 48849 42398
rect 48463 42356 48529 42379
rect 48615 42356 48697 42379
rect 48783 42356 48849 42379
rect 48463 42316 48472 42356
rect 48512 42316 48529 42356
rect 48615 42316 48636 42356
rect 48676 42316 48697 42356
rect 48783 42316 48800 42356
rect 48840 42316 48849 42356
rect 48463 42293 48529 42316
rect 48615 42293 48697 42316
rect 48783 42293 48849 42316
rect 48463 42274 48849 42293
rect 63583 42379 63969 42398
rect 63583 42356 63649 42379
rect 63735 42356 63817 42379
rect 63903 42356 63969 42379
rect 63583 42316 63592 42356
rect 63632 42316 63649 42356
rect 63735 42316 63756 42356
rect 63796 42316 63817 42356
rect 63903 42316 63920 42356
rect 63960 42316 63969 42356
rect 63583 42293 63649 42316
rect 63735 42293 63817 42316
rect 63903 42293 63969 42316
rect 63583 42274 63969 42293
rect 78703 42379 79089 42398
rect 78703 42356 78769 42379
rect 78855 42356 78937 42379
rect 79023 42356 79089 42379
rect 78703 42316 78712 42356
rect 78752 42316 78769 42356
rect 78855 42316 78876 42356
rect 78916 42316 78937 42356
rect 79023 42316 79040 42356
rect 79080 42316 79089 42356
rect 78703 42293 78769 42316
rect 78855 42293 78937 42316
rect 79023 42293 79089 42316
rect 78703 42274 79089 42293
rect 93823 42379 94209 42398
rect 93823 42356 93889 42379
rect 93975 42356 94057 42379
rect 94143 42356 94209 42379
rect 93823 42316 93832 42356
rect 93872 42316 93889 42356
rect 93975 42316 93996 42356
rect 94036 42316 94057 42356
rect 94143 42316 94160 42356
rect 94200 42316 94209 42356
rect 93823 42293 93889 42316
rect 93975 42293 94057 42316
rect 94143 42293 94209 42316
rect 93823 42274 94209 42293
rect 4343 41623 4729 41642
rect 4343 41600 4409 41623
rect 4495 41600 4577 41623
rect 4663 41600 4729 41623
rect 4343 41560 4352 41600
rect 4392 41560 4409 41600
rect 4495 41560 4516 41600
rect 4556 41560 4577 41600
rect 4663 41560 4680 41600
rect 4720 41560 4729 41600
rect 4343 41537 4409 41560
rect 4495 41537 4577 41560
rect 4663 41537 4729 41560
rect 4343 41518 4729 41537
rect 19463 41623 19849 41642
rect 19463 41600 19529 41623
rect 19615 41600 19697 41623
rect 19783 41600 19849 41623
rect 19463 41560 19472 41600
rect 19512 41560 19529 41600
rect 19615 41560 19636 41600
rect 19676 41560 19697 41600
rect 19783 41560 19800 41600
rect 19840 41560 19849 41600
rect 19463 41537 19529 41560
rect 19615 41537 19697 41560
rect 19783 41537 19849 41560
rect 19463 41518 19849 41537
rect 34583 41623 34969 41642
rect 34583 41600 34649 41623
rect 34735 41600 34817 41623
rect 34903 41600 34969 41623
rect 34583 41560 34592 41600
rect 34632 41560 34649 41600
rect 34735 41560 34756 41600
rect 34796 41560 34817 41600
rect 34903 41560 34920 41600
rect 34960 41560 34969 41600
rect 34583 41537 34649 41560
rect 34735 41537 34817 41560
rect 34903 41537 34969 41560
rect 34583 41518 34969 41537
rect 49703 41623 50089 41642
rect 49703 41600 49769 41623
rect 49855 41600 49937 41623
rect 50023 41600 50089 41623
rect 49703 41560 49712 41600
rect 49752 41560 49769 41600
rect 49855 41560 49876 41600
rect 49916 41560 49937 41600
rect 50023 41560 50040 41600
rect 50080 41560 50089 41600
rect 49703 41537 49769 41560
rect 49855 41537 49937 41560
rect 50023 41537 50089 41560
rect 49703 41518 50089 41537
rect 64823 41623 65209 41642
rect 64823 41600 64889 41623
rect 64975 41600 65057 41623
rect 65143 41600 65209 41623
rect 64823 41560 64832 41600
rect 64872 41560 64889 41600
rect 64975 41560 64996 41600
rect 65036 41560 65057 41600
rect 65143 41560 65160 41600
rect 65200 41560 65209 41600
rect 64823 41537 64889 41560
rect 64975 41537 65057 41560
rect 65143 41537 65209 41560
rect 64823 41518 65209 41537
rect 79943 41623 80329 41642
rect 79943 41600 80009 41623
rect 80095 41600 80177 41623
rect 80263 41600 80329 41623
rect 79943 41560 79952 41600
rect 79992 41560 80009 41600
rect 80095 41560 80116 41600
rect 80156 41560 80177 41600
rect 80263 41560 80280 41600
rect 80320 41560 80329 41600
rect 79943 41537 80009 41560
rect 80095 41537 80177 41560
rect 80263 41537 80329 41560
rect 79943 41518 80329 41537
rect 95063 41623 95449 41642
rect 95063 41600 95129 41623
rect 95215 41600 95297 41623
rect 95383 41600 95449 41623
rect 95063 41560 95072 41600
rect 95112 41560 95129 41600
rect 95215 41560 95236 41600
rect 95276 41560 95297 41600
rect 95383 41560 95400 41600
rect 95440 41560 95449 41600
rect 95063 41537 95129 41560
rect 95215 41537 95297 41560
rect 95383 41537 95449 41560
rect 95063 41518 95449 41537
rect 3103 40867 3489 40886
rect 3103 40844 3169 40867
rect 3255 40844 3337 40867
rect 3423 40844 3489 40867
rect 3103 40804 3112 40844
rect 3152 40804 3169 40844
rect 3255 40804 3276 40844
rect 3316 40804 3337 40844
rect 3423 40804 3440 40844
rect 3480 40804 3489 40844
rect 3103 40781 3169 40804
rect 3255 40781 3337 40804
rect 3423 40781 3489 40804
rect 3103 40762 3489 40781
rect 18223 40867 18609 40886
rect 18223 40844 18289 40867
rect 18375 40844 18457 40867
rect 18543 40844 18609 40867
rect 18223 40804 18232 40844
rect 18272 40804 18289 40844
rect 18375 40804 18396 40844
rect 18436 40804 18457 40844
rect 18543 40804 18560 40844
rect 18600 40804 18609 40844
rect 18223 40781 18289 40804
rect 18375 40781 18457 40804
rect 18543 40781 18609 40804
rect 18223 40762 18609 40781
rect 33343 40867 33729 40886
rect 33343 40844 33409 40867
rect 33495 40844 33577 40867
rect 33663 40844 33729 40867
rect 33343 40804 33352 40844
rect 33392 40804 33409 40844
rect 33495 40804 33516 40844
rect 33556 40804 33577 40844
rect 33663 40804 33680 40844
rect 33720 40804 33729 40844
rect 33343 40781 33409 40804
rect 33495 40781 33577 40804
rect 33663 40781 33729 40804
rect 33343 40762 33729 40781
rect 48463 40867 48849 40886
rect 48463 40844 48529 40867
rect 48615 40844 48697 40867
rect 48783 40844 48849 40867
rect 48463 40804 48472 40844
rect 48512 40804 48529 40844
rect 48615 40804 48636 40844
rect 48676 40804 48697 40844
rect 48783 40804 48800 40844
rect 48840 40804 48849 40844
rect 48463 40781 48529 40804
rect 48615 40781 48697 40804
rect 48783 40781 48849 40804
rect 48463 40762 48849 40781
rect 63583 40867 63969 40886
rect 63583 40844 63649 40867
rect 63735 40844 63817 40867
rect 63903 40844 63969 40867
rect 63583 40804 63592 40844
rect 63632 40804 63649 40844
rect 63735 40804 63756 40844
rect 63796 40804 63817 40844
rect 63903 40804 63920 40844
rect 63960 40804 63969 40844
rect 63583 40781 63649 40804
rect 63735 40781 63817 40804
rect 63903 40781 63969 40804
rect 63583 40762 63969 40781
rect 78703 40867 79089 40886
rect 78703 40844 78769 40867
rect 78855 40844 78937 40867
rect 79023 40844 79089 40867
rect 78703 40804 78712 40844
rect 78752 40804 78769 40844
rect 78855 40804 78876 40844
rect 78916 40804 78937 40844
rect 79023 40804 79040 40844
rect 79080 40804 79089 40844
rect 78703 40781 78769 40804
rect 78855 40781 78937 40804
rect 79023 40781 79089 40804
rect 78703 40762 79089 40781
rect 93823 40867 94209 40886
rect 93823 40844 93889 40867
rect 93975 40844 94057 40867
rect 94143 40844 94209 40867
rect 93823 40804 93832 40844
rect 93872 40804 93889 40844
rect 93975 40804 93996 40844
rect 94036 40804 94057 40844
rect 94143 40804 94160 40844
rect 94200 40804 94209 40844
rect 93823 40781 93889 40804
rect 93975 40781 94057 40804
rect 94143 40781 94209 40804
rect 93823 40762 94209 40781
rect 4343 40111 4729 40130
rect 4343 40088 4409 40111
rect 4495 40088 4577 40111
rect 4663 40088 4729 40111
rect 4343 40048 4352 40088
rect 4392 40048 4409 40088
rect 4495 40048 4516 40088
rect 4556 40048 4577 40088
rect 4663 40048 4680 40088
rect 4720 40048 4729 40088
rect 4343 40025 4409 40048
rect 4495 40025 4577 40048
rect 4663 40025 4729 40048
rect 4343 40006 4729 40025
rect 19463 40111 19849 40130
rect 19463 40088 19529 40111
rect 19615 40088 19697 40111
rect 19783 40088 19849 40111
rect 19463 40048 19472 40088
rect 19512 40048 19529 40088
rect 19615 40048 19636 40088
rect 19676 40048 19697 40088
rect 19783 40048 19800 40088
rect 19840 40048 19849 40088
rect 19463 40025 19529 40048
rect 19615 40025 19697 40048
rect 19783 40025 19849 40048
rect 19463 40006 19849 40025
rect 34583 40111 34969 40130
rect 34583 40088 34649 40111
rect 34735 40088 34817 40111
rect 34903 40088 34969 40111
rect 34583 40048 34592 40088
rect 34632 40048 34649 40088
rect 34735 40048 34756 40088
rect 34796 40048 34817 40088
rect 34903 40048 34920 40088
rect 34960 40048 34969 40088
rect 34583 40025 34649 40048
rect 34735 40025 34817 40048
rect 34903 40025 34969 40048
rect 34583 40006 34969 40025
rect 49703 40111 50089 40130
rect 49703 40088 49769 40111
rect 49855 40088 49937 40111
rect 50023 40088 50089 40111
rect 49703 40048 49712 40088
rect 49752 40048 49769 40088
rect 49855 40048 49876 40088
rect 49916 40048 49937 40088
rect 50023 40048 50040 40088
rect 50080 40048 50089 40088
rect 49703 40025 49769 40048
rect 49855 40025 49937 40048
rect 50023 40025 50089 40048
rect 49703 40006 50089 40025
rect 64823 40111 65209 40130
rect 64823 40088 64889 40111
rect 64975 40088 65057 40111
rect 65143 40088 65209 40111
rect 64823 40048 64832 40088
rect 64872 40048 64889 40088
rect 64975 40048 64996 40088
rect 65036 40048 65057 40088
rect 65143 40048 65160 40088
rect 65200 40048 65209 40088
rect 64823 40025 64889 40048
rect 64975 40025 65057 40048
rect 65143 40025 65209 40048
rect 64823 40006 65209 40025
rect 79943 40111 80329 40130
rect 79943 40088 80009 40111
rect 80095 40088 80177 40111
rect 80263 40088 80329 40111
rect 79943 40048 79952 40088
rect 79992 40048 80009 40088
rect 80095 40048 80116 40088
rect 80156 40048 80177 40088
rect 80263 40048 80280 40088
rect 80320 40048 80329 40088
rect 79943 40025 80009 40048
rect 80095 40025 80177 40048
rect 80263 40025 80329 40048
rect 79943 40006 80329 40025
rect 95063 40111 95449 40130
rect 95063 40088 95129 40111
rect 95215 40088 95297 40111
rect 95383 40088 95449 40111
rect 95063 40048 95072 40088
rect 95112 40048 95129 40088
rect 95215 40048 95236 40088
rect 95276 40048 95297 40088
rect 95383 40048 95400 40088
rect 95440 40048 95449 40088
rect 95063 40025 95129 40048
rect 95215 40025 95297 40048
rect 95383 40025 95449 40048
rect 95063 40006 95449 40025
rect 3103 39355 3489 39374
rect 3103 39332 3169 39355
rect 3255 39332 3337 39355
rect 3423 39332 3489 39355
rect 3103 39292 3112 39332
rect 3152 39292 3169 39332
rect 3255 39292 3276 39332
rect 3316 39292 3337 39332
rect 3423 39292 3440 39332
rect 3480 39292 3489 39332
rect 3103 39269 3169 39292
rect 3255 39269 3337 39292
rect 3423 39269 3489 39292
rect 3103 39250 3489 39269
rect 18223 39355 18609 39374
rect 18223 39332 18289 39355
rect 18375 39332 18457 39355
rect 18543 39332 18609 39355
rect 18223 39292 18232 39332
rect 18272 39292 18289 39332
rect 18375 39292 18396 39332
rect 18436 39292 18457 39332
rect 18543 39292 18560 39332
rect 18600 39292 18609 39332
rect 18223 39269 18289 39292
rect 18375 39269 18457 39292
rect 18543 39269 18609 39292
rect 18223 39250 18609 39269
rect 33343 39355 33729 39374
rect 33343 39332 33409 39355
rect 33495 39332 33577 39355
rect 33663 39332 33729 39355
rect 33343 39292 33352 39332
rect 33392 39292 33409 39332
rect 33495 39292 33516 39332
rect 33556 39292 33577 39332
rect 33663 39292 33680 39332
rect 33720 39292 33729 39332
rect 33343 39269 33409 39292
rect 33495 39269 33577 39292
rect 33663 39269 33729 39292
rect 33343 39250 33729 39269
rect 48463 39355 48849 39374
rect 48463 39332 48529 39355
rect 48615 39332 48697 39355
rect 48783 39332 48849 39355
rect 48463 39292 48472 39332
rect 48512 39292 48529 39332
rect 48615 39292 48636 39332
rect 48676 39292 48697 39332
rect 48783 39292 48800 39332
rect 48840 39292 48849 39332
rect 48463 39269 48529 39292
rect 48615 39269 48697 39292
rect 48783 39269 48849 39292
rect 48463 39250 48849 39269
rect 63583 39355 63969 39374
rect 63583 39332 63649 39355
rect 63735 39332 63817 39355
rect 63903 39332 63969 39355
rect 63583 39292 63592 39332
rect 63632 39292 63649 39332
rect 63735 39292 63756 39332
rect 63796 39292 63817 39332
rect 63903 39292 63920 39332
rect 63960 39292 63969 39332
rect 63583 39269 63649 39292
rect 63735 39269 63817 39292
rect 63903 39269 63969 39292
rect 63583 39250 63969 39269
rect 78703 39355 79089 39374
rect 78703 39332 78769 39355
rect 78855 39332 78937 39355
rect 79023 39332 79089 39355
rect 78703 39292 78712 39332
rect 78752 39292 78769 39332
rect 78855 39292 78876 39332
rect 78916 39292 78937 39332
rect 79023 39292 79040 39332
rect 79080 39292 79089 39332
rect 78703 39269 78769 39292
rect 78855 39269 78937 39292
rect 79023 39269 79089 39292
rect 78703 39250 79089 39269
rect 93823 39355 94209 39374
rect 93823 39332 93889 39355
rect 93975 39332 94057 39355
rect 94143 39332 94209 39355
rect 93823 39292 93832 39332
rect 93872 39292 93889 39332
rect 93975 39292 93996 39332
rect 94036 39292 94057 39332
rect 94143 39292 94160 39332
rect 94200 39292 94209 39332
rect 93823 39269 93889 39292
rect 93975 39269 94057 39292
rect 94143 39269 94209 39292
rect 93823 39250 94209 39269
rect 4343 38599 4729 38618
rect 4343 38576 4409 38599
rect 4495 38576 4577 38599
rect 4663 38576 4729 38599
rect 4343 38536 4352 38576
rect 4392 38536 4409 38576
rect 4495 38536 4516 38576
rect 4556 38536 4577 38576
rect 4663 38536 4680 38576
rect 4720 38536 4729 38576
rect 4343 38513 4409 38536
rect 4495 38513 4577 38536
rect 4663 38513 4729 38536
rect 4343 38494 4729 38513
rect 19463 38599 19849 38618
rect 19463 38576 19529 38599
rect 19615 38576 19697 38599
rect 19783 38576 19849 38599
rect 19463 38536 19472 38576
rect 19512 38536 19529 38576
rect 19615 38536 19636 38576
rect 19676 38536 19697 38576
rect 19783 38536 19800 38576
rect 19840 38536 19849 38576
rect 19463 38513 19529 38536
rect 19615 38513 19697 38536
rect 19783 38513 19849 38536
rect 19463 38494 19849 38513
rect 34583 38599 34969 38618
rect 34583 38576 34649 38599
rect 34735 38576 34817 38599
rect 34903 38576 34969 38599
rect 34583 38536 34592 38576
rect 34632 38536 34649 38576
rect 34735 38536 34756 38576
rect 34796 38536 34817 38576
rect 34903 38536 34920 38576
rect 34960 38536 34969 38576
rect 34583 38513 34649 38536
rect 34735 38513 34817 38536
rect 34903 38513 34969 38536
rect 34583 38494 34969 38513
rect 49703 38599 50089 38618
rect 49703 38576 49769 38599
rect 49855 38576 49937 38599
rect 50023 38576 50089 38599
rect 49703 38536 49712 38576
rect 49752 38536 49769 38576
rect 49855 38536 49876 38576
rect 49916 38536 49937 38576
rect 50023 38536 50040 38576
rect 50080 38536 50089 38576
rect 49703 38513 49769 38536
rect 49855 38513 49937 38536
rect 50023 38513 50089 38536
rect 49703 38494 50089 38513
rect 64823 38599 65209 38618
rect 64823 38576 64889 38599
rect 64975 38576 65057 38599
rect 65143 38576 65209 38599
rect 64823 38536 64832 38576
rect 64872 38536 64889 38576
rect 64975 38536 64996 38576
rect 65036 38536 65057 38576
rect 65143 38536 65160 38576
rect 65200 38536 65209 38576
rect 64823 38513 64889 38536
rect 64975 38513 65057 38536
rect 65143 38513 65209 38536
rect 64823 38494 65209 38513
rect 79943 38599 80329 38618
rect 79943 38576 80009 38599
rect 80095 38576 80177 38599
rect 80263 38576 80329 38599
rect 79943 38536 79952 38576
rect 79992 38536 80009 38576
rect 80095 38536 80116 38576
rect 80156 38536 80177 38576
rect 80263 38536 80280 38576
rect 80320 38536 80329 38576
rect 79943 38513 80009 38536
rect 80095 38513 80177 38536
rect 80263 38513 80329 38536
rect 79943 38494 80329 38513
rect 95063 38599 95449 38618
rect 95063 38576 95129 38599
rect 95215 38576 95297 38599
rect 95383 38576 95449 38599
rect 95063 38536 95072 38576
rect 95112 38536 95129 38576
rect 95215 38536 95236 38576
rect 95276 38536 95297 38576
rect 95383 38536 95400 38576
rect 95440 38536 95449 38576
rect 95063 38513 95129 38536
rect 95215 38513 95297 38536
rect 95383 38513 95449 38536
rect 95063 38494 95449 38513
rect 3103 37843 3489 37862
rect 3103 37820 3169 37843
rect 3255 37820 3337 37843
rect 3423 37820 3489 37843
rect 3103 37780 3112 37820
rect 3152 37780 3169 37820
rect 3255 37780 3276 37820
rect 3316 37780 3337 37820
rect 3423 37780 3440 37820
rect 3480 37780 3489 37820
rect 3103 37757 3169 37780
rect 3255 37757 3337 37780
rect 3423 37757 3489 37780
rect 3103 37738 3489 37757
rect 18223 37843 18609 37862
rect 18223 37820 18289 37843
rect 18375 37820 18457 37843
rect 18543 37820 18609 37843
rect 18223 37780 18232 37820
rect 18272 37780 18289 37820
rect 18375 37780 18396 37820
rect 18436 37780 18457 37820
rect 18543 37780 18560 37820
rect 18600 37780 18609 37820
rect 18223 37757 18289 37780
rect 18375 37757 18457 37780
rect 18543 37757 18609 37780
rect 18223 37738 18609 37757
rect 33343 37843 33729 37862
rect 33343 37820 33409 37843
rect 33495 37820 33577 37843
rect 33663 37820 33729 37843
rect 33343 37780 33352 37820
rect 33392 37780 33409 37820
rect 33495 37780 33516 37820
rect 33556 37780 33577 37820
rect 33663 37780 33680 37820
rect 33720 37780 33729 37820
rect 33343 37757 33409 37780
rect 33495 37757 33577 37780
rect 33663 37757 33729 37780
rect 33343 37738 33729 37757
rect 48463 37843 48849 37862
rect 48463 37820 48529 37843
rect 48615 37820 48697 37843
rect 48783 37820 48849 37843
rect 48463 37780 48472 37820
rect 48512 37780 48529 37820
rect 48615 37780 48636 37820
rect 48676 37780 48697 37820
rect 48783 37780 48800 37820
rect 48840 37780 48849 37820
rect 48463 37757 48529 37780
rect 48615 37757 48697 37780
rect 48783 37757 48849 37780
rect 48463 37738 48849 37757
rect 63583 37843 63969 37862
rect 63583 37820 63649 37843
rect 63735 37820 63817 37843
rect 63903 37820 63969 37843
rect 63583 37780 63592 37820
rect 63632 37780 63649 37820
rect 63735 37780 63756 37820
rect 63796 37780 63817 37820
rect 63903 37780 63920 37820
rect 63960 37780 63969 37820
rect 63583 37757 63649 37780
rect 63735 37757 63817 37780
rect 63903 37757 63969 37780
rect 63583 37738 63969 37757
rect 78703 37843 79089 37862
rect 78703 37820 78769 37843
rect 78855 37820 78937 37843
rect 79023 37820 79089 37843
rect 78703 37780 78712 37820
rect 78752 37780 78769 37820
rect 78855 37780 78876 37820
rect 78916 37780 78937 37820
rect 79023 37780 79040 37820
rect 79080 37780 79089 37820
rect 78703 37757 78769 37780
rect 78855 37757 78937 37780
rect 79023 37757 79089 37780
rect 78703 37738 79089 37757
rect 93823 37843 94209 37862
rect 93823 37820 93889 37843
rect 93975 37820 94057 37843
rect 94143 37820 94209 37843
rect 93823 37780 93832 37820
rect 93872 37780 93889 37820
rect 93975 37780 93996 37820
rect 94036 37780 94057 37820
rect 94143 37780 94160 37820
rect 94200 37780 94209 37820
rect 93823 37757 93889 37780
rect 93975 37757 94057 37780
rect 94143 37757 94209 37780
rect 93823 37738 94209 37757
rect 4343 37087 4729 37106
rect 4343 37064 4409 37087
rect 4495 37064 4577 37087
rect 4663 37064 4729 37087
rect 4343 37024 4352 37064
rect 4392 37024 4409 37064
rect 4495 37024 4516 37064
rect 4556 37024 4577 37064
rect 4663 37024 4680 37064
rect 4720 37024 4729 37064
rect 4343 37001 4409 37024
rect 4495 37001 4577 37024
rect 4663 37001 4729 37024
rect 4343 36982 4729 37001
rect 19463 37087 19849 37106
rect 19463 37064 19529 37087
rect 19615 37064 19697 37087
rect 19783 37064 19849 37087
rect 19463 37024 19472 37064
rect 19512 37024 19529 37064
rect 19615 37024 19636 37064
rect 19676 37024 19697 37064
rect 19783 37024 19800 37064
rect 19840 37024 19849 37064
rect 19463 37001 19529 37024
rect 19615 37001 19697 37024
rect 19783 37001 19849 37024
rect 19463 36982 19849 37001
rect 34583 37087 34969 37106
rect 34583 37064 34649 37087
rect 34735 37064 34817 37087
rect 34903 37064 34969 37087
rect 34583 37024 34592 37064
rect 34632 37024 34649 37064
rect 34735 37024 34756 37064
rect 34796 37024 34817 37064
rect 34903 37024 34920 37064
rect 34960 37024 34969 37064
rect 34583 37001 34649 37024
rect 34735 37001 34817 37024
rect 34903 37001 34969 37024
rect 34583 36982 34969 37001
rect 49703 37087 50089 37106
rect 49703 37064 49769 37087
rect 49855 37064 49937 37087
rect 50023 37064 50089 37087
rect 49703 37024 49712 37064
rect 49752 37024 49769 37064
rect 49855 37024 49876 37064
rect 49916 37024 49937 37064
rect 50023 37024 50040 37064
rect 50080 37024 50089 37064
rect 49703 37001 49769 37024
rect 49855 37001 49937 37024
rect 50023 37001 50089 37024
rect 49703 36982 50089 37001
rect 64823 37087 65209 37106
rect 64823 37064 64889 37087
rect 64975 37064 65057 37087
rect 65143 37064 65209 37087
rect 64823 37024 64832 37064
rect 64872 37024 64889 37064
rect 64975 37024 64996 37064
rect 65036 37024 65057 37064
rect 65143 37024 65160 37064
rect 65200 37024 65209 37064
rect 64823 37001 64889 37024
rect 64975 37001 65057 37024
rect 65143 37001 65209 37024
rect 64823 36982 65209 37001
rect 79943 37087 80329 37106
rect 79943 37064 80009 37087
rect 80095 37064 80177 37087
rect 80263 37064 80329 37087
rect 79943 37024 79952 37064
rect 79992 37024 80009 37064
rect 80095 37024 80116 37064
rect 80156 37024 80177 37064
rect 80263 37024 80280 37064
rect 80320 37024 80329 37064
rect 79943 37001 80009 37024
rect 80095 37001 80177 37024
rect 80263 37001 80329 37024
rect 79943 36982 80329 37001
rect 95063 37087 95449 37106
rect 95063 37064 95129 37087
rect 95215 37064 95297 37087
rect 95383 37064 95449 37087
rect 95063 37024 95072 37064
rect 95112 37024 95129 37064
rect 95215 37024 95236 37064
rect 95276 37024 95297 37064
rect 95383 37024 95400 37064
rect 95440 37024 95449 37064
rect 95063 37001 95129 37024
rect 95215 37001 95297 37024
rect 95383 37001 95449 37024
rect 95063 36982 95449 37001
rect 3103 36331 3489 36350
rect 3103 36308 3169 36331
rect 3255 36308 3337 36331
rect 3423 36308 3489 36331
rect 3103 36268 3112 36308
rect 3152 36268 3169 36308
rect 3255 36268 3276 36308
rect 3316 36268 3337 36308
rect 3423 36268 3440 36308
rect 3480 36268 3489 36308
rect 3103 36245 3169 36268
rect 3255 36245 3337 36268
rect 3423 36245 3489 36268
rect 3103 36226 3489 36245
rect 18223 36331 18609 36350
rect 18223 36308 18289 36331
rect 18375 36308 18457 36331
rect 18543 36308 18609 36331
rect 18223 36268 18232 36308
rect 18272 36268 18289 36308
rect 18375 36268 18396 36308
rect 18436 36268 18457 36308
rect 18543 36268 18560 36308
rect 18600 36268 18609 36308
rect 18223 36245 18289 36268
rect 18375 36245 18457 36268
rect 18543 36245 18609 36268
rect 18223 36226 18609 36245
rect 33343 36331 33729 36350
rect 33343 36308 33409 36331
rect 33495 36308 33577 36331
rect 33663 36308 33729 36331
rect 33343 36268 33352 36308
rect 33392 36268 33409 36308
rect 33495 36268 33516 36308
rect 33556 36268 33577 36308
rect 33663 36268 33680 36308
rect 33720 36268 33729 36308
rect 33343 36245 33409 36268
rect 33495 36245 33577 36268
rect 33663 36245 33729 36268
rect 33343 36226 33729 36245
rect 48463 36331 48849 36350
rect 48463 36308 48529 36331
rect 48615 36308 48697 36331
rect 48783 36308 48849 36331
rect 48463 36268 48472 36308
rect 48512 36268 48529 36308
rect 48615 36268 48636 36308
rect 48676 36268 48697 36308
rect 48783 36268 48800 36308
rect 48840 36268 48849 36308
rect 48463 36245 48529 36268
rect 48615 36245 48697 36268
rect 48783 36245 48849 36268
rect 48463 36226 48849 36245
rect 63583 36331 63969 36350
rect 63583 36308 63649 36331
rect 63735 36308 63817 36331
rect 63903 36308 63969 36331
rect 63583 36268 63592 36308
rect 63632 36268 63649 36308
rect 63735 36268 63756 36308
rect 63796 36268 63817 36308
rect 63903 36268 63920 36308
rect 63960 36268 63969 36308
rect 63583 36245 63649 36268
rect 63735 36245 63817 36268
rect 63903 36245 63969 36268
rect 63583 36226 63969 36245
rect 78703 36331 79089 36350
rect 78703 36308 78769 36331
rect 78855 36308 78937 36331
rect 79023 36308 79089 36331
rect 78703 36268 78712 36308
rect 78752 36268 78769 36308
rect 78855 36268 78876 36308
rect 78916 36268 78937 36308
rect 79023 36268 79040 36308
rect 79080 36268 79089 36308
rect 78703 36245 78769 36268
rect 78855 36245 78937 36268
rect 79023 36245 79089 36268
rect 78703 36226 79089 36245
rect 93823 36331 94209 36350
rect 93823 36308 93889 36331
rect 93975 36308 94057 36331
rect 94143 36308 94209 36331
rect 93823 36268 93832 36308
rect 93872 36268 93889 36308
rect 93975 36268 93996 36308
rect 94036 36268 94057 36308
rect 94143 36268 94160 36308
rect 94200 36268 94209 36308
rect 93823 36245 93889 36268
rect 93975 36245 94057 36268
rect 94143 36245 94209 36268
rect 93823 36226 94209 36245
rect 4343 35575 4729 35594
rect 4343 35552 4409 35575
rect 4495 35552 4577 35575
rect 4663 35552 4729 35575
rect 4343 35512 4352 35552
rect 4392 35512 4409 35552
rect 4495 35512 4516 35552
rect 4556 35512 4577 35552
rect 4663 35512 4680 35552
rect 4720 35512 4729 35552
rect 4343 35489 4409 35512
rect 4495 35489 4577 35512
rect 4663 35489 4729 35512
rect 4343 35470 4729 35489
rect 19463 35575 19849 35594
rect 19463 35552 19529 35575
rect 19615 35552 19697 35575
rect 19783 35552 19849 35575
rect 19463 35512 19472 35552
rect 19512 35512 19529 35552
rect 19615 35512 19636 35552
rect 19676 35512 19697 35552
rect 19783 35512 19800 35552
rect 19840 35512 19849 35552
rect 19463 35489 19529 35512
rect 19615 35489 19697 35512
rect 19783 35489 19849 35512
rect 19463 35470 19849 35489
rect 34583 35575 34969 35594
rect 34583 35552 34649 35575
rect 34735 35552 34817 35575
rect 34903 35552 34969 35575
rect 34583 35512 34592 35552
rect 34632 35512 34649 35552
rect 34735 35512 34756 35552
rect 34796 35512 34817 35552
rect 34903 35512 34920 35552
rect 34960 35512 34969 35552
rect 34583 35489 34649 35512
rect 34735 35489 34817 35512
rect 34903 35489 34969 35512
rect 34583 35470 34969 35489
rect 49703 35575 50089 35594
rect 49703 35552 49769 35575
rect 49855 35552 49937 35575
rect 50023 35552 50089 35575
rect 49703 35512 49712 35552
rect 49752 35512 49769 35552
rect 49855 35512 49876 35552
rect 49916 35512 49937 35552
rect 50023 35512 50040 35552
rect 50080 35512 50089 35552
rect 49703 35489 49769 35512
rect 49855 35489 49937 35512
rect 50023 35489 50089 35512
rect 49703 35470 50089 35489
rect 64823 35575 65209 35594
rect 64823 35552 64889 35575
rect 64975 35552 65057 35575
rect 65143 35552 65209 35575
rect 64823 35512 64832 35552
rect 64872 35512 64889 35552
rect 64975 35512 64996 35552
rect 65036 35512 65057 35552
rect 65143 35512 65160 35552
rect 65200 35512 65209 35552
rect 64823 35489 64889 35512
rect 64975 35489 65057 35512
rect 65143 35489 65209 35512
rect 64823 35470 65209 35489
rect 79943 35575 80329 35594
rect 79943 35552 80009 35575
rect 80095 35552 80177 35575
rect 80263 35552 80329 35575
rect 79943 35512 79952 35552
rect 79992 35512 80009 35552
rect 80095 35512 80116 35552
rect 80156 35512 80177 35552
rect 80263 35512 80280 35552
rect 80320 35512 80329 35552
rect 79943 35489 80009 35512
rect 80095 35489 80177 35512
rect 80263 35489 80329 35512
rect 79943 35470 80329 35489
rect 95063 35575 95449 35594
rect 95063 35552 95129 35575
rect 95215 35552 95297 35575
rect 95383 35552 95449 35575
rect 95063 35512 95072 35552
rect 95112 35512 95129 35552
rect 95215 35512 95236 35552
rect 95276 35512 95297 35552
rect 95383 35512 95400 35552
rect 95440 35512 95449 35552
rect 95063 35489 95129 35512
rect 95215 35489 95297 35512
rect 95383 35489 95449 35512
rect 95063 35470 95449 35489
rect 3103 34819 3489 34838
rect 3103 34796 3169 34819
rect 3255 34796 3337 34819
rect 3423 34796 3489 34819
rect 3103 34756 3112 34796
rect 3152 34756 3169 34796
rect 3255 34756 3276 34796
rect 3316 34756 3337 34796
rect 3423 34756 3440 34796
rect 3480 34756 3489 34796
rect 3103 34733 3169 34756
rect 3255 34733 3337 34756
rect 3423 34733 3489 34756
rect 3103 34714 3489 34733
rect 18223 34819 18609 34838
rect 18223 34796 18289 34819
rect 18375 34796 18457 34819
rect 18543 34796 18609 34819
rect 18223 34756 18232 34796
rect 18272 34756 18289 34796
rect 18375 34756 18396 34796
rect 18436 34756 18457 34796
rect 18543 34756 18560 34796
rect 18600 34756 18609 34796
rect 18223 34733 18289 34756
rect 18375 34733 18457 34756
rect 18543 34733 18609 34756
rect 18223 34714 18609 34733
rect 33343 34819 33729 34838
rect 33343 34796 33409 34819
rect 33495 34796 33577 34819
rect 33663 34796 33729 34819
rect 33343 34756 33352 34796
rect 33392 34756 33409 34796
rect 33495 34756 33516 34796
rect 33556 34756 33577 34796
rect 33663 34756 33680 34796
rect 33720 34756 33729 34796
rect 33343 34733 33409 34756
rect 33495 34733 33577 34756
rect 33663 34733 33729 34756
rect 33343 34714 33729 34733
rect 48463 34819 48849 34838
rect 48463 34796 48529 34819
rect 48615 34796 48697 34819
rect 48783 34796 48849 34819
rect 48463 34756 48472 34796
rect 48512 34756 48529 34796
rect 48615 34756 48636 34796
rect 48676 34756 48697 34796
rect 48783 34756 48800 34796
rect 48840 34756 48849 34796
rect 48463 34733 48529 34756
rect 48615 34733 48697 34756
rect 48783 34733 48849 34756
rect 48463 34714 48849 34733
rect 63583 34819 63969 34838
rect 63583 34796 63649 34819
rect 63735 34796 63817 34819
rect 63903 34796 63969 34819
rect 63583 34756 63592 34796
rect 63632 34756 63649 34796
rect 63735 34756 63756 34796
rect 63796 34756 63817 34796
rect 63903 34756 63920 34796
rect 63960 34756 63969 34796
rect 63583 34733 63649 34756
rect 63735 34733 63817 34756
rect 63903 34733 63969 34756
rect 63583 34714 63969 34733
rect 78703 34819 79089 34838
rect 78703 34796 78769 34819
rect 78855 34796 78937 34819
rect 79023 34796 79089 34819
rect 78703 34756 78712 34796
rect 78752 34756 78769 34796
rect 78855 34756 78876 34796
rect 78916 34756 78937 34796
rect 79023 34756 79040 34796
rect 79080 34756 79089 34796
rect 78703 34733 78769 34756
rect 78855 34733 78937 34756
rect 79023 34733 79089 34756
rect 78703 34714 79089 34733
rect 93823 34819 94209 34838
rect 93823 34796 93889 34819
rect 93975 34796 94057 34819
rect 94143 34796 94209 34819
rect 93823 34756 93832 34796
rect 93872 34756 93889 34796
rect 93975 34756 93996 34796
rect 94036 34756 94057 34796
rect 94143 34756 94160 34796
rect 94200 34756 94209 34796
rect 93823 34733 93889 34756
rect 93975 34733 94057 34756
rect 94143 34733 94209 34756
rect 93823 34714 94209 34733
rect 4343 34063 4729 34082
rect 4343 34040 4409 34063
rect 4495 34040 4577 34063
rect 4663 34040 4729 34063
rect 4343 34000 4352 34040
rect 4392 34000 4409 34040
rect 4495 34000 4516 34040
rect 4556 34000 4577 34040
rect 4663 34000 4680 34040
rect 4720 34000 4729 34040
rect 4343 33977 4409 34000
rect 4495 33977 4577 34000
rect 4663 33977 4729 34000
rect 4343 33958 4729 33977
rect 19463 34063 19849 34082
rect 19463 34040 19529 34063
rect 19615 34040 19697 34063
rect 19783 34040 19849 34063
rect 19463 34000 19472 34040
rect 19512 34000 19529 34040
rect 19615 34000 19636 34040
rect 19676 34000 19697 34040
rect 19783 34000 19800 34040
rect 19840 34000 19849 34040
rect 19463 33977 19529 34000
rect 19615 33977 19697 34000
rect 19783 33977 19849 34000
rect 19463 33958 19849 33977
rect 34583 34063 34969 34082
rect 34583 34040 34649 34063
rect 34735 34040 34817 34063
rect 34903 34040 34969 34063
rect 34583 34000 34592 34040
rect 34632 34000 34649 34040
rect 34735 34000 34756 34040
rect 34796 34000 34817 34040
rect 34903 34000 34920 34040
rect 34960 34000 34969 34040
rect 34583 33977 34649 34000
rect 34735 33977 34817 34000
rect 34903 33977 34969 34000
rect 34583 33958 34969 33977
rect 49703 34063 50089 34082
rect 49703 34040 49769 34063
rect 49855 34040 49937 34063
rect 50023 34040 50089 34063
rect 49703 34000 49712 34040
rect 49752 34000 49769 34040
rect 49855 34000 49876 34040
rect 49916 34000 49937 34040
rect 50023 34000 50040 34040
rect 50080 34000 50089 34040
rect 49703 33977 49769 34000
rect 49855 33977 49937 34000
rect 50023 33977 50089 34000
rect 49703 33958 50089 33977
rect 64823 34063 65209 34082
rect 64823 34040 64889 34063
rect 64975 34040 65057 34063
rect 65143 34040 65209 34063
rect 64823 34000 64832 34040
rect 64872 34000 64889 34040
rect 64975 34000 64996 34040
rect 65036 34000 65057 34040
rect 65143 34000 65160 34040
rect 65200 34000 65209 34040
rect 64823 33977 64889 34000
rect 64975 33977 65057 34000
rect 65143 33977 65209 34000
rect 64823 33958 65209 33977
rect 79943 34063 80329 34082
rect 79943 34040 80009 34063
rect 80095 34040 80177 34063
rect 80263 34040 80329 34063
rect 79943 34000 79952 34040
rect 79992 34000 80009 34040
rect 80095 34000 80116 34040
rect 80156 34000 80177 34040
rect 80263 34000 80280 34040
rect 80320 34000 80329 34040
rect 79943 33977 80009 34000
rect 80095 33977 80177 34000
rect 80263 33977 80329 34000
rect 79943 33958 80329 33977
rect 95063 34063 95449 34082
rect 95063 34040 95129 34063
rect 95215 34040 95297 34063
rect 95383 34040 95449 34063
rect 95063 34000 95072 34040
rect 95112 34000 95129 34040
rect 95215 34000 95236 34040
rect 95276 34000 95297 34040
rect 95383 34000 95400 34040
rect 95440 34000 95449 34040
rect 95063 33977 95129 34000
rect 95215 33977 95297 34000
rect 95383 33977 95449 34000
rect 95063 33958 95449 33977
rect 3103 33307 3489 33326
rect 3103 33284 3169 33307
rect 3255 33284 3337 33307
rect 3423 33284 3489 33307
rect 3103 33244 3112 33284
rect 3152 33244 3169 33284
rect 3255 33244 3276 33284
rect 3316 33244 3337 33284
rect 3423 33244 3440 33284
rect 3480 33244 3489 33284
rect 3103 33221 3169 33244
rect 3255 33221 3337 33244
rect 3423 33221 3489 33244
rect 3103 33202 3489 33221
rect 18223 33307 18609 33326
rect 18223 33284 18289 33307
rect 18375 33284 18457 33307
rect 18543 33284 18609 33307
rect 18223 33244 18232 33284
rect 18272 33244 18289 33284
rect 18375 33244 18396 33284
rect 18436 33244 18457 33284
rect 18543 33244 18560 33284
rect 18600 33244 18609 33284
rect 18223 33221 18289 33244
rect 18375 33221 18457 33244
rect 18543 33221 18609 33244
rect 18223 33202 18609 33221
rect 33343 33307 33729 33326
rect 33343 33284 33409 33307
rect 33495 33284 33577 33307
rect 33663 33284 33729 33307
rect 33343 33244 33352 33284
rect 33392 33244 33409 33284
rect 33495 33244 33516 33284
rect 33556 33244 33577 33284
rect 33663 33244 33680 33284
rect 33720 33244 33729 33284
rect 33343 33221 33409 33244
rect 33495 33221 33577 33244
rect 33663 33221 33729 33244
rect 33343 33202 33729 33221
rect 48463 33307 48849 33326
rect 48463 33284 48529 33307
rect 48615 33284 48697 33307
rect 48783 33284 48849 33307
rect 48463 33244 48472 33284
rect 48512 33244 48529 33284
rect 48615 33244 48636 33284
rect 48676 33244 48697 33284
rect 48783 33244 48800 33284
rect 48840 33244 48849 33284
rect 48463 33221 48529 33244
rect 48615 33221 48697 33244
rect 48783 33221 48849 33244
rect 48463 33202 48849 33221
rect 63583 33307 63969 33326
rect 63583 33284 63649 33307
rect 63735 33284 63817 33307
rect 63903 33284 63969 33307
rect 63583 33244 63592 33284
rect 63632 33244 63649 33284
rect 63735 33244 63756 33284
rect 63796 33244 63817 33284
rect 63903 33244 63920 33284
rect 63960 33244 63969 33284
rect 63583 33221 63649 33244
rect 63735 33221 63817 33244
rect 63903 33221 63969 33244
rect 63583 33202 63969 33221
rect 78703 33307 79089 33326
rect 78703 33284 78769 33307
rect 78855 33284 78937 33307
rect 79023 33284 79089 33307
rect 78703 33244 78712 33284
rect 78752 33244 78769 33284
rect 78855 33244 78876 33284
rect 78916 33244 78937 33284
rect 79023 33244 79040 33284
rect 79080 33244 79089 33284
rect 78703 33221 78769 33244
rect 78855 33221 78937 33244
rect 79023 33221 79089 33244
rect 78703 33202 79089 33221
rect 93823 33307 94209 33326
rect 93823 33284 93889 33307
rect 93975 33284 94057 33307
rect 94143 33284 94209 33307
rect 93823 33244 93832 33284
rect 93872 33244 93889 33284
rect 93975 33244 93996 33284
rect 94036 33244 94057 33284
rect 94143 33244 94160 33284
rect 94200 33244 94209 33284
rect 93823 33221 93889 33244
rect 93975 33221 94057 33244
rect 94143 33221 94209 33244
rect 93823 33202 94209 33221
rect 4343 32551 4729 32570
rect 4343 32528 4409 32551
rect 4495 32528 4577 32551
rect 4663 32528 4729 32551
rect 4343 32488 4352 32528
rect 4392 32488 4409 32528
rect 4495 32488 4516 32528
rect 4556 32488 4577 32528
rect 4663 32488 4680 32528
rect 4720 32488 4729 32528
rect 4343 32465 4409 32488
rect 4495 32465 4577 32488
rect 4663 32465 4729 32488
rect 4343 32446 4729 32465
rect 19463 32551 19849 32570
rect 19463 32528 19529 32551
rect 19615 32528 19697 32551
rect 19783 32528 19849 32551
rect 19463 32488 19472 32528
rect 19512 32488 19529 32528
rect 19615 32488 19636 32528
rect 19676 32488 19697 32528
rect 19783 32488 19800 32528
rect 19840 32488 19849 32528
rect 19463 32465 19529 32488
rect 19615 32465 19697 32488
rect 19783 32465 19849 32488
rect 19463 32446 19849 32465
rect 34583 32551 34969 32570
rect 34583 32528 34649 32551
rect 34735 32528 34817 32551
rect 34903 32528 34969 32551
rect 34583 32488 34592 32528
rect 34632 32488 34649 32528
rect 34735 32488 34756 32528
rect 34796 32488 34817 32528
rect 34903 32488 34920 32528
rect 34960 32488 34969 32528
rect 34583 32465 34649 32488
rect 34735 32465 34817 32488
rect 34903 32465 34969 32488
rect 34583 32446 34969 32465
rect 49703 32551 50089 32570
rect 49703 32528 49769 32551
rect 49855 32528 49937 32551
rect 50023 32528 50089 32551
rect 49703 32488 49712 32528
rect 49752 32488 49769 32528
rect 49855 32488 49876 32528
rect 49916 32488 49937 32528
rect 50023 32488 50040 32528
rect 50080 32488 50089 32528
rect 49703 32465 49769 32488
rect 49855 32465 49937 32488
rect 50023 32465 50089 32488
rect 49703 32446 50089 32465
rect 64823 32551 65209 32570
rect 64823 32528 64889 32551
rect 64975 32528 65057 32551
rect 65143 32528 65209 32551
rect 64823 32488 64832 32528
rect 64872 32488 64889 32528
rect 64975 32488 64996 32528
rect 65036 32488 65057 32528
rect 65143 32488 65160 32528
rect 65200 32488 65209 32528
rect 64823 32465 64889 32488
rect 64975 32465 65057 32488
rect 65143 32465 65209 32488
rect 64823 32446 65209 32465
rect 79943 32551 80329 32570
rect 79943 32528 80009 32551
rect 80095 32528 80177 32551
rect 80263 32528 80329 32551
rect 79943 32488 79952 32528
rect 79992 32488 80009 32528
rect 80095 32488 80116 32528
rect 80156 32488 80177 32528
rect 80263 32488 80280 32528
rect 80320 32488 80329 32528
rect 79943 32465 80009 32488
rect 80095 32465 80177 32488
rect 80263 32465 80329 32488
rect 79943 32446 80329 32465
rect 95063 32551 95449 32570
rect 95063 32528 95129 32551
rect 95215 32528 95297 32551
rect 95383 32528 95449 32551
rect 95063 32488 95072 32528
rect 95112 32488 95129 32528
rect 95215 32488 95236 32528
rect 95276 32488 95297 32528
rect 95383 32488 95400 32528
rect 95440 32488 95449 32528
rect 95063 32465 95129 32488
rect 95215 32465 95297 32488
rect 95383 32465 95449 32488
rect 95063 32446 95449 32465
rect 3103 31795 3489 31814
rect 3103 31772 3169 31795
rect 3255 31772 3337 31795
rect 3423 31772 3489 31795
rect 3103 31732 3112 31772
rect 3152 31732 3169 31772
rect 3255 31732 3276 31772
rect 3316 31732 3337 31772
rect 3423 31732 3440 31772
rect 3480 31732 3489 31772
rect 3103 31709 3169 31732
rect 3255 31709 3337 31732
rect 3423 31709 3489 31732
rect 3103 31690 3489 31709
rect 18223 31795 18609 31814
rect 18223 31772 18289 31795
rect 18375 31772 18457 31795
rect 18543 31772 18609 31795
rect 18223 31732 18232 31772
rect 18272 31732 18289 31772
rect 18375 31732 18396 31772
rect 18436 31732 18457 31772
rect 18543 31732 18560 31772
rect 18600 31732 18609 31772
rect 18223 31709 18289 31732
rect 18375 31709 18457 31732
rect 18543 31709 18609 31732
rect 18223 31690 18609 31709
rect 33343 31795 33729 31814
rect 33343 31772 33409 31795
rect 33495 31772 33577 31795
rect 33663 31772 33729 31795
rect 33343 31732 33352 31772
rect 33392 31732 33409 31772
rect 33495 31732 33516 31772
rect 33556 31732 33577 31772
rect 33663 31732 33680 31772
rect 33720 31732 33729 31772
rect 33343 31709 33409 31732
rect 33495 31709 33577 31732
rect 33663 31709 33729 31732
rect 33343 31690 33729 31709
rect 48463 31795 48849 31814
rect 48463 31772 48529 31795
rect 48615 31772 48697 31795
rect 48783 31772 48849 31795
rect 48463 31732 48472 31772
rect 48512 31732 48529 31772
rect 48615 31732 48636 31772
rect 48676 31732 48697 31772
rect 48783 31732 48800 31772
rect 48840 31732 48849 31772
rect 48463 31709 48529 31732
rect 48615 31709 48697 31732
rect 48783 31709 48849 31732
rect 48463 31690 48849 31709
rect 63583 31795 63969 31814
rect 63583 31772 63649 31795
rect 63735 31772 63817 31795
rect 63903 31772 63969 31795
rect 63583 31732 63592 31772
rect 63632 31732 63649 31772
rect 63735 31732 63756 31772
rect 63796 31732 63817 31772
rect 63903 31732 63920 31772
rect 63960 31732 63969 31772
rect 63583 31709 63649 31732
rect 63735 31709 63817 31732
rect 63903 31709 63969 31732
rect 63583 31690 63969 31709
rect 78703 31795 79089 31814
rect 78703 31772 78769 31795
rect 78855 31772 78937 31795
rect 79023 31772 79089 31795
rect 78703 31732 78712 31772
rect 78752 31732 78769 31772
rect 78855 31732 78876 31772
rect 78916 31732 78937 31772
rect 79023 31732 79040 31772
rect 79080 31732 79089 31772
rect 78703 31709 78769 31732
rect 78855 31709 78937 31732
rect 79023 31709 79089 31732
rect 78703 31690 79089 31709
rect 93823 31795 94209 31814
rect 93823 31772 93889 31795
rect 93975 31772 94057 31795
rect 94143 31772 94209 31795
rect 93823 31732 93832 31772
rect 93872 31732 93889 31772
rect 93975 31732 93996 31772
rect 94036 31732 94057 31772
rect 94143 31732 94160 31772
rect 94200 31732 94209 31772
rect 93823 31709 93889 31732
rect 93975 31709 94057 31732
rect 94143 31709 94209 31732
rect 93823 31690 94209 31709
rect 4343 31039 4729 31058
rect 4343 31016 4409 31039
rect 4495 31016 4577 31039
rect 4663 31016 4729 31039
rect 4343 30976 4352 31016
rect 4392 30976 4409 31016
rect 4495 30976 4516 31016
rect 4556 30976 4577 31016
rect 4663 30976 4680 31016
rect 4720 30976 4729 31016
rect 4343 30953 4409 30976
rect 4495 30953 4577 30976
rect 4663 30953 4729 30976
rect 4343 30934 4729 30953
rect 19463 31039 19849 31058
rect 19463 31016 19529 31039
rect 19615 31016 19697 31039
rect 19783 31016 19849 31039
rect 19463 30976 19472 31016
rect 19512 30976 19529 31016
rect 19615 30976 19636 31016
rect 19676 30976 19697 31016
rect 19783 30976 19800 31016
rect 19840 30976 19849 31016
rect 19463 30953 19529 30976
rect 19615 30953 19697 30976
rect 19783 30953 19849 30976
rect 19463 30934 19849 30953
rect 34583 31039 34969 31058
rect 34583 31016 34649 31039
rect 34735 31016 34817 31039
rect 34903 31016 34969 31039
rect 34583 30976 34592 31016
rect 34632 30976 34649 31016
rect 34735 30976 34756 31016
rect 34796 30976 34817 31016
rect 34903 30976 34920 31016
rect 34960 30976 34969 31016
rect 34583 30953 34649 30976
rect 34735 30953 34817 30976
rect 34903 30953 34969 30976
rect 34583 30934 34969 30953
rect 49703 31039 50089 31058
rect 49703 31016 49769 31039
rect 49855 31016 49937 31039
rect 50023 31016 50089 31039
rect 49703 30976 49712 31016
rect 49752 30976 49769 31016
rect 49855 30976 49876 31016
rect 49916 30976 49937 31016
rect 50023 30976 50040 31016
rect 50080 30976 50089 31016
rect 49703 30953 49769 30976
rect 49855 30953 49937 30976
rect 50023 30953 50089 30976
rect 49703 30934 50089 30953
rect 64823 31039 65209 31058
rect 64823 31016 64889 31039
rect 64975 31016 65057 31039
rect 65143 31016 65209 31039
rect 64823 30976 64832 31016
rect 64872 30976 64889 31016
rect 64975 30976 64996 31016
rect 65036 30976 65057 31016
rect 65143 30976 65160 31016
rect 65200 30976 65209 31016
rect 64823 30953 64889 30976
rect 64975 30953 65057 30976
rect 65143 30953 65209 30976
rect 64823 30934 65209 30953
rect 79943 31039 80329 31058
rect 79943 31016 80009 31039
rect 80095 31016 80177 31039
rect 80263 31016 80329 31039
rect 79943 30976 79952 31016
rect 79992 30976 80009 31016
rect 80095 30976 80116 31016
rect 80156 30976 80177 31016
rect 80263 30976 80280 31016
rect 80320 30976 80329 31016
rect 79943 30953 80009 30976
rect 80095 30953 80177 30976
rect 80263 30953 80329 30976
rect 79943 30934 80329 30953
rect 95063 31039 95449 31058
rect 95063 31016 95129 31039
rect 95215 31016 95297 31039
rect 95383 31016 95449 31039
rect 95063 30976 95072 31016
rect 95112 30976 95129 31016
rect 95215 30976 95236 31016
rect 95276 30976 95297 31016
rect 95383 30976 95400 31016
rect 95440 30976 95449 31016
rect 95063 30953 95129 30976
rect 95215 30953 95297 30976
rect 95383 30953 95449 30976
rect 95063 30934 95449 30953
rect 3103 30283 3489 30302
rect 3103 30260 3169 30283
rect 3255 30260 3337 30283
rect 3423 30260 3489 30283
rect 3103 30220 3112 30260
rect 3152 30220 3169 30260
rect 3255 30220 3276 30260
rect 3316 30220 3337 30260
rect 3423 30220 3440 30260
rect 3480 30220 3489 30260
rect 3103 30197 3169 30220
rect 3255 30197 3337 30220
rect 3423 30197 3489 30220
rect 3103 30178 3489 30197
rect 18223 30283 18609 30302
rect 18223 30260 18289 30283
rect 18375 30260 18457 30283
rect 18543 30260 18609 30283
rect 18223 30220 18232 30260
rect 18272 30220 18289 30260
rect 18375 30220 18396 30260
rect 18436 30220 18457 30260
rect 18543 30220 18560 30260
rect 18600 30220 18609 30260
rect 18223 30197 18289 30220
rect 18375 30197 18457 30220
rect 18543 30197 18609 30220
rect 18223 30178 18609 30197
rect 33343 30283 33729 30302
rect 33343 30260 33409 30283
rect 33495 30260 33577 30283
rect 33663 30260 33729 30283
rect 33343 30220 33352 30260
rect 33392 30220 33409 30260
rect 33495 30220 33516 30260
rect 33556 30220 33577 30260
rect 33663 30220 33680 30260
rect 33720 30220 33729 30260
rect 33343 30197 33409 30220
rect 33495 30197 33577 30220
rect 33663 30197 33729 30220
rect 33343 30178 33729 30197
rect 48463 30283 48849 30302
rect 48463 30260 48529 30283
rect 48615 30260 48697 30283
rect 48783 30260 48849 30283
rect 48463 30220 48472 30260
rect 48512 30220 48529 30260
rect 48615 30220 48636 30260
rect 48676 30220 48697 30260
rect 48783 30220 48800 30260
rect 48840 30220 48849 30260
rect 48463 30197 48529 30220
rect 48615 30197 48697 30220
rect 48783 30197 48849 30220
rect 48463 30178 48849 30197
rect 63583 30283 63969 30302
rect 63583 30260 63649 30283
rect 63735 30260 63817 30283
rect 63903 30260 63969 30283
rect 63583 30220 63592 30260
rect 63632 30220 63649 30260
rect 63735 30220 63756 30260
rect 63796 30220 63817 30260
rect 63903 30220 63920 30260
rect 63960 30220 63969 30260
rect 63583 30197 63649 30220
rect 63735 30197 63817 30220
rect 63903 30197 63969 30220
rect 63583 30178 63969 30197
rect 78703 30283 79089 30302
rect 78703 30260 78769 30283
rect 78855 30260 78937 30283
rect 79023 30260 79089 30283
rect 78703 30220 78712 30260
rect 78752 30220 78769 30260
rect 78855 30220 78876 30260
rect 78916 30220 78937 30260
rect 79023 30220 79040 30260
rect 79080 30220 79089 30260
rect 78703 30197 78769 30220
rect 78855 30197 78937 30220
rect 79023 30197 79089 30220
rect 78703 30178 79089 30197
rect 93823 30283 94209 30302
rect 93823 30260 93889 30283
rect 93975 30260 94057 30283
rect 94143 30260 94209 30283
rect 93823 30220 93832 30260
rect 93872 30220 93889 30260
rect 93975 30220 93996 30260
rect 94036 30220 94057 30260
rect 94143 30220 94160 30260
rect 94200 30220 94209 30260
rect 93823 30197 93889 30220
rect 93975 30197 94057 30220
rect 94143 30197 94209 30220
rect 93823 30178 94209 30197
rect 4343 29527 4729 29546
rect 4343 29504 4409 29527
rect 4495 29504 4577 29527
rect 4663 29504 4729 29527
rect 4343 29464 4352 29504
rect 4392 29464 4409 29504
rect 4495 29464 4516 29504
rect 4556 29464 4577 29504
rect 4663 29464 4680 29504
rect 4720 29464 4729 29504
rect 4343 29441 4409 29464
rect 4495 29441 4577 29464
rect 4663 29441 4729 29464
rect 4343 29422 4729 29441
rect 19463 29527 19849 29546
rect 19463 29504 19529 29527
rect 19615 29504 19697 29527
rect 19783 29504 19849 29527
rect 19463 29464 19472 29504
rect 19512 29464 19529 29504
rect 19615 29464 19636 29504
rect 19676 29464 19697 29504
rect 19783 29464 19800 29504
rect 19840 29464 19849 29504
rect 19463 29441 19529 29464
rect 19615 29441 19697 29464
rect 19783 29441 19849 29464
rect 19463 29422 19849 29441
rect 34583 29527 34969 29546
rect 34583 29504 34649 29527
rect 34735 29504 34817 29527
rect 34903 29504 34969 29527
rect 34583 29464 34592 29504
rect 34632 29464 34649 29504
rect 34735 29464 34756 29504
rect 34796 29464 34817 29504
rect 34903 29464 34920 29504
rect 34960 29464 34969 29504
rect 34583 29441 34649 29464
rect 34735 29441 34817 29464
rect 34903 29441 34969 29464
rect 34583 29422 34969 29441
rect 49703 29527 50089 29546
rect 49703 29504 49769 29527
rect 49855 29504 49937 29527
rect 50023 29504 50089 29527
rect 49703 29464 49712 29504
rect 49752 29464 49769 29504
rect 49855 29464 49876 29504
rect 49916 29464 49937 29504
rect 50023 29464 50040 29504
rect 50080 29464 50089 29504
rect 49703 29441 49769 29464
rect 49855 29441 49937 29464
rect 50023 29441 50089 29464
rect 49703 29422 50089 29441
rect 64823 29527 65209 29546
rect 64823 29504 64889 29527
rect 64975 29504 65057 29527
rect 65143 29504 65209 29527
rect 64823 29464 64832 29504
rect 64872 29464 64889 29504
rect 64975 29464 64996 29504
rect 65036 29464 65057 29504
rect 65143 29464 65160 29504
rect 65200 29464 65209 29504
rect 64823 29441 64889 29464
rect 64975 29441 65057 29464
rect 65143 29441 65209 29464
rect 64823 29422 65209 29441
rect 79943 29527 80329 29546
rect 79943 29504 80009 29527
rect 80095 29504 80177 29527
rect 80263 29504 80329 29527
rect 79943 29464 79952 29504
rect 79992 29464 80009 29504
rect 80095 29464 80116 29504
rect 80156 29464 80177 29504
rect 80263 29464 80280 29504
rect 80320 29464 80329 29504
rect 79943 29441 80009 29464
rect 80095 29441 80177 29464
rect 80263 29441 80329 29464
rect 79943 29422 80329 29441
rect 95063 29527 95449 29546
rect 95063 29504 95129 29527
rect 95215 29504 95297 29527
rect 95383 29504 95449 29527
rect 95063 29464 95072 29504
rect 95112 29464 95129 29504
rect 95215 29464 95236 29504
rect 95276 29464 95297 29504
rect 95383 29464 95400 29504
rect 95440 29464 95449 29504
rect 95063 29441 95129 29464
rect 95215 29441 95297 29464
rect 95383 29441 95449 29464
rect 95063 29422 95449 29441
rect 3103 28771 3489 28790
rect 3103 28748 3169 28771
rect 3255 28748 3337 28771
rect 3423 28748 3489 28771
rect 3103 28708 3112 28748
rect 3152 28708 3169 28748
rect 3255 28708 3276 28748
rect 3316 28708 3337 28748
rect 3423 28708 3440 28748
rect 3480 28708 3489 28748
rect 3103 28685 3169 28708
rect 3255 28685 3337 28708
rect 3423 28685 3489 28708
rect 3103 28666 3489 28685
rect 18223 28771 18609 28790
rect 18223 28748 18289 28771
rect 18375 28748 18457 28771
rect 18543 28748 18609 28771
rect 18223 28708 18232 28748
rect 18272 28708 18289 28748
rect 18375 28708 18396 28748
rect 18436 28708 18457 28748
rect 18543 28708 18560 28748
rect 18600 28708 18609 28748
rect 18223 28685 18289 28708
rect 18375 28685 18457 28708
rect 18543 28685 18609 28708
rect 18223 28666 18609 28685
rect 33343 28771 33729 28790
rect 33343 28748 33409 28771
rect 33495 28748 33577 28771
rect 33663 28748 33729 28771
rect 33343 28708 33352 28748
rect 33392 28708 33409 28748
rect 33495 28708 33516 28748
rect 33556 28708 33577 28748
rect 33663 28708 33680 28748
rect 33720 28708 33729 28748
rect 33343 28685 33409 28708
rect 33495 28685 33577 28708
rect 33663 28685 33729 28708
rect 33343 28666 33729 28685
rect 48463 28771 48849 28790
rect 48463 28748 48529 28771
rect 48615 28748 48697 28771
rect 48783 28748 48849 28771
rect 48463 28708 48472 28748
rect 48512 28708 48529 28748
rect 48615 28708 48636 28748
rect 48676 28708 48697 28748
rect 48783 28708 48800 28748
rect 48840 28708 48849 28748
rect 48463 28685 48529 28708
rect 48615 28685 48697 28708
rect 48783 28685 48849 28708
rect 48463 28666 48849 28685
rect 63583 28771 63969 28790
rect 63583 28748 63649 28771
rect 63735 28748 63817 28771
rect 63903 28748 63969 28771
rect 63583 28708 63592 28748
rect 63632 28708 63649 28748
rect 63735 28708 63756 28748
rect 63796 28708 63817 28748
rect 63903 28708 63920 28748
rect 63960 28708 63969 28748
rect 63583 28685 63649 28708
rect 63735 28685 63817 28708
rect 63903 28685 63969 28708
rect 63583 28666 63969 28685
rect 78703 28771 79089 28790
rect 78703 28748 78769 28771
rect 78855 28748 78937 28771
rect 79023 28748 79089 28771
rect 78703 28708 78712 28748
rect 78752 28708 78769 28748
rect 78855 28708 78876 28748
rect 78916 28708 78937 28748
rect 79023 28708 79040 28748
rect 79080 28708 79089 28748
rect 78703 28685 78769 28708
rect 78855 28685 78937 28708
rect 79023 28685 79089 28708
rect 78703 28666 79089 28685
rect 93823 28771 94209 28790
rect 93823 28748 93889 28771
rect 93975 28748 94057 28771
rect 94143 28748 94209 28771
rect 93823 28708 93832 28748
rect 93872 28708 93889 28748
rect 93975 28708 93996 28748
rect 94036 28708 94057 28748
rect 94143 28708 94160 28748
rect 94200 28708 94209 28748
rect 93823 28685 93889 28708
rect 93975 28685 94057 28708
rect 94143 28685 94209 28708
rect 93823 28666 94209 28685
rect 4343 28015 4729 28034
rect 4343 27992 4409 28015
rect 4495 27992 4577 28015
rect 4663 27992 4729 28015
rect 4343 27952 4352 27992
rect 4392 27952 4409 27992
rect 4495 27952 4516 27992
rect 4556 27952 4577 27992
rect 4663 27952 4680 27992
rect 4720 27952 4729 27992
rect 4343 27929 4409 27952
rect 4495 27929 4577 27952
rect 4663 27929 4729 27952
rect 4343 27910 4729 27929
rect 19463 28015 19849 28034
rect 19463 27992 19529 28015
rect 19615 27992 19697 28015
rect 19783 27992 19849 28015
rect 19463 27952 19472 27992
rect 19512 27952 19529 27992
rect 19615 27952 19636 27992
rect 19676 27952 19697 27992
rect 19783 27952 19800 27992
rect 19840 27952 19849 27992
rect 19463 27929 19529 27952
rect 19615 27929 19697 27952
rect 19783 27929 19849 27952
rect 19463 27910 19849 27929
rect 34583 28015 34969 28034
rect 34583 27992 34649 28015
rect 34735 27992 34817 28015
rect 34903 27992 34969 28015
rect 34583 27952 34592 27992
rect 34632 27952 34649 27992
rect 34735 27952 34756 27992
rect 34796 27952 34817 27992
rect 34903 27952 34920 27992
rect 34960 27952 34969 27992
rect 34583 27929 34649 27952
rect 34735 27929 34817 27952
rect 34903 27929 34969 27952
rect 34583 27910 34969 27929
rect 49703 28015 50089 28034
rect 49703 27992 49769 28015
rect 49855 27992 49937 28015
rect 50023 27992 50089 28015
rect 49703 27952 49712 27992
rect 49752 27952 49769 27992
rect 49855 27952 49876 27992
rect 49916 27952 49937 27992
rect 50023 27952 50040 27992
rect 50080 27952 50089 27992
rect 49703 27929 49769 27952
rect 49855 27929 49937 27952
rect 50023 27929 50089 27952
rect 49703 27910 50089 27929
rect 64823 28015 65209 28034
rect 64823 27992 64889 28015
rect 64975 27992 65057 28015
rect 65143 27992 65209 28015
rect 64823 27952 64832 27992
rect 64872 27952 64889 27992
rect 64975 27952 64996 27992
rect 65036 27952 65057 27992
rect 65143 27952 65160 27992
rect 65200 27952 65209 27992
rect 64823 27929 64889 27952
rect 64975 27929 65057 27952
rect 65143 27929 65209 27952
rect 64823 27910 65209 27929
rect 79943 28015 80329 28034
rect 79943 27992 80009 28015
rect 80095 27992 80177 28015
rect 80263 27992 80329 28015
rect 79943 27952 79952 27992
rect 79992 27952 80009 27992
rect 80095 27952 80116 27992
rect 80156 27952 80177 27992
rect 80263 27952 80280 27992
rect 80320 27952 80329 27992
rect 79943 27929 80009 27952
rect 80095 27929 80177 27952
rect 80263 27929 80329 27952
rect 79943 27910 80329 27929
rect 95063 28015 95449 28034
rect 95063 27992 95129 28015
rect 95215 27992 95297 28015
rect 95383 27992 95449 28015
rect 95063 27952 95072 27992
rect 95112 27952 95129 27992
rect 95215 27952 95236 27992
rect 95276 27952 95297 27992
rect 95383 27952 95400 27992
rect 95440 27952 95449 27992
rect 95063 27929 95129 27952
rect 95215 27929 95297 27952
rect 95383 27929 95449 27952
rect 95063 27910 95449 27929
rect 3103 27259 3489 27278
rect 3103 27236 3169 27259
rect 3255 27236 3337 27259
rect 3423 27236 3489 27259
rect 3103 27196 3112 27236
rect 3152 27196 3169 27236
rect 3255 27196 3276 27236
rect 3316 27196 3337 27236
rect 3423 27196 3440 27236
rect 3480 27196 3489 27236
rect 3103 27173 3169 27196
rect 3255 27173 3337 27196
rect 3423 27173 3489 27196
rect 3103 27154 3489 27173
rect 18223 27259 18609 27278
rect 18223 27236 18289 27259
rect 18375 27236 18457 27259
rect 18543 27236 18609 27259
rect 18223 27196 18232 27236
rect 18272 27196 18289 27236
rect 18375 27196 18396 27236
rect 18436 27196 18457 27236
rect 18543 27196 18560 27236
rect 18600 27196 18609 27236
rect 18223 27173 18289 27196
rect 18375 27173 18457 27196
rect 18543 27173 18609 27196
rect 18223 27154 18609 27173
rect 33343 27259 33729 27278
rect 33343 27236 33409 27259
rect 33495 27236 33577 27259
rect 33663 27236 33729 27259
rect 33343 27196 33352 27236
rect 33392 27196 33409 27236
rect 33495 27196 33516 27236
rect 33556 27196 33577 27236
rect 33663 27196 33680 27236
rect 33720 27196 33729 27236
rect 33343 27173 33409 27196
rect 33495 27173 33577 27196
rect 33663 27173 33729 27196
rect 33343 27154 33729 27173
rect 48463 27259 48849 27278
rect 48463 27236 48529 27259
rect 48615 27236 48697 27259
rect 48783 27236 48849 27259
rect 48463 27196 48472 27236
rect 48512 27196 48529 27236
rect 48615 27196 48636 27236
rect 48676 27196 48697 27236
rect 48783 27196 48800 27236
rect 48840 27196 48849 27236
rect 48463 27173 48529 27196
rect 48615 27173 48697 27196
rect 48783 27173 48849 27196
rect 48463 27154 48849 27173
rect 63583 27259 63969 27278
rect 63583 27236 63649 27259
rect 63735 27236 63817 27259
rect 63903 27236 63969 27259
rect 63583 27196 63592 27236
rect 63632 27196 63649 27236
rect 63735 27196 63756 27236
rect 63796 27196 63817 27236
rect 63903 27196 63920 27236
rect 63960 27196 63969 27236
rect 63583 27173 63649 27196
rect 63735 27173 63817 27196
rect 63903 27173 63969 27196
rect 63583 27154 63969 27173
rect 78703 27259 79089 27278
rect 78703 27236 78769 27259
rect 78855 27236 78937 27259
rect 79023 27236 79089 27259
rect 78703 27196 78712 27236
rect 78752 27196 78769 27236
rect 78855 27196 78876 27236
rect 78916 27196 78937 27236
rect 79023 27196 79040 27236
rect 79080 27196 79089 27236
rect 78703 27173 78769 27196
rect 78855 27173 78937 27196
rect 79023 27173 79089 27196
rect 78703 27154 79089 27173
rect 93823 27259 94209 27278
rect 93823 27236 93889 27259
rect 93975 27236 94057 27259
rect 94143 27236 94209 27259
rect 93823 27196 93832 27236
rect 93872 27196 93889 27236
rect 93975 27196 93996 27236
rect 94036 27196 94057 27236
rect 94143 27196 94160 27236
rect 94200 27196 94209 27236
rect 93823 27173 93889 27196
rect 93975 27173 94057 27196
rect 94143 27173 94209 27196
rect 93823 27154 94209 27173
rect 4343 26503 4729 26522
rect 4343 26480 4409 26503
rect 4495 26480 4577 26503
rect 4663 26480 4729 26503
rect 4343 26440 4352 26480
rect 4392 26440 4409 26480
rect 4495 26440 4516 26480
rect 4556 26440 4577 26480
rect 4663 26440 4680 26480
rect 4720 26440 4729 26480
rect 4343 26417 4409 26440
rect 4495 26417 4577 26440
rect 4663 26417 4729 26440
rect 4343 26398 4729 26417
rect 19463 26503 19849 26522
rect 19463 26480 19529 26503
rect 19615 26480 19697 26503
rect 19783 26480 19849 26503
rect 19463 26440 19472 26480
rect 19512 26440 19529 26480
rect 19615 26440 19636 26480
rect 19676 26440 19697 26480
rect 19783 26440 19800 26480
rect 19840 26440 19849 26480
rect 19463 26417 19529 26440
rect 19615 26417 19697 26440
rect 19783 26417 19849 26440
rect 19463 26398 19849 26417
rect 34583 26503 34969 26522
rect 34583 26480 34649 26503
rect 34735 26480 34817 26503
rect 34903 26480 34969 26503
rect 34583 26440 34592 26480
rect 34632 26440 34649 26480
rect 34735 26440 34756 26480
rect 34796 26440 34817 26480
rect 34903 26440 34920 26480
rect 34960 26440 34969 26480
rect 34583 26417 34649 26440
rect 34735 26417 34817 26440
rect 34903 26417 34969 26440
rect 34583 26398 34969 26417
rect 49703 26503 50089 26522
rect 49703 26480 49769 26503
rect 49855 26480 49937 26503
rect 50023 26480 50089 26503
rect 49703 26440 49712 26480
rect 49752 26440 49769 26480
rect 49855 26440 49876 26480
rect 49916 26440 49937 26480
rect 50023 26440 50040 26480
rect 50080 26440 50089 26480
rect 49703 26417 49769 26440
rect 49855 26417 49937 26440
rect 50023 26417 50089 26440
rect 49703 26398 50089 26417
rect 64823 26503 65209 26522
rect 64823 26480 64889 26503
rect 64975 26480 65057 26503
rect 65143 26480 65209 26503
rect 64823 26440 64832 26480
rect 64872 26440 64889 26480
rect 64975 26440 64996 26480
rect 65036 26440 65057 26480
rect 65143 26440 65160 26480
rect 65200 26440 65209 26480
rect 64823 26417 64889 26440
rect 64975 26417 65057 26440
rect 65143 26417 65209 26440
rect 64823 26398 65209 26417
rect 79943 26503 80329 26522
rect 79943 26480 80009 26503
rect 80095 26480 80177 26503
rect 80263 26480 80329 26503
rect 79943 26440 79952 26480
rect 79992 26440 80009 26480
rect 80095 26440 80116 26480
rect 80156 26440 80177 26480
rect 80263 26440 80280 26480
rect 80320 26440 80329 26480
rect 79943 26417 80009 26440
rect 80095 26417 80177 26440
rect 80263 26417 80329 26440
rect 79943 26398 80329 26417
rect 95063 26503 95449 26522
rect 95063 26480 95129 26503
rect 95215 26480 95297 26503
rect 95383 26480 95449 26503
rect 95063 26440 95072 26480
rect 95112 26440 95129 26480
rect 95215 26440 95236 26480
rect 95276 26440 95297 26480
rect 95383 26440 95400 26480
rect 95440 26440 95449 26480
rect 95063 26417 95129 26440
rect 95215 26417 95297 26440
rect 95383 26417 95449 26440
rect 95063 26398 95449 26417
rect 3103 25747 3489 25766
rect 3103 25724 3169 25747
rect 3255 25724 3337 25747
rect 3423 25724 3489 25747
rect 3103 25684 3112 25724
rect 3152 25684 3169 25724
rect 3255 25684 3276 25724
rect 3316 25684 3337 25724
rect 3423 25684 3440 25724
rect 3480 25684 3489 25724
rect 3103 25661 3169 25684
rect 3255 25661 3337 25684
rect 3423 25661 3489 25684
rect 3103 25642 3489 25661
rect 18223 25747 18609 25766
rect 18223 25724 18289 25747
rect 18375 25724 18457 25747
rect 18543 25724 18609 25747
rect 18223 25684 18232 25724
rect 18272 25684 18289 25724
rect 18375 25684 18396 25724
rect 18436 25684 18457 25724
rect 18543 25684 18560 25724
rect 18600 25684 18609 25724
rect 18223 25661 18289 25684
rect 18375 25661 18457 25684
rect 18543 25661 18609 25684
rect 18223 25642 18609 25661
rect 33343 25747 33729 25766
rect 33343 25724 33409 25747
rect 33495 25724 33577 25747
rect 33663 25724 33729 25747
rect 33343 25684 33352 25724
rect 33392 25684 33409 25724
rect 33495 25684 33516 25724
rect 33556 25684 33577 25724
rect 33663 25684 33680 25724
rect 33720 25684 33729 25724
rect 33343 25661 33409 25684
rect 33495 25661 33577 25684
rect 33663 25661 33729 25684
rect 33343 25642 33729 25661
rect 48463 25747 48849 25766
rect 48463 25724 48529 25747
rect 48615 25724 48697 25747
rect 48783 25724 48849 25747
rect 48463 25684 48472 25724
rect 48512 25684 48529 25724
rect 48615 25684 48636 25724
rect 48676 25684 48697 25724
rect 48783 25684 48800 25724
rect 48840 25684 48849 25724
rect 48463 25661 48529 25684
rect 48615 25661 48697 25684
rect 48783 25661 48849 25684
rect 48463 25642 48849 25661
rect 63583 25747 63969 25766
rect 63583 25724 63649 25747
rect 63735 25724 63817 25747
rect 63903 25724 63969 25747
rect 63583 25684 63592 25724
rect 63632 25684 63649 25724
rect 63735 25684 63756 25724
rect 63796 25684 63817 25724
rect 63903 25684 63920 25724
rect 63960 25684 63969 25724
rect 63583 25661 63649 25684
rect 63735 25661 63817 25684
rect 63903 25661 63969 25684
rect 63583 25642 63969 25661
rect 78703 25747 79089 25766
rect 78703 25724 78769 25747
rect 78855 25724 78937 25747
rect 79023 25724 79089 25747
rect 78703 25684 78712 25724
rect 78752 25684 78769 25724
rect 78855 25684 78876 25724
rect 78916 25684 78937 25724
rect 79023 25684 79040 25724
rect 79080 25684 79089 25724
rect 78703 25661 78769 25684
rect 78855 25661 78937 25684
rect 79023 25661 79089 25684
rect 78703 25642 79089 25661
rect 93823 25747 94209 25766
rect 93823 25724 93889 25747
rect 93975 25724 94057 25747
rect 94143 25724 94209 25747
rect 93823 25684 93832 25724
rect 93872 25684 93889 25724
rect 93975 25684 93996 25724
rect 94036 25684 94057 25724
rect 94143 25684 94160 25724
rect 94200 25684 94209 25724
rect 93823 25661 93889 25684
rect 93975 25661 94057 25684
rect 94143 25661 94209 25684
rect 93823 25642 94209 25661
rect 4343 24991 4729 25010
rect 4343 24968 4409 24991
rect 4495 24968 4577 24991
rect 4663 24968 4729 24991
rect 4343 24928 4352 24968
rect 4392 24928 4409 24968
rect 4495 24928 4516 24968
rect 4556 24928 4577 24968
rect 4663 24928 4680 24968
rect 4720 24928 4729 24968
rect 4343 24905 4409 24928
rect 4495 24905 4577 24928
rect 4663 24905 4729 24928
rect 4343 24886 4729 24905
rect 19463 24991 19849 25010
rect 19463 24968 19529 24991
rect 19615 24968 19697 24991
rect 19783 24968 19849 24991
rect 19463 24928 19472 24968
rect 19512 24928 19529 24968
rect 19615 24928 19636 24968
rect 19676 24928 19697 24968
rect 19783 24928 19800 24968
rect 19840 24928 19849 24968
rect 19463 24905 19529 24928
rect 19615 24905 19697 24928
rect 19783 24905 19849 24928
rect 19463 24886 19849 24905
rect 34583 24991 34969 25010
rect 34583 24968 34649 24991
rect 34735 24968 34817 24991
rect 34903 24968 34969 24991
rect 34583 24928 34592 24968
rect 34632 24928 34649 24968
rect 34735 24928 34756 24968
rect 34796 24928 34817 24968
rect 34903 24928 34920 24968
rect 34960 24928 34969 24968
rect 34583 24905 34649 24928
rect 34735 24905 34817 24928
rect 34903 24905 34969 24928
rect 34583 24886 34969 24905
rect 49703 24991 50089 25010
rect 49703 24968 49769 24991
rect 49855 24968 49937 24991
rect 50023 24968 50089 24991
rect 49703 24928 49712 24968
rect 49752 24928 49769 24968
rect 49855 24928 49876 24968
rect 49916 24928 49937 24968
rect 50023 24928 50040 24968
rect 50080 24928 50089 24968
rect 49703 24905 49769 24928
rect 49855 24905 49937 24928
rect 50023 24905 50089 24928
rect 49703 24886 50089 24905
rect 64823 24991 65209 25010
rect 64823 24968 64889 24991
rect 64975 24968 65057 24991
rect 65143 24968 65209 24991
rect 64823 24928 64832 24968
rect 64872 24928 64889 24968
rect 64975 24928 64996 24968
rect 65036 24928 65057 24968
rect 65143 24928 65160 24968
rect 65200 24928 65209 24968
rect 64823 24905 64889 24928
rect 64975 24905 65057 24928
rect 65143 24905 65209 24928
rect 64823 24886 65209 24905
rect 79943 24991 80329 25010
rect 79943 24968 80009 24991
rect 80095 24968 80177 24991
rect 80263 24968 80329 24991
rect 79943 24928 79952 24968
rect 79992 24928 80009 24968
rect 80095 24928 80116 24968
rect 80156 24928 80177 24968
rect 80263 24928 80280 24968
rect 80320 24928 80329 24968
rect 79943 24905 80009 24928
rect 80095 24905 80177 24928
rect 80263 24905 80329 24928
rect 79943 24886 80329 24905
rect 95063 24991 95449 25010
rect 95063 24968 95129 24991
rect 95215 24968 95297 24991
rect 95383 24968 95449 24991
rect 95063 24928 95072 24968
rect 95112 24928 95129 24968
rect 95215 24928 95236 24968
rect 95276 24928 95297 24968
rect 95383 24928 95400 24968
rect 95440 24928 95449 24968
rect 95063 24905 95129 24928
rect 95215 24905 95297 24928
rect 95383 24905 95449 24928
rect 95063 24886 95449 24905
rect 3103 24235 3489 24254
rect 3103 24212 3169 24235
rect 3255 24212 3337 24235
rect 3423 24212 3489 24235
rect 3103 24172 3112 24212
rect 3152 24172 3169 24212
rect 3255 24172 3276 24212
rect 3316 24172 3337 24212
rect 3423 24172 3440 24212
rect 3480 24172 3489 24212
rect 3103 24149 3169 24172
rect 3255 24149 3337 24172
rect 3423 24149 3489 24172
rect 3103 24130 3489 24149
rect 18223 24235 18609 24254
rect 18223 24212 18289 24235
rect 18375 24212 18457 24235
rect 18543 24212 18609 24235
rect 18223 24172 18232 24212
rect 18272 24172 18289 24212
rect 18375 24172 18396 24212
rect 18436 24172 18457 24212
rect 18543 24172 18560 24212
rect 18600 24172 18609 24212
rect 18223 24149 18289 24172
rect 18375 24149 18457 24172
rect 18543 24149 18609 24172
rect 18223 24130 18609 24149
rect 33343 24235 33729 24254
rect 33343 24212 33409 24235
rect 33495 24212 33577 24235
rect 33663 24212 33729 24235
rect 33343 24172 33352 24212
rect 33392 24172 33409 24212
rect 33495 24172 33516 24212
rect 33556 24172 33577 24212
rect 33663 24172 33680 24212
rect 33720 24172 33729 24212
rect 33343 24149 33409 24172
rect 33495 24149 33577 24172
rect 33663 24149 33729 24172
rect 33343 24130 33729 24149
rect 48463 24235 48849 24254
rect 48463 24212 48529 24235
rect 48615 24212 48697 24235
rect 48783 24212 48849 24235
rect 48463 24172 48472 24212
rect 48512 24172 48529 24212
rect 48615 24172 48636 24212
rect 48676 24172 48697 24212
rect 48783 24172 48800 24212
rect 48840 24172 48849 24212
rect 48463 24149 48529 24172
rect 48615 24149 48697 24172
rect 48783 24149 48849 24172
rect 48463 24130 48849 24149
rect 63583 24235 63969 24254
rect 63583 24212 63649 24235
rect 63735 24212 63817 24235
rect 63903 24212 63969 24235
rect 63583 24172 63592 24212
rect 63632 24172 63649 24212
rect 63735 24172 63756 24212
rect 63796 24172 63817 24212
rect 63903 24172 63920 24212
rect 63960 24172 63969 24212
rect 63583 24149 63649 24172
rect 63735 24149 63817 24172
rect 63903 24149 63969 24172
rect 63583 24130 63969 24149
rect 78703 24235 79089 24254
rect 78703 24212 78769 24235
rect 78855 24212 78937 24235
rect 79023 24212 79089 24235
rect 78703 24172 78712 24212
rect 78752 24172 78769 24212
rect 78855 24172 78876 24212
rect 78916 24172 78937 24212
rect 79023 24172 79040 24212
rect 79080 24172 79089 24212
rect 78703 24149 78769 24172
rect 78855 24149 78937 24172
rect 79023 24149 79089 24172
rect 78703 24130 79089 24149
rect 93823 24235 94209 24254
rect 93823 24212 93889 24235
rect 93975 24212 94057 24235
rect 94143 24212 94209 24235
rect 93823 24172 93832 24212
rect 93872 24172 93889 24212
rect 93975 24172 93996 24212
rect 94036 24172 94057 24212
rect 94143 24172 94160 24212
rect 94200 24172 94209 24212
rect 93823 24149 93889 24172
rect 93975 24149 94057 24172
rect 94143 24149 94209 24172
rect 93823 24130 94209 24149
rect 4343 23479 4729 23498
rect 4343 23456 4409 23479
rect 4495 23456 4577 23479
rect 4663 23456 4729 23479
rect 4343 23416 4352 23456
rect 4392 23416 4409 23456
rect 4495 23416 4516 23456
rect 4556 23416 4577 23456
rect 4663 23416 4680 23456
rect 4720 23416 4729 23456
rect 4343 23393 4409 23416
rect 4495 23393 4577 23416
rect 4663 23393 4729 23416
rect 4343 23374 4729 23393
rect 19463 23479 19849 23498
rect 19463 23456 19529 23479
rect 19615 23456 19697 23479
rect 19783 23456 19849 23479
rect 19463 23416 19472 23456
rect 19512 23416 19529 23456
rect 19615 23416 19636 23456
rect 19676 23416 19697 23456
rect 19783 23416 19800 23456
rect 19840 23416 19849 23456
rect 19463 23393 19529 23416
rect 19615 23393 19697 23416
rect 19783 23393 19849 23416
rect 19463 23374 19849 23393
rect 34583 23479 34969 23498
rect 34583 23456 34649 23479
rect 34735 23456 34817 23479
rect 34903 23456 34969 23479
rect 34583 23416 34592 23456
rect 34632 23416 34649 23456
rect 34735 23416 34756 23456
rect 34796 23416 34817 23456
rect 34903 23416 34920 23456
rect 34960 23416 34969 23456
rect 34583 23393 34649 23416
rect 34735 23393 34817 23416
rect 34903 23393 34969 23416
rect 34583 23374 34969 23393
rect 49703 23479 50089 23498
rect 49703 23456 49769 23479
rect 49855 23456 49937 23479
rect 50023 23456 50089 23479
rect 49703 23416 49712 23456
rect 49752 23416 49769 23456
rect 49855 23416 49876 23456
rect 49916 23416 49937 23456
rect 50023 23416 50040 23456
rect 50080 23416 50089 23456
rect 49703 23393 49769 23416
rect 49855 23393 49937 23416
rect 50023 23393 50089 23416
rect 49703 23374 50089 23393
rect 64823 23479 65209 23498
rect 64823 23456 64889 23479
rect 64975 23456 65057 23479
rect 65143 23456 65209 23479
rect 64823 23416 64832 23456
rect 64872 23416 64889 23456
rect 64975 23416 64996 23456
rect 65036 23416 65057 23456
rect 65143 23416 65160 23456
rect 65200 23416 65209 23456
rect 64823 23393 64889 23416
rect 64975 23393 65057 23416
rect 65143 23393 65209 23416
rect 64823 23374 65209 23393
rect 79943 23479 80329 23498
rect 79943 23456 80009 23479
rect 80095 23456 80177 23479
rect 80263 23456 80329 23479
rect 79943 23416 79952 23456
rect 79992 23416 80009 23456
rect 80095 23416 80116 23456
rect 80156 23416 80177 23456
rect 80263 23416 80280 23456
rect 80320 23416 80329 23456
rect 79943 23393 80009 23416
rect 80095 23393 80177 23416
rect 80263 23393 80329 23416
rect 79943 23374 80329 23393
rect 95063 23479 95449 23498
rect 95063 23456 95129 23479
rect 95215 23456 95297 23479
rect 95383 23456 95449 23479
rect 95063 23416 95072 23456
rect 95112 23416 95129 23456
rect 95215 23416 95236 23456
rect 95276 23416 95297 23456
rect 95383 23416 95400 23456
rect 95440 23416 95449 23456
rect 95063 23393 95129 23416
rect 95215 23393 95297 23416
rect 95383 23393 95449 23416
rect 95063 23374 95449 23393
rect 3103 22723 3489 22742
rect 3103 22700 3169 22723
rect 3255 22700 3337 22723
rect 3423 22700 3489 22723
rect 3103 22660 3112 22700
rect 3152 22660 3169 22700
rect 3255 22660 3276 22700
rect 3316 22660 3337 22700
rect 3423 22660 3440 22700
rect 3480 22660 3489 22700
rect 3103 22637 3169 22660
rect 3255 22637 3337 22660
rect 3423 22637 3489 22660
rect 3103 22618 3489 22637
rect 18223 22723 18609 22742
rect 18223 22700 18289 22723
rect 18375 22700 18457 22723
rect 18543 22700 18609 22723
rect 18223 22660 18232 22700
rect 18272 22660 18289 22700
rect 18375 22660 18396 22700
rect 18436 22660 18457 22700
rect 18543 22660 18560 22700
rect 18600 22660 18609 22700
rect 18223 22637 18289 22660
rect 18375 22637 18457 22660
rect 18543 22637 18609 22660
rect 18223 22618 18609 22637
rect 33343 22723 33729 22742
rect 33343 22700 33409 22723
rect 33495 22700 33577 22723
rect 33663 22700 33729 22723
rect 33343 22660 33352 22700
rect 33392 22660 33409 22700
rect 33495 22660 33516 22700
rect 33556 22660 33577 22700
rect 33663 22660 33680 22700
rect 33720 22660 33729 22700
rect 33343 22637 33409 22660
rect 33495 22637 33577 22660
rect 33663 22637 33729 22660
rect 33343 22618 33729 22637
rect 48463 22723 48849 22742
rect 48463 22700 48529 22723
rect 48615 22700 48697 22723
rect 48783 22700 48849 22723
rect 48463 22660 48472 22700
rect 48512 22660 48529 22700
rect 48615 22660 48636 22700
rect 48676 22660 48697 22700
rect 48783 22660 48800 22700
rect 48840 22660 48849 22700
rect 48463 22637 48529 22660
rect 48615 22637 48697 22660
rect 48783 22637 48849 22660
rect 48463 22618 48849 22637
rect 63583 22723 63969 22742
rect 63583 22700 63649 22723
rect 63735 22700 63817 22723
rect 63903 22700 63969 22723
rect 63583 22660 63592 22700
rect 63632 22660 63649 22700
rect 63735 22660 63756 22700
rect 63796 22660 63817 22700
rect 63903 22660 63920 22700
rect 63960 22660 63969 22700
rect 63583 22637 63649 22660
rect 63735 22637 63817 22660
rect 63903 22637 63969 22660
rect 63583 22618 63969 22637
rect 78703 22723 79089 22742
rect 78703 22700 78769 22723
rect 78855 22700 78937 22723
rect 79023 22700 79089 22723
rect 78703 22660 78712 22700
rect 78752 22660 78769 22700
rect 78855 22660 78876 22700
rect 78916 22660 78937 22700
rect 79023 22660 79040 22700
rect 79080 22660 79089 22700
rect 78703 22637 78769 22660
rect 78855 22637 78937 22660
rect 79023 22637 79089 22660
rect 78703 22618 79089 22637
rect 93823 22723 94209 22742
rect 93823 22700 93889 22723
rect 93975 22700 94057 22723
rect 94143 22700 94209 22723
rect 93823 22660 93832 22700
rect 93872 22660 93889 22700
rect 93975 22660 93996 22700
rect 94036 22660 94057 22700
rect 94143 22660 94160 22700
rect 94200 22660 94209 22700
rect 93823 22637 93889 22660
rect 93975 22637 94057 22660
rect 94143 22637 94209 22660
rect 93823 22618 94209 22637
rect 4343 21967 4729 21986
rect 4343 21944 4409 21967
rect 4495 21944 4577 21967
rect 4663 21944 4729 21967
rect 4343 21904 4352 21944
rect 4392 21904 4409 21944
rect 4495 21904 4516 21944
rect 4556 21904 4577 21944
rect 4663 21904 4680 21944
rect 4720 21904 4729 21944
rect 4343 21881 4409 21904
rect 4495 21881 4577 21904
rect 4663 21881 4729 21904
rect 4343 21862 4729 21881
rect 19463 21967 19849 21986
rect 19463 21944 19529 21967
rect 19615 21944 19697 21967
rect 19783 21944 19849 21967
rect 19463 21904 19472 21944
rect 19512 21904 19529 21944
rect 19615 21904 19636 21944
rect 19676 21904 19697 21944
rect 19783 21904 19800 21944
rect 19840 21904 19849 21944
rect 19463 21881 19529 21904
rect 19615 21881 19697 21904
rect 19783 21881 19849 21904
rect 19463 21862 19849 21881
rect 34583 21967 34969 21986
rect 34583 21944 34649 21967
rect 34735 21944 34817 21967
rect 34903 21944 34969 21967
rect 34583 21904 34592 21944
rect 34632 21904 34649 21944
rect 34735 21904 34756 21944
rect 34796 21904 34817 21944
rect 34903 21904 34920 21944
rect 34960 21904 34969 21944
rect 34583 21881 34649 21904
rect 34735 21881 34817 21904
rect 34903 21881 34969 21904
rect 34583 21862 34969 21881
rect 49703 21967 50089 21986
rect 49703 21944 49769 21967
rect 49855 21944 49937 21967
rect 50023 21944 50089 21967
rect 49703 21904 49712 21944
rect 49752 21904 49769 21944
rect 49855 21904 49876 21944
rect 49916 21904 49937 21944
rect 50023 21904 50040 21944
rect 50080 21904 50089 21944
rect 49703 21881 49769 21904
rect 49855 21881 49937 21904
rect 50023 21881 50089 21904
rect 49703 21862 50089 21881
rect 64823 21967 65209 21986
rect 64823 21944 64889 21967
rect 64975 21944 65057 21967
rect 65143 21944 65209 21967
rect 64823 21904 64832 21944
rect 64872 21904 64889 21944
rect 64975 21904 64996 21944
rect 65036 21904 65057 21944
rect 65143 21904 65160 21944
rect 65200 21904 65209 21944
rect 64823 21881 64889 21904
rect 64975 21881 65057 21904
rect 65143 21881 65209 21904
rect 64823 21862 65209 21881
rect 79943 21967 80329 21986
rect 79943 21944 80009 21967
rect 80095 21944 80177 21967
rect 80263 21944 80329 21967
rect 79943 21904 79952 21944
rect 79992 21904 80009 21944
rect 80095 21904 80116 21944
rect 80156 21904 80177 21944
rect 80263 21904 80280 21944
rect 80320 21904 80329 21944
rect 79943 21881 80009 21904
rect 80095 21881 80177 21904
rect 80263 21881 80329 21904
rect 79943 21862 80329 21881
rect 95063 21967 95449 21986
rect 95063 21944 95129 21967
rect 95215 21944 95297 21967
rect 95383 21944 95449 21967
rect 95063 21904 95072 21944
rect 95112 21904 95129 21944
rect 95215 21904 95236 21944
rect 95276 21904 95297 21944
rect 95383 21904 95400 21944
rect 95440 21904 95449 21944
rect 95063 21881 95129 21904
rect 95215 21881 95297 21904
rect 95383 21881 95449 21904
rect 95063 21862 95449 21881
rect 3103 21211 3489 21230
rect 3103 21188 3169 21211
rect 3255 21188 3337 21211
rect 3423 21188 3489 21211
rect 3103 21148 3112 21188
rect 3152 21148 3169 21188
rect 3255 21148 3276 21188
rect 3316 21148 3337 21188
rect 3423 21148 3440 21188
rect 3480 21148 3489 21188
rect 3103 21125 3169 21148
rect 3255 21125 3337 21148
rect 3423 21125 3489 21148
rect 3103 21106 3489 21125
rect 18223 21211 18609 21230
rect 18223 21188 18289 21211
rect 18375 21188 18457 21211
rect 18543 21188 18609 21211
rect 18223 21148 18232 21188
rect 18272 21148 18289 21188
rect 18375 21148 18396 21188
rect 18436 21148 18457 21188
rect 18543 21148 18560 21188
rect 18600 21148 18609 21188
rect 18223 21125 18289 21148
rect 18375 21125 18457 21148
rect 18543 21125 18609 21148
rect 18223 21106 18609 21125
rect 33343 21211 33729 21230
rect 33343 21188 33409 21211
rect 33495 21188 33577 21211
rect 33663 21188 33729 21211
rect 33343 21148 33352 21188
rect 33392 21148 33409 21188
rect 33495 21148 33516 21188
rect 33556 21148 33577 21188
rect 33663 21148 33680 21188
rect 33720 21148 33729 21188
rect 33343 21125 33409 21148
rect 33495 21125 33577 21148
rect 33663 21125 33729 21148
rect 33343 21106 33729 21125
rect 48463 21211 48849 21230
rect 48463 21188 48529 21211
rect 48615 21188 48697 21211
rect 48783 21188 48849 21211
rect 48463 21148 48472 21188
rect 48512 21148 48529 21188
rect 48615 21148 48636 21188
rect 48676 21148 48697 21188
rect 48783 21148 48800 21188
rect 48840 21148 48849 21188
rect 48463 21125 48529 21148
rect 48615 21125 48697 21148
rect 48783 21125 48849 21148
rect 48463 21106 48849 21125
rect 63583 21211 63969 21230
rect 63583 21188 63649 21211
rect 63735 21188 63817 21211
rect 63903 21188 63969 21211
rect 63583 21148 63592 21188
rect 63632 21148 63649 21188
rect 63735 21148 63756 21188
rect 63796 21148 63817 21188
rect 63903 21148 63920 21188
rect 63960 21148 63969 21188
rect 63583 21125 63649 21148
rect 63735 21125 63817 21148
rect 63903 21125 63969 21148
rect 63583 21106 63969 21125
rect 78703 21211 79089 21230
rect 78703 21188 78769 21211
rect 78855 21188 78937 21211
rect 79023 21188 79089 21211
rect 78703 21148 78712 21188
rect 78752 21148 78769 21188
rect 78855 21148 78876 21188
rect 78916 21148 78937 21188
rect 79023 21148 79040 21188
rect 79080 21148 79089 21188
rect 78703 21125 78769 21148
rect 78855 21125 78937 21148
rect 79023 21125 79089 21148
rect 78703 21106 79089 21125
rect 93823 21211 94209 21230
rect 93823 21188 93889 21211
rect 93975 21188 94057 21211
rect 94143 21188 94209 21211
rect 93823 21148 93832 21188
rect 93872 21148 93889 21188
rect 93975 21148 93996 21188
rect 94036 21148 94057 21188
rect 94143 21148 94160 21188
rect 94200 21148 94209 21188
rect 93823 21125 93889 21148
rect 93975 21125 94057 21148
rect 94143 21125 94209 21148
rect 93823 21106 94209 21125
rect 4343 20455 4729 20474
rect 4343 20432 4409 20455
rect 4495 20432 4577 20455
rect 4663 20432 4729 20455
rect 4343 20392 4352 20432
rect 4392 20392 4409 20432
rect 4495 20392 4516 20432
rect 4556 20392 4577 20432
rect 4663 20392 4680 20432
rect 4720 20392 4729 20432
rect 4343 20369 4409 20392
rect 4495 20369 4577 20392
rect 4663 20369 4729 20392
rect 4343 20350 4729 20369
rect 19463 20455 19849 20474
rect 19463 20432 19529 20455
rect 19615 20432 19697 20455
rect 19783 20432 19849 20455
rect 19463 20392 19472 20432
rect 19512 20392 19529 20432
rect 19615 20392 19636 20432
rect 19676 20392 19697 20432
rect 19783 20392 19800 20432
rect 19840 20392 19849 20432
rect 19463 20369 19529 20392
rect 19615 20369 19697 20392
rect 19783 20369 19849 20392
rect 19463 20350 19849 20369
rect 34583 20455 34969 20474
rect 34583 20432 34649 20455
rect 34735 20432 34817 20455
rect 34903 20432 34969 20455
rect 34583 20392 34592 20432
rect 34632 20392 34649 20432
rect 34735 20392 34756 20432
rect 34796 20392 34817 20432
rect 34903 20392 34920 20432
rect 34960 20392 34969 20432
rect 34583 20369 34649 20392
rect 34735 20369 34817 20392
rect 34903 20369 34969 20392
rect 34583 20350 34969 20369
rect 49703 20455 50089 20474
rect 49703 20432 49769 20455
rect 49855 20432 49937 20455
rect 50023 20432 50089 20455
rect 49703 20392 49712 20432
rect 49752 20392 49769 20432
rect 49855 20392 49876 20432
rect 49916 20392 49937 20432
rect 50023 20392 50040 20432
rect 50080 20392 50089 20432
rect 49703 20369 49769 20392
rect 49855 20369 49937 20392
rect 50023 20369 50089 20392
rect 49703 20350 50089 20369
rect 64823 20455 65209 20474
rect 64823 20432 64889 20455
rect 64975 20432 65057 20455
rect 65143 20432 65209 20455
rect 64823 20392 64832 20432
rect 64872 20392 64889 20432
rect 64975 20392 64996 20432
rect 65036 20392 65057 20432
rect 65143 20392 65160 20432
rect 65200 20392 65209 20432
rect 64823 20369 64889 20392
rect 64975 20369 65057 20392
rect 65143 20369 65209 20392
rect 64823 20350 65209 20369
rect 79943 20455 80329 20474
rect 79943 20432 80009 20455
rect 80095 20432 80177 20455
rect 80263 20432 80329 20455
rect 79943 20392 79952 20432
rect 79992 20392 80009 20432
rect 80095 20392 80116 20432
rect 80156 20392 80177 20432
rect 80263 20392 80280 20432
rect 80320 20392 80329 20432
rect 79943 20369 80009 20392
rect 80095 20369 80177 20392
rect 80263 20369 80329 20392
rect 79943 20350 80329 20369
rect 95063 20455 95449 20474
rect 95063 20432 95129 20455
rect 95215 20432 95297 20455
rect 95383 20432 95449 20455
rect 95063 20392 95072 20432
rect 95112 20392 95129 20432
rect 95215 20392 95236 20432
rect 95276 20392 95297 20432
rect 95383 20392 95400 20432
rect 95440 20392 95449 20432
rect 95063 20369 95129 20392
rect 95215 20369 95297 20392
rect 95383 20369 95449 20392
rect 95063 20350 95449 20369
rect 3103 19699 3489 19718
rect 3103 19676 3169 19699
rect 3255 19676 3337 19699
rect 3423 19676 3489 19699
rect 3103 19636 3112 19676
rect 3152 19636 3169 19676
rect 3255 19636 3276 19676
rect 3316 19636 3337 19676
rect 3423 19636 3440 19676
rect 3480 19636 3489 19676
rect 3103 19613 3169 19636
rect 3255 19613 3337 19636
rect 3423 19613 3489 19636
rect 3103 19594 3489 19613
rect 18223 19699 18609 19718
rect 18223 19676 18289 19699
rect 18375 19676 18457 19699
rect 18543 19676 18609 19699
rect 18223 19636 18232 19676
rect 18272 19636 18289 19676
rect 18375 19636 18396 19676
rect 18436 19636 18457 19676
rect 18543 19636 18560 19676
rect 18600 19636 18609 19676
rect 18223 19613 18289 19636
rect 18375 19613 18457 19636
rect 18543 19613 18609 19636
rect 18223 19594 18609 19613
rect 33343 19699 33729 19718
rect 33343 19676 33409 19699
rect 33495 19676 33577 19699
rect 33663 19676 33729 19699
rect 33343 19636 33352 19676
rect 33392 19636 33409 19676
rect 33495 19636 33516 19676
rect 33556 19636 33577 19676
rect 33663 19636 33680 19676
rect 33720 19636 33729 19676
rect 33343 19613 33409 19636
rect 33495 19613 33577 19636
rect 33663 19613 33729 19636
rect 33343 19594 33729 19613
rect 48463 19699 48849 19718
rect 48463 19676 48529 19699
rect 48615 19676 48697 19699
rect 48783 19676 48849 19699
rect 48463 19636 48472 19676
rect 48512 19636 48529 19676
rect 48615 19636 48636 19676
rect 48676 19636 48697 19676
rect 48783 19636 48800 19676
rect 48840 19636 48849 19676
rect 48463 19613 48529 19636
rect 48615 19613 48697 19636
rect 48783 19613 48849 19636
rect 48463 19594 48849 19613
rect 63583 19699 63969 19718
rect 63583 19676 63649 19699
rect 63735 19676 63817 19699
rect 63903 19676 63969 19699
rect 63583 19636 63592 19676
rect 63632 19636 63649 19676
rect 63735 19636 63756 19676
rect 63796 19636 63817 19676
rect 63903 19636 63920 19676
rect 63960 19636 63969 19676
rect 63583 19613 63649 19636
rect 63735 19613 63817 19636
rect 63903 19613 63969 19636
rect 63583 19594 63969 19613
rect 78703 19699 79089 19718
rect 78703 19676 78769 19699
rect 78855 19676 78937 19699
rect 79023 19676 79089 19699
rect 78703 19636 78712 19676
rect 78752 19636 78769 19676
rect 78855 19636 78876 19676
rect 78916 19636 78937 19676
rect 79023 19636 79040 19676
rect 79080 19636 79089 19676
rect 78703 19613 78769 19636
rect 78855 19613 78937 19636
rect 79023 19613 79089 19636
rect 78703 19594 79089 19613
rect 93823 19699 94209 19718
rect 93823 19676 93889 19699
rect 93975 19676 94057 19699
rect 94143 19676 94209 19699
rect 93823 19636 93832 19676
rect 93872 19636 93889 19676
rect 93975 19636 93996 19676
rect 94036 19636 94057 19676
rect 94143 19636 94160 19676
rect 94200 19636 94209 19676
rect 93823 19613 93889 19636
rect 93975 19613 94057 19636
rect 94143 19613 94209 19636
rect 93823 19594 94209 19613
rect 4343 18943 4729 18962
rect 4343 18920 4409 18943
rect 4495 18920 4577 18943
rect 4663 18920 4729 18943
rect 4343 18880 4352 18920
rect 4392 18880 4409 18920
rect 4495 18880 4516 18920
rect 4556 18880 4577 18920
rect 4663 18880 4680 18920
rect 4720 18880 4729 18920
rect 4343 18857 4409 18880
rect 4495 18857 4577 18880
rect 4663 18857 4729 18880
rect 4343 18838 4729 18857
rect 19463 18943 19849 18962
rect 19463 18920 19529 18943
rect 19615 18920 19697 18943
rect 19783 18920 19849 18943
rect 19463 18880 19472 18920
rect 19512 18880 19529 18920
rect 19615 18880 19636 18920
rect 19676 18880 19697 18920
rect 19783 18880 19800 18920
rect 19840 18880 19849 18920
rect 19463 18857 19529 18880
rect 19615 18857 19697 18880
rect 19783 18857 19849 18880
rect 19463 18838 19849 18857
rect 34583 18943 34969 18962
rect 34583 18920 34649 18943
rect 34735 18920 34817 18943
rect 34903 18920 34969 18943
rect 34583 18880 34592 18920
rect 34632 18880 34649 18920
rect 34735 18880 34756 18920
rect 34796 18880 34817 18920
rect 34903 18880 34920 18920
rect 34960 18880 34969 18920
rect 34583 18857 34649 18880
rect 34735 18857 34817 18880
rect 34903 18857 34969 18880
rect 34583 18838 34969 18857
rect 49703 18943 50089 18962
rect 49703 18920 49769 18943
rect 49855 18920 49937 18943
rect 50023 18920 50089 18943
rect 49703 18880 49712 18920
rect 49752 18880 49769 18920
rect 49855 18880 49876 18920
rect 49916 18880 49937 18920
rect 50023 18880 50040 18920
rect 50080 18880 50089 18920
rect 49703 18857 49769 18880
rect 49855 18857 49937 18880
rect 50023 18857 50089 18880
rect 49703 18838 50089 18857
rect 64823 18943 65209 18962
rect 64823 18920 64889 18943
rect 64975 18920 65057 18943
rect 65143 18920 65209 18943
rect 64823 18880 64832 18920
rect 64872 18880 64889 18920
rect 64975 18880 64996 18920
rect 65036 18880 65057 18920
rect 65143 18880 65160 18920
rect 65200 18880 65209 18920
rect 64823 18857 64889 18880
rect 64975 18857 65057 18880
rect 65143 18857 65209 18880
rect 64823 18838 65209 18857
rect 79943 18943 80329 18962
rect 79943 18920 80009 18943
rect 80095 18920 80177 18943
rect 80263 18920 80329 18943
rect 79943 18880 79952 18920
rect 79992 18880 80009 18920
rect 80095 18880 80116 18920
rect 80156 18880 80177 18920
rect 80263 18880 80280 18920
rect 80320 18880 80329 18920
rect 79943 18857 80009 18880
rect 80095 18857 80177 18880
rect 80263 18857 80329 18880
rect 79943 18838 80329 18857
rect 95063 18943 95449 18962
rect 95063 18920 95129 18943
rect 95215 18920 95297 18943
rect 95383 18920 95449 18943
rect 95063 18880 95072 18920
rect 95112 18880 95129 18920
rect 95215 18880 95236 18920
rect 95276 18880 95297 18920
rect 95383 18880 95400 18920
rect 95440 18880 95449 18920
rect 95063 18857 95129 18880
rect 95215 18857 95297 18880
rect 95383 18857 95449 18880
rect 95063 18838 95449 18857
rect 3103 18187 3489 18206
rect 3103 18164 3169 18187
rect 3255 18164 3337 18187
rect 3423 18164 3489 18187
rect 3103 18124 3112 18164
rect 3152 18124 3169 18164
rect 3255 18124 3276 18164
rect 3316 18124 3337 18164
rect 3423 18124 3440 18164
rect 3480 18124 3489 18164
rect 3103 18101 3169 18124
rect 3255 18101 3337 18124
rect 3423 18101 3489 18124
rect 3103 18082 3489 18101
rect 18223 18187 18609 18206
rect 18223 18164 18289 18187
rect 18375 18164 18457 18187
rect 18543 18164 18609 18187
rect 18223 18124 18232 18164
rect 18272 18124 18289 18164
rect 18375 18124 18396 18164
rect 18436 18124 18457 18164
rect 18543 18124 18560 18164
rect 18600 18124 18609 18164
rect 18223 18101 18289 18124
rect 18375 18101 18457 18124
rect 18543 18101 18609 18124
rect 18223 18082 18609 18101
rect 33343 18187 33729 18206
rect 33343 18164 33409 18187
rect 33495 18164 33577 18187
rect 33663 18164 33729 18187
rect 33343 18124 33352 18164
rect 33392 18124 33409 18164
rect 33495 18124 33516 18164
rect 33556 18124 33577 18164
rect 33663 18124 33680 18164
rect 33720 18124 33729 18164
rect 33343 18101 33409 18124
rect 33495 18101 33577 18124
rect 33663 18101 33729 18124
rect 33343 18082 33729 18101
rect 48463 18187 48849 18206
rect 48463 18164 48529 18187
rect 48615 18164 48697 18187
rect 48783 18164 48849 18187
rect 48463 18124 48472 18164
rect 48512 18124 48529 18164
rect 48615 18124 48636 18164
rect 48676 18124 48697 18164
rect 48783 18124 48800 18164
rect 48840 18124 48849 18164
rect 48463 18101 48529 18124
rect 48615 18101 48697 18124
rect 48783 18101 48849 18124
rect 48463 18082 48849 18101
rect 63583 18187 63969 18206
rect 63583 18164 63649 18187
rect 63735 18164 63817 18187
rect 63903 18164 63969 18187
rect 63583 18124 63592 18164
rect 63632 18124 63649 18164
rect 63735 18124 63756 18164
rect 63796 18124 63817 18164
rect 63903 18124 63920 18164
rect 63960 18124 63969 18164
rect 63583 18101 63649 18124
rect 63735 18101 63817 18124
rect 63903 18101 63969 18124
rect 63583 18082 63969 18101
rect 78703 18187 79089 18206
rect 78703 18164 78769 18187
rect 78855 18164 78937 18187
rect 79023 18164 79089 18187
rect 78703 18124 78712 18164
rect 78752 18124 78769 18164
rect 78855 18124 78876 18164
rect 78916 18124 78937 18164
rect 79023 18124 79040 18164
rect 79080 18124 79089 18164
rect 78703 18101 78769 18124
rect 78855 18101 78937 18124
rect 79023 18101 79089 18124
rect 78703 18082 79089 18101
rect 93823 18187 94209 18206
rect 93823 18164 93889 18187
rect 93975 18164 94057 18187
rect 94143 18164 94209 18187
rect 93823 18124 93832 18164
rect 93872 18124 93889 18164
rect 93975 18124 93996 18164
rect 94036 18124 94057 18164
rect 94143 18124 94160 18164
rect 94200 18124 94209 18164
rect 93823 18101 93889 18124
rect 93975 18101 94057 18124
rect 94143 18101 94209 18124
rect 93823 18082 94209 18101
rect 4343 17431 4729 17450
rect 4343 17408 4409 17431
rect 4495 17408 4577 17431
rect 4663 17408 4729 17431
rect 4343 17368 4352 17408
rect 4392 17368 4409 17408
rect 4495 17368 4516 17408
rect 4556 17368 4577 17408
rect 4663 17368 4680 17408
rect 4720 17368 4729 17408
rect 4343 17345 4409 17368
rect 4495 17345 4577 17368
rect 4663 17345 4729 17368
rect 4343 17326 4729 17345
rect 19463 17431 19849 17450
rect 19463 17408 19529 17431
rect 19615 17408 19697 17431
rect 19783 17408 19849 17431
rect 19463 17368 19472 17408
rect 19512 17368 19529 17408
rect 19615 17368 19636 17408
rect 19676 17368 19697 17408
rect 19783 17368 19800 17408
rect 19840 17368 19849 17408
rect 19463 17345 19529 17368
rect 19615 17345 19697 17368
rect 19783 17345 19849 17368
rect 19463 17326 19849 17345
rect 34583 17431 34969 17450
rect 34583 17408 34649 17431
rect 34735 17408 34817 17431
rect 34903 17408 34969 17431
rect 34583 17368 34592 17408
rect 34632 17368 34649 17408
rect 34735 17368 34756 17408
rect 34796 17368 34817 17408
rect 34903 17368 34920 17408
rect 34960 17368 34969 17408
rect 34583 17345 34649 17368
rect 34735 17345 34817 17368
rect 34903 17345 34969 17368
rect 34583 17326 34969 17345
rect 49703 17431 50089 17450
rect 49703 17408 49769 17431
rect 49855 17408 49937 17431
rect 50023 17408 50089 17431
rect 49703 17368 49712 17408
rect 49752 17368 49769 17408
rect 49855 17368 49876 17408
rect 49916 17368 49937 17408
rect 50023 17368 50040 17408
rect 50080 17368 50089 17408
rect 49703 17345 49769 17368
rect 49855 17345 49937 17368
rect 50023 17345 50089 17368
rect 49703 17326 50089 17345
rect 64823 17431 65209 17450
rect 64823 17408 64889 17431
rect 64975 17408 65057 17431
rect 65143 17408 65209 17431
rect 64823 17368 64832 17408
rect 64872 17368 64889 17408
rect 64975 17368 64996 17408
rect 65036 17368 65057 17408
rect 65143 17368 65160 17408
rect 65200 17368 65209 17408
rect 64823 17345 64889 17368
rect 64975 17345 65057 17368
rect 65143 17345 65209 17368
rect 64823 17326 65209 17345
rect 79943 17431 80329 17450
rect 79943 17408 80009 17431
rect 80095 17408 80177 17431
rect 80263 17408 80329 17431
rect 79943 17368 79952 17408
rect 79992 17368 80009 17408
rect 80095 17368 80116 17408
rect 80156 17368 80177 17408
rect 80263 17368 80280 17408
rect 80320 17368 80329 17408
rect 79943 17345 80009 17368
rect 80095 17345 80177 17368
rect 80263 17345 80329 17368
rect 79943 17326 80329 17345
rect 95063 17431 95449 17450
rect 95063 17408 95129 17431
rect 95215 17408 95297 17431
rect 95383 17408 95449 17431
rect 95063 17368 95072 17408
rect 95112 17368 95129 17408
rect 95215 17368 95236 17408
rect 95276 17368 95297 17408
rect 95383 17368 95400 17408
rect 95440 17368 95449 17408
rect 95063 17345 95129 17368
rect 95215 17345 95297 17368
rect 95383 17345 95449 17368
rect 95063 17326 95449 17345
rect 3103 16675 3489 16694
rect 3103 16652 3169 16675
rect 3255 16652 3337 16675
rect 3423 16652 3489 16675
rect 3103 16612 3112 16652
rect 3152 16612 3169 16652
rect 3255 16612 3276 16652
rect 3316 16612 3337 16652
rect 3423 16612 3440 16652
rect 3480 16612 3489 16652
rect 3103 16589 3169 16612
rect 3255 16589 3337 16612
rect 3423 16589 3489 16612
rect 3103 16570 3489 16589
rect 18223 16675 18609 16694
rect 18223 16652 18289 16675
rect 18375 16652 18457 16675
rect 18543 16652 18609 16675
rect 18223 16612 18232 16652
rect 18272 16612 18289 16652
rect 18375 16612 18396 16652
rect 18436 16612 18457 16652
rect 18543 16612 18560 16652
rect 18600 16612 18609 16652
rect 18223 16589 18289 16612
rect 18375 16589 18457 16612
rect 18543 16589 18609 16612
rect 18223 16570 18609 16589
rect 33343 16675 33729 16694
rect 33343 16652 33409 16675
rect 33495 16652 33577 16675
rect 33663 16652 33729 16675
rect 33343 16612 33352 16652
rect 33392 16612 33409 16652
rect 33495 16612 33516 16652
rect 33556 16612 33577 16652
rect 33663 16612 33680 16652
rect 33720 16612 33729 16652
rect 33343 16589 33409 16612
rect 33495 16589 33577 16612
rect 33663 16589 33729 16612
rect 33343 16570 33729 16589
rect 48463 16675 48849 16694
rect 48463 16652 48529 16675
rect 48615 16652 48697 16675
rect 48783 16652 48849 16675
rect 48463 16612 48472 16652
rect 48512 16612 48529 16652
rect 48615 16612 48636 16652
rect 48676 16612 48697 16652
rect 48783 16612 48800 16652
rect 48840 16612 48849 16652
rect 48463 16589 48529 16612
rect 48615 16589 48697 16612
rect 48783 16589 48849 16612
rect 48463 16570 48849 16589
rect 63583 16675 63969 16694
rect 63583 16652 63649 16675
rect 63735 16652 63817 16675
rect 63903 16652 63969 16675
rect 63583 16612 63592 16652
rect 63632 16612 63649 16652
rect 63735 16612 63756 16652
rect 63796 16612 63817 16652
rect 63903 16612 63920 16652
rect 63960 16612 63969 16652
rect 63583 16589 63649 16612
rect 63735 16589 63817 16612
rect 63903 16589 63969 16612
rect 63583 16570 63969 16589
rect 78703 16675 79089 16694
rect 78703 16652 78769 16675
rect 78855 16652 78937 16675
rect 79023 16652 79089 16675
rect 78703 16612 78712 16652
rect 78752 16612 78769 16652
rect 78855 16612 78876 16652
rect 78916 16612 78937 16652
rect 79023 16612 79040 16652
rect 79080 16612 79089 16652
rect 78703 16589 78769 16612
rect 78855 16589 78937 16612
rect 79023 16589 79089 16612
rect 78703 16570 79089 16589
rect 93823 16675 94209 16694
rect 93823 16652 93889 16675
rect 93975 16652 94057 16675
rect 94143 16652 94209 16675
rect 93823 16612 93832 16652
rect 93872 16612 93889 16652
rect 93975 16612 93996 16652
rect 94036 16612 94057 16652
rect 94143 16612 94160 16652
rect 94200 16612 94209 16652
rect 93823 16589 93889 16612
rect 93975 16589 94057 16612
rect 94143 16589 94209 16612
rect 93823 16570 94209 16589
rect 4343 15919 4729 15938
rect 4343 15896 4409 15919
rect 4495 15896 4577 15919
rect 4663 15896 4729 15919
rect 4343 15856 4352 15896
rect 4392 15856 4409 15896
rect 4495 15856 4516 15896
rect 4556 15856 4577 15896
rect 4663 15856 4680 15896
rect 4720 15856 4729 15896
rect 4343 15833 4409 15856
rect 4495 15833 4577 15856
rect 4663 15833 4729 15856
rect 4343 15814 4729 15833
rect 19463 15919 19849 15938
rect 19463 15896 19529 15919
rect 19615 15896 19697 15919
rect 19783 15896 19849 15919
rect 19463 15856 19472 15896
rect 19512 15856 19529 15896
rect 19615 15856 19636 15896
rect 19676 15856 19697 15896
rect 19783 15856 19800 15896
rect 19840 15856 19849 15896
rect 19463 15833 19529 15856
rect 19615 15833 19697 15856
rect 19783 15833 19849 15856
rect 19463 15814 19849 15833
rect 34583 15919 34969 15938
rect 34583 15896 34649 15919
rect 34735 15896 34817 15919
rect 34903 15896 34969 15919
rect 34583 15856 34592 15896
rect 34632 15856 34649 15896
rect 34735 15856 34756 15896
rect 34796 15856 34817 15896
rect 34903 15856 34920 15896
rect 34960 15856 34969 15896
rect 34583 15833 34649 15856
rect 34735 15833 34817 15856
rect 34903 15833 34969 15856
rect 34583 15814 34969 15833
rect 49703 15919 50089 15938
rect 49703 15896 49769 15919
rect 49855 15896 49937 15919
rect 50023 15896 50089 15919
rect 49703 15856 49712 15896
rect 49752 15856 49769 15896
rect 49855 15856 49876 15896
rect 49916 15856 49937 15896
rect 50023 15856 50040 15896
rect 50080 15856 50089 15896
rect 49703 15833 49769 15856
rect 49855 15833 49937 15856
rect 50023 15833 50089 15856
rect 49703 15814 50089 15833
rect 64823 15919 65209 15938
rect 64823 15896 64889 15919
rect 64975 15896 65057 15919
rect 65143 15896 65209 15919
rect 64823 15856 64832 15896
rect 64872 15856 64889 15896
rect 64975 15856 64996 15896
rect 65036 15856 65057 15896
rect 65143 15856 65160 15896
rect 65200 15856 65209 15896
rect 64823 15833 64889 15856
rect 64975 15833 65057 15856
rect 65143 15833 65209 15856
rect 64823 15814 65209 15833
rect 79943 15919 80329 15938
rect 79943 15896 80009 15919
rect 80095 15896 80177 15919
rect 80263 15896 80329 15919
rect 79943 15856 79952 15896
rect 79992 15856 80009 15896
rect 80095 15856 80116 15896
rect 80156 15856 80177 15896
rect 80263 15856 80280 15896
rect 80320 15856 80329 15896
rect 79943 15833 80009 15856
rect 80095 15833 80177 15856
rect 80263 15833 80329 15856
rect 79943 15814 80329 15833
rect 95063 15919 95449 15938
rect 95063 15896 95129 15919
rect 95215 15896 95297 15919
rect 95383 15896 95449 15919
rect 95063 15856 95072 15896
rect 95112 15856 95129 15896
rect 95215 15856 95236 15896
rect 95276 15856 95297 15896
rect 95383 15856 95400 15896
rect 95440 15856 95449 15896
rect 95063 15833 95129 15856
rect 95215 15833 95297 15856
rect 95383 15833 95449 15856
rect 95063 15814 95449 15833
rect 3103 15163 3489 15182
rect 3103 15140 3169 15163
rect 3255 15140 3337 15163
rect 3423 15140 3489 15163
rect 3103 15100 3112 15140
rect 3152 15100 3169 15140
rect 3255 15100 3276 15140
rect 3316 15100 3337 15140
rect 3423 15100 3440 15140
rect 3480 15100 3489 15140
rect 3103 15077 3169 15100
rect 3255 15077 3337 15100
rect 3423 15077 3489 15100
rect 3103 15058 3489 15077
rect 18223 15163 18609 15182
rect 18223 15140 18289 15163
rect 18375 15140 18457 15163
rect 18543 15140 18609 15163
rect 18223 15100 18232 15140
rect 18272 15100 18289 15140
rect 18375 15100 18396 15140
rect 18436 15100 18457 15140
rect 18543 15100 18560 15140
rect 18600 15100 18609 15140
rect 18223 15077 18289 15100
rect 18375 15077 18457 15100
rect 18543 15077 18609 15100
rect 18223 15058 18609 15077
rect 33343 15163 33729 15182
rect 33343 15140 33409 15163
rect 33495 15140 33577 15163
rect 33663 15140 33729 15163
rect 33343 15100 33352 15140
rect 33392 15100 33409 15140
rect 33495 15100 33516 15140
rect 33556 15100 33577 15140
rect 33663 15100 33680 15140
rect 33720 15100 33729 15140
rect 33343 15077 33409 15100
rect 33495 15077 33577 15100
rect 33663 15077 33729 15100
rect 33343 15058 33729 15077
rect 48463 15163 48849 15182
rect 48463 15140 48529 15163
rect 48615 15140 48697 15163
rect 48783 15140 48849 15163
rect 48463 15100 48472 15140
rect 48512 15100 48529 15140
rect 48615 15100 48636 15140
rect 48676 15100 48697 15140
rect 48783 15100 48800 15140
rect 48840 15100 48849 15140
rect 48463 15077 48529 15100
rect 48615 15077 48697 15100
rect 48783 15077 48849 15100
rect 48463 15058 48849 15077
rect 63583 15163 63969 15182
rect 63583 15140 63649 15163
rect 63735 15140 63817 15163
rect 63903 15140 63969 15163
rect 63583 15100 63592 15140
rect 63632 15100 63649 15140
rect 63735 15100 63756 15140
rect 63796 15100 63817 15140
rect 63903 15100 63920 15140
rect 63960 15100 63969 15140
rect 63583 15077 63649 15100
rect 63735 15077 63817 15100
rect 63903 15077 63969 15100
rect 63583 15058 63969 15077
rect 78703 15163 79089 15182
rect 78703 15140 78769 15163
rect 78855 15140 78937 15163
rect 79023 15140 79089 15163
rect 78703 15100 78712 15140
rect 78752 15100 78769 15140
rect 78855 15100 78876 15140
rect 78916 15100 78937 15140
rect 79023 15100 79040 15140
rect 79080 15100 79089 15140
rect 78703 15077 78769 15100
rect 78855 15077 78937 15100
rect 79023 15077 79089 15100
rect 78703 15058 79089 15077
rect 93823 15163 94209 15182
rect 93823 15140 93889 15163
rect 93975 15140 94057 15163
rect 94143 15140 94209 15163
rect 93823 15100 93832 15140
rect 93872 15100 93889 15140
rect 93975 15100 93996 15140
rect 94036 15100 94057 15140
rect 94143 15100 94160 15140
rect 94200 15100 94209 15140
rect 93823 15077 93889 15100
rect 93975 15077 94057 15100
rect 94143 15077 94209 15100
rect 93823 15058 94209 15077
rect 4343 14407 4729 14426
rect 4343 14384 4409 14407
rect 4495 14384 4577 14407
rect 4663 14384 4729 14407
rect 4343 14344 4352 14384
rect 4392 14344 4409 14384
rect 4495 14344 4516 14384
rect 4556 14344 4577 14384
rect 4663 14344 4680 14384
rect 4720 14344 4729 14384
rect 4343 14321 4409 14344
rect 4495 14321 4577 14344
rect 4663 14321 4729 14344
rect 4343 14302 4729 14321
rect 19463 14407 19849 14426
rect 19463 14384 19529 14407
rect 19615 14384 19697 14407
rect 19783 14384 19849 14407
rect 19463 14344 19472 14384
rect 19512 14344 19529 14384
rect 19615 14344 19636 14384
rect 19676 14344 19697 14384
rect 19783 14344 19800 14384
rect 19840 14344 19849 14384
rect 19463 14321 19529 14344
rect 19615 14321 19697 14344
rect 19783 14321 19849 14344
rect 19463 14302 19849 14321
rect 34583 14407 34969 14426
rect 34583 14384 34649 14407
rect 34735 14384 34817 14407
rect 34903 14384 34969 14407
rect 34583 14344 34592 14384
rect 34632 14344 34649 14384
rect 34735 14344 34756 14384
rect 34796 14344 34817 14384
rect 34903 14344 34920 14384
rect 34960 14344 34969 14384
rect 34583 14321 34649 14344
rect 34735 14321 34817 14344
rect 34903 14321 34969 14344
rect 34583 14302 34969 14321
rect 49703 14407 50089 14426
rect 49703 14384 49769 14407
rect 49855 14384 49937 14407
rect 50023 14384 50089 14407
rect 49703 14344 49712 14384
rect 49752 14344 49769 14384
rect 49855 14344 49876 14384
rect 49916 14344 49937 14384
rect 50023 14344 50040 14384
rect 50080 14344 50089 14384
rect 49703 14321 49769 14344
rect 49855 14321 49937 14344
rect 50023 14321 50089 14344
rect 49703 14302 50089 14321
rect 64823 14407 65209 14426
rect 64823 14384 64889 14407
rect 64975 14384 65057 14407
rect 65143 14384 65209 14407
rect 64823 14344 64832 14384
rect 64872 14344 64889 14384
rect 64975 14344 64996 14384
rect 65036 14344 65057 14384
rect 65143 14344 65160 14384
rect 65200 14344 65209 14384
rect 64823 14321 64889 14344
rect 64975 14321 65057 14344
rect 65143 14321 65209 14344
rect 64823 14302 65209 14321
rect 79943 14407 80329 14426
rect 79943 14384 80009 14407
rect 80095 14384 80177 14407
rect 80263 14384 80329 14407
rect 79943 14344 79952 14384
rect 79992 14344 80009 14384
rect 80095 14344 80116 14384
rect 80156 14344 80177 14384
rect 80263 14344 80280 14384
rect 80320 14344 80329 14384
rect 79943 14321 80009 14344
rect 80095 14321 80177 14344
rect 80263 14321 80329 14344
rect 79943 14302 80329 14321
rect 95063 14407 95449 14426
rect 95063 14384 95129 14407
rect 95215 14384 95297 14407
rect 95383 14384 95449 14407
rect 95063 14344 95072 14384
rect 95112 14344 95129 14384
rect 95215 14344 95236 14384
rect 95276 14344 95297 14384
rect 95383 14344 95400 14384
rect 95440 14344 95449 14384
rect 95063 14321 95129 14344
rect 95215 14321 95297 14344
rect 95383 14321 95449 14344
rect 95063 14302 95449 14321
rect 3103 13651 3489 13670
rect 3103 13628 3169 13651
rect 3255 13628 3337 13651
rect 3423 13628 3489 13651
rect 3103 13588 3112 13628
rect 3152 13588 3169 13628
rect 3255 13588 3276 13628
rect 3316 13588 3337 13628
rect 3423 13588 3440 13628
rect 3480 13588 3489 13628
rect 3103 13565 3169 13588
rect 3255 13565 3337 13588
rect 3423 13565 3489 13588
rect 3103 13546 3489 13565
rect 18223 13651 18609 13670
rect 18223 13628 18289 13651
rect 18375 13628 18457 13651
rect 18543 13628 18609 13651
rect 18223 13588 18232 13628
rect 18272 13588 18289 13628
rect 18375 13588 18396 13628
rect 18436 13588 18457 13628
rect 18543 13588 18560 13628
rect 18600 13588 18609 13628
rect 18223 13565 18289 13588
rect 18375 13565 18457 13588
rect 18543 13565 18609 13588
rect 18223 13546 18609 13565
rect 33343 13651 33729 13670
rect 33343 13628 33409 13651
rect 33495 13628 33577 13651
rect 33663 13628 33729 13651
rect 33343 13588 33352 13628
rect 33392 13588 33409 13628
rect 33495 13588 33516 13628
rect 33556 13588 33577 13628
rect 33663 13588 33680 13628
rect 33720 13588 33729 13628
rect 33343 13565 33409 13588
rect 33495 13565 33577 13588
rect 33663 13565 33729 13588
rect 33343 13546 33729 13565
rect 48463 13651 48849 13670
rect 48463 13628 48529 13651
rect 48615 13628 48697 13651
rect 48783 13628 48849 13651
rect 48463 13588 48472 13628
rect 48512 13588 48529 13628
rect 48615 13588 48636 13628
rect 48676 13588 48697 13628
rect 48783 13588 48800 13628
rect 48840 13588 48849 13628
rect 48463 13565 48529 13588
rect 48615 13565 48697 13588
rect 48783 13565 48849 13588
rect 48463 13546 48849 13565
rect 63583 13651 63969 13670
rect 63583 13628 63649 13651
rect 63735 13628 63817 13651
rect 63903 13628 63969 13651
rect 63583 13588 63592 13628
rect 63632 13588 63649 13628
rect 63735 13588 63756 13628
rect 63796 13588 63817 13628
rect 63903 13588 63920 13628
rect 63960 13588 63969 13628
rect 63583 13565 63649 13588
rect 63735 13565 63817 13588
rect 63903 13565 63969 13588
rect 63583 13546 63969 13565
rect 78703 13651 79089 13670
rect 78703 13628 78769 13651
rect 78855 13628 78937 13651
rect 79023 13628 79089 13651
rect 78703 13588 78712 13628
rect 78752 13588 78769 13628
rect 78855 13588 78876 13628
rect 78916 13588 78937 13628
rect 79023 13588 79040 13628
rect 79080 13588 79089 13628
rect 78703 13565 78769 13588
rect 78855 13565 78937 13588
rect 79023 13565 79089 13588
rect 78703 13546 79089 13565
rect 93823 13651 94209 13670
rect 93823 13628 93889 13651
rect 93975 13628 94057 13651
rect 94143 13628 94209 13651
rect 93823 13588 93832 13628
rect 93872 13588 93889 13628
rect 93975 13588 93996 13628
rect 94036 13588 94057 13628
rect 94143 13588 94160 13628
rect 94200 13588 94209 13628
rect 93823 13565 93889 13588
rect 93975 13565 94057 13588
rect 94143 13565 94209 13588
rect 93823 13546 94209 13565
rect 4343 12895 4729 12914
rect 4343 12872 4409 12895
rect 4495 12872 4577 12895
rect 4663 12872 4729 12895
rect 4343 12832 4352 12872
rect 4392 12832 4409 12872
rect 4495 12832 4516 12872
rect 4556 12832 4577 12872
rect 4663 12832 4680 12872
rect 4720 12832 4729 12872
rect 4343 12809 4409 12832
rect 4495 12809 4577 12832
rect 4663 12809 4729 12832
rect 4343 12790 4729 12809
rect 19463 12895 19849 12914
rect 19463 12872 19529 12895
rect 19615 12872 19697 12895
rect 19783 12872 19849 12895
rect 19463 12832 19472 12872
rect 19512 12832 19529 12872
rect 19615 12832 19636 12872
rect 19676 12832 19697 12872
rect 19783 12832 19800 12872
rect 19840 12832 19849 12872
rect 19463 12809 19529 12832
rect 19615 12809 19697 12832
rect 19783 12809 19849 12832
rect 19463 12790 19849 12809
rect 34583 12895 34969 12914
rect 34583 12872 34649 12895
rect 34735 12872 34817 12895
rect 34903 12872 34969 12895
rect 34583 12832 34592 12872
rect 34632 12832 34649 12872
rect 34735 12832 34756 12872
rect 34796 12832 34817 12872
rect 34903 12832 34920 12872
rect 34960 12832 34969 12872
rect 34583 12809 34649 12832
rect 34735 12809 34817 12832
rect 34903 12809 34969 12832
rect 34583 12790 34969 12809
rect 49703 12895 50089 12914
rect 49703 12872 49769 12895
rect 49855 12872 49937 12895
rect 50023 12872 50089 12895
rect 49703 12832 49712 12872
rect 49752 12832 49769 12872
rect 49855 12832 49876 12872
rect 49916 12832 49937 12872
rect 50023 12832 50040 12872
rect 50080 12832 50089 12872
rect 49703 12809 49769 12832
rect 49855 12809 49937 12832
rect 50023 12809 50089 12832
rect 49703 12790 50089 12809
rect 64823 12895 65209 12914
rect 64823 12872 64889 12895
rect 64975 12872 65057 12895
rect 65143 12872 65209 12895
rect 64823 12832 64832 12872
rect 64872 12832 64889 12872
rect 64975 12832 64996 12872
rect 65036 12832 65057 12872
rect 65143 12832 65160 12872
rect 65200 12832 65209 12872
rect 64823 12809 64889 12832
rect 64975 12809 65057 12832
rect 65143 12809 65209 12832
rect 64823 12790 65209 12809
rect 79943 12895 80329 12914
rect 79943 12872 80009 12895
rect 80095 12872 80177 12895
rect 80263 12872 80329 12895
rect 79943 12832 79952 12872
rect 79992 12832 80009 12872
rect 80095 12832 80116 12872
rect 80156 12832 80177 12872
rect 80263 12832 80280 12872
rect 80320 12832 80329 12872
rect 79943 12809 80009 12832
rect 80095 12809 80177 12832
rect 80263 12809 80329 12832
rect 79943 12790 80329 12809
rect 95063 12895 95449 12914
rect 95063 12872 95129 12895
rect 95215 12872 95297 12895
rect 95383 12872 95449 12895
rect 95063 12832 95072 12872
rect 95112 12832 95129 12872
rect 95215 12832 95236 12872
rect 95276 12832 95297 12872
rect 95383 12832 95400 12872
rect 95440 12832 95449 12872
rect 95063 12809 95129 12832
rect 95215 12809 95297 12832
rect 95383 12809 95449 12832
rect 95063 12790 95449 12809
rect 3103 12139 3489 12158
rect 3103 12116 3169 12139
rect 3255 12116 3337 12139
rect 3423 12116 3489 12139
rect 3103 12076 3112 12116
rect 3152 12076 3169 12116
rect 3255 12076 3276 12116
rect 3316 12076 3337 12116
rect 3423 12076 3440 12116
rect 3480 12076 3489 12116
rect 3103 12053 3169 12076
rect 3255 12053 3337 12076
rect 3423 12053 3489 12076
rect 3103 12034 3489 12053
rect 18223 12139 18609 12158
rect 18223 12116 18289 12139
rect 18375 12116 18457 12139
rect 18543 12116 18609 12139
rect 18223 12076 18232 12116
rect 18272 12076 18289 12116
rect 18375 12076 18396 12116
rect 18436 12076 18457 12116
rect 18543 12076 18560 12116
rect 18600 12076 18609 12116
rect 18223 12053 18289 12076
rect 18375 12053 18457 12076
rect 18543 12053 18609 12076
rect 18223 12034 18609 12053
rect 33343 12139 33729 12158
rect 33343 12116 33409 12139
rect 33495 12116 33577 12139
rect 33663 12116 33729 12139
rect 33343 12076 33352 12116
rect 33392 12076 33409 12116
rect 33495 12076 33516 12116
rect 33556 12076 33577 12116
rect 33663 12076 33680 12116
rect 33720 12076 33729 12116
rect 33343 12053 33409 12076
rect 33495 12053 33577 12076
rect 33663 12053 33729 12076
rect 33343 12034 33729 12053
rect 48463 12139 48849 12158
rect 48463 12116 48529 12139
rect 48615 12116 48697 12139
rect 48783 12116 48849 12139
rect 48463 12076 48472 12116
rect 48512 12076 48529 12116
rect 48615 12076 48636 12116
rect 48676 12076 48697 12116
rect 48783 12076 48800 12116
rect 48840 12076 48849 12116
rect 48463 12053 48529 12076
rect 48615 12053 48697 12076
rect 48783 12053 48849 12076
rect 48463 12034 48849 12053
rect 63583 12139 63969 12158
rect 63583 12116 63649 12139
rect 63735 12116 63817 12139
rect 63903 12116 63969 12139
rect 63583 12076 63592 12116
rect 63632 12076 63649 12116
rect 63735 12076 63756 12116
rect 63796 12076 63817 12116
rect 63903 12076 63920 12116
rect 63960 12076 63969 12116
rect 63583 12053 63649 12076
rect 63735 12053 63817 12076
rect 63903 12053 63969 12076
rect 63583 12034 63969 12053
rect 78703 12139 79089 12158
rect 78703 12116 78769 12139
rect 78855 12116 78937 12139
rect 79023 12116 79089 12139
rect 78703 12076 78712 12116
rect 78752 12076 78769 12116
rect 78855 12076 78876 12116
rect 78916 12076 78937 12116
rect 79023 12076 79040 12116
rect 79080 12076 79089 12116
rect 78703 12053 78769 12076
rect 78855 12053 78937 12076
rect 79023 12053 79089 12076
rect 78703 12034 79089 12053
rect 93823 12139 94209 12158
rect 93823 12116 93889 12139
rect 93975 12116 94057 12139
rect 94143 12116 94209 12139
rect 93823 12076 93832 12116
rect 93872 12076 93889 12116
rect 93975 12076 93996 12116
rect 94036 12076 94057 12116
rect 94143 12076 94160 12116
rect 94200 12076 94209 12116
rect 93823 12053 93889 12076
rect 93975 12053 94057 12076
rect 94143 12053 94209 12076
rect 93823 12034 94209 12053
rect 4343 11383 4729 11402
rect 4343 11360 4409 11383
rect 4495 11360 4577 11383
rect 4663 11360 4729 11383
rect 4343 11320 4352 11360
rect 4392 11320 4409 11360
rect 4495 11320 4516 11360
rect 4556 11320 4577 11360
rect 4663 11320 4680 11360
rect 4720 11320 4729 11360
rect 4343 11297 4409 11320
rect 4495 11297 4577 11320
rect 4663 11297 4729 11320
rect 4343 11278 4729 11297
rect 19463 11383 19849 11402
rect 19463 11360 19529 11383
rect 19615 11360 19697 11383
rect 19783 11360 19849 11383
rect 19463 11320 19472 11360
rect 19512 11320 19529 11360
rect 19615 11320 19636 11360
rect 19676 11320 19697 11360
rect 19783 11320 19800 11360
rect 19840 11320 19849 11360
rect 19463 11297 19529 11320
rect 19615 11297 19697 11320
rect 19783 11297 19849 11320
rect 19463 11278 19849 11297
rect 34583 11383 34969 11402
rect 34583 11360 34649 11383
rect 34735 11360 34817 11383
rect 34903 11360 34969 11383
rect 34583 11320 34592 11360
rect 34632 11320 34649 11360
rect 34735 11320 34756 11360
rect 34796 11320 34817 11360
rect 34903 11320 34920 11360
rect 34960 11320 34969 11360
rect 34583 11297 34649 11320
rect 34735 11297 34817 11320
rect 34903 11297 34969 11320
rect 34583 11278 34969 11297
rect 49703 11383 50089 11402
rect 49703 11360 49769 11383
rect 49855 11360 49937 11383
rect 50023 11360 50089 11383
rect 49703 11320 49712 11360
rect 49752 11320 49769 11360
rect 49855 11320 49876 11360
rect 49916 11320 49937 11360
rect 50023 11320 50040 11360
rect 50080 11320 50089 11360
rect 49703 11297 49769 11320
rect 49855 11297 49937 11320
rect 50023 11297 50089 11320
rect 49703 11278 50089 11297
rect 64823 11383 65209 11402
rect 64823 11360 64889 11383
rect 64975 11360 65057 11383
rect 65143 11360 65209 11383
rect 64823 11320 64832 11360
rect 64872 11320 64889 11360
rect 64975 11320 64996 11360
rect 65036 11320 65057 11360
rect 65143 11320 65160 11360
rect 65200 11320 65209 11360
rect 64823 11297 64889 11320
rect 64975 11297 65057 11320
rect 65143 11297 65209 11320
rect 64823 11278 65209 11297
rect 79943 11383 80329 11402
rect 79943 11360 80009 11383
rect 80095 11360 80177 11383
rect 80263 11360 80329 11383
rect 79943 11320 79952 11360
rect 79992 11320 80009 11360
rect 80095 11320 80116 11360
rect 80156 11320 80177 11360
rect 80263 11320 80280 11360
rect 80320 11320 80329 11360
rect 79943 11297 80009 11320
rect 80095 11297 80177 11320
rect 80263 11297 80329 11320
rect 79943 11278 80329 11297
rect 95063 11383 95449 11402
rect 95063 11360 95129 11383
rect 95215 11360 95297 11383
rect 95383 11360 95449 11383
rect 95063 11320 95072 11360
rect 95112 11320 95129 11360
rect 95215 11320 95236 11360
rect 95276 11320 95297 11360
rect 95383 11320 95400 11360
rect 95440 11320 95449 11360
rect 95063 11297 95129 11320
rect 95215 11297 95297 11320
rect 95383 11297 95449 11320
rect 95063 11278 95449 11297
rect 3103 10627 3489 10646
rect 3103 10604 3169 10627
rect 3255 10604 3337 10627
rect 3423 10604 3489 10627
rect 3103 10564 3112 10604
rect 3152 10564 3169 10604
rect 3255 10564 3276 10604
rect 3316 10564 3337 10604
rect 3423 10564 3440 10604
rect 3480 10564 3489 10604
rect 3103 10541 3169 10564
rect 3255 10541 3337 10564
rect 3423 10541 3489 10564
rect 3103 10522 3489 10541
rect 18223 10627 18609 10646
rect 18223 10604 18289 10627
rect 18375 10604 18457 10627
rect 18543 10604 18609 10627
rect 18223 10564 18232 10604
rect 18272 10564 18289 10604
rect 18375 10564 18396 10604
rect 18436 10564 18457 10604
rect 18543 10564 18560 10604
rect 18600 10564 18609 10604
rect 18223 10541 18289 10564
rect 18375 10541 18457 10564
rect 18543 10541 18609 10564
rect 18223 10522 18609 10541
rect 33343 10627 33729 10646
rect 33343 10604 33409 10627
rect 33495 10604 33577 10627
rect 33663 10604 33729 10627
rect 33343 10564 33352 10604
rect 33392 10564 33409 10604
rect 33495 10564 33516 10604
rect 33556 10564 33577 10604
rect 33663 10564 33680 10604
rect 33720 10564 33729 10604
rect 33343 10541 33409 10564
rect 33495 10541 33577 10564
rect 33663 10541 33729 10564
rect 33343 10522 33729 10541
rect 48463 10627 48849 10646
rect 48463 10604 48529 10627
rect 48615 10604 48697 10627
rect 48783 10604 48849 10627
rect 48463 10564 48472 10604
rect 48512 10564 48529 10604
rect 48615 10564 48636 10604
rect 48676 10564 48697 10604
rect 48783 10564 48800 10604
rect 48840 10564 48849 10604
rect 48463 10541 48529 10564
rect 48615 10541 48697 10564
rect 48783 10541 48849 10564
rect 48463 10522 48849 10541
rect 63583 10627 63969 10646
rect 63583 10604 63649 10627
rect 63735 10604 63817 10627
rect 63903 10604 63969 10627
rect 63583 10564 63592 10604
rect 63632 10564 63649 10604
rect 63735 10564 63756 10604
rect 63796 10564 63817 10604
rect 63903 10564 63920 10604
rect 63960 10564 63969 10604
rect 63583 10541 63649 10564
rect 63735 10541 63817 10564
rect 63903 10541 63969 10564
rect 63583 10522 63969 10541
rect 78703 10627 79089 10646
rect 78703 10604 78769 10627
rect 78855 10604 78937 10627
rect 79023 10604 79089 10627
rect 78703 10564 78712 10604
rect 78752 10564 78769 10604
rect 78855 10564 78876 10604
rect 78916 10564 78937 10604
rect 79023 10564 79040 10604
rect 79080 10564 79089 10604
rect 78703 10541 78769 10564
rect 78855 10541 78937 10564
rect 79023 10541 79089 10564
rect 78703 10522 79089 10541
rect 93823 10627 94209 10646
rect 93823 10604 93889 10627
rect 93975 10604 94057 10627
rect 94143 10604 94209 10627
rect 93823 10564 93832 10604
rect 93872 10564 93889 10604
rect 93975 10564 93996 10604
rect 94036 10564 94057 10604
rect 94143 10564 94160 10604
rect 94200 10564 94209 10604
rect 93823 10541 93889 10564
rect 93975 10541 94057 10564
rect 94143 10541 94209 10564
rect 93823 10522 94209 10541
rect 4343 9871 4729 9890
rect 4343 9848 4409 9871
rect 4495 9848 4577 9871
rect 4663 9848 4729 9871
rect 4343 9808 4352 9848
rect 4392 9808 4409 9848
rect 4495 9808 4516 9848
rect 4556 9808 4577 9848
rect 4663 9808 4680 9848
rect 4720 9808 4729 9848
rect 4343 9785 4409 9808
rect 4495 9785 4577 9808
rect 4663 9785 4729 9808
rect 4343 9766 4729 9785
rect 19463 9871 19849 9890
rect 19463 9848 19529 9871
rect 19615 9848 19697 9871
rect 19783 9848 19849 9871
rect 19463 9808 19472 9848
rect 19512 9808 19529 9848
rect 19615 9808 19636 9848
rect 19676 9808 19697 9848
rect 19783 9808 19800 9848
rect 19840 9808 19849 9848
rect 19463 9785 19529 9808
rect 19615 9785 19697 9808
rect 19783 9785 19849 9808
rect 19463 9766 19849 9785
rect 34583 9871 34969 9890
rect 34583 9848 34649 9871
rect 34735 9848 34817 9871
rect 34903 9848 34969 9871
rect 34583 9808 34592 9848
rect 34632 9808 34649 9848
rect 34735 9808 34756 9848
rect 34796 9808 34817 9848
rect 34903 9808 34920 9848
rect 34960 9808 34969 9848
rect 34583 9785 34649 9808
rect 34735 9785 34817 9808
rect 34903 9785 34969 9808
rect 34583 9766 34969 9785
rect 49703 9871 50089 9890
rect 49703 9848 49769 9871
rect 49855 9848 49937 9871
rect 50023 9848 50089 9871
rect 49703 9808 49712 9848
rect 49752 9808 49769 9848
rect 49855 9808 49876 9848
rect 49916 9808 49937 9848
rect 50023 9808 50040 9848
rect 50080 9808 50089 9848
rect 49703 9785 49769 9808
rect 49855 9785 49937 9808
rect 50023 9785 50089 9808
rect 49703 9766 50089 9785
rect 64823 9871 65209 9890
rect 64823 9848 64889 9871
rect 64975 9848 65057 9871
rect 65143 9848 65209 9871
rect 64823 9808 64832 9848
rect 64872 9808 64889 9848
rect 64975 9808 64996 9848
rect 65036 9808 65057 9848
rect 65143 9808 65160 9848
rect 65200 9808 65209 9848
rect 64823 9785 64889 9808
rect 64975 9785 65057 9808
rect 65143 9785 65209 9808
rect 64823 9766 65209 9785
rect 79943 9871 80329 9890
rect 79943 9848 80009 9871
rect 80095 9848 80177 9871
rect 80263 9848 80329 9871
rect 79943 9808 79952 9848
rect 79992 9808 80009 9848
rect 80095 9808 80116 9848
rect 80156 9808 80177 9848
rect 80263 9808 80280 9848
rect 80320 9808 80329 9848
rect 79943 9785 80009 9808
rect 80095 9785 80177 9808
rect 80263 9785 80329 9808
rect 79943 9766 80329 9785
rect 95063 9871 95449 9890
rect 95063 9848 95129 9871
rect 95215 9848 95297 9871
rect 95383 9848 95449 9871
rect 95063 9808 95072 9848
rect 95112 9808 95129 9848
rect 95215 9808 95236 9848
rect 95276 9808 95297 9848
rect 95383 9808 95400 9848
rect 95440 9808 95449 9848
rect 95063 9785 95129 9808
rect 95215 9785 95297 9808
rect 95383 9785 95449 9808
rect 95063 9766 95449 9785
rect 3103 9115 3489 9134
rect 3103 9092 3169 9115
rect 3255 9092 3337 9115
rect 3423 9092 3489 9115
rect 3103 9052 3112 9092
rect 3152 9052 3169 9092
rect 3255 9052 3276 9092
rect 3316 9052 3337 9092
rect 3423 9052 3440 9092
rect 3480 9052 3489 9092
rect 3103 9029 3169 9052
rect 3255 9029 3337 9052
rect 3423 9029 3489 9052
rect 3103 9010 3489 9029
rect 18223 9115 18609 9134
rect 18223 9092 18289 9115
rect 18375 9092 18457 9115
rect 18543 9092 18609 9115
rect 18223 9052 18232 9092
rect 18272 9052 18289 9092
rect 18375 9052 18396 9092
rect 18436 9052 18457 9092
rect 18543 9052 18560 9092
rect 18600 9052 18609 9092
rect 18223 9029 18289 9052
rect 18375 9029 18457 9052
rect 18543 9029 18609 9052
rect 18223 9010 18609 9029
rect 33343 9115 33729 9134
rect 33343 9092 33409 9115
rect 33495 9092 33577 9115
rect 33663 9092 33729 9115
rect 33343 9052 33352 9092
rect 33392 9052 33409 9092
rect 33495 9052 33516 9092
rect 33556 9052 33577 9092
rect 33663 9052 33680 9092
rect 33720 9052 33729 9092
rect 33343 9029 33409 9052
rect 33495 9029 33577 9052
rect 33663 9029 33729 9052
rect 33343 9010 33729 9029
rect 48463 9115 48849 9134
rect 48463 9092 48529 9115
rect 48615 9092 48697 9115
rect 48783 9092 48849 9115
rect 48463 9052 48472 9092
rect 48512 9052 48529 9092
rect 48615 9052 48636 9092
rect 48676 9052 48697 9092
rect 48783 9052 48800 9092
rect 48840 9052 48849 9092
rect 48463 9029 48529 9052
rect 48615 9029 48697 9052
rect 48783 9029 48849 9052
rect 48463 9010 48849 9029
rect 63583 9115 63969 9134
rect 63583 9092 63649 9115
rect 63735 9092 63817 9115
rect 63903 9092 63969 9115
rect 63583 9052 63592 9092
rect 63632 9052 63649 9092
rect 63735 9052 63756 9092
rect 63796 9052 63817 9092
rect 63903 9052 63920 9092
rect 63960 9052 63969 9092
rect 63583 9029 63649 9052
rect 63735 9029 63817 9052
rect 63903 9029 63969 9052
rect 63583 9010 63969 9029
rect 78703 9115 79089 9134
rect 78703 9092 78769 9115
rect 78855 9092 78937 9115
rect 79023 9092 79089 9115
rect 78703 9052 78712 9092
rect 78752 9052 78769 9092
rect 78855 9052 78876 9092
rect 78916 9052 78937 9092
rect 79023 9052 79040 9092
rect 79080 9052 79089 9092
rect 78703 9029 78769 9052
rect 78855 9029 78937 9052
rect 79023 9029 79089 9052
rect 78703 9010 79089 9029
rect 93823 9115 94209 9134
rect 93823 9092 93889 9115
rect 93975 9092 94057 9115
rect 94143 9092 94209 9115
rect 93823 9052 93832 9092
rect 93872 9052 93889 9092
rect 93975 9052 93996 9092
rect 94036 9052 94057 9092
rect 94143 9052 94160 9092
rect 94200 9052 94209 9092
rect 93823 9029 93889 9052
rect 93975 9029 94057 9052
rect 94143 9029 94209 9052
rect 93823 9010 94209 9029
rect 4343 8359 4729 8378
rect 4343 8336 4409 8359
rect 4495 8336 4577 8359
rect 4663 8336 4729 8359
rect 4343 8296 4352 8336
rect 4392 8296 4409 8336
rect 4495 8296 4516 8336
rect 4556 8296 4577 8336
rect 4663 8296 4680 8336
rect 4720 8296 4729 8336
rect 4343 8273 4409 8296
rect 4495 8273 4577 8296
rect 4663 8273 4729 8296
rect 4343 8254 4729 8273
rect 19463 8359 19849 8378
rect 19463 8336 19529 8359
rect 19615 8336 19697 8359
rect 19783 8336 19849 8359
rect 19463 8296 19472 8336
rect 19512 8296 19529 8336
rect 19615 8296 19636 8336
rect 19676 8296 19697 8336
rect 19783 8296 19800 8336
rect 19840 8296 19849 8336
rect 19463 8273 19529 8296
rect 19615 8273 19697 8296
rect 19783 8273 19849 8296
rect 19463 8254 19849 8273
rect 34583 8359 34969 8378
rect 34583 8336 34649 8359
rect 34735 8336 34817 8359
rect 34903 8336 34969 8359
rect 34583 8296 34592 8336
rect 34632 8296 34649 8336
rect 34735 8296 34756 8336
rect 34796 8296 34817 8336
rect 34903 8296 34920 8336
rect 34960 8296 34969 8336
rect 34583 8273 34649 8296
rect 34735 8273 34817 8296
rect 34903 8273 34969 8296
rect 34583 8254 34969 8273
rect 49703 8359 50089 8378
rect 49703 8336 49769 8359
rect 49855 8336 49937 8359
rect 50023 8336 50089 8359
rect 49703 8296 49712 8336
rect 49752 8296 49769 8336
rect 49855 8296 49876 8336
rect 49916 8296 49937 8336
rect 50023 8296 50040 8336
rect 50080 8296 50089 8336
rect 49703 8273 49769 8296
rect 49855 8273 49937 8296
rect 50023 8273 50089 8296
rect 49703 8254 50089 8273
rect 64823 8359 65209 8378
rect 64823 8336 64889 8359
rect 64975 8336 65057 8359
rect 65143 8336 65209 8359
rect 64823 8296 64832 8336
rect 64872 8296 64889 8336
rect 64975 8296 64996 8336
rect 65036 8296 65057 8336
rect 65143 8296 65160 8336
rect 65200 8296 65209 8336
rect 64823 8273 64889 8296
rect 64975 8273 65057 8296
rect 65143 8273 65209 8296
rect 64823 8254 65209 8273
rect 79943 8359 80329 8378
rect 79943 8336 80009 8359
rect 80095 8336 80177 8359
rect 80263 8336 80329 8359
rect 79943 8296 79952 8336
rect 79992 8296 80009 8336
rect 80095 8296 80116 8336
rect 80156 8296 80177 8336
rect 80263 8296 80280 8336
rect 80320 8296 80329 8336
rect 79943 8273 80009 8296
rect 80095 8273 80177 8296
rect 80263 8273 80329 8296
rect 79943 8254 80329 8273
rect 95063 8359 95449 8378
rect 95063 8336 95129 8359
rect 95215 8336 95297 8359
rect 95383 8336 95449 8359
rect 95063 8296 95072 8336
rect 95112 8296 95129 8336
rect 95215 8296 95236 8336
rect 95276 8296 95297 8336
rect 95383 8296 95400 8336
rect 95440 8296 95449 8336
rect 95063 8273 95129 8296
rect 95215 8273 95297 8296
rect 95383 8273 95449 8296
rect 95063 8254 95449 8273
rect 3103 7603 3489 7622
rect 3103 7580 3169 7603
rect 3255 7580 3337 7603
rect 3423 7580 3489 7603
rect 3103 7540 3112 7580
rect 3152 7540 3169 7580
rect 3255 7540 3276 7580
rect 3316 7540 3337 7580
rect 3423 7540 3440 7580
rect 3480 7540 3489 7580
rect 3103 7517 3169 7540
rect 3255 7517 3337 7540
rect 3423 7517 3489 7540
rect 3103 7498 3489 7517
rect 18223 7603 18609 7622
rect 18223 7580 18289 7603
rect 18375 7580 18457 7603
rect 18543 7580 18609 7603
rect 18223 7540 18232 7580
rect 18272 7540 18289 7580
rect 18375 7540 18396 7580
rect 18436 7540 18457 7580
rect 18543 7540 18560 7580
rect 18600 7540 18609 7580
rect 18223 7517 18289 7540
rect 18375 7517 18457 7540
rect 18543 7517 18609 7540
rect 18223 7498 18609 7517
rect 33343 7603 33729 7622
rect 33343 7580 33409 7603
rect 33495 7580 33577 7603
rect 33663 7580 33729 7603
rect 33343 7540 33352 7580
rect 33392 7540 33409 7580
rect 33495 7540 33516 7580
rect 33556 7540 33577 7580
rect 33663 7540 33680 7580
rect 33720 7540 33729 7580
rect 33343 7517 33409 7540
rect 33495 7517 33577 7540
rect 33663 7517 33729 7540
rect 33343 7498 33729 7517
rect 48463 7603 48849 7622
rect 48463 7580 48529 7603
rect 48615 7580 48697 7603
rect 48783 7580 48849 7603
rect 48463 7540 48472 7580
rect 48512 7540 48529 7580
rect 48615 7540 48636 7580
rect 48676 7540 48697 7580
rect 48783 7540 48800 7580
rect 48840 7540 48849 7580
rect 48463 7517 48529 7540
rect 48615 7517 48697 7540
rect 48783 7517 48849 7540
rect 48463 7498 48849 7517
rect 63583 7603 63969 7622
rect 63583 7580 63649 7603
rect 63735 7580 63817 7603
rect 63903 7580 63969 7603
rect 63583 7540 63592 7580
rect 63632 7540 63649 7580
rect 63735 7540 63756 7580
rect 63796 7540 63817 7580
rect 63903 7540 63920 7580
rect 63960 7540 63969 7580
rect 63583 7517 63649 7540
rect 63735 7517 63817 7540
rect 63903 7517 63969 7540
rect 63583 7498 63969 7517
rect 78703 7603 79089 7622
rect 78703 7580 78769 7603
rect 78855 7580 78937 7603
rect 79023 7580 79089 7603
rect 78703 7540 78712 7580
rect 78752 7540 78769 7580
rect 78855 7540 78876 7580
rect 78916 7540 78937 7580
rect 79023 7540 79040 7580
rect 79080 7540 79089 7580
rect 78703 7517 78769 7540
rect 78855 7517 78937 7540
rect 79023 7517 79089 7540
rect 78703 7498 79089 7517
rect 93823 7603 94209 7622
rect 93823 7580 93889 7603
rect 93975 7580 94057 7603
rect 94143 7580 94209 7603
rect 93823 7540 93832 7580
rect 93872 7540 93889 7580
rect 93975 7540 93996 7580
rect 94036 7540 94057 7580
rect 94143 7540 94160 7580
rect 94200 7540 94209 7580
rect 93823 7517 93889 7540
rect 93975 7517 94057 7540
rect 94143 7517 94209 7540
rect 93823 7498 94209 7517
rect 4343 6847 4729 6866
rect 4343 6824 4409 6847
rect 4495 6824 4577 6847
rect 4663 6824 4729 6847
rect 4343 6784 4352 6824
rect 4392 6784 4409 6824
rect 4495 6784 4516 6824
rect 4556 6784 4577 6824
rect 4663 6784 4680 6824
rect 4720 6784 4729 6824
rect 4343 6761 4409 6784
rect 4495 6761 4577 6784
rect 4663 6761 4729 6784
rect 4343 6742 4729 6761
rect 19463 6847 19849 6866
rect 19463 6824 19529 6847
rect 19615 6824 19697 6847
rect 19783 6824 19849 6847
rect 19463 6784 19472 6824
rect 19512 6784 19529 6824
rect 19615 6784 19636 6824
rect 19676 6784 19697 6824
rect 19783 6784 19800 6824
rect 19840 6784 19849 6824
rect 19463 6761 19529 6784
rect 19615 6761 19697 6784
rect 19783 6761 19849 6784
rect 19463 6742 19849 6761
rect 34583 6847 34969 6866
rect 34583 6824 34649 6847
rect 34735 6824 34817 6847
rect 34903 6824 34969 6847
rect 34583 6784 34592 6824
rect 34632 6784 34649 6824
rect 34735 6784 34756 6824
rect 34796 6784 34817 6824
rect 34903 6784 34920 6824
rect 34960 6784 34969 6824
rect 34583 6761 34649 6784
rect 34735 6761 34817 6784
rect 34903 6761 34969 6784
rect 34583 6742 34969 6761
rect 49703 6847 50089 6866
rect 49703 6824 49769 6847
rect 49855 6824 49937 6847
rect 50023 6824 50089 6847
rect 49703 6784 49712 6824
rect 49752 6784 49769 6824
rect 49855 6784 49876 6824
rect 49916 6784 49937 6824
rect 50023 6784 50040 6824
rect 50080 6784 50089 6824
rect 49703 6761 49769 6784
rect 49855 6761 49937 6784
rect 50023 6761 50089 6784
rect 49703 6742 50089 6761
rect 64823 6847 65209 6866
rect 64823 6824 64889 6847
rect 64975 6824 65057 6847
rect 65143 6824 65209 6847
rect 64823 6784 64832 6824
rect 64872 6784 64889 6824
rect 64975 6784 64996 6824
rect 65036 6784 65057 6824
rect 65143 6784 65160 6824
rect 65200 6784 65209 6824
rect 64823 6761 64889 6784
rect 64975 6761 65057 6784
rect 65143 6761 65209 6784
rect 64823 6742 65209 6761
rect 79943 6847 80329 6866
rect 79943 6824 80009 6847
rect 80095 6824 80177 6847
rect 80263 6824 80329 6847
rect 79943 6784 79952 6824
rect 79992 6784 80009 6824
rect 80095 6784 80116 6824
rect 80156 6784 80177 6824
rect 80263 6784 80280 6824
rect 80320 6784 80329 6824
rect 79943 6761 80009 6784
rect 80095 6761 80177 6784
rect 80263 6761 80329 6784
rect 79943 6742 80329 6761
rect 95063 6847 95449 6866
rect 95063 6824 95129 6847
rect 95215 6824 95297 6847
rect 95383 6824 95449 6847
rect 95063 6784 95072 6824
rect 95112 6784 95129 6824
rect 95215 6784 95236 6824
rect 95276 6784 95297 6824
rect 95383 6784 95400 6824
rect 95440 6784 95449 6824
rect 95063 6761 95129 6784
rect 95215 6761 95297 6784
rect 95383 6761 95449 6784
rect 95063 6742 95449 6761
rect 3103 6091 3489 6110
rect 3103 6068 3169 6091
rect 3255 6068 3337 6091
rect 3423 6068 3489 6091
rect 3103 6028 3112 6068
rect 3152 6028 3169 6068
rect 3255 6028 3276 6068
rect 3316 6028 3337 6068
rect 3423 6028 3440 6068
rect 3480 6028 3489 6068
rect 3103 6005 3169 6028
rect 3255 6005 3337 6028
rect 3423 6005 3489 6028
rect 3103 5986 3489 6005
rect 18223 6091 18609 6110
rect 18223 6068 18289 6091
rect 18375 6068 18457 6091
rect 18543 6068 18609 6091
rect 18223 6028 18232 6068
rect 18272 6028 18289 6068
rect 18375 6028 18396 6068
rect 18436 6028 18457 6068
rect 18543 6028 18560 6068
rect 18600 6028 18609 6068
rect 18223 6005 18289 6028
rect 18375 6005 18457 6028
rect 18543 6005 18609 6028
rect 18223 5986 18609 6005
rect 33343 6091 33729 6110
rect 33343 6068 33409 6091
rect 33495 6068 33577 6091
rect 33663 6068 33729 6091
rect 33343 6028 33352 6068
rect 33392 6028 33409 6068
rect 33495 6028 33516 6068
rect 33556 6028 33577 6068
rect 33663 6028 33680 6068
rect 33720 6028 33729 6068
rect 33343 6005 33409 6028
rect 33495 6005 33577 6028
rect 33663 6005 33729 6028
rect 33343 5986 33729 6005
rect 48463 6091 48849 6110
rect 48463 6068 48529 6091
rect 48615 6068 48697 6091
rect 48783 6068 48849 6091
rect 48463 6028 48472 6068
rect 48512 6028 48529 6068
rect 48615 6028 48636 6068
rect 48676 6028 48697 6068
rect 48783 6028 48800 6068
rect 48840 6028 48849 6068
rect 48463 6005 48529 6028
rect 48615 6005 48697 6028
rect 48783 6005 48849 6028
rect 48463 5986 48849 6005
rect 63583 6091 63969 6110
rect 63583 6068 63649 6091
rect 63735 6068 63817 6091
rect 63903 6068 63969 6091
rect 63583 6028 63592 6068
rect 63632 6028 63649 6068
rect 63735 6028 63756 6068
rect 63796 6028 63817 6068
rect 63903 6028 63920 6068
rect 63960 6028 63969 6068
rect 63583 6005 63649 6028
rect 63735 6005 63817 6028
rect 63903 6005 63969 6028
rect 63583 5986 63969 6005
rect 78703 6091 79089 6110
rect 78703 6068 78769 6091
rect 78855 6068 78937 6091
rect 79023 6068 79089 6091
rect 78703 6028 78712 6068
rect 78752 6028 78769 6068
rect 78855 6028 78876 6068
rect 78916 6028 78937 6068
rect 79023 6028 79040 6068
rect 79080 6028 79089 6068
rect 78703 6005 78769 6028
rect 78855 6005 78937 6028
rect 79023 6005 79089 6028
rect 78703 5986 79089 6005
rect 93823 6091 94209 6110
rect 93823 6068 93889 6091
rect 93975 6068 94057 6091
rect 94143 6068 94209 6091
rect 93823 6028 93832 6068
rect 93872 6028 93889 6068
rect 93975 6028 93996 6068
rect 94036 6028 94057 6068
rect 94143 6028 94160 6068
rect 94200 6028 94209 6068
rect 93823 6005 93889 6028
rect 93975 6005 94057 6028
rect 94143 6005 94209 6028
rect 93823 5986 94209 6005
rect 4343 5335 4729 5354
rect 4343 5312 4409 5335
rect 4495 5312 4577 5335
rect 4663 5312 4729 5335
rect 4343 5272 4352 5312
rect 4392 5272 4409 5312
rect 4495 5272 4516 5312
rect 4556 5272 4577 5312
rect 4663 5272 4680 5312
rect 4720 5272 4729 5312
rect 4343 5249 4409 5272
rect 4495 5249 4577 5272
rect 4663 5249 4729 5272
rect 4343 5230 4729 5249
rect 19463 5335 19849 5354
rect 19463 5312 19529 5335
rect 19615 5312 19697 5335
rect 19783 5312 19849 5335
rect 19463 5272 19472 5312
rect 19512 5272 19529 5312
rect 19615 5272 19636 5312
rect 19676 5272 19697 5312
rect 19783 5272 19800 5312
rect 19840 5272 19849 5312
rect 19463 5249 19529 5272
rect 19615 5249 19697 5272
rect 19783 5249 19849 5272
rect 19463 5230 19849 5249
rect 34583 5335 34969 5354
rect 34583 5312 34649 5335
rect 34735 5312 34817 5335
rect 34903 5312 34969 5335
rect 34583 5272 34592 5312
rect 34632 5272 34649 5312
rect 34735 5272 34756 5312
rect 34796 5272 34817 5312
rect 34903 5272 34920 5312
rect 34960 5272 34969 5312
rect 34583 5249 34649 5272
rect 34735 5249 34817 5272
rect 34903 5249 34969 5272
rect 34583 5230 34969 5249
rect 49703 5335 50089 5354
rect 49703 5312 49769 5335
rect 49855 5312 49937 5335
rect 50023 5312 50089 5335
rect 49703 5272 49712 5312
rect 49752 5272 49769 5312
rect 49855 5272 49876 5312
rect 49916 5272 49937 5312
rect 50023 5272 50040 5312
rect 50080 5272 50089 5312
rect 49703 5249 49769 5272
rect 49855 5249 49937 5272
rect 50023 5249 50089 5272
rect 49703 5230 50089 5249
rect 64823 5335 65209 5354
rect 64823 5312 64889 5335
rect 64975 5312 65057 5335
rect 65143 5312 65209 5335
rect 64823 5272 64832 5312
rect 64872 5272 64889 5312
rect 64975 5272 64996 5312
rect 65036 5272 65057 5312
rect 65143 5272 65160 5312
rect 65200 5272 65209 5312
rect 64823 5249 64889 5272
rect 64975 5249 65057 5272
rect 65143 5249 65209 5272
rect 64823 5230 65209 5249
rect 79943 5335 80329 5354
rect 79943 5312 80009 5335
rect 80095 5312 80177 5335
rect 80263 5312 80329 5335
rect 79943 5272 79952 5312
rect 79992 5272 80009 5312
rect 80095 5272 80116 5312
rect 80156 5272 80177 5312
rect 80263 5272 80280 5312
rect 80320 5272 80329 5312
rect 79943 5249 80009 5272
rect 80095 5249 80177 5272
rect 80263 5249 80329 5272
rect 79943 5230 80329 5249
rect 95063 5335 95449 5354
rect 95063 5312 95129 5335
rect 95215 5312 95297 5335
rect 95383 5312 95449 5335
rect 95063 5272 95072 5312
rect 95112 5272 95129 5312
rect 95215 5272 95236 5312
rect 95276 5272 95297 5312
rect 95383 5272 95400 5312
rect 95440 5272 95449 5312
rect 95063 5249 95129 5272
rect 95215 5249 95297 5272
rect 95383 5249 95449 5272
rect 95063 5230 95449 5249
rect 3103 4579 3489 4598
rect 3103 4556 3169 4579
rect 3255 4556 3337 4579
rect 3423 4556 3489 4579
rect 3103 4516 3112 4556
rect 3152 4516 3169 4556
rect 3255 4516 3276 4556
rect 3316 4516 3337 4556
rect 3423 4516 3440 4556
rect 3480 4516 3489 4556
rect 3103 4493 3169 4516
rect 3255 4493 3337 4516
rect 3423 4493 3489 4516
rect 3103 4474 3489 4493
rect 18223 4579 18609 4598
rect 18223 4556 18289 4579
rect 18375 4556 18457 4579
rect 18543 4556 18609 4579
rect 18223 4516 18232 4556
rect 18272 4516 18289 4556
rect 18375 4516 18396 4556
rect 18436 4516 18457 4556
rect 18543 4516 18560 4556
rect 18600 4516 18609 4556
rect 18223 4493 18289 4516
rect 18375 4493 18457 4516
rect 18543 4493 18609 4516
rect 18223 4474 18609 4493
rect 33343 4579 33729 4598
rect 33343 4556 33409 4579
rect 33495 4556 33577 4579
rect 33663 4556 33729 4579
rect 33343 4516 33352 4556
rect 33392 4516 33409 4556
rect 33495 4516 33516 4556
rect 33556 4516 33577 4556
rect 33663 4516 33680 4556
rect 33720 4516 33729 4556
rect 33343 4493 33409 4516
rect 33495 4493 33577 4516
rect 33663 4493 33729 4516
rect 33343 4474 33729 4493
rect 48463 4579 48849 4598
rect 48463 4556 48529 4579
rect 48615 4556 48697 4579
rect 48783 4556 48849 4579
rect 48463 4516 48472 4556
rect 48512 4516 48529 4556
rect 48615 4516 48636 4556
rect 48676 4516 48697 4556
rect 48783 4516 48800 4556
rect 48840 4516 48849 4556
rect 48463 4493 48529 4516
rect 48615 4493 48697 4516
rect 48783 4493 48849 4516
rect 48463 4474 48849 4493
rect 63583 4579 63969 4598
rect 63583 4556 63649 4579
rect 63735 4556 63817 4579
rect 63903 4556 63969 4579
rect 63583 4516 63592 4556
rect 63632 4516 63649 4556
rect 63735 4516 63756 4556
rect 63796 4516 63817 4556
rect 63903 4516 63920 4556
rect 63960 4516 63969 4556
rect 63583 4493 63649 4516
rect 63735 4493 63817 4516
rect 63903 4493 63969 4516
rect 63583 4474 63969 4493
rect 78703 4579 79089 4598
rect 78703 4556 78769 4579
rect 78855 4556 78937 4579
rect 79023 4556 79089 4579
rect 78703 4516 78712 4556
rect 78752 4516 78769 4556
rect 78855 4516 78876 4556
rect 78916 4516 78937 4556
rect 79023 4516 79040 4556
rect 79080 4516 79089 4556
rect 78703 4493 78769 4516
rect 78855 4493 78937 4516
rect 79023 4493 79089 4516
rect 78703 4474 79089 4493
rect 93823 4579 94209 4598
rect 93823 4556 93889 4579
rect 93975 4556 94057 4579
rect 94143 4556 94209 4579
rect 93823 4516 93832 4556
rect 93872 4516 93889 4556
rect 93975 4516 93996 4556
rect 94036 4516 94057 4556
rect 94143 4516 94160 4556
rect 94200 4516 94209 4556
rect 93823 4493 93889 4516
rect 93975 4493 94057 4516
rect 94143 4493 94209 4516
rect 93823 4474 94209 4493
rect 4343 3823 4729 3842
rect 4343 3800 4409 3823
rect 4495 3800 4577 3823
rect 4663 3800 4729 3823
rect 4343 3760 4352 3800
rect 4392 3760 4409 3800
rect 4495 3760 4516 3800
rect 4556 3760 4577 3800
rect 4663 3760 4680 3800
rect 4720 3760 4729 3800
rect 4343 3737 4409 3760
rect 4495 3737 4577 3760
rect 4663 3737 4729 3760
rect 4343 3718 4729 3737
rect 19463 3823 19849 3842
rect 19463 3800 19529 3823
rect 19615 3800 19697 3823
rect 19783 3800 19849 3823
rect 19463 3760 19472 3800
rect 19512 3760 19529 3800
rect 19615 3760 19636 3800
rect 19676 3760 19697 3800
rect 19783 3760 19800 3800
rect 19840 3760 19849 3800
rect 19463 3737 19529 3760
rect 19615 3737 19697 3760
rect 19783 3737 19849 3760
rect 19463 3718 19849 3737
rect 34583 3823 34969 3842
rect 34583 3800 34649 3823
rect 34735 3800 34817 3823
rect 34903 3800 34969 3823
rect 34583 3760 34592 3800
rect 34632 3760 34649 3800
rect 34735 3760 34756 3800
rect 34796 3760 34817 3800
rect 34903 3760 34920 3800
rect 34960 3760 34969 3800
rect 34583 3737 34649 3760
rect 34735 3737 34817 3760
rect 34903 3737 34969 3760
rect 34583 3718 34969 3737
rect 49703 3823 50089 3842
rect 49703 3800 49769 3823
rect 49855 3800 49937 3823
rect 50023 3800 50089 3823
rect 49703 3760 49712 3800
rect 49752 3760 49769 3800
rect 49855 3760 49876 3800
rect 49916 3760 49937 3800
rect 50023 3760 50040 3800
rect 50080 3760 50089 3800
rect 49703 3737 49769 3760
rect 49855 3737 49937 3760
rect 50023 3737 50089 3760
rect 49703 3718 50089 3737
rect 64823 3823 65209 3842
rect 64823 3800 64889 3823
rect 64975 3800 65057 3823
rect 65143 3800 65209 3823
rect 64823 3760 64832 3800
rect 64872 3760 64889 3800
rect 64975 3760 64996 3800
rect 65036 3760 65057 3800
rect 65143 3760 65160 3800
rect 65200 3760 65209 3800
rect 64823 3737 64889 3760
rect 64975 3737 65057 3760
rect 65143 3737 65209 3760
rect 64823 3718 65209 3737
rect 79943 3823 80329 3842
rect 79943 3800 80009 3823
rect 80095 3800 80177 3823
rect 80263 3800 80329 3823
rect 79943 3760 79952 3800
rect 79992 3760 80009 3800
rect 80095 3760 80116 3800
rect 80156 3760 80177 3800
rect 80263 3760 80280 3800
rect 80320 3760 80329 3800
rect 79943 3737 80009 3760
rect 80095 3737 80177 3760
rect 80263 3737 80329 3760
rect 79943 3718 80329 3737
rect 95063 3823 95449 3842
rect 95063 3800 95129 3823
rect 95215 3800 95297 3823
rect 95383 3800 95449 3823
rect 95063 3760 95072 3800
rect 95112 3760 95129 3800
rect 95215 3760 95236 3800
rect 95276 3760 95297 3800
rect 95383 3760 95400 3800
rect 95440 3760 95449 3800
rect 95063 3737 95129 3760
rect 95215 3737 95297 3760
rect 95383 3737 95449 3760
rect 95063 3718 95449 3737
rect 3103 3067 3489 3086
rect 3103 3044 3169 3067
rect 3255 3044 3337 3067
rect 3423 3044 3489 3067
rect 3103 3004 3112 3044
rect 3152 3004 3169 3044
rect 3255 3004 3276 3044
rect 3316 3004 3337 3044
rect 3423 3004 3440 3044
rect 3480 3004 3489 3044
rect 3103 2981 3169 3004
rect 3255 2981 3337 3004
rect 3423 2981 3489 3004
rect 3103 2962 3489 2981
rect 18223 3067 18609 3086
rect 18223 3044 18289 3067
rect 18375 3044 18457 3067
rect 18543 3044 18609 3067
rect 18223 3004 18232 3044
rect 18272 3004 18289 3044
rect 18375 3004 18396 3044
rect 18436 3004 18457 3044
rect 18543 3004 18560 3044
rect 18600 3004 18609 3044
rect 18223 2981 18289 3004
rect 18375 2981 18457 3004
rect 18543 2981 18609 3004
rect 18223 2962 18609 2981
rect 33343 3067 33729 3086
rect 33343 3044 33409 3067
rect 33495 3044 33577 3067
rect 33663 3044 33729 3067
rect 33343 3004 33352 3044
rect 33392 3004 33409 3044
rect 33495 3004 33516 3044
rect 33556 3004 33577 3044
rect 33663 3004 33680 3044
rect 33720 3004 33729 3044
rect 33343 2981 33409 3004
rect 33495 2981 33577 3004
rect 33663 2981 33729 3004
rect 33343 2962 33729 2981
rect 48463 3067 48849 3086
rect 48463 3044 48529 3067
rect 48615 3044 48697 3067
rect 48783 3044 48849 3067
rect 48463 3004 48472 3044
rect 48512 3004 48529 3044
rect 48615 3004 48636 3044
rect 48676 3004 48697 3044
rect 48783 3004 48800 3044
rect 48840 3004 48849 3044
rect 48463 2981 48529 3004
rect 48615 2981 48697 3004
rect 48783 2981 48849 3004
rect 48463 2962 48849 2981
rect 63583 3067 63969 3086
rect 63583 3044 63649 3067
rect 63735 3044 63817 3067
rect 63903 3044 63969 3067
rect 63583 3004 63592 3044
rect 63632 3004 63649 3044
rect 63735 3004 63756 3044
rect 63796 3004 63817 3044
rect 63903 3004 63920 3044
rect 63960 3004 63969 3044
rect 63583 2981 63649 3004
rect 63735 2981 63817 3004
rect 63903 2981 63969 3004
rect 63583 2962 63969 2981
rect 78703 3067 79089 3086
rect 78703 3044 78769 3067
rect 78855 3044 78937 3067
rect 79023 3044 79089 3067
rect 78703 3004 78712 3044
rect 78752 3004 78769 3044
rect 78855 3004 78876 3044
rect 78916 3004 78937 3044
rect 79023 3004 79040 3044
rect 79080 3004 79089 3044
rect 78703 2981 78769 3004
rect 78855 2981 78937 3004
rect 79023 2981 79089 3004
rect 78703 2962 79089 2981
rect 93823 3067 94209 3086
rect 93823 3044 93889 3067
rect 93975 3044 94057 3067
rect 94143 3044 94209 3067
rect 93823 3004 93832 3044
rect 93872 3004 93889 3044
rect 93975 3004 93996 3044
rect 94036 3004 94057 3044
rect 94143 3004 94160 3044
rect 94200 3004 94209 3044
rect 93823 2981 93889 3004
rect 93975 2981 94057 3004
rect 94143 2981 94209 3004
rect 93823 2962 94209 2981
rect 4343 2311 4729 2330
rect 4343 2288 4409 2311
rect 4495 2288 4577 2311
rect 4663 2288 4729 2311
rect 4343 2248 4352 2288
rect 4392 2248 4409 2288
rect 4495 2248 4516 2288
rect 4556 2248 4577 2288
rect 4663 2248 4680 2288
rect 4720 2248 4729 2288
rect 4343 2225 4409 2248
rect 4495 2225 4577 2248
rect 4663 2225 4729 2248
rect 4343 2206 4729 2225
rect 19463 2311 19849 2330
rect 19463 2288 19529 2311
rect 19615 2288 19697 2311
rect 19783 2288 19849 2311
rect 19463 2248 19472 2288
rect 19512 2248 19529 2288
rect 19615 2248 19636 2288
rect 19676 2248 19697 2288
rect 19783 2248 19800 2288
rect 19840 2248 19849 2288
rect 19463 2225 19529 2248
rect 19615 2225 19697 2248
rect 19783 2225 19849 2248
rect 19463 2206 19849 2225
rect 34583 2311 34969 2330
rect 34583 2288 34649 2311
rect 34735 2288 34817 2311
rect 34903 2288 34969 2311
rect 34583 2248 34592 2288
rect 34632 2248 34649 2288
rect 34735 2248 34756 2288
rect 34796 2248 34817 2288
rect 34903 2248 34920 2288
rect 34960 2248 34969 2288
rect 34583 2225 34649 2248
rect 34735 2225 34817 2248
rect 34903 2225 34969 2248
rect 34583 2206 34969 2225
rect 49703 2311 50089 2330
rect 49703 2288 49769 2311
rect 49855 2288 49937 2311
rect 50023 2288 50089 2311
rect 49703 2248 49712 2288
rect 49752 2248 49769 2288
rect 49855 2248 49876 2288
rect 49916 2248 49937 2288
rect 50023 2248 50040 2288
rect 50080 2248 50089 2288
rect 49703 2225 49769 2248
rect 49855 2225 49937 2248
rect 50023 2225 50089 2248
rect 49703 2206 50089 2225
rect 64823 2311 65209 2330
rect 64823 2288 64889 2311
rect 64975 2288 65057 2311
rect 65143 2288 65209 2311
rect 64823 2248 64832 2288
rect 64872 2248 64889 2288
rect 64975 2248 64996 2288
rect 65036 2248 65057 2288
rect 65143 2248 65160 2288
rect 65200 2248 65209 2288
rect 64823 2225 64889 2248
rect 64975 2225 65057 2248
rect 65143 2225 65209 2248
rect 64823 2206 65209 2225
rect 79943 2311 80329 2330
rect 79943 2288 80009 2311
rect 80095 2288 80177 2311
rect 80263 2288 80329 2311
rect 79943 2248 79952 2288
rect 79992 2248 80009 2288
rect 80095 2248 80116 2288
rect 80156 2248 80177 2288
rect 80263 2248 80280 2288
rect 80320 2248 80329 2288
rect 79943 2225 80009 2248
rect 80095 2225 80177 2248
rect 80263 2225 80329 2248
rect 79943 2206 80329 2225
rect 95063 2311 95449 2330
rect 95063 2288 95129 2311
rect 95215 2288 95297 2311
rect 95383 2288 95449 2311
rect 95063 2248 95072 2288
rect 95112 2248 95129 2288
rect 95215 2248 95236 2288
rect 95276 2248 95297 2288
rect 95383 2248 95400 2288
rect 95440 2248 95449 2288
rect 95063 2225 95129 2248
rect 95215 2225 95297 2248
rect 95383 2225 95449 2248
rect 95063 2206 95449 2225
rect 3103 1555 3489 1574
rect 3103 1532 3169 1555
rect 3255 1532 3337 1555
rect 3423 1532 3489 1555
rect 3103 1492 3112 1532
rect 3152 1492 3169 1532
rect 3255 1492 3276 1532
rect 3316 1492 3337 1532
rect 3423 1492 3440 1532
rect 3480 1492 3489 1532
rect 3103 1469 3169 1492
rect 3255 1469 3337 1492
rect 3423 1469 3489 1492
rect 3103 1450 3489 1469
rect 18223 1555 18609 1574
rect 18223 1532 18289 1555
rect 18375 1532 18457 1555
rect 18543 1532 18609 1555
rect 18223 1492 18232 1532
rect 18272 1492 18289 1532
rect 18375 1492 18396 1532
rect 18436 1492 18457 1532
rect 18543 1492 18560 1532
rect 18600 1492 18609 1532
rect 18223 1469 18289 1492
rect 18375 1469 18457 1492
rect 18543 1469 18609 1492
rect 18223 1450 18609 1469
rect 33343 1555 33729 1574
rect 33343 1532 33409 1555
rect 33495 1532 33577 1555
rect 33663 1532 33729 1555
rect 33343 1492 33352 1532
rect 33392 1492 33409 1532
rect 33495 1492 33516 1532
rect 33556 1492 33577 1532
rect 33663 1492 33680 1532
rect 33720 1492 33729 1532
rect 33343 1469 33409 1492
rect 33495 1469 33577 1492
rect 33663 1469 33729 1492
rect 33343 1450 33729 1469
rect 48463 1555 48849 1574
rect 48463 1532 48529 1555
rect 48615 1532 48697 1555
rect 48783 1532 48849 1555
rect 48463 1492 48472 1532
rect 48512 1492 48529 1532
rect 48615 1492 48636 1532
rect 48676 1492 48697 1532
rect 48783 1492 48800 1532
rect 48840 1492 48849 1532
rect 48463 1469 48529 1492
rect 48615 1469 48697 1492
rect 48783 1469 48849 1492
rect 48463 1450 48849 1469
rect 63583 1555 63969 1574
rect 63583 1532 63649 1555
rect 63735 1532 63817 1555
rect 63903 1532 63969 1555
rect 63583 1492 63592 1532
rect 63632 1492 63649 1532
rect 63735 1492 63756 1532
rect 63796 1492 63817 1532
rect 63903 1492 63920 1532
rect 63960 1492 63969 1532
rect 63583 1469 63649 1492
rect 63735 1469 63817 1492
rect 63903 1469 63969 1492
rect 63583 1450 63969 1469
rect 78703 1555 79089 1574
rect 78703 1532 78769 1555
rect 78855 1532 78937 1555
rect 79023 1532 79089 1555
rect 78703 1492 78712 1532
rect 78752 1492 78769 1532
rect 78855 1492 78876 1532
rect 78916 1492 78937 1532
rect 79023 1492 79040 1532
rect 79080 1492 79089 1532
rect 78703 1469 78769 1492
rect 78855 1469 78937 1492
rect 79023 1469 79089 1492
rect 78703 1450 79089 1469
rect 93823 1555 94209 1574
rect 93823 1532 93889 1555
rect 93975 1532 94057 1555
rect 94143 1532 94209 1555
rect 93823 1492 93832 1532
rect 93872 1492 93889 1532
rect 93975 1492 93996 1532
rect 94036 1492 94057 1532
rect 94143 1492 94160 1532
rect 94200 1492 94209 1532
rect 93823 1469 93889 1492
rect 93975 1469 94057 1492
rect 94143 1469 94209 1492
rect 93823 1450 94209 1469
rect 4343 799 4729 818
rect 4343 776 4409 799
rect 4495 776 4577 799
rect 4663 776 4729 799
rect 4343 736 4352 776
rect 4392 736 4409 776
rect 4495 736 4516 776
rect 4556 736 4577 776
rect 4663 736 4680 776
rect 4720 736 4729 776
rect 4343 713 4409 736
rect 4495 713 4577 736
rect 4663 713 4729 736
rect 4343 694 4729 713
rect 19463 799 19849 818
rect 19463 776 19529 799
rect 19615 776 19697 799
rect 19783 776 19849 799
rect 19463 736 19472 776
rect 19512 736 19529 776
rect 19615 736 19636 776
rect 19676 736 19697 776
rect 19783 736 19800 776
rect 19840 736 19849 776
rect 19463 713 19529 736
rect 19615 713 19697 736
rect 19783 713 19849 736
rect 19463 694 19849 713
rect 34583 799 34969 818
rect 34583 776 34649 799
rect 34735 776 34817 799
rect 34903 776 34969 799
rect 34583 736 34592 776
rect 34632 736 34649 776
rect 34735 736 34756 776
rect 34796 736 34817 776
rect 34903 736 34920 776
rect 34960 736 34969 776
rect 34583 713 34649 736
rect 34735 713 34817 736
rect 34903 713 34969 736
rect 34583 694 34969 713
rect 49703 799 50089 818
rect 49703 776 49769 799
rect 49855 776 49937 799
rect 50023 776 50089 799
rect 49703 736 49712 776
rect 49752 736 49769 776
rect 49855 736 49876 776
rect 49916 736 49937 776
rect 50023 736 50040 776
rect 50080 736 50089 776
rect 49703 713 49769 736
rect 49855 713 49937 736
rect 50023 713 50089 736
rect 49703 694 50089 713
rect 64823 799 65209 818
rect 64823 776 64889 799
rect 64975 776 65057 799
rect 65143 776 65209 799
rect 64823 736 64832 776
rect 64872 736 64889 776
rect 64975 736 64996 776
rect 65036 736 65057 776
rect 65143 736 65160 776
rect 65200 736 65209 776
rect 64823 713 64889 736
rect 64975 713 65057 736
rect 65143 713 65209 736
rect 64823 694 65209 713
rect 79943 799 80329 818
rect 79943 776 80009 799
rect 80095 776 80177 799
rect 80263 776 80329 799
rect 79943 736 79952 776
rect 79992 736 80009 776
rect 80095 736 80116 776
rect 80156 736 80177 776
rect 80263 736 80280 776
rect 80320 736 80329 776
rect 79943 713 80009 736
rect 80095 713 80177 736
rect 80263 713 80329 736
rect 79943 694 80329 713
rect 95063 799 95449 818
rect 95063 776 95129 799
rect 95215 776 95297 799
rect 95383 776 95449 799
rect 95063 736 95072 776
rect 95112 736 95129 776
rect 95215 736 95236 776
rect 95276 736 95297 776
rect 95383 736 95400 776
rect 95440 736 95449 776
rect 95063 713 95129 736
rect 95215 713 95297 736
rect 95383 713 95449 736
rect 95063 694 95449 713
<< via5 >>
rect 3169 81668 3255 81691
rect 3337 81668 3423 81691
rect 3169 81628 3194 81668
rect 3194 81628 3234 81668
rect 3234 81628 3255 81668
rect 3337 81628 3358 81668
rect 3358 81628 3398 81668
rect 3398 81628 3423 81668
rect 3169 81605 3255 81628
rect 3337 81605 3423 81628
rect 18289 81668 18375 81691
rect 18457 81668 18543 81691
rect 18289 81628 18314 81668
rect 18314 81628 18354 81668
rect 18354 81628 18375 81668
rect 18457 81628 18478 81668
rect 18478 81628 18518 81668
rect 18518 81628 18543 81668
rect 18289 81605 18375 81628
rect 18457 81605 18543 81628
rect 33409 81668 33495 81691
rect 33577 81668 33663 81691
rect 33409 81628 33434 81668
rect 33434 81628 33474 81668
rect 33474 81628 33495 81668
rect 33577 81628 33598 81668
rect 33598 81628 33638 81668
rect 33638 81628 33663 81668
rect 33409 81605 33495 81628
rect 33577 81605 33663 81628
rect 48529 81668 48615 81691
rect 48697 81668 48783 81691
rect 48529 81628 48554 81668
rect 48554 81628 48594 81668
rect 48594 81628 48615 81668
rect 48697 81628 48718 81668
rect 48718 81628 48758 81668
rect 48758 81628 48783 81668
rect 48529 81605 48615 81628
rect 48697 81605 48783 81628
rect 63649 81668 63735 81691
rect 63817 81668 63903 81691
rect 63649 81628 63674 81668
rect 63674 81628 63714 81668
rect 63714 81628 63735 81668
rect 63817 81628 63838 81668
rect 63838 81628 63878 81668
rect 63878 81628 63903 81668
rect 63649 81605 63735 81628
rect 63817 81605 63903 81628
rect 78769 81668 78855 81691
rect 78937 81668 79023 81691
rect 78769 81628 78794 81668
rect 78794 81628 78834 81668
rect 78834 81628 78855 81668
rect 78937 81628 78958 81668
rect 78958 81628 78998 81668
rect 78998 81628 79023 81668
rect 78769 81605 78855 81628
rect 78937 81605 79023 81628
rect 93889 81668 93975 81691
rect 94057 81668 94143 81691
rect 93889 81628 93914 81668
rect 93914 81628 93954 81668
rect 93954 81628 93975 81668
rect 94057 81628 94078 81668
rect 94078 81628 94118 81668
rect 94118 81628 94143 81668
rect 93889 81605 93975 81628
rect 94057 81605 94143 81628
rect 4409 80912 4495 80935
rect 4577 80912 4663 80935
rect 4409 80872 4434 80912
rect 4434 80872 4474 80912
rect 4474 80872 4495 80912
rect 4577 80872 4598 80912
rect 4598 80872 4638 80912
rect 4638 80872 4663 80912
rect 4409 80849 4495 80872
rect 4577 80849 4663 80872
rect 19529 80912 19615 80935
rect 19697 80912 19783 80935
rect 19529 80872 19554 80912
rect 19554 80872 19594 80912
rect 19594 80872 19615 80912
rect 19697 80872 19718 80912
rect 19718 80872 19758 80912
rect 19758 80872 19783 80912
rect 19529 80849 19615 80872
rect 19697 80849 19783 80872
rect 34649 80912 34735 80935
rect 34817 80912 34903 80935
rect 34649 80872 34674 80912
rect 34674 80872 34714 80912
rect 34714 80872 34735 80912
rect 34817 80872 34838 80912
rect 34838 80872 34878 80912
rect 34878 80872 34903 80912
rect 34649 80849 34735 80872
rect 34817 80849 34903 80872
rect 49769 80912 49855 80935
rect 49937 80912 50023 80935
rect 49769 80872 49794 80912
rect 49794 80872 49834 80912
rect 49834 80872 49855 80912
rect 49937 80872 49958 80912
rect 49958 80872 49998 80912
rect 49998 80872 50023 80912
rect 49769 80849 49855 80872
rect 49937 80849 50023 80872
rect 64889 80912 64975 80935
rect 65057 80912 65143 80935
rect 64889 80872 64914 80912
rect 64914 80872 64954 80912
rect 64954 80872 64975 80912
rect 65057 80872 65078 80912
rect 65078 80872 65118 80912
rect 65118 80872 65143 80912
rect 64889 80849 64975 80872
rect 65057 80849 65143 80872
rect 80009 80912 80095 80935
rect 80177 80912 80263 80935
rect 80009 80872 80034 80912
rect 80034 80872 80074 80912
rect 80074 80872 80095 80912
rect 80177 80872 80198 80912
rect 80198 80872 80238 80912
rect 80238 80872 80263 80912
rect 80009 80849 80095 80872
rect 80177 80849 80263 80872
rect 95129 80912 95215 80935
rect 95297 80912 95383 80935
rect 95129 80872 95154 80912
rect 95154 80872 95194 80912
rect 95194 80872 95215 80912
rect 95297 80872 95318 80912
rect 95318 80872 95358 80912
rect 95358 80872 95383 80912
rect 95129 80849 95215 80872
rect 95297 80849 95383 80872
rect 3169 80156 3255 80179
rect 3337 80156 3423 80179
rect 3169 80116 3194 80156
rect 3194 80116 3234 80156
rect 3234 80116 3255 80156
rect 3337 80116 3358 80156
rect 3358 80116 3398 80156
rect 3398 80116 3423 80156
rect 3169 80093 3255 80116
rect 3337 80093 3423 80116
rect 18289 80156 18375 80179
rect 18457 80156 18543 80179
rect 18289 80116 18314 80156
rect 18314 80116 18354 80156
rect 18354 80116 18375 80156
rect 18457 80116 18478 80156
rect 18478 80116 18518 80156
rect 18518 80116 18543 80156
rect 18289 80093 18375 80116
rect 18457 80093 18543 80116
rect 33409 80156 33495 80179
rect 33577 80156 33663 80179
rect 33409 80116 33434 80156
rect 33434 80116 33474 80156
rect 33474 80116 33495 80156
rect 33577 80116 33598 80156
rect 33598 80116 33638 80156
rect 33638 80116 33663 80156
rect 33409 80093 33495 80116
rect 33577 80093 33663 80116
rect 48529 80156 48615 80179
rect 48697 80156 48783 80179
rect 48529 80116 48554 80156
rect 48554 80116 48594 80156
rect 48594 80116 48615 80156
rect 48697 80116 48718 80156
rect 48718 80116 48758 80156
rect 48758 80116 48783 80156
rect 48529 80093 48615 80116
rect 48697 80093 48783 80116
rect 63649 80156 63735 80179
rect 63817 80156 63903 80179
rect 63649 80116 63674 80156
rect 63674 80116 63714 80156
rect 63714 80116 63735 80156
rect 63817 80116 63838 80156
rect 63838 80116 63878 80156
rect 63878 80116 63903 80156
rect 63649 80093 63735 80116
rect 63817 80093 63903 80116
rect 78769 80156 78855 80179
rect 78937 80156 79023 80179
rect 78769 80116 78794 80156
rect 78794 80116 78834 80156
rect 78834 80116 78855 80156
rect 78937 80116 78958 80156
rect 78958 80116 78998 80156
rect 78998 80116 79023 80156
rect 78769 80093 78855 80116
rect 78937 80093 79023 80116
rect 93889 80156 93975 80179
rect 94057 80156 94143 80179
rect 93889 80116 93914 80156
rect 93914 80116 93954 80156
rect 93954 80116 93975 80156
rect 94057 80116 94078 80156
rect 94078 80116 94118 80156
rect 94118 80116 94143 80156
rect 93889 80093 93975 80116
rect 94057 80093 94143 80116
rect 4409 79400 4495 79423
rect 4577 79400 4663 79423
rect 4409 79360 4434 79400
rect 4434 79360 4474 79400
rect 4474 79360 4495 79400
rect 4577 79360 4598 79400
rect 4598 79360 4638 79400
rect 4638 79360 4663 79400
rect 4409 79337 4495 79360
rect 4577 79337 4663 79360
rect 19529 79400 19615 79423
rect 19697 79400 19783 79423
rect 19529 79360 19554 79400
rect 19554 79360 19594 79400
rect 19594 79360 19615 79400
rect 19697 79360 19718 79400
rect 19718 79360 19758 79400
rect 19758 79360 19783 79400
rect 19529 79337 19615 79360
rect 19697 79337 19783 79360
rect 34649 79400 34735 79423
rect 34817 79400 34903 79423
rect 34649 79360 34674 79400
rect 34674 79360 34714 79400
rect 34714 79360 34735 79400
rect 34817 79360 34838 79400
rect 34838 79360 34878 79400
rect 34878 79360 34903 79400
rect 34649 79337 34735 79360
rect 34817 79337 34903 79360
rect 49769 79400 49855 79423
rect 49937 79400 50023 79423
rect 49769 79360 49794 79400
rect 49794 79360 49834 79400
rect 49834 79360 49855 79400
rect 49937 79360 49958 79400
rect 49958 79360 49998 79400
rect 49998 79360 50023 79400
rect 49769 79337 49855 79360
rect 49937 79337 50023 79360
rect 64889 79400 64975 79423
rect 65057 79400 65143 79423
rect 64889 79360 64914 79400
rect 64914 79360 64954 79400
rect 64954 79360 64975 79400
rect 65057 79360 65078 79400
rect 65078 79360 65118 79400
rect 65118 79360 65143 79400
rect 64889 79337 64975 79360
rect 65057 79337 65143 79360
rect 80009 79400 80095 79423
rect 80177 79400 80263 79423
rect 80009 79360 80034 79400
rect 80034 79360 80074 79400
rect 80074 79360 80095 79400
rect 80177 79360 80198 79400
rect 80198 79360 80238 79400
rect 80238 79360 80263 79400
rect 80009 79337 80095 79360
rect 80177 79337 80263 79360
rect 95129 79400 95215 79423
rect 95297 79400 95383 79423
rect 95129 79360 95154 79400
rect 95154 79360 95194 79400
rect 95194 79360 95215 79400
rect 95297 79360 95318 79400
rect 95318 79360 95358 79400
rect 95358 79360 95383 79400
rect 95129 79337 95215 79360
rect 95297 79337 95383 79360
rect 3169 78644 3255 78667
rect 3337 78644 3423 78667
rect 3169 78604 3194 78644
rect 3194 78604 3234 78644
rect 3234 78604 3255 78644
rect 3337 78604 3358 78644
rect 3358 78604 3398 78644
rect 3398 78604 3423 78644
rect 3169 78581 3255 78604
rect 3337 78581 3423 78604
rect 18289 78644 18375 78667
rect 18457 78644 18543 78667
rect 18289 78604 18314 78644
rect 18314 78604 18354 78644
rect 18354 78604 18375 78644
rect 18457 78604 18478 78644
rect 18478 78604 18518 78644
rect 18518 78604 18543 78644
rect 18289 78581 18375 78604
rect 18457 78581 18543 78604
rect 33409 78644 33495 78667
rect 33577 78644 33663 78667
rect 33409 78604 33434 78644
rect 33434 78604 33474 78644
rect 33474 78604 33495 78644
rect 33577 78604 33598 78644
rect 33598 78604 33638 78644
rect 33638 78604 33663 78644
rect 33409 78581 33495 78604
rect 33577 78581 33663 78604
rect 48529 78644 48615 78667
rect 48697 78644 48783 78667
rect 48529 78604 48554 78644
rect 48554 78604 48594 78644
rect 48594 78604 48615 78644
rect 48697 78604 48718 78644
rect 48718 78604 48758 78644
rect 48758 78604 48783 78644
rect 48529 78581 48615 78604
rect 48697 78581 48783 78604
rect 63649 78644 63735 78667
rect 63817 78644 63903 78667
rect 63649 78604 63674 78644
rect 63674 78604 63714 78644
rect 63714 78604 63735 78644
rect 63817 78604 63838 78644
rect 63838 78604 63878 78644
rect 63878 78604 63903 78644
rect 63649 78581 63735 78604
rect 63817 78581 63903 78604
rect 78769 78644 78855 78667
rect 78937 78644 79023 78667
rect 78769 78604 78794 78644
rect 78794 78604 78834 78644
rect 78834 78604 78855 78644
rect 78937 78604 78958 78644
rect 78958 78604 78998 78644
rect 78998 78604 79023 78644
rect 78769 78581 78855 78604
rect 78937 78581 79023 78604
rect 93889 78644 93975 78667
rect 94057 78644 94143 78667
rect 93889 78604 93914 78644
rect 93914 78604 93954 78644
rect 93954 78604 93975 78644
rect 94057 78604 94078 78644
rect 94078 78604 94118 78644
rect 94118 78604 94143 78644
rect 93889 78581 93975 78604
rect 94057 78581 94143 78604
rect 4409 77888 4495 77911
rect 4577 77888 4663 77911
rect 4409 77848 4434 77888
rect 4434 77848 4474 77888
rect 4474 77848 4495 77888
rect 4577 77848 4598 77888
rect 4598 77848 4638 77888
rect 4638 77848 4663 77888
rect 4409 77825 4495 77848
rect 4577 77825 4663 77848
rect 19529 77888 19615 77911
rect 19697 77888 19783 77911
rect 19529 77848 19554 77888
rect 19554 77848 19594 77888
rect 19594 77848 19615 77888
rect 19697 77848 19718 77888
rect 19718 77848 19758 77888
rect 19758 77848 19783 77888
rect 19529 77825 19615 77848
rect 19697 77825 19783 77848
rect 34649 77888 34735 77911
rect 34817 77888 34903 77911
rect 34649 77848 34674 77888
rect 34674 77848 34714 77888
rect 34714 77848 34735 77888
rect 34817 77848 34838 77888
rect 34838 77848 34878 77888
rect 34878 77848 34903 77888
rect 34649 77825 34735 77848
rect 34817 77825 34903 77848
rect 49769 77888 49855 77911
rect 49937 77888 50023 77911
rect 49769 77848 49794 77888
rect 49794 77848 49834 77888
rect 49834 77848 49855 77888
rect 49937 77848 49958 77888
rect 49958 77848 49998 77888
rect 49998 77848 50023 77888
rect 49769 77825 49855 77848
rect 49937 77825 50023 77848
rect 64889 77888 64975 77911
rect 65057 77888 65143 77911
rect 64889 77848 64914 77888
rect 64914 77848 64954 77888
rect 64954 77848 64975 77888
rect 65057 77848 65078 77888
rect 65078 77848 65118 77888
rect 65118 77848 65143 77888
rect 64889 77825 64975 77848
rect 65057 77825 65143 77848
rect 80009 77888 80095 77911
rect 80177 77888 80263 77911
rect 80009 77848 80034 77888
rect 80034 77848 80074 77888
rect 80074 77848 80095 77888
rect 80177 77848 80198 77888
rect 80198 77848 80238 77888
rect 80238 77848 80263 77888
rect 80009 77825 80095 77848
rect 80177 77825 80263 77848
rect 95129 77888 95215 77911
rect 95297 77888 95383 77911
rect 95129 77848 95154 77888
rect 95154 77848 95194 77888
rect 95194 77848 95215 77888
rect 95297 77848 95318 77888
rect 95318 77848 95358 77888
rect 95358 77848 95383 77888
rect 95129 77825 95215 77848
rect 95297 77825 95383 77848
rect 3169 77132 3255 77155
rect 3337 77132 3423 77155
rect 3169 77092 3194 77132
rect 3194 77092 3234 77132
rect 3234 77092 3255 77132
rect 3337 77092 3358 77132
rect 3358 77092 3398 77132
rect 3398 77092 3423 77132
rect 3169 77069 3255 77092
rect 3337 77069 3423 77092
rect 18289 77132 18375 77155
rect 18457 77132 18543 77155
rect 18289 77092 18314 77132
rect 18314 77092 18354 77132
rect 18354 77092 18375 77132
rect 18457 77092 18478 77132
rect 18478 77092 18518 77132
rect 18518 77092 18543 77132
rect 18289 77069 18375 77092
rect 18457 77069 18543 77092
rect 33409 77132 33495 77155
rect 33577 77132 33663 77155
rect 33409 77092 33434 77132
rect 33434 77092 33474 77132
rect 33474 77092 33495 77132
rect 33577 77092 33598 77132
rect 33598 77092 33638 77132
rect 33638 77092 33663 77132
rect 33409 77069 33495 77092
rect 33577 77069 33663 77092
rect 48529 77132 48615 77155
rect 48697 77132 48783 77155
rect 48529 77092 48554 77132
rect 48554 77092 48594 77132
rect 48594 77092 48615 77132
rect 48697 77092 48718 77132
rect 48718 77092 48758 77132
rect 48758 77092 48783 77132
rect 48529 77069 48615 77092
rect 48697 77069 48783 77092
rect 63649 77132 63735 77155
rect 63817 77132 63903 77155
rect 63649 77092 63674 77132
rect 63674 77092 63714 77132
rect 63714 77092 63735 77132
rect 63817 77092 63838 77132
rect 63838 77092 63878 77132
rect 63878 77092 63903 77132
rect 63649 77069 63735 77092
rect 63817 77069 63903 77092
rect 78769 77132 78855 77155
rect 78937 77132 79023 77155
rect 78769 77092 78794 77132
rect 78794 77092 78834 77132
rect 78834 77092 78855 77132
rect 78937 77092 78958 77132
rect 78958 77092 78998 77132
rect 78998 77092 79023 77132
rect 78769 77069 78855 77092
rect 78937 77069 79023 77092
rect 93889 77132 93975 77155
rect 94057 77132 94143 77155
rect 93889 77092 93914 77132
rect 93914 77092 93954 77132
rect 93954 77092 93975 77132
rect 94057 77092 94078 77132
rect 94078 77092 94118 77132
rect 94118 77092 94143 77132
rect 93889 77069 93975 77092
rect 94057 77069 94143 77092
rect 4409 76376 4495 76399
rect 4577 76376 4663 76399
rect 4409 76336 4434 76376
rect 4434 76336 4474 76376
rect 4474 76336 4495 76376
rect 4577 76336 4598 76376
rect 4598 76336 4638 76376
rect 4638 76336 4663 76376
rect 4409 76313 4495 76336
rect 4577 76313 4663 76336
rect 19529 76376 19615 76399
rect 19697 76376 19783 76399
rect 19529 76336 19554 76376
rect 19554 76336 19594 76376
rect 19594 76336 19615 76376
rect 19697 76336 19718 76376
rect 19718 76336 19758 76376
rect 19758 76336 19783 76376
rect 19529 76313 19615 76336
rect 19697 76313 19783 76336
rect 34649 76376 34735 76399
rect 34817 76376 34903 76399
rect 34649 76336 34674 76376
rect 34674 76336 34714 76376
rect 34714 76336 34735 76376
rect 34817 76336 34838 76376
rect 34838 76336 34878 76376
rect 34878 76336 34903 76376
rect 34649 76313 34735 76336
rect 34817 76313 34903 76336
rect 49769 76376 49855 76399
rect 49937 76376 50023 76399
rect 49769 76336 49794 76376
rect 49794 76336 49834 76376
rect 49834 76336 49855 76376
rect 49937 76336 49958 76376
rect 49958 76336 49998 76376
rect 49998 76336 50023 76376
rect 49769 76313 49855 76336
rect 49937 76313 50023 76336
rect 64889 76376 64975 76399
rect 65057 76376 65143 76399
rect 64889 76336 64914 76376
rect 64914 76336 64954 76376
rect 64954 76336 64975 76376
rect 65057 76336 65078 76376
rect 65078 76336 65118 76376
rect 65118 76336 65143 76376
rect 64889 76313 64975 76336
rect 65057 76313 65143 76336
rect 80009 76376 80095 76399
rect 80177 76376 80263 76399
rect 80009 76336 80034 76376
rect 80034 76336 80074 76376
rect 80074 76336 80095 76376
rect 80177 76336 80198 76376
rect 80198 76336 80238 76376
rect 80238 76336 80263 76376
rect 80009 76313 80095 76336
rect 80177 76313 80263 76336
rect 95129 76376 95215 76399
rect 95297 76376 95383 76399
rect 95129 76336 95154 76376
rect 95154 76336 95194 76376
rect 95194 76336 95215 76376
rect 95297 76336 95318 76376
rect 95318 76336 95358 76376
rect 95358 76336 95383 76376
rect 95129 76313 95215 76336
rect 95297 76313 95383 76336
rect 3169 75620 3255 75643
rect 3337 75620 3423 75643
rect 3169 75580 3194 75620
rect 3194 75580 3234 75620
rect 3234 75580 3255 75620
rect 3337 75580 3358 75620
rect 3358 75580 3398 75620
rect 3398 75580 3423 75620
rect 3169 75557 3255 75580
rect 3337 75557 3423 75580
rect 18289 75620 18375 75643
rect 18457 75620 18543 75643
rect 18289 75580 18314 75620
rect 18314 75580 18354 75620
rect 18354 75580 18375 75620
rect 18457 75580 18478 75620
rect 18478 75580 18518 75620
rect 18518 75580 18543 75620
rect 18289 75557 18375 75580
rect 18457 75557 18543 75580
rect 33409 75620 33495 75643
rect 33577 75620 33663 75643
rect 33409 75580 33434 75620
rect 33434 75580 33474 75620
rect 33474 75580 33495 75620
rect 33577 75580 33598 75620
rect 33598 75580 33638 75620
rect 33638 75580 33663 75620
rect 33409 75557 33495 75580
rect 33577 75557 33663 75580
rect 48529 75620 48615 75643
rect 48697 75620 48783 75643
rect 48529 75580 48554 75620
rect 48554 75580 48594 75620
rect 48594 75580 48615 75620
rect 48697 75580 48718 75620
rect 48718 75580 48758 75620
rect 48758 75580 48783 75620
rect 48529 75557 48615 75580
rect 48697 75557 48783 75580
rect 63649 75620 63735 75643
rect 63817 75620 63903 75643
rect 63649 75580 63674 75620
rect 63674 75580 63714 75620
rect 63714 75580 63735 75620
rect 63817 75580 63838 75620
rect 63838 75580 63878 75620
rect 63878 75580 63903 75620
rect 63649 75557 63735 75580
rect 63817 75557 63903 75580
rect 78769 75620 78855 75643
rect 78937 75620 79023 75643
rect 78769 75580 78794 75620
rect 78794 75580 78834 75620
rect 78834 75580 78855 75620
rect 78937 75580 78958 75620
rect 78958 75580 78998 75620
rect 78998 75580 79023 75620
rect 78769 75557 78855 75580
rect 78937 75557 79023 75580
rect 93889 75620 93975 75643
rect 94057 75620 94143 75643
rect 93889 75580 93914 75620
rect 93914 75580 93954 75620
rect 93954 75580 93975 75620
rect 94057 75580 94078 75620
rect 94078 75580 94118 75620
rect 94118 75580 94143 75620
rect 93889 75557 93975 75580
rect 94057 75557 94143 75580
rect 4409 74864 4495 74887
rect 4577 74864 4663 74887
rect 4409 74824 4434 74864
rect 4434 74824 4474 74864
rect 4474 74824 4495 74864
rect 4577 74824 4598 74864
rect 4598 74824 4638 74864
rect 4638 74824 4663 74864
rect 4409 74801 4495 74824
rect 4577 74801 4663 74824
rect 19529 74864 19615 74887
rect 19697 74864 19783 74887
rect 19529 74824 19554 74864
rect 19554 74824 19594 74864
rect 19594 74824 19615 74864
rect 19697 74824 19718 74864
rect 19718 74824 19758 74864
rect 19758 74824 19783 74864
rect 19529 74801 19615 74824
rect 19697 74801 19783 74824
rect 34649 74864 34735 74887
rect 34817 74864 34903 74887
rect 34649 74824 34674 74864
rect 34674 74824 34714 74864
rect 34714 74824 34735 74864
rect 34817 74824 34838 74864
rect 34838 74824 34878 74864
rect 34878 74824 34903 74864
rect 34649 74801 34735 74824
rect 34817 74801 34903 74824
rect 49769 74864 49855 74887
rect 49937 74864 50023 74887
rect 49769 74824 49794 74864
rect 49794 74824 49834 74864
rect 49834 74824 49855 74864
rect 49937 74824 49958 74864
rect 49958 74824 49998 74864
rect 49998 74824 50023 74864
rect 49769 74801 49855 74824
rect 49937 74801 50023 74824
rect 64889 74864 64975 74887
rect 65057 74864 65143 74887
rect 64889 74824 64914 74864
rect 64914 74824 64954 74864
rect 64954 74824 64975 74864
rect 65057 74824 65078 74864
rect 65078 74824 65118 74864
rect 65118 74824 65143 74864
rect 64889 74801 64975 74824
rect 65057 74801 65143 74824
rect 80009 74864 80095 74887
rect 80177 74864 80263 74887
rect 80009 74824 80034 74864
rect 80034 74824 80074 74864
rect 80074 74824 80095 74864
rect 80177 74824 80198 74864
rect 80198 74824 80238 74864
rect 80238 74824 80263 74864
rect 80009 74801 80095 74824
rect 80177 74801 80263 74824
rect 95129 74864 95215 74887
rect 95297 74864 95383 74887
rect 95129 74824 95154 74864
rect 95154 74824 95194 74864
rect 95194 74824 95215 74864
rect 95297 74824 95318 74864
rect 95318 74824 95358 74864
rect 95358 74824 95383 74864
rect 95129 74801 95215 74824
rect 95297 74801 95383 74824
rect 3169 74108 3255 74131
rect 3337 74108 3423 74131
rect 3169 74068 3194 74108
rect 3194 74068 3234 74108
rect 3234 74068 3255 74108
rect 3337 74068 3358 74108
rect 3358 74068 3398 74108
rect 3398 74068 3423 74108
rect 3169 74045 3255 74068
rect 3337 74045 3423 74068
rect 18289 74108 18375 74131
rect 18457 74108 18543 74131
rect 18289 74068 18314 74108
rect 18314 74068 18354 74108
rect 18354 74068 18375 74108
rect 18457 74068 18478 74108
rect 18478 74068 18518 74108
rect 18518 74068 18543 74108
rect 18289 74045 18375 74068
rect 18457 74045 18543 74068
rect 33409 74108 33495 74131
rect 33577 74108 33663 74131
rect 33409 74068 33434 74108
rect 33434 74068 33474 74108
rect 33474 74068 33495 74108
rect 33577 74068 33598 74108
rect 33598 74068 33638 74108
rect 33638 74068 33663 74108
rect 33409 74045 33495 74068
rect 33577 74045 33663 74068
rect 48529 74108 48615 74131
rect 48697 74108 48783 74131
rect 48529 74068 48554 74108
rect 48554 74068 48594 74108
rect 48594 74068 48615 74108
rect 48697 74068 48718 74108
rect 48718 74068 48758 74108
rect 48758 74068 48783 74108
rect 48529 74045 48615 74068
rect 48697 74045 48783 74068
rect 63649 74108 63735 74131
rect 63817 74108 63903 74131
rect 63649 74068 63674 74108
rect 63674 74068 63714 74108
rect 63714 74068 63735 74108
rect 63817 74068 63838 74108
rect 63838 74068 63878 74108
rect 63878 74068 63903 74108
rect 63649 74045 63735 74068
rect 63817 74045 63903 74068
rect 78769 74108 78855 74131
rect 78937 74108 79023 74131
rect 78769 74068 78794 74108
rect 78794 74068 78834 74108
rect 78834 74068 78855 74108
rect 78937 74068 78958 74108
rect 78958 74068 78998 74108
rect 78998 74068 79023 74108
rect 78769 74045 78855 74068
rect 78937 74045 79023 74068
rect 93889 74108 93975 74131
rect 94057 74108 94143 74131
rect 93889 74068 93914 74108
rect 93914 74068 93954 74108
rect 93954 74068 93975 74108
rect 94057 74068 94078 74108
rect 94078 74068 94118 74108
rect 94118 74068 94143 74108
rect 93889 74045 93975 74068
rect 94057 74045 94143 74068
rect 4409 73352 4495 73375
rect 4577 73352 4663 73375
rect 4409 73312 4434 73352
rect 4434 73312 4474 73352
rect 4474 73312 4495 73352
rect 4577 73312 4598 73352
rect 4598 73312 4638 73352
rect 4638 73312 4663 73352
rect 4409 73289 4495 73312
rect 4577 73289 4663 73312
rect 19529 73352 19615 73375
rect 19697 73352 19783 73375
rect 19529 73312 19554 73352
rect 19554 73312 19594 73352
rect 19594 73312 19615 73352
rect 19697 73312 19718 73352
rect 19718 73312 19758 73352
rect 19758 73312 19783 73352
rect 19529 73289 19615 73312
rect 19697 73289 19783 73312
rect 34649 73352 34735 73375
rect 34817 73352 34903 73375
rect 34649 73312 34674 73352
rect 34674 73312 34714 73352
rect 34714 73312 34735 73352
rect 34817 73312 34838 73352
rect 34838 73312 34878 73352
rect 34878 73312 34903 73352
rect 34649 73289 34735 73312
rect 34817 73289 34903 73312
rect 49769 73352 49855 73375
rect 49937 73352 50023 73375
rect 49769 73312 49794 73352
rect 49794 73312 49834 73352
rect 49834 73312 49855 73352
rect 49937 73312 49958 73352
rect 49958 73312 49998 73352
rect 49998 73312 50023 73352
rect 49769 73289 49855 73312
rect 49937 73289 50023 73312
rect 64889 73352 64975 73375
rect 65057 73352 65143 73375
rect 64889 73312 64914 73352
rect 64914 73312 64954 73352
rect 64954 73312 64975 73352
rect 65057 73312 65078 73352
rect 65078 73312 65118 73352
rect 65118 73312 65143 73352
rect 64889 73289 64975 73312
rect 65057 73289 65143 73312
rect 80009 73352 80095 73375
rect 80177 73352 80263 73375
rect 80009 73312 80034 73352
rect 80034 73312 80074 73352
rect 80074 73312 80095 73352
rect 80177 73312 80198 73352
rect 80198 73312 80238 73352
rect 80238 73312 80263 73352
rect 80009 73289 80095 73312
rect 80177 73289 80263 73312
rect 95129 73352 95215 73375
rect 95297 73352 95383 73375
rect 95129 73312 95154 73352
rect 95154 73312 95194 73352
rect 95194 73312 95215 73352
rect 95297 73312 95318 73352
rect 95318 73312 95358 73352
rect 95358 73312 95383 73352
rect 95129 73289 95215 73312
rect 95297 73289 95383 73312
rect 3169 72596 3255 72619
rect 3337 72596 3423 72619
rect 3169 72556 3194 72596
rect 3194 72556 3234 72596
rect 3234 72556 3255 72596
rect 3337 72556 3358 72596
rect 3358 72556 3398 72596
rect 3398 72556 3423 72596
rect 3169 72533 3255 72556
rect 3337 72533 3423 72556
rect 18289 72596 18375 72619
rect 18457 72596 18543 72619
rect 18289 72556 18314 72596
rect 18314 72556 18354 72596
rect 18354 72556 18375 72596
rect 18457 72556 18478 72596
rect 18478 72556 18518 72596
rect 18518 72556 18543 72596
rect 18289 72533 18375 72556
rect 18457 72533 18543 72556
rect 33409 72596 33495 72619
rect 33577 72596 33663 72619
rect 33409 72556 33434 72596
rect 33434 72556 33474 72596
rect 33474 72556 33495 72596
rect 33577 72556 33598 72596
rect 33598 72556 33638 72596
rect 33638 72556 33663 72596
rect 33409 72533 33495 72556
rect 33577 72533 33663 72556
rect 48529 72596 48615 72619
rect 48697 72596 48783 72619
rect 48529 72556 48554 72596
rect 48554 72556 48594 72596
rect 48594 72556 48615 72596
rect 48697 72556 48718 72596
rect 48718 72556 48758 72596
rect 48758 72556 48783 72596
rect 48529 72533 48615 72556
rect 48697 72533 48783 72556
rect 63649 72596 63735 72619
rect 63817 72596 63903 72619
rect 63649 72556 63674 72596
rect 63674 72556 63714 72596
rect 63714 72556 63735 72596
rect 63817 72556 63838 72596
rect 63838 72556 63878 72596
rect 63878 72556 63903 72596
rect 63649 72533 63735 72556
rect 63817 72533 63903 72556
rect 78769 72596 78855 72619
rect 78937 72596 79023 72619
rect 78769 72556 78794 72596
rect 78794 72556 78834 72596
rect 78834 72556 78855 72596
rect 78937 72556 78958 72596
rect 78958 72556 78998 72596
rect 78998 72556 79023 72596
rect 78769 72533 78855 72556
rect 78937 72533 79023 72556
rect 93889 72596 93975 72619
rect 94057 72596 94143 72619
rect 93889 72556 93914 72596
rect 93914 72556 93954 72596
rect 93954 72556 93975 72596
rect 94057 72556 94078 72596
rect 94078 72556 94118 72596
rect 94118 72556 94143 72596
rect 93889 72533 93975 72556
rect 94057 72533 94143 72556
rect 4409 71840 4495 71863
rect 4577 71840 4663 71863
rect 4409 71800 4434 71840
rect 4434 71800 4474 71840
rect 4474 71800 4495 71840
rect 4577 71800 4598 71840
rect 4598 71800 4638 71840
rect 4638 71800 4663 71840
rect 4409 71777 4495 71800
rect 4577 71777 4663 71800
rect 19529 71840 19615 71863
rect 19697 71840 19783 71863
rect 19529 71800 19554 71840
rect 19554 71800 19594 71840
rect 19594 71800 19615 71840
rect 19697 71800 19718 71840
rect 19718 71800 19758 71840
rect 19758 71800 19783 71840
rect 19529 71777 19615 71800
rect 19697 71777 19783 71800
rect 34649 71840 34735 71863
rect 34817 71840 34903 71863
rect 34649 71800 34674 71840
rect 34674 71800 34714 71840
rect 34714 71800 34735 71840
rect 34817 71800 34838 71840
rect 34838 71800 34878 71840
rect 34878 71800 34903 71840
rect 34649 71777 34735 71800
rect 34817 71777 34903 71800
rect 49769 71840 49855 71863
rect 49937 71840 50023 71863
rect 49769 71800 49794 71840
rect 49794 71800 49834 71840
rect 49834 71800 49855 71840
rect 49937 71800 49958 71840
rect 49958 71800 49998 71840
rect 49998 71800 50023 71840
rect 49769 71777 49855 71800
rect 49937 71777 50023 71800
rect 64889 71840 64975 71863
rect 65057 71840 65143 71863
rect 64889 71800 64914 71840
rect 64914 71800 64954 71840
rect 64954 71800 64975 71840
rect 65057 71800 65078 71840
rect 65078 71800 65118 71840
rect 65118 71800 65143 71840
rect 64889 71777 64975 71800
rect 65057 71777 65143 71800
rect 80009 71840 80095 71863
rect 80177 71840 80263 71863
rect 80009 71800 80034 71840
rect 80034 71800 80074 71840
rect 80074 71800 80095 71840
rect 80177 71800 80198 71840
rect 80198 71800 80238 71840
rect 80238 71800 80263 71840
rect 80009 71777 80095 71800
rect 80177 71777 80263 71800
rect 95129 71840 95215 71863
rect 95297 71840 95383 71863
rect 95129 71800 95154 71840
rect 95154 71800 95194 71840
rect 95194 71800 95215 71840
rect 95297 71800 95318 71840
rect 95318 71800 95358 71840
rect 95358 71800 95383 71840
rect 95129 71777 95215 71800
rect 95297 71777 95383 71800
rect 3169 71084 3255 71107
rect 3337 71084 3423 71107
rect 3169 71044 3194 71084
rect 3194 71044 3234 71084
rect 3234 71044 3255 71084
rect 3337 71044 3358 71084
rect 3358 71044 3398 71084
rect 3398 71044 3423 71084
rect 3169 71021 3255 71044
rect 3337 71021 3423 71044
rect 18289 71084 18375 71107
rect 18457 71084 18543 71107
rect 18289 71044 18314 71084
rect 18314 71044 18354 71084
rect 18354 71044 18375 71084
rect 18457 71044 18478 71084
rect 18478 71044 18518 71084
rect 18518 71044 18543 71084
rect 18289 71021 18375 71044
rect 18457 71021 18543 71044
rect 33409 71084 33495 71107
rect 33577 71084 33663 71107
rect 33409 71044 33434 71084
rect 33434 71044 33474 71084
rect 33474 71044 33495 71084
rect 33577 71044 33598 71084
rect 33598 71044 33638 71084
rect 33638 71044 33663 71084
rect 33409 71021 33495 71044
rect 33577 71021 33663 71044
rect 48529 71084 48615 71107
rect 48697 71084 48783 71107
rect 48529 71044 48554 71084
rect 48554 71044 48594 71084
rect 48594 71044 48615 71084
rect 48697 71044 48718 71084
rect 48718 71044 48758 71084
rect 48758 71044 48783 71084
rect 48529 71021 48615 71044
rect 48697 71021 48783 71044
rect 63649 71084 63735 71107
rect 63817 71084 63903 71107
rect 63649 71044 63674 71084
rect 63674 71044 63714 71084
rect 63714 71044 63735 71084
rect 63817 71044 63838 71084
rect 63838 71044 63878 71084
rect 63878 71044 63903 71084
rect 63649 71021 63735 71044
rect 63817 71021 63903 71044
rect 78769 71084 78855 71107
rect 78937 71084 79023 71107
rect 78769 71044 78794 71084
rect 78794 71044 78834 71084
rect 78834 71044 78855 71084
rect 78937 71044 78958 71084
rect 78958 71044 78998 71084
rect 78998 71044 79023 71084
rect 78769 71021 78855 71044
rect 78937 71021 79023 71044
rect 93889 71084 93975 71107
rect 94057 71084 94143 71107
rect 93889 71044 93914 71084
rect 93914 71044 93954 71084
rect 93954 71044 93975 71084
rect 94057 71044 94078 71084
rect 94078 71044 94118 71084
rect 94118 71044 94143 71084
rect 93889 71021 93975 71044
rect 94057 71021 94143 71044
rect 4409 70328 4495 70351
rect 4577 70328 4663 70351
rect 4409 70288 4434 70328
rect 4434 70288 4474 70328
rect 4474 70288 4495 70328
rect 4577 70288 4598 70328
rect 4598 70288 4638 70328
rect 4638 70288 4663 70328
rect 4409 70265 4495 70288
rect 4577 70265 4663 70288
rect 19529 70328 19615 70351
rect 19697 70328 19783 70351
rect 19529 70288 19554 70328
rect 19554 70288 19594 70328
rect 19594 70288 19615 70328
rect 19697 70288 19718 70328
rect 19718 70288 19758 70328
rect 19758 70288 19783 70328
rect 19529 70265 19615 70288
rect 19697 70265 19783 70288
rect 34649 70328 34735 70351
rect 34817 70328 34903 70351
rect 34649 70288 34674 70328
rect 34674 70288 34714 70328
rect 34714 70288 34735 70328
rect 34817 70288 34838 70328
rect 34838 70288 34878 70328
rect 34878 70288 34903 70328
rect 34649 70265 34735 70288
rect 34817 70265 34903 70288
rect 49769 70328 49855 70351
rect 49937 70328 50023 70351
rect 49769 70288 49794 70328
rect 49794 70288 49834 70328
rect 49834 70288 49855 70328
rect 49937 70288 49958 70328
rect 49958 70288 49998 70328
rect 49998 70288 50023 70328
rect 49769 70265 49855 70288
rect 49937 70265 50023 70288
rect 64889 70328 64975 70351
rect 65057 70328 65143 70351
rect 64889 70288 64914 70328
rect 64914 70288 64954 70328
rect 64954 70288 64975 70328
rect 65057 70288 65078 70328
rect 65078 70288 65118 70328
rect 65118 70288 65143 70328
rect 64889 70265 64975 70288
rect 65057 70265 65143 70288
rect 80009 70328 80095 70351
rect 80177 70328 80263 70351
rect 80009 70288 80034 70328
rect 80034 70288 80074 70328
rect 80074 70288 80095 70328
rect 80177 70288 80198 70328
rect 80198 70288 80238 70328
rect 80238 70288 80263 70328
rect 80009 70265 80095 70288
rect 80177 70265 80263 70288
rect 95129 70328 95215 70351
rect 95297 70328 95383 70351
rect 95129 70288 95154 70328
rect 95154 70288 95194 70328
rect 95194 70288 95215 70328
rect 95297 70288 95318 70328
rect 95318 70288 95358 70328
rect 95358 70288 95383 70328
rect 95129 70265 95215 70288
rect 95297 70265 95383 70288
rect 3169 69572 3255 69595
rect 3337 69572 3423 69595
rect 3169 69532 3194 69572
rect 3194 69532 3234 69572
rect 3234 69532 3255 69572
rect 3337 69532 3358 69572
rect 3358 69532 3398 69572
rect 3398 69532 3423 69572
rect 3169 69509 3255 69532
rect 3337 69509 3423 69532
rect 18289 69572 18375 69595
rect 18457 69572 18543 69595
rect 18289 69532 18314 69572
rect 18314 69532 18354 69572
rect 18354 69532 18375 69572
rect 18457 69532 18478 69572
rect 18478 69532 18518 69572
rect 18518 69532 18543 69572
rect 18289 69509 18375 69532
rect 18457 69509 18543 69532
rect 33409 69572 33495 69595
rect 33577 69572 33663 69595
rect 33409 69532 33434 69572
rect 33434 69532 33474 69572
rect 33474 69532 33495 69572
rect 33577 69532 33598 69572
rect 33598 69532 33638 69572
rect 33638 69532 33663 69572
rect 33409 69509 33495 69532
rect 33577 69509 33663 69532
rect 48529 69572 48615 69595
rect 48697 69572 48783 69595
rect 48529 69532 48554 69572
rect 48554 69532 48594 69572
rect 48594 69532 48615 69572
rect 48697 69532 48718 69572
rect 48718 69532 48758 69572
rect 48758 69532 48783 69572
rect 48529 69509 48615 69532
rect 48697 69509 48783 69532
rect 63649 69572 63735 69595
rect 63817 69572 63903 69595
rect 63649 69532 63674 69572
rect 63674 69532 63714 69572
rect 63714 69532 63735 69572
rect 63817 69532 63838 69572
rect 63838 69532 63878 69572
rect 63878 69532 63903 69572
rect 63649 69509 63735 69532
rect 63817 69509 63903 69532
rect 78769 69572 78855 69595
rect 78937 69572 79023 69595
rect 78769 69532 78794 69572
rect 78794 69532 78834 69572
rect 78834 69532 78855 69572
rect 78937 69532 78958 69572
rect 78958 69532 78998 69572
rect 78998 69532 79023 69572
rect 78769 69509 78855 69532
rect 78937 69509 79023 69532
rect 93889 69572 93975 69595
rect 94057 69572 94143 69595
rect 93889 69532 93914 69572
rect 93914 69532 93954 69572
rect 93954 69532 93975 69572
rect 94057 69532 94078 69572
rect 94078 69532 94118 69572
rect 94118 69532 94143 69572
rect 93889 69509 93975 69532
rect 94057 69509 94143 69532
rect 4409 68816 4495 68839
rect 4577 68816 4663 68839
rect 4409 68776 4434 68816
rect 4434 68776 4474 68816
rect 4474 68776 4495 68816
rect 4577 68776 4598 68816
rect 4598 68776 4638 68816
rect 4638 68776 4663 68816
rect 4409 68753 4495 68776
rect 4577 68753 4663 68776
rect 19529 68816 19615 68839
rect 19697 68816 19783 68839
rect 19529 68776 19554 68816
rect 19554 68776 19594 68816
rect 19594 68776 19615 68816
rect 19697 68776 19718 68816
rect 19718 68776 19758 68816
rect 19758 68776 19783 68816
rect 19529 68753 19615 68776
rect 19697 68753 19783 68776
rect 34649 68816 34735 68839
rect 34817 68816 34903 68839
rect 34649 68776 34674 68816
rect 34674 68776 34714 68816
rect 34714 68776 34735 68816
rect 34817 68776 34838 68816
rect 34838 68776 34878 68816
rect 34878 68776 34903 68816
rect 34649 68753 34735 68776
rect 34817 68753 34903 68776
rect 49769 68816 49855 68839
rect 49937 68816 50023 68839
rect 49769 68776 49794 68816
rect 49794 68776 49834 68816
rect 49834 68776 49855 68816
rect 49937 68776 49958 68816
rect 49958 68776 49998 68816
rect 49998 68776 50023 68816
rect 49769 68753 49855 68776
rect 49937 68753 50023 68776
rect 64889 68816 64975 68839
rect 65057 68816 65143 68839
rect 64889 68776 64914 68816
rect 64914 68776 64954 68816
rect 64954 68776 64975 68816
rect 65057 68776 65078 68816
rect 65078 68776 65118 68816
rect 65118 68776 65143 68816
rect 64889 68753 64975 68776
rect 65057 68753 65143 68776
rect 80009 68816 80095 68839
rect 80177 68816 80263 68839
rect 80009 68776 80034 68816
rect 80034 68776 80074 68816
rect 80074 68776 80095 68816
rect 80177 68776 80198 68816
rect 80198 68776 80238 68816
rect 80238 68776 80263 68816
rect 80009 68753 80095 68776
rect 80177 68753 80263 68776
rect 95129 68816 95215 68839
rect 95297 68816 95383 68839
rect 95129 68776 95154 68816
rect 95154 68776 95194 68816
rect 95194 68776 95215 68816
rect 95297 68776 95318 68816
rect 95318 68776 95358 68816
rect 95358 68776 95383 68816
rect 95129 68753 95215 68776
rect 95297 68753 95383 68776
rect 3169 68060 3255 68083
rect 3337 68060 3423 68083
rect 3169 68020 3194 68060
rect 3194 68020 3234 68060
rect 3234 68020 3255 68060
rect 3337 68020 3358 68060
rect 3358 68020 3398 68060
rect 3398 68020 3423 68060
rect 3169 67997 3255 68020
rect 3337 67997 3423 68020
rect 18289 68060 18375 68083
rect 18457 68060 18543 68083
rect 18289 68020 18314 68060
rect 18314 68020 18354 68060
rect 18354 68020 18375 68060
rect 18457 68020 18478 68060
rect 18478 68020 18518 68060
rect 18518 68020 18543 68060
rect 18289 67997 18375 68020
rect 18457 67997 18543 68020
rect 33409 68060 33495 68083
rect 33577 68060 33663 68083
rect 33409 68020 33434 68060
rect 33434 68020 33474 68060
rect 33474 68020 33495 68060
rect 33577 68020 33598 68060
rect 33598 68020 33638 68060
rect 33638 68020 33663 68060
rect 33409 67997 33495 68020
rect 33577 67997 33663 68020
rect 48529 68060 48615 68083
rect 48697 68060 48783 68083
rect 48529 68020 48554 68060
rect 48554 68020 48594 68060
rect 48594 68020 48615 68060
rect 48697 68020 48718 68060
rect 48718 68020 48758 68060
rect 48758 68020 48783 68060
rect 48529 67997 48615 68020
rect 48697 67997 48783 68020
rect 63649 68060 63735 68083
rect 63817 68060 63903 68083
rect 63649 68020 63674 68060
rect 63674 68020 63714 68060
rect 63714 68020 63735 68060
rect 63817 68020 63838 68060
rect 63838 68020 63878 68060
rect 63878 68020 63903 68060
rect 63649 67997 63735 68020
rect 63817 67997 63903 68020
rect 78769 68060 78855 68083
rect 78937 68060 79023 68083
rect 78769 68020 78794 68060
rect 78794 68020 78834 68060
rect 78834 68020 78855 68060
rect 78937 68020 78958 68060
rect 78958 68020 78998 68060
rect 78998 68020 79023 68060
rect 78769 67997 78855 68020
rect 78937 67997 79023 68020
rect 93889 68060 93975 68083
rect 94057 68060 94143 68083
rect 93889 68020 93914 68060
rect 93914 68020 93954 68060
rect 93954 68020 93975 68060
rect 94057 68020 94078 68060
rect 94078 68020 94118 68060
rect 94118 68020 94143 68060
rect 93889 67997 93975 68020
rect 94057 67997 94143 68020
rect 4409 67304 4495 67327
rect 4577 67304 4663 67327
rect 4409 67264 4434 67304
rect 4434 67264 4474 67304
rect 4474 67264 4495 67304
rect 4577 67264 4598 67304
rect 4598 67264 4638 67304
rect 4638 67264 4663 67304
rect 4409 67241 4495 67264
rect 4577 67241 4663 67264
rect 19529 67304 19615 67327
rect 19697 67304 19783 67327
rect 19529 67264 19554 67304
rect 19554 67264 19594 67304
rect 19594 67264 19615 67304
rect 19697 67264 19718 67304
rect 19718 67264 19758 67304
rect 19758 67264 19783 67304
rect 19529 67241 19615 67264
rect 19697 67241 19783 67264
rect 34649 67304 34735 67327
rect 34817 67304 34903 67327
rect 34649 67264 34674 67304
rect 34674 67264 34714 67304
rect 34714 67264 34735 67304
rect 34817 67264 34838 67304
rect 34838 67264 34878 67304
rect 34878 67264 34903 67304
rect 34649 67241 34735 67264
rect 34817 67241 34903 67264
rect 49769 67304 49855 67327
rect 49937 67304 50023 67327
rect 49769 67264 49794 67304
rect 49794 67264 49834 67304
rect 49834 67264 49855 67304
rect 49937 67264 49958 67304
rect 49958 67264 49998 67304
rect 49998 67264 50023 67304
rect 49769 67241 49855 67264
rect 49937 67241 50023 67264
rect 64889 67304 64975 67327
rect 65057 67304 65143 67327
rect 64889 67264 64914 67304
rect 64914 67264 64954 67304
rect 64954 67264 64975 67304
rect 65057 67264 65078 67304
rect 65078 67264 65118 67304
rect 65118 67264 65143 67304
rect 64889 67241 64975 67264
rect 65057 67241 65143 67264
rect 80009 67304 80095 67327
rect 80177 67304 80263 67327
rect 80009 67264 80034 67304
rect 80034 67264 80074 67304
rect 80074 67264 80095 67304
rect 80177 67264 80198 67304
rect 80198 67264 80238 67304
rect 80238 67264 80263 67304
rect 80009 67241 80095 67264
rect 80177 67241 80263 67264
rect 95129 67304 95215 67327
rect 95297 67304 95383 67327
rect 95129 67264 95154 67304
rect 95154 67264 95194 67304
rect 95194 67264 95215 67304
rect 95297 67264 95318 67304
rect 95318 67264 95358 67304
rect 95358 67264 95383 67304
rect 95129 67241 95215 67264
rect 95297 67241 95383 67264
rect 3169 66548 3255 66571
rect 3337 66548 3423 66571
rect 3169 66508 3194 66548
rect 3194 66508 3234 66548
rect 3234 66508 3255 66548
rect 3337 66508 3358 66548
rect 3358 66508 3398 66548
rect 3398 66508 3423 66548
rect 3169 66485 3255 66508
rect 3337 66485 3423 66508
rect 18289 66548 18375 66571
rect 18457 66548 18543 66571
rect 18289 66508 18314 66548
rect 18314 66508 18354 66548
rect 18354 66508 18375 66548
rect 18457 66508 18478 66548
rect 18478 66508 18518 66548
rect 18518 66508 18543 66548
rect 18289 66485 18375 66508
rect 18457 66485 18543 66508
rect 33409 66548 33495 66571
rect 33577 66548 33663 66571
rect 33409 66508 33434 66548
rect 33434 66508 33474 66548
rect 33474 66508 33495 66548
rect 33577 66508 33598 66548
rect 33598 66508 33638 66548
rect 33638 66508 33663 66548
rect 33409 66485 33495 66508
rect 33577 66485 33663 66508
rect 48529 66548 48615 66571
rect 48697 66548 48783 66571
rect 48529 66508 48554 66548
rect 48554 66508 48594 66548
rect 48594 66508 48615 66548
rect 48697 66508 48718 66548
rect 48718 66508 48758 66548
rect 48758 66508 48783 66548
rect 48529 66485 48615 66508
rect 48697 66485 48783 66508
rect 63649 66548 63735 66571
rect 63817 66548 63903 66571
rect 63649 66508 63674 66548
rect 63674 66508 63714 66548
rect 63714 66508 63735 66548
rect 63817 66508 63838 66548
rect 63838 66508 63878 66548
rect 63878 66508 63903 66548
rect 63649 66485 63735 66508
rect 63817 66485 63903 66508
rect 78769 66548 78855 66571
rect 78937 66548 79023 66571
rect 78769 66508 78794 66548
rect 78794 66508 78834 66548
rect 78834 66508 78855 66548
rect 78937 66508 78958 66548
rect 78958 66508 78998 66548
rect 78998 66508 79023 66548
rect 78769 66485 78855 66508
rect 78937 66485 79023 66508
rect 93889 66548 93975 66571
rect 94057 66548 94143 66571
rect 93889 66508 93914 66548
rect 93914 66508 93954 66548
rect 93954 66508 93975 66548
rect 94057 66508 94078 66548
rect 94078 66508 94118 66548
rect 94118 66508 94143 66548
rect 93889 66485 93975 66508
rect 94057 66485 94143 66508
rect 4409 65792 4495 65815
rect 4577 65792 4663 65815
rect 4409 65752 4434 65792
rect 4434 65752 4474 65792
rect 4474 65752 4495 65792
rect 4577 65752 4598 65792
rect 4598 65752 4638 65792
rect 4638 65752 4663 65792
rect 4409 65729 4495 65752
rect 4577 65729 4663 65752
rect 19529 65792 19615 65815
rect 19697 65792 19783 65815
rect 19529 65752 19554 65792
rect 19554 65752 19594 65792
rect 19594 65752 19615 65792
rect 19697 65752 19718 65792
rect 19718 65752 19758 65792
rect 19758 65752 19783 65792
rect 19529 65729 19615 65752
rect 19697 65729 19783 65752
rect 34649 65792 34735 65815
rect 34817 65792 34903 65815
rect 34649 65752 34674 65792
rect 34674 65752 34714 65792
rect 34714 65752 34735 65792
rect 34817 65752 34838 65792
rect 34838 65752 34878 65792
rect 34878 65752 34903 65792
rect 34649 65729 34735 65752
rect 34817 65729 34903 65752
rect 49769 65792 49855 65815
rect 49937 65792 50023 65815
rect 49769 65752 49794 65792
rect 49794 65752 49834 65792
rect 49834 65752 49855 65792
rect 49937 65752 49958 65792
rect 49958 65752 49998 65792
rect 49998 65752 50023 65792
rect 49769 65729 49855 65752
rect 49937 65729 50023 65752
rect 64889 65792 64975 65815
rect 65057 65792 65143 65815
rect 64889 65752 64914 65792
rect 64914 65752 64954 65792
rect 64954 65752 64975 65792
rect 65057 65752 65078 65792
rect 65078 65752 65118 65792
rect 65118 65752 65143 65792
rect 64889 65729 64975 65752
rect 65057 65729 65143 65752
rect 80009 65792 80095 65815
rect 80177 65792 80263 65815
rect 80009 65752 80034 65792
rect 80034 65752 80074 65792
rect 80074 65752 80095 65792
rect 80177 65752 80198 65792
rect 80198 65752 80238 65792
rect 80238 65752 80263 65792
rect 80009 65729 80095 65752
rect 80177 65729 80263 65752
rect 95129 65792 95215 65815
rect 95297 65792 95383 65815
rect 95129 65752 95154 65792
rect 95154 65752 95194 65792
rect 95194 65752 95215 65792
rect 95297 65752 95318 65792
rect 95318 65752 95358 65792
rect 95358 65752 95383 65792
rect 95129 65729 95215 65752
rect 95297 65729 95383 65752
rect 3169 65036 3255 65059
rect 3337 65036 3423 65059
rect 3169 64996 3194 65036
rect 3194 64996 3234 65036
rect 3234 64996 3255 65036
rect 3337 64996 3358 65036
rect 3358 64996 3398 65036
rect 3398 64996 3423 65036
rect 3169 64973 3255 64996
rect 3337 64973 3423 64996
rect 18289 65036 18375 65059
rect 18457 65036 18543 65059
rect 18289 64996 18314 65036
rect 18314 64996 18354 65036
rect 18354 64996 18375 65036
rect 18457 64996 18478 65036
rect 18478 64996 18518 65036
rect 18518 64996 18543 65036
rect 18289 64973 18375 64996
rect 18457 64973 18543 64996
rect 33409 65036 33495 65059
rect 33577 65036 33663 65059
rect 33409 64996 33434 65036
rect 33434 64996 33474 65036
rect 33474 64996 33495 65036
rect 33577 64996 33598 65036
rect 33598 64996 33638 65036
rect 33638 64996 33663 65036
rect 33409 64973 33495 64996
rect 33577 64973 33663 64996
rect 48529 65036 48615 65059
rect 48697 65036 48783 65059
rect 48529 64996 48554 65036
rect 48554 64996 48594 65036
rect 48594 64996 48615 65036
rect 48697 64996 48718 65036
rect 48718 64996 48758 65036
rect 48758 64996 48783 65036
rect 48529 64973 48615 64996
rect 48697 64973 48783 64996
rect 63649 65036 63735 65059
rect 63817 65036 63903 65059
rect 63649 64996 63674 65036
rect 63674 64996 63714 65036
rect 63714 64996 63735 65036
rect 63817 64996 63838 65036
rect 63838 64996 63878 65036
rect 63878 64996 63903 65036
rect 63649 64973 63735 64996
rect 63817 64973 63903 64996
rect 78769 65036 78855 65059
rect 78937 65036 79023 65059
rect 78769 64996 78794 65036
rect 78794 64996 78834 65036
rect 78834 64996 78855 65036
rect 78937 64996 78958 65036
rect 78958 64996 78998 65036
rect 78998 64996 79023 65036
rect 78769 64973 78855 64996
rect 78937 64973 79023 64996
rect 93889 65036 93975 65059
rect 94057 65036 94143 65059
rect 93889 64996 93914 65036
rect 93914 64996 93954 65036
rect 93954 64996 93975 65036
rect 94057 64996 94078 65036
rect 94078 64996 94118 65036
rect 94118 64996 94143 65036
rect 93889 64973 93975 64996
rect 94057 64973 94143 64996
rect 4409 64280 4495 64303
rect 4577 64280 4663 64303
rect 4409 64240 4434 64280
rect 4434 64240 4474 64280
rect 4474 64240 4495 64280
rect 4577 64240 4598 64280
rect 4598 64240 4638 64280
rect 4638 64240 4663 64280
rect 4409 64217 4495 64240
rect 4577 64217 4663 64240
rect 19529 64280 19615 64303
rect 19697 64280 19783 64303
rect 19529 64240 19554 64280
rect 19554 64240 19594 64280
rect 19594 64240 19615 64280
rect 19697 64240 19718 64280
rect 19718 64240 19758 64280
rect 19758 64240 19783 64280
rect 19529 64217 19615 64240
rect 19697 64217 19783 64240
rect 34649 64280 34735 64303
rect 34817 64280 34903 64303
rect 34649 64240 34674 64280
rect 34674 64240 34714 64280
rect 34714 64240 34735 64280
rect 34817 64240 34838 64280
rect 34838 64240 34878 64280
rect 34878 64240 34903 64280
rect 34649 64217 34735 64240
rect 34817 64217 34903 64240
rect 49769 64280 49855 64303
rect 49937 64280 50023 64303
rect 49769 64240 49794 64280
rect 49794 64240 49834 64280
rect 49834 64240 49855 64280
rect 49937 64240 49958 64280
rect 49958 64240 49998 64280
rect 49998 64240 50023 64280
rect 49769 64217 49855 64240
rect 49937 64217 50023 64240
rect 64889 64280 64975 64303
rect 65057 64280 65143 64303
rect 64889 64240 64914 64280
rect 64914 64240 64954 64280
rect 64954 64240 64975 64280
rect 65057 64240 65078 64280
rect 65078 64240 65118 64280
rect 65118 64240 65143 64280
rect 64889 64217 64975 64240
rect 65057 64217 65143 64240
rect 80009 64280 80095 64303
rect 80177 64280 80263 64303
rect 80009 64240 80034 64280
rect 80034 64240 80074 64280
rect 80074 64240 80095 64280
rect 80177 64240 80198 64280
rect 80198 64240 80238 64280
rect 80238 64240 80263 64280
rect 80009 64217 80095 64240
rect 80177 64217 80263 64240
rect 95129 64280 95215 64303
rect 95297 64280 95383 64303
rect 95129 64240 95154 64280
rect 95154 64240 95194 64280
rect 95194 64240 95215 64280
rect 95297 64240 95318 64280
rect 95318 64240 95358 64280
rect 95358 64240 95383 64280
rect 95129 64217 95215 64240
rect 95297 64217 95383 64240
rect 3169 63524 3255 63547
rect 3337 63524 3423 63547
rect 3169 63484 3194 63524
rect 3194 63484 3234 63524
rect 3234 63484 3255 63524
rect 3337 63484 3358 63524
rect 3358 63484 3398 63524
rect 3398 63484 3423 63524
rect 3169 63461 3255 63484
rect 3337 63461 3423 63484
rect 18289 63524 18375 63547
rect 18457 63524 18543 63547
rect 18289 63484 18314 63524
rect 18314 63484 18354 63524
rect 18354 63484 18375 63524
rect 18457 63484 18478 63524
rect 18478 63484 18518 63524
rect 18518 63484 18543 63524
rect 18289 63461 18375 63484
rect 18457 63461 18543 63484
rect 33409 63524 33495 63547
rect 33577 63524 33663 63547
rect 33409 63484 33434 63524
rect 33434 63484 33474 63524
rect 33474 63484 33495 63524
rect 33577 63484 33598 63524
rect 33598 63484 33638 63524
rect 33638 63484 33663 63524
rect 33409 63461 33495 63484
rect 33577 63461 33663 63484
rect 48529 63524 48615 63547
rect 48697 63524 48783 63547
rect 48529 63484 48554 63524
rect 48554 63484 48594 63524
rect 48594 63484 48615 63524
rect 48697 63484 48718 63524
rect 48718 63484 48758 63524
rect 48758 63484 48783 63524
rect 48529 63461 48615 63484
rect 48697 63461 48783 63484
rect 63649 63524 63735 63547
rect 63817 63524 63903 63547
rect 63649 63484 63674 63524
rect 63674 63484 63714 63524
rect 63714 63484 63735 63524
rect 63817 63484 63838 63524
rect 63838 63484 63878 63524
rect 63878 63484 63903 63524
rect 63649 63461 63735 63484
rect 63817 63461 63903 63484
rect 78769 63524 78855 63547
rect 78937 63524 79023 63547
rect 78769 63484 78794 63524
rect 78794 63484 78834 63524
rect 78834 63484 78855 63524
rect 78937 63484 78958 63524
rect 78958 63484 78998 63524
rect 78998 63484 79023 63524
rect 78769 63461 78855 63484
rect 78937 63461 79023 63484
rect 93889 63524 93975 63547
rect 94057 63524 94143 63547
rect 93889 63484 93914 63524
rect 93914 63484 93954 63524
rect 93954 63484 93975 63524
rect 94057 63484 94078 63524
rect 94078 63484 94118 63524
rect 94118 63484 94143 63524
rect 93889 63461 93975 63484
rect 94057 63461 94143 63484
rect 4409 62768 4495 62791
rect 4577 62768 4663 62791
rect 4409 62728 4434 62768
rect 4434 62728 4474 62768
rect 4474 62728 4495 62768
rect 4577 62728 4598 62768
rect 4598 62728 4638 62768
rect 4638 62728 4663 62768
rect 4409 62705 4495 62728
rect 4577 62705 4663 62728
rect 19529 62768 19615 62791
rect 19697 62768 19783 62791
rect 19529 62728 19554 62768
rect 19554 62728 19594 62768
rect 19594 62728 19615 62768
rect 19697 62728 19718 62768
rect 19718 62728 19758 62768
rect 19758 62728 19783 62768
rect 19529 62705 19615 62728
rect 19697 62705 19783 62728
rect 34649 62768 34735 62791
rect 34817 62768 34903 62791
rect 34649 62728 34674 62768
rect 34674 62728 34714 62768
rect 34714 62728 34735 62768
rect 34817 62728 34838 62768
rect 34838 62728 34878 62768
rect 34878 62728 34903 62768
rect 34649 62705 34735 62728
rect 34817 62705 34903 62728
rect 49769 62768 49855 62791
rect 49937 62768 50023 62791
rect 49769 62728 49794 62768
rect 49794 62728 49834 62768
rect 49834 62728 49855 62768
rect 49937 62728 49958 62768
rect 49958 62728 49998 62768
rect 49998 62728 50023 62768
rect 49769 62705 49855 62728
rect 49937 62705 50023 62728
rect 64889 62768 64975 62791
rect 65057 62768 65143 62791
rect 64889 62728 64914 62768
rect 64914 62728 64954 62768
rect 64954 62728 64975 62768
rect 65057 62728 65078 62768
rect 65078 62728 65118 62768
rect 65118 62728 65143 62768
rect 64889 62705 64975 62728
rect 65057 62705 65143 62728
rect 80009 62768 80095 62791
rect 80177 62768 80263 62791
rect 80009 62728 80034 62768
rect 80034 62728 80074 62768
rect 80074 62728 80095 62768
rect 80177 62728 80198 62768
rect 80198 62728 80238 62768
rect 80238 62728 80263 62768
rect 80009 62705 80095 62728
rect 80177 62705 80263 62728
rect 95129 62768 95215 62791
rect 95297 62768 95383 62791
rect 95129 62728 95154 62768
rect 95154 62728 95194 62768
rect 95194 62728 95215 62768
rect 95297 62728 95318 62768
rect 95318 62728 95358 62768
rect 95358 62728 95383 62768
rect 95129 62705 95215 62728
rect 95297 62705 95383 62728
rect 3169 62012 3255 62035
rect 3337 62012 3423 62035
rect 3169 61972 3194 62012
rect 3194 61972 3234 62012
rect 3234 61972 3255 62012
rect 3337 61972 3358 62012
rect 3358 61972 3398 62012
rect 3398 61972 3423 62012
rect 3169 61949 3255 61972
rect 3337 61949 3423 61972
rect 18289 62012 18375 62035
rect 18457 62012 18543 62035
rect 18289 61972 18314 62012
rect 18314 61972 18354 62012
rect 18354 61972 18375 62012
rect 18457 61972 18478 62012
rect 18478 61972 18518 62012
rect 18518 61972 18543 62012
rect 18289 61949 18375 61972
rect 18457 61949 18543 61972
rect 33409 62012 33495 62035
rect 33577 62012 33663 62035
rect 33409 61972 33434 62012
rect 33434 61972 33474 62012
rect 33474 61972 33495 62012
rect 33577 61972 33598 62012
rect 33598 61972 33638 62012
rect 33638 61972 33663 62012
rect 33409 61949 33495 61972
rect 33577 61949 33663 61972
rect 48529 62012 48615 62035
rect 48697 62012 48783 62035
rect 48529 61972 48554 62012
rect 48554 61972 48594 62012
rect 48594 61972 48615 62012
rect 48697 61972 48718 62012
rect 48718 61972 48758 62012
rect 48758 61972 48783 62012
rect 48529 61949 48615 61972
rect 48697 61949 48783 61972
rect 63649 62012 63735 62035
rect 63817 62012 63903 62035
rect 63649 61972 63674 62012
rect 63674 61972 63714 62012
rect 63714 61972 63735 62012
rect 63817 61972 63838 62012
rect 63838 61972 63878 62012
rect 63878 61972 63903 62012
rect 63649 61949 63735 61972
rect 63817 61949 63903 61972
rect 78769 62012 78855 62035
rect 78937 62012 79023 62035
rect 78769 61972 78794 62012
rect 78794 61972 78834 62012
rect 78834 61972 78855 62012
rect 78937 61972 78958 62012
rect 78958 61972 78998 62012
rect 78998 61972 79023 62012
rect 78769 61949 78855 61972
rect 78937 61949 79023 61972
rect 93889 62012 93975 62035
rect 94057 62012 94143 62035
rect 93889 61972 93914 62012
rect 93914 61972 93954 62012
rect 93954 61972 93975 62012
rect 94057 61972 94078 62012
rect 94078 61972 94118 62012
rect 94118 61972 94143 62012
rect 93889 61949 93975 61972
rect 94057 61949 94143 61972
rect 4409 61256 4495 61279
rect 4577 61256 4663 61279
rect 4409 61216 4434 61256
rect 4434 61216 4474 61256
rect 4474 61216 4495 61256
rect 4577 61216 4598 61256
rect 4598 61216 4638 61256
rect 4638 61216 4663 61256
rect 4409 61193 4495 61216
rect 4577 61193 4663 61216
rect 19529 61256 19615 61279
rect 19697 61256 19783 61279
rect 19529 61216 19554 61256
rect 19554 61216 19594 61256
rect 19594 61216 19615 61256
rect 19697 61216 19718 61256
rect 19718 61216 19758 61256
rect 19758 61216 19783 61256
rect 19529 61193 19615 61216
rect 19697 61193 19783 61216
rect 34649 61256 34735 61279
rect 34817 61256 34903 61279
rect 34649 61216 34674 61256
rect 34674 61216 34714 61256
rect 34714 61216 34735 61256
rect 34817 61216 34838 61256
rect 34838 61216 34878 61256
rect 34878 61216 34903 61256
rect 34649 61193 34735 61216
rect 34817 61193 34903 61216
rect 49769 61256 49855 61279
rect 49937 61256 50023 61279
rect 49769 61216 49794 61256
rect 49794 61216 49834 61256
rect 49834 61216 49855 61256
rect 49937 61216 49958 61256
rect 49958 61216 49998 61256
rect 49998 61216 50023 61256
rect 49769 61193 49855 61216
rect 49937 61193 50023 61216
rect 64889 61256 64975 61279
rect 65057 61256 65143 61279
rect 64889 61216 64914 61256
rect 64914 61216 64954 61256
rect 64954 61216 64975 61256
rect 65057 61216 65078 61256
rect 65078 61216 65118 61256
rect 65118 61216 65143 61256
rect 64889 61193 64975 61216
rect 65057 61193 65143 61216
rect 80009 61256 80095 61279
rect 80177 61256 80263 61279
rect 80009 61216 80034 61256
rect 80034 61216 80074 61256
rect 80074 61216 80095 61256
rect 80177 61216 80198 61256
rect 80198 61216 80238 61256
rect 80238 61216 80263 61256
rect 80009 61193 80095 61216
rect 80177 61193 80263 61216
rect 95129 61256 95215 61279
rect 95297 61256 95383 61279
rect 95129 61216 95154 61256
rect 95154 61216 95194 61256
rect 95194 61216 95215 61256
rect 95297 61216 95318 61256
rect 95318 61216 95358 61256
rect 95358 61216 95383 61256
rect 95129 61193 95215 61216
rect 95297 61193 95383 61216
rect 3169 60500 3255 60523
rect 3337 60500 3423 60523
rect 3169 60460 3194 60500
rect 3194 60460 3234 60500
rect 3234 60460 3255 60500
rect 3337 60460 3358 60500
rect 3358 60460 3398 60500
rect 3398 60460 3423 60500
rect 3169 60437 3255 60460
rect 3337 60437 3423 60460
rect 18289 60500 18375 60523
rect 18457 60500 18543 60523
rect 18289 60460 18314 60500
rect 18314 60460 18354 60500
rect 18354 60460 18375 60500
rect 18457 60460 18478 60500
rect 18478 60460 18518 60500
rect 18518 60460 18543 60500
rect 18289 60437 18375 60460
rect 18457 60437 18543 60460
rect 33409 60500 33495 60523
rect 33577 60500 33663 60523
rect 33409 60460 33434 60500
rect 33434 60460 33474 60500
rect 33474 60460 33495 60500
rect 33577 60460 33598 60500
rect 33598 60460 33638 60500
rect 33638 60460 33663 60500
rect 33409 60437 33495 60460
rect 33577 60437 33663 60460
rect 48529 60500 48615 60523
rect 48697 60500 48783 60523
rect 48529 60460 48554 60500
rect 48554 60460 48594 60500
rect 48594 60460 48615 60500
rect 48697 60460 48718 60500
rect 48718 60460 48758 60500
rect 48758 60460 48783 60500
rect 48529 60437 48615 60460
rect 48697 60437 48783 60460
rect 63649 60500 63735 60523
rect 63817 60500 63903 60523
rect 63649 60460 63674 60500
rect 63674 60460 63714 60500
rect 63714 60460 63735 60500
rect 63817 60460 63838 60500
rect 63838 60460 63878 60500
rect 63878 60460 63903 60500
rect 63649 60437 63735 60460
rect 63817 60437 63903 60460
rect 78769 60500 78855 60523
rect 78937 60500 79023 60523
rect 78769 60460 78794 60500
rect 78794 60460 78834 60500
rect 78834 60460 78855 60500
rect 78937 60460 78958 60500
rect 78958 60460 78998 60500
rect 78998 60460 79023 60500
rect 78769 60437 78855 60460
rect 78937 60437 79023 60460
rect 93889 60500 93975 60523
rect 94057 60500 94143 60523
rect 93889 60460 93914 60500
rect 93914 60460 93954 60500
rect 93954 60460 93975 60500
rect 94057 60460 94078 60500
rect 94078 60460 94118 60500
rect 94118 60460 94143 60500
rect 93889 60437 93975 60460
rect 94057 60437 94143 60460
rect 4409 59744 4495 59767
rect 4577 59744 4663 59767
rect 4409 59704 4434 59744
rect 4434 59704 4474 59744
rect 4474 59704 4495 59744
rect 4577 59704 4598 59744
rect 4598 59704 4638 59744
rect 4638 59704 4663 59744
rect 4409 59681 4495 59704
rect 4577 59681 4663 59704
rect 19529 59744 19615 59767
rect 19697 59744 19783 59767
rect 19529 59704 19554 59744
rect 19554 59704 19594 59744
rect 19594 59704 19615 59744
rect 19697 59704 19718 59744
rect 19718 59704 19758 59744
rect 19758 59704 19783 59744
rect 19529 59681 19615 59704
rect 19697 59681 19783 59704
rect 34649 59744 34735 59767
rect 34817 59744 34903 59767
rect 34649 59704 34674 59744
rect 34674 59704 34714 59744
rect 34714 59704 34735 59744
rect 34817 59704 34838 59744
rect 34838 59704 34878 59744
rect 34878 59704 34903 59744
rect 34649 59681 34735 59704
rect 34817 59681 34903 59704
rect 49769 59744 49855 59767
rect 49937 59744 50023 59767
rect 49769 59704 49794 59744
rect 49794 59704 49834 59744
rect 49834 59704 49855 59744
rect 49937 59704 49958 59744
rect 49958 59704 49998 59744
rect 49998 59704 50023 59744
rect 49769 59681 49855 59704
rect 49937 59681 50023 59704
rect 64889 59744 64975 59767
rect 65057 59744 65143 59767
rect 64889 59704 64914 59744
rect 64914 59704 64954 59744
rect 64954 59704 64975 59744
rect 65057 59704 65078 59744
rect 65078 59704 65118 59744
rect 65118 59704 65143 59744
rect 64889 59681 64975 59704
rect 65057 59681 65143 59704
rect 80009 59744 80095 59767
rect 80177 59744 80263 59767
rect 80009 59704 80034 59744
rect 80034 59704 80074 59744
rect 80074 59704 80095 59744
rect 80177 59704 80198 59744
rect 80198 59704 80238 59744
rect 80238 59704 80263 59744
rect 80009 59681 80095 59704
rect 80177 59681 80263 59704
rect 95129 59744 95215 59767
rect 95297 59744 95383 59767
rect 95129 59704 95154 59744
rect 95154 59704 95194 59744
rect 95194 59704 95215 59744
rect 95297 59704 95318 59744
rect 95318 59704 95358 59744
rect 95358 59704 95383 59744
rect 95129 59681 95215 59704
rect 95297 59681 95383 59704
rect 3169 58988 3255 59011
rect 3337 58988 3423 59011
rect 3169 58948 3194 58988
rect 3194 58948 3234 58988
rect 3234 58948 3255 58988
rect 3337 58948 3358 58988
rect 3358 58948 3398 58988
rect 3398 58948 3423 58988
rect 3169 58925 3255 58948
rect 3337 58925 3423 58948
rect 18289 58988 18375 59011
rect 18457 58988 18543 59011
rect 18289 58948 18314 58988
rect 18314 58948 18354 58988
rect 18354 58948 18375 58988
rect 18457 58948 18478 58988
rect 18478 58948 18518 58988
rect 18518 58948 18543 58988
rect 18289 58925 18375 58948
rect 18457 58925 18543 58948
rect 33409 58988 33495 59011
rect 33577 58988 33663 59011
rect 33409 58948 33434 58988
rect 33434 58948 33474 58988
rect 33474 58948 33495 58988
rect 33577 58948 33598 58988
rect 33598 58948 33638 58988
rect 33638 58948 33663 58988
rect 33409 58925 33495 58948
rect 33577 58925 33663 58948
rect 48529 58988 48615 59011
rect 48697 58988 48783 59011
rect 48529 58948 48554 58988
rect 48554 58948 48594 58988
rect 48594 58948 48615 58988
rect 48697 58948 48718 58988
rect 48718 58948 48758 58988
rect 48758 58948 48783 58988
rect 48529 58925 48615 58948
rect 48697 58925 48783 58948
rect 63649 58988 63735 59011
rect 63817 58988 63903 59011
rect 63649 58948 63674 58988
rect 63674 58948 63714 58988
rect 63714 58948 63735 58988
rect 63817 58948 63838 58988
rect 63838 58948 63878 58988
rect 63878 58948 63903 58988
rect 63649 58925 63735 58948
rect 63817 58925 63903 58948
rect 78769 58988 78855 59011
rect 78937 58988 79023 59011
rect 78769 58948 78794 58988
rect 78794 58948 78834 58988
rect 78834 58948 78855 58988
rect 78937 58948 78958 58988
rect 78958 58948 78998 58988
rect 78998 58948 79023 58988
rect 78769 58925 78855 58948
rect 78937 58925 79023 58948
rect 93889 58988 93975 59011
rect 94057 58988 94143 59011
rect 93889 58948 93914 58988
rect 93914 58948 93954 58988
rect 93954 58948 93975 58988
rect 94057 58948 94078 58988
rect 94078 58948 94118 58988
rect 94118 58948 94143 58988
rect 93889 58925 93975 58948
rect 94057 58925 94143 58948
rect 4409 58232 4495 58255
rect 4577 58232 4663 58255
rect 4409 58192 4434 58232
rect 4434 58192 4474 58232
rect 4474 58192 4495 58232
rect 4577 58192 4598 58232
rect 4598 58192 4638 58232
rect 4638 58192 4663 58232
rect 4409 58169 4495 58192
rect 4577 58169 4663 58192
rect 19529 58232 19615 58255
rect 19697 58232 19783 58255
rect 19529 58192 19554 58232
rect 19554 58192 19594 58232
rect 19594 58192 19615 58232
rect 19697 58192 19718 58232
rect 19718 58192 19758 58232
rect 19758 58192 19783 58232
rect 19529 58169 19615 58192
rect 19697 58169 19783 58192
rect 34649 58232 34735 58255
rect 34817 58232 34903 58255
rect 34649 58192 34674 58232
rect 34674 58192 34714 58232
rect 34714 58192 34735 58232
rect 34817 58192 34838 58232
rect 34838 58192 34878 58232
rect 34878 58192 34903 58232
rect 34649 58169 34735 58192
rect 34817 58169 34903 58192
rect 49769 58232 49855 58255
rect 49937 58232 50023 58255
rect 49769 58192 49794 58232
rect 49794 58192 49834 58232
rect 49834 58192 49855 58232
rect 49937 58192 49958 58232
rect 49958 58192 49998 58232
rect 49998 58192 50023 58232
rect 49769 58169 49855 58192
rect 49937 58169 50023 58192
rect 64889 58232 64975 58255
rect 65057 58232 65143 58255
rect 64889 58192 64914 58232
rect 64914 58192 64954 58232
rect 64954 58192 64975 58232
rect 65057 58192 65078 58232
rect 65078 58192 65118 58232
rect 65118 58192 65143 58232
rect 64889 58169 64975 58192
rect 65057 58169 65143 58192
rect 80009 58232 80095 58255
rect 80177 58232 80263 58255
rect 80009 58192 80034 58232
rect 80034 58192 80074 58232
rect 80074 58192 80095 58232
rect 80177 58192 80198 58232
rect 80198 58192 80238 58232
rect 80238 58192 80263 58232
rect 80009 58169 80095 58192
rect 80177 58169 80263 58192
rect 95129 58232 95215 58255
rect 95297 58232 95383 58255
rect 95129 58192 95154 58232
rect 95154 58192 95194 58232
rect 95194 58192 95215 58232
rect 95297 58192 95318 58232
rect 95318 58192 95358 58232
rect 95358 58192 95383 58232
rect 95129 58169 95215 58192
rect 95297 58169 95383 58192
rect 3169 57476 3255 57499
rect 3337 57476 3423 57499
rect 3169 57436 3194 57476
rect 3194 57436 3234 57476
rect 3234 57436 3255 57476
rect 3337 57436 3358 57476
rect 3358 57436 3398 57476
rect 3398 57436 3423 57476
rect 3169 57413 3255 57436
rect 3337 57413 3423 57436
rect 18289 57476 18375 57499
rect 18457 57476 18543 57499
rect 18289 57436 18314 57476
rect 18314 57436 18354 57476
rect 18354 57436 18375 57476
rect 18457 57436 18478 57476
rect 18478 57436 18518 57476
rect 18518 57436 18543 57476
rect 18289 57413 18375 57436
rect 18457 57413 18543 57436
rect 33409 57476 33495 57499
rect 33577 57476 33663 57499
rect 33409 57436 33434 57476
rect 33434 57436 33474 57476
rect 33474 57436 33495 57476
rect 33577 57436 33598 57476
rect 33598 57436 33638 57476
rect 33638 57436 33663 57476
rect 33409 57413 33495 57436
rect 33577 57413 33663 57436
rect 48529 57476 48615 57499
rect 48697 57476 48783 57499
rect 48529 57436 48554 57476
rect 48554 57436 48594 57476
rect 48594 57436 48615 57476
rect 48697 57436 48718 57476
rect 48718 57436 48758 57476
rect 48758 57436 48783 57476
rect 48529 57413 48615 57436
rect 48697 57413 48783 57436
rect 63649 57476 63735 57499
rect 63817 57476 63903 57499
rect 63649 57436 63674 57476
rect 63674 57436 63714 57476
rect 63714 57436 63735 57476
rect 63817 57436 63838 57476
rect 63838 57436 63878 57476
rect 63878 57436 63903 57476
rect 63649 57413 63735 57436
rect 63817 57413 63903 57436
rect 78769 57476 78855 57499
rect 78937 57476 79023 57499
rect 78769 57436 78794 57476
rect 78794 57436 78834 57476
rect 78834 57436 78855 57476
rect 78937 57436 78958 57476
rect 78958 57436 78998 57476
rect 78998 57436 79023 57476
rect 78769 57413 78855 57436
rect 78937 57413 79023 57436
rect 93889 57476 93975 57499
rect 94057 57476 94143 57499
rect 93889 57436 93914 57476
rect 93914 57436 93954 57476
rect 93954 57436 93975 57476
rect 94057 57436 94078 57476
rect 94078 57436 94118 57476
rect 94118 57436 94143 57476
rect 93889 57413 93975 57436
rect 94057 57413 94143 57436
rect 4409 56720 4495 56743
rect 4577 56720 4663 56743
rect 4409 56680 4434 56720
rect 4434 56680 4474 56720
rect 4474 56680 4495 56720
rect 4577 56680 4598 56720
rect 4598 56680 4638 56720
rect 4638 56680 4663 56720
rect 4409 56657 4495 56680
rect 4577 56657 4663 56680
rect 19529 56720 19615 56743
rect 19697 56720 19783 56743
rect 19529 56680 19554 56720
rect 19554 56680 19594 56720
rect 19594 56680 19615 56720
rect 19697 56680 19718 56720
rect 19718 56680 19758 56720
rect 19758 56680 19783 56720
rect 19529 56657 19615 56680
rect 19697 56657 19783 56680
rect 34649 56720 34735 56743
rect 34817 56720 34903 56743
rect 34649 56680 34674 56720
rect 34674 56680 34714 56720
rect 34714 56680 34735 56720
rect 34817 56680 34838 56720
rect 34838 56680 34878 56720
rect 34878 56680 34903 56720
rect 34649 56657 34735 56680
rect 34817 56657 34903 56680
rect 49769 56720 49855 56743
rect 49937 56720 50023 56743
rect 49769 56680 49794 56720
rect 49794 56680 49834 56720
rect 49834 56680 49855 56720
rect 49937 56680 49958 56720
rect 49958 56680 49998 56720
rect 49998 56680 50023 56720
rect 49769 56657 49855 56680
rect 49937 56657 50023 56680
rect 64889 56720 64975 56743
rect 65057 56720 65143 56743
rect 64889 56680 64914 56720
rect 64914 56680 64954 56720
rect 64954 56680 64975 56720
rect 65057 56680 65078 56720
rect 65078 56680 65118 56720
rect 65118 56680 65143 56720
rect 64889 56657 64975 56680
rect 65057 56657 65143 56680
rect 80009 56720 80095 56743
rect 80177 56720 80263 56743
rect 80009 56680 80034 56720
rect 80034 56680 80074 56720
rect 80074 56680 80095 56720
rect 80177 56680 80198 56720
rect 80198 56680 80238 56720
rect 80238 56680 80263 56720
rect 80009 56657 80095 56680
rect 80177 56657 80263 56680
rect 95129 56720 95215 56743
rect 95297 56720 95383 56743
rect 95129 56680 95154 56720
rect 95154 56680 95194 56720
rect 95194 56680 95215 56720
rect 95297 56680 95318 56720
rect 95318 56680 95358 56720
rect 95358 56680 95383 56720
rect 95129 56657 95215 56680
rect 95297 56657 95383 56680
rect 3169 55964 3255 55987
rect 3337 55964 3423 55987
rect 3169 55924 3194 55964
rect 3194 55924 3234 55964
rect 3234 55924 3255 55964
rect 3337 55924 3358 55964
rect 3358 55924 3398 55964
rect 3398 55924 3423 55964
rect 3169 55901 3255 55924
rect 3337 55901 3423 55924
rect 18289 55964 18375 55987
rect 18457 55964 18543 55987
rect 18289 55924 18314 55964
rect 18314 55924 18354 55964
rect 18354 55924 18375 55964
rect 18457 55924 18478 55964
rect 18478 55924 18518 55964
rect 18518 55924 18543 55964
rect 18289 55901 18375 55924
rect 18457 55901 18543 55924
rect 33409 55964 33495 55987
rect 33577 55964 33663 55987
rect 33409 55924 33434 55964
rect 33434 55924 33474 55964
rect 33474 55924 33495 55964
rect 33577 55924 33598 55964
rect 33598 55924 33638 55964
rect 33638 55924 33663 55964
rect 33409 55901 33495 55924
rect 33577 55901 33663 55924
rect 48529 55964 48615 55987
rect 48697 55964 48783 55987
rect 48529 55924 48554 55964
rect 48554 55924 48594 55964
rect 48594 55924 48615 55964
rect 48697 55924 48718 55964
rect 48718 55924 48758 55964
rect 48758 55924 48783 55964
rect 48529 55901 48615 55924
rect 48697 55901 48783 55924
rect 63649 55964 63735 55987
rect 63817 55964 63903 55987
rect 63649 55924 63674 55964
rect 63674 55924 63714 55964
rect 63714 55924 63735 55964
rect 63817 55924 63838 55964
rect 63838 55924 63878 55964
rect 63878 55924 63903 55964
rect 63649 55901 63735 55924
rect 63817 55901 63903 55924
rect 78769 55964 78855 55987
rect 78937 55964 79023 55987
rect 78769 55924 78794 55964
rect 78794 55924 78834 55964
rect 78834 55924 78855 55964
rect 78937 55924 78958 55964
rect 78958 55924 78998 55964
rect 78998 55924 79023 55964
rect 78769 55901 78855 55924
rect 78937 55901 79023 55924
rect 93889 55964 93975 55987
rect 94057 55964 94143 55987
rect 93889 55924 93914 55964
rect 93914 55924 93954 55964
rect 93954 55924 93975 55964
rect 94057 55924 94078 55964
rect 94078 55924 94118 55964
rect 94118 55924 94143 55964
rect 93889 55901 93975 55924
rect 94057 55901 94143 55924
rect 4409 55208 4495 55231
rect 4577 55208 4663 55231
rect 4409 55168 4434 55208
rect 4434 55168 4474 55208
rect 4474 55168 4495 55208
rect 4577 55168 4598 55208
rect 4598 55168 4638 55208
rect 4638 55168 4663 55208
rect 4409 55145 4495 55168
rect 4577 55145 4663 55168
rect 19529 55208 19615 55231
rect 19697 55208 19783 55231
rect 19529 55168 19554 55208
rect 19554 55168 19594 55208
rect 19594 55168 19615 55208
rect 19697 55168 19718 55208
rect 19718 55168 19758 55208
rect 19758 55168 19783 55208
rect 19529 55145 19615 55168
rect 19697 55145 19783 55168
rect 34649 55208 34735 55231
rect 34817 55208 34903 55231
rect 34649 55168 34674 55208
rect 34674 55168 34714 55208
rect 34714 55168 34735 55208
rect 34817 55168 34838 55208
rect 34838 55168 34878 55208
rect 34878 55168 34903 55208
rect 34649 55145 34735 55168
rect 34817 55145 34903 55168
rect 49769 55208 49855 55231
rect 49937 55208 50023 55231
rect 49769 55168 49794 55208
rect 49794 55168 49834 55208
rect 49834 55168 49855 55208
rect 49937 55168 49958 55208
rect 49958 55168 49998 55208
rect 49998 55168 50023 55208
rect 49769 55145 49855 55168
rect 49937 55145 50023 55168
rect 64889 55208 64975 55231
rect 65057 55208 65143 55231
rect 64889 55168 64914 55208
rect 64914 55168 64954 55208
rect 64954 55168 64975 55208
rect 65057 55168 65078 55208
rect 65078 55168 65118 55208
rect 65118 55168 65143 55208
rect 64889 55145 64975 55168
rect 65057 55145 65143 55168
rect 80009 55208 80095 55231
rect 80177 55208 80263 55231
rect 80009 55168 80034 55208
rect 80034 55168 80074 55208
rect 80074 55168 80095 55208
rect 80177 55168 80198 55208
rect 80198 55168 80238 55208
rect 80238 55168 80263 55208
rect 80009 55145 80095 55168
rect 80177 55145 80263 55168
rect 95129 55208 95215 55231
rect 95297 55208 95383 55231
rect 95129 55168 95154 55208
rect 95154 55168 95194 55208
rect 95194 55168 95215 55208
rect 95297 55168 95318 55208
rect 95318 55168 95358 55208
rect 95358 55168 95383 55208
rect 95129 55145 95215 55168
rect 95297 55145 95383 55168
rect 3169 54452 3255 54475
rect 3337 54452 3423 54475
rect 3169 54412 3194 54452
rect 3194 54412 3234 54452
rect 3234 54412 3255 54452
rect 3337 54412 3358 54452
rect 3358 54412 3398 54452
rect 3398 54412 3423 54452
rect 3169 54389 3255 54412
rect 3337 54389 3423 54412
rect 18289 54452 18375 54475
rect 18457 54452 18543 54475
rect 18289 54412 18314 54452
rect 18314 54412 18354 54452
rect 18354 54412 18375 54452
rect 18457 54412 18478 54452
rect 18478 54412 18518 54452
rect 18518 54412 18543 54452
rect 18289 54389 18375 54412
rect 18457 54389 18543 54412
rect 33409 54452 33495 54475
rect 33577 54452 33663 54475
rect 33409 54412 33434 54452
rect 33434 54412 33474 54452
rect 33474 54412 33495 54452
rect 33577 54412 33598 54452
rect 33598 54412 33638 54452
rect 33638 54412 33663 54452
rect 33409 54389 33495 54412
rect 33577 54389 33663 54412
rect 48529 54452 48615 54475
rect 48697 54452 48783 54475
rect 48529 54412 48554 54452
rect 48554 54412 48594 54452
rect 48594 54412 48615 54452
rect 48697 54412 48718 54452
rect 48718 54412 48758 54452
rect 48758 54412 48783 54452
rect 48529 54389 48615 54412
rect 48697 54389 48783 54412
rect 63649 54452 63735 54475
rect 63817 54452 63903 54475
rect 63649 54412 63674 54452
rect 63674 54412 63714 54452
rect 63714 54412 63735 54452
rect 63817 54412 63838 54452
rect 63838 54412 63878 54452
rect 63878 54412 63903 54452
rect 63649 54389 63735 54412
rect 63817 54389 63903 54412
rect 78769 54452 78855 54475
rect 78937 54452 79023 54475
rect 78769 54412 78794 54452
rect 78794 54412 78834 54452
rect 78834 54412 78855 54452
rect 78937 54412 78958 54452
rect 78958 54412 78998 54452
rect 78998 54412 79023 54452
rect 78769 54389 78855 54412
rect 78937 54389 79023 54412
rect 93889 54452 93975 54475
rect 94057 54452 94143 54475
rect 93889 54412 93914 54452
rect 93914 54412 93954 54452
rect 93954 54412 93975 54452
rect 94057 54412 94078 54452
rect 94078 54412 94118 54452
rect 94118 54412 94143 54452
rect 93889 54389 93975 54412
rect 94057 54389 94143 54412
rect 4409 53696 4495 53719
rect 4577 53696 4663 53719
rect 4409 53656 4434 53696
rect 4434 53656 4474 53696
rect 4474 53656 4495 53696
rect 4577 53656 4598 53696
rect 4598 53656 4638 53696
rect 4638 53656 4663 53696
rect 4409 53633 4495 53656
rect 4577 53633 4663 53656
rect 19529 53696 19615 53719
rect 19697 53696 19783 53719
rect 19529 53656 19554 53696
rect 19554 53656 19594 53696
rect 19594 53656 19615 53696
rect 19697 53656 19718 53696
rect 19718 53656 19758 53696
rect 19758 53656 19783 53696
rect 19529 53633 19615 53656
rect 19697 53633 19783 53656
rect 34649 53696 34735 53719
rect 34817 53696 34903 53719
rect 34649 53656 34674 53696
rect 34674 53656 34714 53696
rect 34714 53656 34735 53696
rect 34817 53656 34838 53696
rect 34838 53656 34878 53696
rect 34878 53656 34903 53696
rect 34649 53633 34735 53656
rect 34817 53633 34903 53656
rect 49769 53696 49855 53719
rect 49937 53696 50023 53719
rect 49769 53656 49794 53696
rect 49794 53656 49834 53696
rect 49834 53656 49855 53696
rect 49937 53656 49958 53696
rect 49958 53656 49998 53696
rect 49998 53656 50023 53696
rect 49769 53633 49855 53656
rect 49937 53633 50023 53656
rect 64889 53696 64975 53719
rect 65057 53696 65143 53719
rect 64889 53656 64914 53696
rect 64914 53656 64954 53696
rect 64954 53656 64975 53696
rect 65057 53656 65078 53696
rect 65078 53656 65118 53696
rect 65118 53656 65143 53696
rect 64889 53633 64975 53656
rect 65057 53633 65143 53656
rect 80009 53696 80095 53719
rect 80177 53696 80263 53719
rect 80009 53656 80034 53696
rect 80034 53656 80074 53696
rect 80074 53656 80095 53696
rect 80177 53656 80198 53696
rect 80198 53656 80238 53696
rect 80238 53656 80263 53696
rect 80009 53633 80095 53656
rect 80177 53633 80263 53656
rect 95129 53696 95215 53719
rect 95297 53696 95383 53719
rect 95129 53656 95154 53696
rect 95154 53656 95194 53696
rect 95194 53656 95215 53696
rect 95297 53656 95318 53696
rect 95318 53656 95358 53696
rect 95358 53656 95383 53696
rect 95129 53633 95215 53656
rect 95297 53633 95383 53656
rect 3169 52940 3255 52963
rect 3337 52940 3423 52963
rect 3169 52900 3194 52940
rect 3194 52900 3234 52940
rect 3234 52900 3255 52940
rect 3337 52900 3358 52940
rect 3358 52900 3398 52940
rect 3398 52900 3423 52940
rect 3169 52877 3255 52900
rect 3337 52877 3423 52900
rect 18289 52940 18375 52963
rect 18457 52940 18543 52963
rect 18289 52900 18314 52940
rect 18314 52900 18354 52940
rect 18354 52900 18375 52940
rect 18457 52900 18478 52940
rect 18478 52900 18518 52940
rect 18518 52900 18543 52940
rect 18289 52877 18375 52900
rect 18457 52877 18543 52900
rect 33409 52940 33495 52963
rect 33577 52940 33663 52963
rect 33409 52900 33434 52940
rect 33434 52900 33474 52940
rect 33474 52900 33495 52940
rect 33577 52900 33598 52940
rect 33598 52900 33638 52940
rect 33638 52900 33663 52940
rect 33409 52877 33495 52900
rect 33577 52877 33663 52900
rect 48529 52940 48615 52963
rect 48697 52940 48783 52963
rect 48529 52900 48554 52940
rect 48554 52900 48594 52940
rect 48594 52900 48615 52940
rect 48697 52900 48718 52940
rect 48718 52900 48758 52940
rect 48758 52900 48783 52940
rect 48529 52877 48615 52900
rect 48697 52877 48783 52900
rect 63649 52940 63735 52963
rect 63817 52940 63903 52963
rect 63649 52900 63674 52940
rect 63674 52900 63714 52940
rect 63714 52900 63735 52940
rect 63817 52900 63838 52940
rect 63838 52900 63878 52940
rect 63878 52900 63903 52940
rect 63649 52877 63735 52900
rect 63817 52877 63903 52900
rect 78769 52940 78855 52963
rect 78937 52940 79023 52963
rect 78769 52900 78794 52940
rect 78794 52900 78834 52940
rect 78834 52900 78855 52940
rect 78937 52900 78958 52940
rect 78958 52900 78998 52940
rect 78998 52900 79023 52940
rect 78769 52877 78855 52900
rect 78937 52877 79023 52900
rect 93889 52940 93975 52963
rect 94057 52940 94143 52963
rect 93889 52900 93914 52940
rect 93914 52900 93954 52940
rect 93954 52900 93975 52940
rect 94057 52900 94078 52940
rect 94078 52900 94118 52940
rect 94118 52900 94143 52940
rect 93889 52877 93975 52900
rect 94057 52877 94143 52900
rect 4409 52184 4495 52207
rect 4577 52184 4663 52207
rect 4409 52144 4434 52184
rect 4434 52144 4474 52184
rect 4474 52144 4495 52184
rect 4577 52144 4598 52184
rect 4598 52144 4638 52184
rect 4638 52144 4663 52184
rect 4409 52121 4495 52144
rect 4577 52121 4663 52144
rect 19529 52184 19615 52207
rect 19697 52184 19783 52207
rect 19529 52144 19554 52184
rect 19554 52144 19594 52184
rect 19594 52144 19615 52184
rect 19697 52144 19718 52184
rect 19718 52144 19758 52184
rect 19758 52144 19783 52184
rect 19529 52121 19615 52144
rect 19697 52121 19783 52144
rect 34649 52184 34735 52207
rect 34817 52184 34903 52207
rect 34649 52144 34674 52184
rect 34674 52144 34714 52184
rect 34714 52144 34735 52184
rect 34817 52144 34838 52184
rect 34838 52144 34878 52184
rect 34878 52144 34903 52184
rect 34649 52121 34735 52144
rect 34817 52121 34903 52144
rect 49769 52184 49855 52207
rect 49937 52184 50023 52207
rect 49769 52144 49794 52184
rect 49794 52144 49834 52184
rect 49834 52144 49855 52184
rect 49937 52144 49958 52184
rect 49958 52144 49998 52184
rect 49998 52144 50023 52184
rect 49769 52121 49855 52144
rect 49937 52121 50023 52144
rect 64889 52184 64975 52207
rect 65057 52184 65143 52207
rect 64889 52144 64914 52184
rect 64914 52144 64954 52184
rect 64954 52144 64975 52184
rect 65057 52144 65078 52184
rect 65078 52144 65118 52184
rect 65118 52144 65143 52184
rect 64889 52121 64975 52144
rect 65057 52121 65143 52144
rect 80009 52184 80095 52207
rect 80177 52184 80263 52207
rect 80009 52144 80034 52184
rect 80034 52144 80074 52184
rect 80074 52144 80095 52184
rect 80177 52144 80198 52184
rect 80198 52144 80238 52184
rect 80238 52144 80263 52184
rect 80009 52121 80095 52144
rect 80177 52121 80263 52144
rect 95129 52184 95215 52207
rect 95297 52184 95383 52207
rect 95129 52144 95154 52184
rect 95154 52144 95194 52184
rect 95194 52144 95215 52184
rect 95297 52144 95318 52184
rect 95318 52144 95358 52184
rect 95358 52144 95383 52184
rect 95129 52121 95215 52144
rect 95297 52121 95383 52144
rect 3169 51428 3255 51451
rect 3337 51428 3423 51451
rect 3169 51388 3194 51428
rect 3194 51388 3234 51428
rect 3234 51388 3255 51428
rect 3337 51388 3358 51428
rect 3358 51388 3398 51428
rect 3398 51388 3423 51428
rect 3169 51365 3255 51388
rect 3337 51365 3423 51388
rect 18289 51428 18375 51451
rect 18457 51428 18543 51451
rect 18289 51388 18314 51428
rect 18314 51388 18354 51428
rect 18354 51388 18375 51428
rect 18457 51388 18478 51428
rect 18478 51388 18518 51428
rect 18518 51388 18543 51428
rect 18289 51365 18375 51388
rect 18457 51365 18543 51388
rect 33409 51428 33495 51451
rect 33577 51428 33663 51451
rect 33409 51388 33434 51428
rect 33434 51388 33474 51428
rect 33474 51388 33495 51428
rect 33577 51388 33598 51428
rect 33598 51388 33638 51428
rect 33638 51388 33663 51428
rect 33409 51365 33495 51388
rect 33577 51365 33663 51388
rect 48529 51428 48615 51451
rect 48697 51428 48783 51451
rect 48529 51388 48554 51428
rect 48554 51388 48594 51428
rect 48594 51388 48615 51428
rect 48697 51388 48718 51428
rect 48718 51388 48758 51428
rect 48758 51388 48783 51428
rect 48529 51365 48615 51388
rect 48697 51365 48783 51388
rect 63649 51428 63735 51451
rect 63817 51428 63903 51451
rect 63649 51388 63674 51428
rect 63674 51388 63714 51428
rect 63714 51388 63735 51428
rect 63817 51388 63838 51428
rect 63838 51388 63878 51428
rect 63878 51388 63903 51428
rect 63649 51365 63735 51388
rect 63817 51365 63903 51388
rect 78769 51428 78855 51451
rect 78937 51428 79023 51451
rect 78769 51388 78794 51428
rect 78794 51388 78834 51428
rect 78834 51388 78855 51428
rect 78937 51388 78958 51428
rect 78958 51388 78998 51428
rect 78998 51388 79023 51428
rect 78769 51365 78855 51388
rect 78937 51365 79023 51388
rect 93889 51428 93975 51451
rect 94057 51428 94143 51451
rect 93889 51388 93914 51428
rect 93914 51388 93954 51428
rect 93954 51388 93975 51428
rect 94057 51388 94078 51428
rect 94078 51388 94118 51428
rect 94118 51388 94143 51428
rect 93889 51365 93975 51388
rect 94057 51365 94143 51388
rect 4409 50672 4495 50695
rect 4577 50672 4663 50695
rect 4409 50632 4434 50672
rect 4434 50632 4474 50672
rect 4474 50632 4495 50672
rect 4577 50632 4598 50672
rect 4598 50632 4638 50672
rect 4638 50632 4663 50672
rect 4409 50609 4495 50632
rect 4577 50609 4663 50632
rect 19529 50672 19615 50695
rect 19697 50672 19783 50695
rect 19529 50632 19554 50672
rect 19554 50632 19594 50672
rect 19594 50632 19615 50672
rect 19697 50632 19718 50672
rect 19718 50632 19758 50672
rect 19758 50632 19783 50672
rect 19529 50609 19615 50632
rect 19697 50609 19783 50632
rect 34649 50672 34735 50695
rect 34817 50672 34903 50695
rect 34649 50632 34674 50672
rect 34674 50632 34714 50672
rect 34714 50632 34735 50672
rect 34817 50632 34838 50672
rect 34838 50632 34878 50672
rect 34878 50632 34903 50672
rect 34649 50609 34735 50632
rect 34817 50609 34903 50632
rect 49769 50672 49855 50695
rect 49937 50672 50023 50695
rect 49769 50632 49794 50672
rect 49794 50632 49834 50672
rect 49834 50632 49855 50672
rect 49937 50632 49958 50672
rect 49958 50632 49998 50672
rect 49998 50632 50023 50672
rect 49769 50609 49855 50632
rect 49937 50609 50023 50632
rect 64889 50672 64975 50695
rect 65057 50672 65143 50695
rect 64889 50632 64914 50672
rect 64914 50632 64954 50672
rect 64954 50632 64975 50672
rect 65057 50632 65078 50672
rect 65078 50632 65118 50672
rect 65118 50632 65143 50672
rect 64889 50609 64975 50632
rect 65057 50609 65143 50632
rect 80009 50672 80095 50695
rect 80177 50672 80263 50695
rect 80009 50632 80034 50672
rect 80034 50632 80074 50672
rect 80074 50632 80095 50672
rect 80177 50632 80198 50672
rect 80198 50632 80238 50672
rect 80238 50632 80263 50672
rect 80009 50609 80095 50632
rect 80177 50609 80263 50632
rect 95129 50672 95215 50695
rect 95297 50672 95383 50695
rect 95129 50632 95154 50672
rect 95154 50632 95194 50672
rect 95194 50632 95215 50672
rect 95297 50632 95318 50672
rect 95318 50632 95358 50672
rect 95358 50632 95383 50672
rect 95129 50609 95215 50632
rect 95297 50609 95383 50632
rect 3169 49916 3255 49939
rect 3337 49916 3423 49939
rect 3169 49876 3194 49916
rect 3194 49876 3234 49916
rect 3234 49876 3255 49916
rect 3337 49876 3358 49916
rect 3358 49876 3398 49916
rect 3398 49876 3423 49916
rect 3169 49853 3255 49876
rect 3337 49853 3423 49876
rect 18289 49916 18375 49939
rect 18457 49916 18543 49939
rect 18289 49876 18314 49916
rect 18314 49876 18354 49916
rect 18354 49876 18375 49916
rect 18457 49876 18478 49916
rect 18478 49876 18518 49916
rect 18518 49876 18543 49916
rect 18289 49853 18375 49876
rect 18457 49853 18543 49876
rect 33409 49916 33495 49939
rect 33577 49916 33663 49939
rect 33409 49876 33434 49916
rect 33434 49876 33474 49916
rect 33474 49876 33495 49916
rect 33577 49876 33598 49916
rect 33598 49876 33638 49916
rect 33638 49876 33663 49916
rect 33409 49853 33495 49876
rect 33577 49853 33663 49876
rect 48529 49916 48615 49939
rect 48697 49916 48783 49939
rect 48529 49876 48554 49916
rect 48554 49876 48594 49916
rect 48594 49876 48615 49916
rect 48697 49876 48718 49916
rect 48718 49876 48758 49916
rect 48758 49876 48783 49916
rect 48529 49853 48615 49876
rect 48697 49853 48783 49876
rect 63649 49916 63735 49939
rect 63817 49916 63903 49939
rect 63649 49876 63674 49916
rect 63674 49876 63714 49916
rect 63714 49876 63735 49916
rect 63817 49876 63838 49916
rect 63838 49876 63878 49916
rect 63878 49876 63903 49916
rect 63649 49853 63735 49876
rect 63817 49853 63903 49876
rect 78769 49916 78855 49939
rect 78937 49916 79023 49939
rect 78769 49876 78794 49916
rect 78794 49876 78834 49916
rect 78834 49876 78855 49916
rect 78937 49876 78958 49916
rect 78958 49876 78998 49916
rect 78998 49876 79023 49916
rect 78769 49853 78855 49876
rect 78937 49853 79023 49876
rect 93889 49916 93975 49939
rect 94057 49916 94143 49939
rect 93889 49876 93914 49916
rect 93914 49876 93954 49916
rect 93954 49876 93975 49916
rect 94057 49876 94078 49916
rect 94078 49876 94118 49916
rect 94118 49876 94143 49916
rect 93889 49853 93975 49876
rect 94057 49853 94143 49876
rect 4409 49160 4495 49183
rect 4577 49160 4663 49183
rect 4409 49120 4434 49160
rect 4434 49120 4474 49160
rect 4474 49120 4495 49160
rect 4577 49120 4598 49160
rect 4598 49120 4638 49160
rect 4638 49120 4663 49160
rect 4409 49097 4495 49120
rect 4577 49097 4663 49120
rect 19529 49160 19615 49183
rect 19697 49160 19783 49183
rect 19529 49120 19554 49160
rect 19554 49120 19594 49160
rect 19594 49120 19615 49160
rect 19697 49120 19718 49160
rect 19718 49120 19758 49160
rect 19758 49120 19783 49160
rect 19529 49097 19615 49120
rect 19697 49097 19783 49120
rect 34649 49160 34735 49183
rect 34817 49160 34903 49183
rect 34649 49120 34674 49160
rect 34674 49120 34714 49160
rect 34714 49120 34735 49160
rect 34817 49120 34838 49160
rect 34838 49120 34878 49160
rect 34878 49120 34903 49160
rect 34649 49097 34735 49120
rect 34817 49097 34903 49120
rect 49769 49160 49855 49183
rect 49937 49160 50023 49183
rect 49769 49120 49794 49160
rect 49794 49120 49834 49160
rect 49834 49120 49855 49160
rect 49937 49120 49958 49160
rect 49958 49120 49998 49160
rect 49998 49120 50023 49160
rect 49769 49097 49855 49120
rect 49937 49097 50023 49120
rect 64889 49160 64975 49183
rect 65057 49160 65143 49183
rect 64889 49120 64914 49160
rect 64914 49120 64954 49160
rect 64954 49120 64975 49160
rect 65057 49120 65078 49160
rect 65078 49120 65118 49160
rect 65118 49120 65143 49160
rect 64889 49097 64975 49120
rect 65057 49097 65143 49120
rect 80009 49160 80095 49183
rect 80177 49160 80263 49183
rect 80009 49120 80034 49160
rect 80034 49120 80074 49160
rect 80074 49120 80095 49160
rect 80177 49120 80198 49160
rect 80198 49120 80238 49160
rect 80238 49120 80263 49160
rect 80009 49097 80095 49120
rect 80177 49097 80263 49120
rect 95129 49160 95215 49183
rect 95297 49160 95383 49183
rect 95129 49120 95154 49160
rect 95154 49120 95194 49160
rect 95194 49120 95215 49160
rect 95297 49120 95318 49160
rect 95318 49120 95358 49160
rect 95358 49120 95383 49160
rect 95129 49097 95215 49120
rect 95297 49097 95383 49120
rect 3169 48404 3255 48427
rect 3337 48404 3423 48427
rect 3169 48364 3194 48404
rect 3194 48364 3234 48404
rect 3234 48364 3255 48404
rect 3337 48364 3358 48404
rect 3358 48364 3398 48404
rect 3398 48364 3423 48404
rect 3169 48341 3255 48364
rect 3337 48341 3423 48364
rect 18289 48404 18375 48427
rect 18457 48404 18543 48427
rect 18289 48364 18314 48404
rect 18314 48364 18354 48404
rect 18354 48364 18375 48404
rect 18457 48364 18478 48404
rect 18478 48364 18518 48404
rect 18518 48364 18543 48404
rect 18289 48341 18375 48364
rect 18457 48341 18543 48364
rect 33409 48404 33495 48427
rect 33577 48404 33663 48427
rect 33409 48364 33434 48404
rect 33434 48364 33474 48404
rect 33474 48364 33495 48404
rect 33577 48364 33598 48404
rect 33598 48364 33638 48404
rect 33638 48364 33663 48404
rect 33409 48341 33495 48364
rect 33577 48341 33663 48364
rect 48529 48404 48615 48427
rect 48697 48404 48783 48427
rect 48529 48364 48554 48404
rect 48554 48364 48594 48404
rect 48594 48364 48615 48404
rect 48697 48364 48718 48404
rect 48718 48364 48758 48404
rect 48758 48364 48783 48404
rect 48529 48341 48615 48364
rect 48697 48341 48783 48364
rect 63649 48404 63735 48427
rect 63817 48404 63903 48427
rect 63649 48364 63674 48404
rect 63674 48364 63714 48404
rect 63714 48364 63735 48404
rect 63817 48364 63838 48404
rect 63838 48364 63878 48404
rect 63878 48364 63903 48404
rect 63649 48341 63735 48364
rect 63817 48341 63903 48364
rect 78769 48404 78855 48427
rect 78937 48404 79023 48427
rect 78769 48364 78794 48404
rect 78794 48364 78834 48404
rect 78834 48364 78855 48404
rect 78937 48364 78958 48404
rect 78958 48364 78998 48404
rect 78998 48364 79023 48404
rect 78769 48341 78855 48364
rect 78937 48341 79023 48364
rect 93889 48404 93975 48427
rect 94057 48404 94143 48427
rect 93889 48364 93914 48404
rect 93914 48364 93954 48404
rect 93954 48364 93975 48404
rect 94057 48364 94078 48404
rect 94078 48364 94118 48404
rect 94118 48364 94143 48404
rect 93889 48341 93975 48364
rect 94057 48341 94143 48364
rect 4409 47648 4495 47671
rect 4577 47648 4663 47671
rect 4409 47608 4434 47648
rect 4434 47608 4474 47648
rect 4474 47608 4495 47648
rect 4577 47608 4598 47648
rect 4598 47608 4638 47648
rect 4638 47608 4663 47648
rect 4409 47585 4495 47608
rect 4577 47585 4663 47608
rect 19529 47648 19615 47671
rect 19697 47648 19783 47671
rect 19529 47608 19554 47648
rect 19554 47608 19594 47648
rect 19594 47608 19615 47648
rect 19697 47608 19718 47648
rect 19718 47608 19758 47648
rect 19758 47608 19783 47648
rect 19529 47585 19615 47608
rect 19697 47585 19783 47608
rect 34649 47648 34735 47671
rect 34817 47648 34903 47671
rect 34649 47608 34674 47648
rect 34674 47608 34714 47648
rect 34714 47608 34735 47648
rect 34817 47608 34838 47648
rect 34838 47608 34878 47648
rect 34878 47608 34903 47648
rect 34649 47585 34735 47608
rect 34817 47585 34903 47608
rect 49769 47648 49855 47671
rect 49937 47648 50023 47671
rect 49769 47608 49794 47648
rect 49794 47608 49834 47648
rect 49834 47608 49855 47648
rect 49937 47608 49958 47648
rect 49958 47608 49998 47648
rect 49998 47608 50023 47648
rect 49769 47585 49855 47608
rect 49937 47585 50023 47608
rect 64889 47648 64975 47671
rect 65057 47648 65143 47671
rect 64889 47608 64914 47648
rect 64914 47608 64954 47648
rect 64954 47608 64975 47648
rect 65057 47608 65078 47648
rect 65078 47608 65118 47648
rect 65118 47608 65143 47648
rect 64889 47585 64975 47608
rect 65057 47585 65143 47608
rect 80009 47648 80095 47671
rect 80177 47648 80263 47671
rect 80009 47608 80034 47648
rect 80034 47608 80074 47648
rect 80074 47608 80095 47648
rect 80177 47608 80198 47648
rect 80198 47608 80238 47648
rect 80238 47608 80263 47648
rect 80009 47585 80095 47608
rect 80177 47585 80263 47608
rect 95129 47648 95215 47671
rect 95297 47648 95383 47671
rect 95129 47608 95154 47648
rect 95154 47608 95194 47648
rect 95194 47608 95215 47648
rect 95297 47608 95318 47648
rect 95318 47608 95358 47648
rect 95358 47608 95383 47648
rect 95129 47585 95215 47608
rect 95297 47585 95383 47608
rect 3169 46892 3255 46915
rect 3337 46892 3423 46915
rect 3169 46852 3194 46892
rect 3194 46852 3234 46892
rect 3234 46852 3255 46892
rect 3337 46852 3358 46892
rect 3358 46852 3398 46892
rect 3398 46852 3423 46892
rect 3169 46829 3255 46852
rect 3337 46829 3423 46852
rect 18289 46892 18375 46915
rect 18457 46892 18543 46915
rect 18289 46852 18314 46892
rect 18314 46852 18354 46892
rect 18354 46852 18375 46892
rect 18457 46852 18478 46892
rect 18478 46852 18518 46892
rect 18518 46852 18543 46892
rect 18289 46829 18375 46852
rect 18457 46829 18543 46852
rect 33409 46892 33495 46915
rect 33577 46892 33663 46915
rect 33409 46852 33434 46892
rect 33434 46852 33474 46892
rect 33474 46852 33495 46892
rect 33577 46852 33598 46892
rect 33598 46852 33638 46892
rect 33638 46852 33663 46892
rect 33409 46829 33495 46852
rect 33577 46829 33663 46852
rect 48529 46892 48615 46915
rect 48697 46892 48783 46915
rect 48529 46852 48554 46892
rect 48554 46852 48594 46892
rect 48594 46852 48615 46892
rect 48697 46852 48718 46892
rect 48718 46852 48758 46892
rect 48758 46852 48783 46892
rect 48529 46829 48615 46852
rect 48697 46829 48783 46852
rect 63649 46892 63735 46915
rect 63817 46892 63903 46915
rect 63649 46852 63674 46892
rect 63674 46852 63714 46892
rect 63714 46852 63735 46892
rect 63817 46852 63838 46892
rect 63838 46852 63878 46892
rect 63878 46852 63903 46892
rect 63649 46829 63735 46852
rect 63817 46829 63903 46852
rect 78769 46892 78855 46915
rect 78937 46892 79023 46915
rect 78769 46852 78794 46892
rect 78794 46852 78834 46892
rect 78834 46852 78855 46892
rect 78937 46852 78958 46892
rect 78958 46852 78998 46892
rect 78998 46852 79023 46892
rect 78769 46829 78855 46852
rect 78937 46829 79023 46852
rect 93889 46892 93975 46915
rect 94057 46892 94143 46915
rect 93889 46852 93914 46892
rect 93914 46852 93954 46892
rect 93954 46852 93975 46892
rect 94057 46852 94078 46892
rect 94078 46852 94118 46892
rect 94118 46852 94143 46892
rect 93889 46829 93975 46852
rect 94057 46829 94143 46852
rect 4409 46136 4495 46159
rect 4577 46136 4663 46159
rect 4409 46096 4434 46136
rect 4434 46096 4474 46136
rect 4474 46096 4495 46136
rect 4577 46096 4598 46136
rect 4598 46096 4638 46136
rect 4638 46096 4663 46136
rect 4409 46073 4495 46096
rect 4577 46073 4663 46096
rect 19529 46136 19615 46159
rect 19697 46136 19783 46159
rect 19529 46096 19554 46136
rect 19554 46096 19594 46136
rect 19594 46096 19615 46136
rect 19697 46096 19718 46136
rect 19718 46096 19758 46136
rect 19758 46096 19783 46136
rect 19529 46073 19615 46096
rect 19697 46073 19783 46096
rect 34649 46136 34735 46159
rect 34817 46136 34903 46159
rect 34649 46096 34674 46136
rect 34674 46096 34714 46136
rect 34714 46096 34735 46136
rect 34817 46096 34838 46136
rect 34838 46096 34878 46136
rect 34878 46096 34903 46136
rect 34649 46073 34735 46096
rect 34817 46073 34903 46096
rect 49769 46136 49855 46159
rect 49937 46136 50023 46159
rect 49769 46096 49794 46136
rect 49794 46096 49834 46136
rect 49834 46096 49855 46136
rect 49937 46096 49958 46136
rect 49958 46096 49998 46136
rect 49998 46096 50023 46136
rect 49769 46073 49855 46096
rect 49937 46073 50023 46096
rect 64889 46136 64975 46159
rect 65057 46136 65143 46159
rect 64889 46096 64914 46136
rect 64914 46096 64954 46136
rect 64954 46096 64975 46136
rect 65057 46096 65078 46136
rect 65078 46096 65118 46136
rect 65118 46096 65143 46136
rect 64889 46073 64975 46096
rect 65057 46073 65143 46096
rect 80009 46136 80095 46159
rect 80177 46136 80263 46159
rect 80009 46096 80034 46136
rect 80034 46096 80074 46136
rect 80074 46096 80095 46136
rect 80177 46096 80198 46136
rect 80198 46096 80238 46136
rect 80238 46096 80263 46136
rect 80009 46073 80095 46096
rect 80177 46073 80263 46096
rect 95129 46136 95215 46159
rect 95297 46136 95383 46159
rect 95129 46096 95154 46136
rect 95154 46096 95194 46136
rect 95194 46096 95215 46136
rect 95297 46096 95318 46136
rect 95318 46096 95358 46136
rect 95358 46096 95383 46136
rect 95129 46073 95215 46096
rect 95297 46073 95383 46096
rect 3169 45380 3255 45403
rect 3337 45380 3423 45403
rect 3169 45340 3194 45380
rect 3194 45340 3234 45380
rect 3234 45340 3255 45380
rect 3337 45340 3358 45380
rect 3358 45340 3398 45380
rect 3398 45340 3423 45380
rect 3169 45317 3255 45340
rect 3337 45317 3423 45340
rect 18289 45380 18375 45403
rect 18457 45380 18543 45403
rect 18289 45340 18314 45380
rect 18314 45340 18354 45380
rect 18354 45340 18375 45380
rect 18457 45340 18478 45380
rect 18478 45340 18518 45380
rect 18518 45340 18543 45380
rect 18289 45317 18375 45340
rect 18457 45317 18543 45340
rect 33409 45380 33495 45403
rect 33577 45380 33663 45403
rect 33409 45340 33434 45380
rect 33434 45340 33474 45380
rect 33474 45340 33495 45380
rect 33577 45340 33598 45380
rect 33598 45340 33638 45380
rect 33638 45340 33663 45380
rect 33409 45317 33495 45340
rect 33577 45317 33663 45340
rect 48529 45380 48615 45403
rect 48697 45380 48783 45403
rect 48529 45340 48554 45380
rect 48554 45340 48594 45380
rect 48594 45340 48615 45380
rect 48697 45340 48718 45380
rect 48718 45340 48758 45380
rect 48758 45340 48783 45380
rect 48529 45317 48615 45340
rect 48697 45317 48783 45340
rect 63649 45380 63735 45403
rect 63817 45380 63903 45403
rect 63649 45340 63674 45380
rect 63674 45340 63714 45380
rect 63714 45340 63735 45380
rect 63817 45340 63838 45380
rect 63838 45340 63878 45380
rect 63878 45340 63903 45380
rect 63649 45317 63735 45340
rect 63817 45317 63903 45340
rect 78769 45380 78855 45403
rect 78937 45380 79023 45403
rect 78769 45340 78794 45380
rect 78794 45340 78834 45380
rect 78834 45340 78855 45380
rect 78937 45340 78958 45380
rect 78958 45340 78998 45380
rect 78998 45340 79023 45380
rect 78769 45317 78855 45340
rect 78937 45317 79023 45340
rect 93889 45380 93975 45403
rect 94057 45380 94143 45403
rect 93889 45340 93914 45380
rect 93914 45340 93954 45380
rect 93954 45340 93975 45380
rect 94057 45340 94078 45380
rect 94078 45340 94118 45380
rect 94118 45340 94143 45380
rect 93889 45317 93975 45340
rect 94057 45317 94143 45340
rect 4409 44624 4495 44647
rect 4577 44624 4663 44647
rect 4409 44584 4434 44624
rect 4434 44584 4474 44624
rect 4474 44584 4495 44624
rect 4577 44584 4598 44624
rect 4598 44584 4638 44624
rect 4638 44584 4663 44624
rect 4409 44561 4495 44584
rect 4577 44561 4663 44584
rect 19529 44624 19615 44647
rect 19697 44624 19783 44647
rect 19529 44584 19554 44624
rect 19554 44584 19594 44624
rect 19594 44584 19615 44624
rect 19697 44584 19718 44624
rect 19718 44584 19758 44624
rect 19758 44584 19783 44624
rect 19529 44561 19615 44584
rect 19697 44561 19783 44584
rect 34649 44624 34735 44647
rect 34817 44624 34903 44647
rect 34649 44584 34674 44624
rect 34674 44584 34714 44624
rect 34714 44584 34735 44624
rect 34817 44584 34838 44624
rect 34838 44584 34878 44624
rect 34878 44584 34903 44624
rect 34649 44561 34735 44584
rect 34817 44561 34903 44584
rect 49769 44624 49855 44647
rect 49937 44624 50023 44647
rect 49769 44584 49794 44624
rect 49794 44584 49834 44624
rect 49834 44584 49855 44624
rect 49937 44584 49958 44624
rect 49958 44584 49998 44624
rect 49998 44584 50023 44624
rect 49769 44561 49855 44584
rect 49937 44561 50023 44584
rect 64889 44624 64975 44647
rect 65057 44624 65143 44647
rect 64889 44584 64914 44624
rect 64914 44584 64954 44624
rect 64954 44584 64975 44624
rect 65057 44584 65078 44624
rect 65078 44584 65118 44624
rect 65118 44584 65143 44624
rect 64889 44561 64975 44584
rect 65057 44561 65143 44584
rect 80009 44624 80095 44647
rect 80177 44624 80263 44647
rect 80009 44584 80034 44624
rect 80034 44584 80074 44624
rect 80074 44584 80095 44624
rect 80177 44584 80198 44624
rect 80198 44584 80238 44624
rect 80238 44584 80263 44624
rect 80009 44561 80095 44584
rect 80177 44561 80263 44584
rect 95129 44624 95215 44647
rect 95297 44624 95383 44647
rect 95129 44584 95154 44624
rect 95154 44584 95194 44624
rect 95194 44584 95215 44624
rect 95297 44584 95318 44624
rect 95318 44584 95358 44624
rect 95358 44584 95383 44624
rect 95129 44561 95215 44584
rect 95297 44561 95383 44584
rect 3169 43868 3255 43891
rect 3337 43868 3423 43891
rect 3169 43828 3194 43868
rect 3194 43828 3234 43868
rect 3234 43828 3255 43868
rect 3337 43828 3358 43868
rect 3358 43828 3398 43868
rect 3398 43828 3423 43868
rect 3169 43805 3255 43828
rect 3337 43805 3423 43828
rect 18289 43868 18375 43891
rect 18457 43868 18543 43891
rect 18289 43828 18314 43868
rect 18314 43828 18354 43868
rect 18354 43828 18375 43868
rect 18457 43828 18478 43868
rect 18478 43828 18518 43868
rect 18518 43828 18543 43868
rect 18289 43805 18375 43828
rect 18457 43805 18543 43828
rect 33409 43868 33495 43891
rect 33577 43868 33663 43891
rect 33409 43828 33434 43868
rect 33434 43828 33474 43868
rect 33474 43828 33495 43868
rect 33577 43828 33598 43868
rect 33598 43828 33638 43868
rect 33638 43828 33663 43868
rect 33409 43805 33495 43828
rect 33577 43805 33663 43828
rect 48529 43868 48615 43891
rect 48697 43868 48783 43891
rect 48529 43828 48554 43868
rect 48554 43828 48594 43868
rect 48594 43828 48615 43868
rect 48697 43828 48718 43868
rect 48718 43828 48758 43868
rect 48758 43828 48783 43868
rect 48529 43805 48615 43828
rect 48697 43805 48783 43828
rect 63649 43868 63735 43891
rect 63817 43868 63903 43891
rect 63649 43828 63674 43868
rect 63674 43828 63714 43868
rect 63714 43828 63735 43868
rect 63817 43828 63838 43868
rect 63838 43828 63878 43868
rect 63878 43828 63903 43868
rect 63649 43805 63735 43828
rect 63817 43805 63903 43828
rect 78769 43868 78855 43891
rect 78937 43868 79023 43891
rect 78769 43828 78794 43868
rect 78794 43828 78834 43868
rect 78834 43828 78855 43868
rect 78937 43828 78958 43868
rect 78958 43828 78998 43868
rect 78998 43828 79023 43868
rect 78769 43805 78855 43828
rect 78937 43805 79023 43828
rect 93889 43868 93975 43891
rect 94057 43868 94143 43891
rect 93889 43828 93914 43868
rect 93914 43828 93954 43868
rect 93954 43828 93975 43868
rect 94057 43828 94078 43868
rect 94078 43828 94118 43868
rect 94118 43828 94143 43868
rect 93889 43805 93975 43828
rect 94057 43805 94143 43828
rect 4409 43112 4495 43135
rect 4577 43112 4663 43135
rect 4409 43072 4434 43112
rect 4434 43072 4474 43112
rect 4474 43072 4495 43112
rect 4577 43072 4598 43112
rect 4598 43072 4638 43112
rect 4638 43072 4663 43112
rect 4409 43049 4495 43072
rect 4577 43049 4663 43072
rect 19529 43112 19615 43135
rect 19697 43112 19783 43135
rect 19529 43072 19554 43112
rect 19554 43072 19594 43112
rect 19594 43072 19615 43112
rect 19697 43072 19718 43112
rect 19718 43072 19758 43112
rect 19758 43072 19783 43112
rect 19529 43049 19615 43072
rect 19697 43049 19783 43072
rect 34649 43112 34735 43135
rect 34817 43112 34903 43135
rect 34649 43072 34674 43112
rect 34674 43072 34714 43112
rect 34714 43072 34735 43112
rect 34817 43072 34838 43112
rect 34838 43072 34878 43112
rect 34878 43072 34903 43112
rect 34649 43049 34735 43072
rect 34817 43049 34903 43072
rect 49769 43112 49855 43135
rect 49937 43112 50023 43135
rect 49769 43072 49794 43112
rect 49794 43072 49834 43112
rect 49834 43072 49855 43112
rect 49937 43072 49958 43112
rect 49958 43072 49998 43112
rect 49998 43072 50023 43112
rect 49769 43049 49855 43072
rect 49937 43049 50023 43072
rect 64889 43112 64975 43135
rect 65057 43112 65143 43135
rect 64889 43072 64914 43112
rect 64914 43072 64954 43112
rect 64954 43072 64975 43112
rect 65057 43072 65078 43112
rect 65078 43072 65118 43112
rect 65118 43072 65143 43112
rect 64889 43049 64975 43072
rect 65057 43049 65143 43072
rect 80009 43112 80095 43135
rect 80177 43112 80263 43135
rect 80009 43072 80034 43112
rect 80034 43072 80074 43112
rect 80074 43072 80095 43112
rect 80177 43072 80198 43112
rect 80198 43072 80238 43112
rect 80238 43072 80263 43112
rect 80009 43049 80095 43072
rect 80177 43049 80263 43072
rect 95129 43112 95215 43135
rect 95297 43112 95383 43135
rect 95129 43072 95154 43112
rect 95154 43072 95194 43112
rect 95194 43072 95215 43112
rect 95297 43072 95318 43112
rect 95318 43072 95358 43112
rect 95358 43072 95383 43112
rect 95129 43049 95215 43072
rect 95297 43049 95383 43072
rect 3169 42356 3255 42379
rect 3337 42356 3423 42379
rect 3169 42316 3194 42356
rect 3194 42316 3234 42356
rect 3234 42316 3255 42356
rect 3337 42316 3358 42356
rect 3358 42316 3398 42356
rect 3398 42316 3423 42356
rect 3169 42293 3255 42316
rect 3337 42293 3423 42316
rect 18289 42356 18375 42379
rect 18457 42356 18543 42379
rect 18289 42316 18314 42356
rect 18314 42316 18354 42356
rect 18354 42316 18375 42356
rect 18457 42316 18478 42356
rect 18478 42316 18518 42356
rect 18518 42316 18543 42356
rect 18289 42293 18375 42316
rect 18457 42293 18543 42316
rect 33409 42356 33495 42379
rect 33577 42356 33663 42379
rect 33409 42316 33434 42356
rect 33434 42316 33474 42356
rect 33474 42316 33495 42356
rect 33577 42316 33598 42356
rect 33598 42316 33638 42356
rect 33638 42316 33663 42356
rect 33409 42293 33495 42316
rect 33577 42293 33663 42316
rect 48529 42356 48615 42379
rect 48697 42356 48783 42379
rect 48529 42316 48554 42356
rect 48554 42316 48594 42356
rect 48594 42316 48615 42356
rect 48697 42316 48718 42356
rect 48718 42316 48758 42356
rect 48758 42316 48783 42356
rect 48529 42293 48615 42316
rect 48697 42293 48783 42316
rect 63649 42356 63735 42379
rect 63817 42356 63903 42379
rect 63649 42316 63674 42356
rect 63674 42316 63714 42356
rect 63714 42316 63735 42356
rect 63817 42316 63838 42356
rect 63838 42316 63878 42356
rect 63878 42316 63903 42356
rect 63649 42293 63735 42316
rect 63817 42293 63903 42316
rect 78769 42356 78855 42379
rect 78937 42356 79023 42379
rect 78769 42316 78794 42356
rect 78794 42316 78834 42356
rect 78834 42316 78855 42356
rect 78937 42316 78958 42356
rect 78958 42316 78998 42356
rect 78998 42316 79023 42356
rect 78769 42293 78855 42316
rect 78937 42293 79023 42316
rect 93889 42356 93975 42379
rect 94057 42356 94143 42379
rect 93889 42316 93914 42356
rect 93914 42316 93954 42356
rect 93954 42316 93975 42356
rect 94057 42316 94078 42356
rect 94078 42316 94118 42356
rect 94118 42316 94143 42356
rect 93889 42293 93975 42316
rect 94057 42293 94143 42316
rect 4409 41600 4495 41623
rect 4577 41600 4663 41623
rect 4409 41560 4434 41600
rect 4434 41560 4474 41600
rect 4474 41560 4495 41600
rect 4577 41560 4598 41600
rect 4598 41560 4638 41600
rect 4638 41560 4663 41600
rect 4409 41537 4495 41560
rect 4577 41537 4663 41560
rect 19529 41600 19615 41623
rect 19697 41600 19783 41623
rect 19529 41560 19554 41600
rect 19554 41560 19594 41600
rect 19594 41560 19615 41600
rect 19697 41560 19718 41600
rect 19718 41560 19758 41600
rect 19758 41560 19783 41600
rect 19529 41537 19615 41560
rect 19697 41537 19783 41560
rect 34649 41600 34735 41623
rect 34817 41600 34903 41623
rect 34649 41560 34674 41600
rect 34674 41560 34714 41600
rect 34714 41560 34735 41600
rect 34817 41560 34838 41600
rect 34838 41560 34878 41600
rect 34878 41560 34903 41600
rect 34649 41537 34735 41560
rect 34817 41537 34903 41560
rect 49769 41600 49855 41623
rect 49937 41600 50023 41623
rect 49769 41560 49794 41600
rect 49794 41560 49834 41600
rect 49834 41560 49855 41600
rect 49937 41560 49958 41600
rect 49958 41560 49998 41600
rect 49998 41560 50023 41600
rect 49769 41537 49855 41560
rect 49937 41537 50023 41560
rect 64889 41600 64975 41623
rect 65057 41600 65143 41623
rect 64889 41560 64914 41600
rect 64914 41560 64954 41600
rect 64954 41560 64975 41600
rect 65057 41560 65078 41600
rect 65078 41560 65118 41600
rect 65118 41560 65143 41600
rect 64889 41537 64975 41560
rect 65057 41537 65143 41560
rect 80009 41600 80095 41623
rect 80177 41600 80263 41623
rect 80009 41560 80034 41600
rect 80034 41560 80074 41600
rect 80074 41560 80095 41600
rect 80177 41560 80198 41600
rect 80198 41560 80238 41600
rect 80238 41560 80263 41600
rect 80009 41537 80095 41560
rect 80177 41537 80263 41560
rect 95129 41600 95215 41623
rect 95297 41600 95383 41623
rect 95129 41560 95154 41600
rect 95154 41560 95194 41600
rect 95194 41560 95215 41600
rect 95297 41560 95318 41600
rect 95318 41560 95358 41600
rect 95358 41560 95383 41600
rect 95129 41537 95215 41560
rect 95297 41537 95383 41560
rect 3169 40844 3255 40867
rect 3337 40844 3423 40867
rect 3169 40804 3194 40844
rect 3194 40804 3234 40844
rect 3234 40804 3255 40844
rect 3337 40804 3358 40844
rect 3358 40804 3398 40844
rect 3398 40804 3423 40844
rect 3169 40781 3255 40804
rect 3337 40781 3423 40804
rect 18289 40844 18375 40867
rect 18457 40844 18543 40867
rect 18289 40804 18314 40844
rect 18314 40804 18354 40844
rect 18354 40804 18375 40844
rect 18457 40804 18478 40844
rect 18478 40804 18518 40844
rect 18518 40804 18543 40844
rect 18289 40781 18375 40804
rect 18457 40781 18543 40804
rect 33409 40844 33495 40867
rect 33577 40844 33663 40867
rect 33409 40804 33434 40844
rect 33434 40804 33474 40844
rect 33474 40804 33495 40844
rect 33577 40804 33598 40844
rect 33598 40804 33638 40844
rect 33638 40804 33663 40844
rect 33409 40781 33495 40804
rect 33577 40781 33663 40804
rect 48529 40844 48615 40867
rect 48697 40844 48783 40867
rect 48529 40804 48554 40844
rect 48554 40804 48594 40844
rect 48594 40804 48615 40844
rect 48697 40804 48718 40844
rect 48718 40804 48758 40844
rect 48758 40804 48783 40844
rect 48529 40781 48615 40804
rect 48697 40781 48783 40804
rect 63649 40844 63735 40867
rect 63817 40844 63903 40867
rect 63649 40804 63674 40844
rect 63674 40804 63714 40844
rect 63714 40804 63735 40844
rect 63817 40804 63838 40844
rect 63838 40804 63878 40844
rect 63878 40804 63903 40844
rect 63649 40781 63735 40804
rect 63817 40781 63903 40804
rect 78769 40844 78855 40867
rect 78937 40844 79023 40867
rect 78769 40804 78794 40844
rect 78794 40804 78834 40844
rect 78834 40804 78855 40844
rect 78937 40804 78958 40844
rect 78958 40804 78998 40844
rect 78998 40804 79023 40844
rect 78769 40781 78855 40804
rect 78937 40781 79023 40804
rect 93889 40844 93975 40867
rect 94057 40844 94143 40867
rect 93889 40804 93914 40844
rect 93914 40804 93954 40844
rect 93954 40804 93975 40844
rect 94057 40804 94078 40844
rect 94078 40804 94118 40844
rect 94118 40804 94143 40844
rect 93889 40781 93975 40804
rect 94057 40781 94143 40804
rect 4409 40088 4495 40111
rect 4577 40088 4663 40111
rect 4409 40048 4434 40088
rect 4434 40048 4474 40088
rect 4474 40048 4495 40088
rect 4577 40048 4598 40088
rect 4598 40048 4638 40088
rect 4638 40048 4663 40088
rect 4409 40025 4495 40048
rect 4577 40025 4663 40048
rect 19529 40088 19615 40111
rect 19697 40088 19783 40111
rect 19529 40048 19554 40088
rect 19554 40048 19594 40088
rect 19594 40048 19615 40088
rect 19697 40048 19718 40088
rect 19718 40048 19758 40088
rect 19758 40048 19783 40088
rect 19529 40025 19615 40048
rect 19697 40025 19783 40048
rect 34649 40088 34735 40111
rect 34817 40088 34903 40111
rect 34649 40048 34674 40088
rect 34674 40048 34714 40088
rect 34714 40048 34735 40088
rect 34817 40048 34838 40088
rect 34838 40048 34878 40088
rect 34878 40048 34903 40088
rect 34649 40025 34735 40048
rect 34817 40025 34903 40048
rect 49769 40088 49855 40111
rect 49937 40088 50023 40111
rect 49769 40048 49794 40088
rect 49794 40048 49834 40088
rect 49834 40048 49855 40088
rect 49937 40048 49958 40088
rect 49958 40048 49998 40088
rect 49998 40048 50023 40088
rect 49769 40025 49855 40048
rect 49937 40025 50023 40048
rect 64889 40088 64975 40111
rect 65057 40088 65143 40111
rect 64889 40048 64914 40088
rect 64914 40048 64954 40088
rect 64954 40048 64975 40088
rect 65057 40048 65078 40088
rect 65078 40048 65118 40088
rect 65118 40048 65143 40088
rect 64889 40025 64975 40048
rect 65057 40025 65143 40048
rect 80009 40088 80095 40111
rect 80177 40088 80263 40111
rect 80009 40048 80034 40088
rect 80034 40048 80074 40088
rect 80074 40048 80095 40088
rect 80177 40048 80198 40088
rect 80198 40048 80238 40088
rect 80238 40048 80263 40088
rect 80009 40025 80095 40048
rect 80177 40025 80263 40048
rect 95129 40088 95215 40111
rect 95297 40088 95383 40111
rect 95129 40048 95154 40088
rect 95154 40048 95194 40088
rect 95194 40048 95215 40088
rect 95297 40048 95318 40088
rect 95318 40048 95358 40088
rect 95358 40048 95383 40088
rect 95129 40025 95215 40048
rect 95297 40025 95383 40048
rect 3169 39332 3255 39355
rect 3337 39332 3423 39355
rect 3169 39292 3194 39332
rect 3194 39292 3234 39332
rect 3234 39292 3255 39332
rect 3337 39292 3358 39332
rect 3358 39292 3398 39332
rect 3398 39292 3423 39332
rect 3169 39269 3255 39292
rect 3337 39269 3423 39292
rect 18289 39332 18375 39355
rect 18457 39332 18543 39355
rect 18289 39292 18314 39332
rect 18314 39292 18354 39332
rect 18354 39292 18375 39332
rect 18457 39292 18478 39332
rect 18478 39292 18518 39332
rect 18518 39292 18543 39332
rect 18289 39269 18375 39292
rect 18457 39269 18543 39292
rect 33409 39332 33495 39355
rect 33577 39332 33663 39355
rect 33409 39292 33434 39332
rect 33434 39292 33474 39332
rect 33474 39292 33495 39332
rect 33577 39292 33598 39332
rect 33598 39292 33638 39332
rect 33638 39292 33663 39332
rect 33409 39269 33495 39292
rect 33577 39269 33663 39292
rect 48529 39332 48615 39355
rect 48697 39332 48783 39355
rect 48529 39292 48554 39332
rect 48554 39292 48594 39332
rect 48594 39292 48615 39332
rect 48697 39292 48718 39332
rect 48718 39292 48758 39332
rect 48758 39292 48783 39332
rect 48529 39269 48615 39292
rect 48697 39269 48783 39292
rect 63649 39332 63735 39355
rect 63817 39332 63903 39355
rect 63649 39292 63674 39332
rect 63674 39292 63714 39332
rect 63714 39292 63735 39332
rect 63817 39292 63838 39332
rect 63838 39292 63878 39332
rect 63878 39292 63903 39332
rect 63649 39269 63735 39292
rect 63817 39269 63903 39292
rect 78769 39332 78855 39355
rect 78937 39332 79023 39355
rect 78769 39292 78794 39332
rect 78794 39292 78834 39332
rect 78834 39292 78855 39332
rect 78937 39292 78958 39332
rect 78958 39292 78998 39332
rect 78998 39292 79023 39332
rect 78769 39269 78855 39292
rect 78937 39269 79023 39292
rect 93889 39332 93975 39355
rect 94057 39332 94143 39355
rect 93889 39292 93914 39332
rect 93914 39292 93954 39332
rect 93954 39292 93975 39332
rect 94057 39292 94078 39332
rect 94078 39292 94118 39332
rect 94118 39292 94143 39332
rect 93889 39269 93975 39292
rect 94057 39269 94143 39292
rect 4409 38576 4495 38599
rect 4577 38576 4663 38599
rect 4409 38536 4434 38576
rect 4434 38536 4474 38576
rect 4474 38536 4495 38576
rect 4577 38536 4598 38576
rect 4598 38536 4638 38576
rect 4638 38536 4663 38576
rect 4409 38513 4495 38536
rect 4577 38513 4663 38536
rect 19529 38576 19615 38599
rect 19697 38576 19783 38599
rect 19529 38536 19554 38576
rect 19554 38536 19594 38576
rect 19594 38536 19615 38576
rect 19697 38536 19718 38576
rect 19718 38536 19758 38576
rect 19758 38536 19783 38576
rect 19529 38513 19615 38536
rect 19697 38513 19783 38536
rect 34649 38576 34735 38599
rect 34817 38576 34903 38599
rect 34649 38536 34674 38576
rect 34674 38536 34714 38576
rect 34714 38536 34735 38576
rect 34817 38536 34838 38576
rect 34838 38536 34878 38576
rect 34878 38536 34903 38576
rect 34649 38513 34735 38536
rect 34817 38513 34903 38536
rect 49769 38576 49855 38599
rect 49937 38576 50023 38599
rect 49769 38536 49794 38576
rect 49794 38536 49834 38576
rect 49834 38536 49855 38576
rect 49937 38536 49958 38576
rect 49958 38536 49998 38576
rect 49998 38536 50023 38576
rect 49769 38513 49855 38536
rect 49937 38513 50023 38536
rect 64889 38576 64975 38599
rect 65057 38576 65143 38599
rect 64889 38536 64914 38576
rect 64914 38536 64954 38576
rect 64954 38536 64975 38576
rect 65057 38536 65078 38576
rect 65078 38536 65118 38576
rect 65118 38536 65143 38576
rect 64889 38513 64975 38536
rect 65057 38513 65143 38536
rect 80009 38576 80095 38599
rect 80177 38576 80263 38599
rect 80009 38536 80034 38576
rect 80034 38536 80074 38576
rect 80074 38536 80095 38576
rect 80177 38536 80198 38576
rect 80198 38536 80238 38576
rect 80238 38536 80263 38576
rect 80009 38513 80095 38536
rect 80177 38513 80263 38536
rect 95129 38576 95215 38599
rect 95297 38576 95383 38599
rect 95129 38536 95154 38576
rect 95154 38536 95194 38576
rect 95194 38536 95215 38576
rect 95297 38536 95318 38576
rect 95318 38536 95358 38576
rect 95358 38536 95383 38576
rect 95129 38513 95215 38536
rect 95297 38513 95383 38536
rect 3169 37820 3255 37843
rect 3337 37820 3423 37843
rect 3169 37780 3194 37820
rect 3194 37780 3234 37820
rect 3234 37780 3255 37820
rect 3337 37780 3358 37820
rect 3358 37780 3398 37820
rect 3398 37780 3423 37820
rect 3169 37757 3255 37780
rect 3337 37757 3423 37780
rect 18289 37820 18375 37843
rect 18457 37820 18543 37843
rect 18289 37780 18314 37820
rect 18314 37780 18354 37820
rect 18354 37780 18375 37820
rect 18457 37780 18478 37820
rect 18478 37780 18518 37820
rect 18518 37780 18543 37820
rect 18289 37757 18375 37780
rect 18457 37757 18543 37780
rect 33409 37820 33495 37843
rect 33577 37820 33663 37843
rect 33409 37780 33434 37820
rect 33434 37780 33474 37820
rect 33474 37780 33495 37820
rect 33577 37780 33598 37820
rect 33598 37780 33638 37820
rect 33638 37780 33663 37820
rect 33409 37757 33495 37780
rect 33577 37757 33663 37780
rect 48529 37820 48615 37843
rect 48697 37820 48783 37843
rect 48529 37780 48554 37820
rect 48554 37780 48594 37820
rect 48594 37780 48615 37820
rect 48697 37780 48718 37820
rect 48718 37780 48758 37820
rect 48758 37780 48783 37820
rect 48529 37757 48615 37780
rect 48697 37757 48783 37780
rect 63649 37820 63735 37843
rect 63817 37820 63903 37843
rect 63649 37780 63674 37820
rect 63674 37780 63714 37820
rect 63714 37780 63735 37820
rect 63817 37780 63838 37820
rect 63838 37780 63878 37820
rect 63878 37780 63903 37820
rect 63649 37757 63735 37780
rect 63817 37757 63903 37780
rect 78769 37820 78855 37843
rect 78937 37820 79023 37843
rect 78769 37780 78794 37820
rect 78794 37780 78834 37820
rect 78834 37780 78855 37820
rect 78937 37780 78958 37820
rect 78958 37780 78998 37820
rect 78998 37780 79023 37820
rect 78769 37757 78855 37780
rect 78937 37757 79023 37780
rect 93889 37820 93975 37843
rect 94057 37820 94143 37843
rect 93889 37780 93914 37820
rect 93914 37780 93954 37820
rect 93954 37780 93975 37820
rect 94057 37780 94078 37820
rect 94078 37780 94118 37820
rect 94118 37780 94143 37820
rect 93889 37757 93975 37780
rect 94057 37757 94143 37780
rect 4409 37064 4495 37087
rect 4577 37064 4663 37087
rect 4409 37024 4434 37064
rect 4434 37024 4474 37064
rect 4474 37024 4495 37064
rect 4577 37024 4598 37064
rect 4598 37024 4638 37064
rect 4638 37024 4663 37064
rect 4409 37001 4495 37024
rect 4577 37001 4663 37024
rect 19529 37064 19615 37087
rect 19697 37064 19783 37087
rect 19529 37024 19554 37064
rect 19554 37024 19594 37064
rect 19594 37024 19615 37064
rect 19697 37024 19718 37064
rect 19718 37024 19758 37064
rect 19758 37024 19783 37064
rect 19529 37001 19615 37024
rect 19697 37001 19783 37024
rect 34649 37064 34735 37087
rect 34817 37064 34903 37087
rect 34649 37024 34674 37064
rect 34674 37024 34714 37064
rect 34714 37024 34735 37064
rect 34817 37024 34838 37064
rect 34838 37024 34878 37064
rect 34878 37024 34903 37064
rect 34649 37001 34735 37024
rect 34817 37001 34903 37024
rect 49769 37064 49855 37087
rect 49937 37064 50023 37087
rect 49769 37024 49794 37064
rect 49794 37024 49834 37064
rect 49834 37024 49855 37064
rect 49937 37024 49958 37064
rect 49958 37024 49998 37064
rect 49998 37024 50023 37064
rect 49769 37001 49855 37024
rect 49937 37001 50023 37024
rect 64889 37064 64975 37087
rect 65057 37064 65143 37087
rect 64889 37024 64914 37064
rect 64914 37024 64954 37064
rect 64954 37024 64975 37064
rect 65057 37024 65078 37064
rect 65078 37024 65118 37064
rect 65118 37024 65143 37064
rect 64889 37001 64975 37024
rect 65057 37001 65143 37024
rect 80009 37064 80095 37087
rect 80177 37064 80263 37087
rect 80009 37024 80034 37064
rect 80034 37024 80074 37064
rect 80074 37024 80095 37064
rect 80177 37024 80198 37064
rect 80198 37024 80238 37064
rect 80238 37024 80263 37064
rect 80009 37001 80095 37024
rect 80177 37001 80263 37024
rect 95129 37064 95215 37087
rect 95297 37064 95383 37087
rect 95129 37024 95154 37064
rect 95154 37024 95194 37064
rect 95194 37024 95215 37064
rect 95297 37024 95318 37064
rect 95318 37024 95358 37064
rect 95358 37024 95383 37064
rect 95129 37001 95215 37024
rect 95297 37001 95383 37024
rect 3169 36308 3255 36331
rect 3337 36308 3423 36331
rect 3169 36268 3194 36308
rect 3194 36268 3234 36308
rect 3234 36268 3255 36308
rect 3337 36268 3358 36308
rect 3358 36268 3398 36308
rect 3398 36268 3423 36308
rect 3169 36245 3255 36268
rect 3337 36245 3423 36268
rect 18289 36308 18375 36331
rect 18457 36308 18543 36331
rect 18289 36268 18314 36308
rect 18314 36268 18354 36308
rect 18354 36268 18375 36308
rect 18457 36268 18478 36308
rect 18478 36268 18518 36308
rect 18518 36268 18543 36308
rect 18289 36245 18375 36268
rect 18457 36245 18543 36268
rect 33409 36308 33495 36331
rect 33577 36308 33663 36331
rect 33409 36268 33434 36308
rect 33434 36268 33474 36308
rect 33474 36268 33495 36308
rect 33577 36268 33598 36308
rect 33598 36268 33638 36308
rect 33638 36268 33663 36308
rect 33409 36245 33495 36268
rect 33577 36245 33663 36268
rect 48529 36308 48615 36331
rect 48697 36308 48783 36331
rect 48529 36268 48554 36308
rect 48554 36268 48594 36308
rect 48594 36268 48615 36308
rect 48697 36268 48718 36308
rect 48718 36268 48758 36308
rect 48758 36268 48783 36308
rect 48529 36245 48615 36268
rect 48697 36245 48783 36268
rect 63649 36308 63735 36331
rect 63817 36308 63903 36331
rect 63649 36268 63674 36308
rect 63674 36268 63714 36308
rect 63714 36268 63735 36308
rect 63817 36268 63838 36308
rect 63838 36268 63878 36308
rect 63878 36268 63903 36308
rect 63649 36245 63735 36268
rect 63817 36245 63903 36268
rect 78769 36308 78855 36331
rect 78937 36308 79023 36331
rect 78769 36268 78794 36308
rect 78794 36268 78834 36308
rect 78834 36268 78855 36308
rect 78937 36268 78958 36308
rect 78958 36268 78998 36308
rect 78998 36268 79023 36308
rect 78769 36245 78855 36268
rect 78937 36245 79023 36268
rect 93889 36308 93975 36331
rect 94057 36308 94143 36331
rect 93889 36268 93914 36308
rect 93914 36268 93954 36308
rect 93954 36268 93975 36308
rect 94057 36268 94078 36308
rect 94078 36268 94118 36308
rect 94118 36268 94143 36308
rect 93889 36245 93975 36268
rect 94057 36245 94143 36268
rect 4409 35552 4495 35575
rect 4577 35552 4663 35575
rect 4409 35512 4434 35552
rect 4434 35512 4474 35552
rect 4474 35512 4495 35552
rect 4577 35512 4598 35552
rect 4598 35512 4638 35552
rect 4638 35512 4663 35552
rect 4409 35489 4495 35512
rect 4577 35489 4663 35512
rect 19529 35552 19615 35575
rect 19697 35552 19783 35575
rect 19529 35512 19554 35552
rect 19554 35512 19594 35552
rect 19594 35512 19615 35552
rect 19697 35512 19718 35552
rect 19718 35512 19758 35552
rect 19758 35512 19783 35552
rect 19529 35489 19615 35512
rect 19697 35489 19783 35512
rect 34649 35552 34735 35575
rect 34817 35552 34903 35575
rect 34649 35512 34674 35552
rect 34674 35512 34714 35552
rect 34714 35512 34735 35552
rect 34817 35512 34838 35552
rect 34838 35512 34878 35552
rect 34878 35512 34903 35552
rect 34649 35489 34735 35512
rect 34817 35489 34903 35512
rect 49769 35552 49855 35575
rect 49937 35552 50023 35575
rect 49769 35512 49794 35552
rect 49794 35512 49834 35552
rect 49834 35512 49855 35552
rect 49937 35512 49958 35552
rect 49958 35512 49998 35552
rect 49998 35512 50023 35552
rect 49769 35489 49855 35512
rect 49937 35489 50023 35512
rect 64889 35552 64975 35575
rect 65057 35552 65143 35575
rect 64889 35512 64914 35552
rect 64914 35512 64954 35552
rect 64954 35512 64975 35552
rect 65057 35512 65078 35552
rect 65078 35512 65118 35552
rect 65118 35512 65143 35552
rect 64889 35489 64975 35512
rect 65057 35489 65143 35512
rect 80009 35552 80095 35575
rect 80177 35552 80263 35575
rect 80009 35512 80034 35552
rect 80034 35512 80074 35552
rect 80074 35512 80095 35552
rect 80177 35512 80198 35552
rect 80198 35512 80238 35552
rect 80238 35512 80263 35552
rect 80009 35489 80095 35512
rect 80177 35489 80263 35512
rect 95129 35552 95215 35575
rect 95297 35552 95383 35575
rect 95129 35512 95154 35552
rect 95154 35512 95194 35552
rect 95194 35512 95215 35552
rect 95297 35512 95318 35552
rect 95318 35512 95358 35552
rect 95358 35512 95383 35552
rect 95129 35489 95215 35512
rect 95297 35489 95383 35512
rect 3169 34796 3255 34819
rect 3337 34796 3423 34819
rect 3169 34756 3194 34796
rect 3194 34756 3234 34796
rect 3234 34756 3255 34796
rect 3337 34756 3358 34796
rect 3358 34756 3398 34796
rect 3398 34756 3423 34796
rect 3169 34733 3255 34756
rect 3337 34733 3423 34756
rect 18289 34796 18375 34819
rect 18457 34796 18543 34819
rect 18289 34756 18314 34796
rect 18314 34756 18354 34796
rect 18354 34756 18375 34796
rect 18457 34756 18478 34796
rect 18478 34756 18518 34796
rect 18518 34756 18543 34796
rect 18289 34733 18375 34756
rect 18457 34733 18543 34756
rect 33409 34796 33495 34819
rect 33577 34796 33663 34819
rect 33409 34756 33434 34796
rect 33434 34756 33474 34796
rect 33474 34756 33495 34796
rect 33577 34756 33598 34796
rect 33598 34756 33638 34796
rect 33638 34756 33663 34796
rect 33409 34733 33495 34756
rect 33577 34733 33663 34756
rect 48529 34796 48615 34819
rect 48697 34796 48783 34819
rect 48529 34756 48554 34796
rect 48554 34756 48594 34796
rect 48594 34756 48615 34796
rect 48697 34756 48718 34796
rect 48718 34756 48758 34796
rect 48758 34756 48783 34796
rect 48529 34733 48615 34756
rect 48697 34733 48783 34756
rect 63649 34796 63735 34819
rect 63817 34796 63903 34819
rect 63649 34756 63674 34796
rect 63674 34756 63714 34796
rect 63714 34756 63735 34796
rect 63817 34756 63838 34796
rect 63838 34756 63878 34796
rect 63878 34756 63903 34796
rect 63649 34733 63735 34756
rect 63817 34733 63903 34756
rect 78769 34796 78855 34819
rect 78937 34796 79023 34819
rect 78769 34756 78794 34796
rect 78794 34756 78834 34796
rect 78834 34756 78855 34796
rect 78937 34756 78958 34796
rect 78958 34756 78998 34796
rect 78998 34756 79023 34796
rect 78769 34733 78855 34756
rect 78937 34733 79023 34756
rect 93889 34796 93975 34819
rect 94057 34796 94143 34819
rect 93889 34756 93914 34796
rect 93914 34756 93954 34796
rect 93954 34756 93975 34796
rect 94057 34756 94078 34796
rect 94078 34756 94118 34796
rect 94118 34756 94143 34796
rect 93889 34733 93975 34756
rect 94057 34733 94143 34756
rect 4409 34040 4495 34063
rect 4577 34040 4663 34063
rect 4409 34000 4434 34040
rect 4434 34000 4474 34040
rect 4474 34000 4495 34040
rect 4577 34000 4598 34040
rect 4598 34000 4638 34040
rect 4638 34000 4663 34040
rect 4409 33977 4495 34000
rect 4577 33977 4663 34000
rect 19529 34040 19615 34063
rect 19697 34040 19783 34063
rect 19529 34000 19554 34040
rect 19554 34000 19594 34040
rect 19594 34000 19615 34040
rect 19697 34000 19718 34040
rect 19718 34000 19758 34040
rect 19758 34000 19783 34040
rect 19529 33977 19615 34000
rect 19697 33977 19783 34000
rect 34649 34040 34735 34063
rect 34817 34040 34903 34063
rect 34649 34000 34674 34040
rect 34674 34000 34714 34040
rect 34714 34000 34735 34040
rect 34817 34000 34838 34040
rect 34838 34000 34878 34040
rect 34878 34000 34903 34040
rect 34649 33977 34735 34000
rect 34817 33977 34903 34000
rect 49769 34040 49855 34063
rect 49937 34040 50023 34063
rect 49769 34000 49794 34040
rect 49794 34000 49834 34040
rect 49834 34000 49855 34040
rect 49937 34000 49958 34040
rect 49958 34000 49998 34040
rect 49998 34000 50023 34040
rect 49769 33977 49855 34000
rect 49937 33977 50023 34000
rect 64889 34040 64975 34063
rect 65057 34040 65143 34063
rect 64889 34000 64914 34040
rect 64914 34000 64954 34040
rect 64954 34000 64975 34040
rect 65057 34000 65078 34040
rect 65078 34000 65118 34040
rect 65118 34000 65143 34040
rect 64889 33977 64975 34000
rect 65057 33977 65143 34000
rect 80009 34040 80095 34063
rect 80177 34040 80263 34063
rect 80009 34000 80034 34040
rect 80034 34000 80074 34040
rect 80074 34000 80095 34040
rect 80177 34000 80198 34040
rect 80198 34000 80238 34040
rect 80238 34000 80263 34040
rect 80009 33977 80095 34000
rect 80177 33977 80263 34000
rect 95129 34040 95215 34063
rect 95297 34040 95383 34063
rect 95129 34000 95154 34040
rect 95154 34000 95194 34040
rect 95194 34000 95215 34040
rect 95297 34000 95318 34040
rect 95318 34000 95358 34040
rect 95358 34000 95383 34040
rect 95129 33977 95215 34000
rect 95297 33977 95383 34000
rect 3169 33284 3255 33307
rect 3337 33284 3423 33307
rect 3169 33244 3194 33284
rect 3194 33244 3234 33284
rect 3234 33244 3255 33284
rect 3337 33244 3358 33284
rect 3358 33244 3398 33284
rect 3398 33244 3423 33284
rect 3169 33221 3255 33244
rect 3337 33221 3423 33244
rect 18289 33284 18375 33307
rect 18457 33284 18543 33307
rect 18289 33244 18314 33284
rect 18314 33244 18354 33284
rect 18354 33244 18375 33284
rect 18457 33244 18478 33284
rect 18478 33244 18518 33284
rect 18518 33244 18543 33284
rect 18289 33221 18375 33244
rect 18457 33221 18543 33244
rect 33409 33284 33495 33307
rect 33577 33284 33663 33307
rect 33409 33244 33434 33284
rect 33434 33244 33474 33284
rect 33474 33244 33495 33284
rect 33577 33244 33598 33284
rect 33598 33244 33638 33284
rect 33638 33244 33663 33284
rect 33409 33221 33495 33244
rect 33577 33221 33663 33244
rect 48529 33284 48615 33307
rect 48697 33284 48783 33307
rect 48529 33244 48554 33284
rect 48554 33244 48594 33284
rect 48594 33244 48615 33284
rect 48697 33244 48718 33284
rect 48718 33244 48758 33284
rect 48758 33244 48783 33284
rect 48529 33221 48615 33244
rect 48697 33221 48783 33244
rect 63649 33284 63735 33307
rect 63817 33284 63903 33307
rect 63649 33244 63674 33284
rect 63674 33244 63714 33284
rect 63714 33244 63735 33284
rect 63817 33244 63838 33284
rect 63838 33244 63878 33284
rect 63878 33244 63903 33284
rect 63649 33221 63735 33244
rect 63817 33221 63903 33244
rect 78769 33284 78855 33307
rect 78937 33284 79023 33307
rect 78769 33244 78794 33284
rect 78794 33244 78834 33284
rect 78834 33244 78855 33284
rect 78937 33244 78958 33284
rect 78958 33244 78998 33284
rect 78998 33244 79023 33284
rect 78769 33221 78855 33244
rect 78937 33221 79023 33244
rect 93889 33284 93975 33307
rect 94057 33284 94143 33307
rect 93889 33244 93914 33284
rect 93914 33244 93954 33284
rect 93954 33244 93975 33284
rect 94057 33244 94078 33284
rect 94078 33244 94118 33284
rect 94118 33244 94143 33284
rect 93889 33221 93975 33244
rect 94057 33221 94143 33244
rect 4409 32528 4495 32551
rect 4577 32528 4663 32551
rect 4409 32488 4434 32528
rect 4434 32488 4474 32528
rect 4474 32488 4495 32528
rect 4577 32488 4598 32528
rect 4598 32488 4638 32528
rect 4638 32488 4663 32528
rect 4409 32465 4495 32488
rect 4577 32465 4663 32488
rect 19529 32528 19615 32551
rect 19697 32528 19783 32551
rect 19529 32488 19554 32528
rect 19554 32488 19594 32528
rect 19594 32488 19615 32528
rect 19697 32488 19718 32528
rect 19718 32488 19758 32528
rect 19758 32488 19783 32528
rect 19529 32465 19615 32488
rect 19697 32465 19783 32488
rect 34649 32528 34735 32551
rect 34817 32528 34903 32551
rect 34649 32488 34674 32528
rect 34674 32488 34714 32528
rect 34714 32488 34735 32528
rect 34817 32488 34838 32528
rect 34838 32488 34878 32528
rect 34878 32488 34903 32528
rect 34649 32465 34735 32488
rect 34817 32465 34903 32488
rect 49769 32528 49855 32551
rect 49937 32528 50023 32551
rect 49769 32488 49794 32528
rect 49794 32488 49834 32528
rect 49834 32488 49855 32528
rect 49937 32488 49958 32528
rect 49958 32488 49998 32528
rect 49998 32488 50023 32528
rect 49769 32465 49855 32488
rect 49937 32465 50023 32488
rect 64889 32528 64975 32551
rect 65057 32528 65143 32551
rect 64889 32488 64914 32528
rect 64914 32488 64954 32528
rect 64954 32488 64975 32528
rect 65057 32488 65078 32528
rect 65078 32488 65118 32528
rect 65118 32488 65143 32528
rect 64889 32465 64975 32488
rect 65057 32465 65143 32488
rect 80009 32528 80095 32551
rect 80177 32528 80263 32551
rect 80009 32488 80034 32528
rect 80034 32488 80074 32528
rect 80074 32488 80095 32528
rect 80177 32488 80198 32528
rect 80198 32488 80238 32528
rect 80238 32488 80263 32528
rect 80009 32465 80095 32488
rect 80177 32465 80263 32488
rect 95129 32528 95215 32551
rect 95297 32528 95383 32551
rect 95129 32488 95154 32528
rect 95154 32488 95194 32528
rect 95194 32488 95215 32528
rect 95297 32488 95318 32528
rect 95318 32488 95358 32528
rect 95358 32488 95383 32528
rect 95129 32465 95215 32488
rect 95297 32465 95383 32488
rect 3169 31772 3255 31795
rect 3337 31772 3423 31795
rect 3169 31732 3194 31772
rect 3194 31732 3234 31772
rect 3234 31732 3255 31772
rect 3337 31732 3358 31772
rect 3358 31732 3398 31772
rect 3398 31732 3423 31772
rect 3169 31709 3255 31732
rect 3337 31709 3423 31732
rect 18289 31772 18375 31795
rect 18457 31772 18543 31795
rect 18289 31732 18314 31772
rect 18314 31732 18354 31772
rect 18354 31732 18375 31772
rect 18457 31732 18478 31772
rect 18478 31732 18518 31772
rect 18518 31732 18543 31772
rect 18289 31709 18375 31732
rect 18457 31709 18543 31732
rect 33409 31772 33495 31795
rect 33577 31772 33663 31795
rect 33409 31732 33434 31772
rect 33434 31732 33474 31772
rect 33474 31732 33495 31772
rect 33577 31732 33598 31772
rect 33598 31732 33638 31772
rect 33638 31732 33663 31772
rect 33409 31709 33495 31732
rect 33577 31709 33663 31732
rect 48529 31772 48615 31795
rect 48697 31772 48783 31795
rect 48529 31732 48554 31772
rect 48554 31732 48594 31772
rect 48594 31732 48615 31772
rect 48697 31732 48718 31772
rect 48718 31732 48758 31772
rect 48758 31732 48783 31772
rect 48529 31709 48615 31732
rect 48697 31709 48783 31732
rect 63649 31772 63735 31795
rect 63817 31772 63903 31795
rect 63649 31732 63674 31772
rect 63674 31732 63714 31772
rect 63714 31732 63735 31772
rect 63817 31732 63838 31772
rect 63838 31732 63878 31772
rect 63878 31732 63903 31772
rect 63649 31709 63735 31732
rect 63817 31709 63903 31732
rect 78769 31772 78855 31795
rect 78937 31772 79023 31795
rect 78769 31732 78794 31772
rect 78794 31732 78834 31772
rect 78834 31732 78855 31772
rect 78937 31732 78958 31772
rect 78958 31732 78998 31772
rect 78998 31732 79023 31772
rect 78769 31709 78855 31732
rect 78937 31709 79023 31732
rect 93889 31772 93975 31795
rect 94057 31772 94143 31795
rect 93889 31732 93914 31772
rect 93914 31732 93954 31772
rect 93954 31732 93975 31772
rect 94057 31732 94078 31772
rect 94078 31732 94118 31772
rect 94118 31732 94143 31772
rect 93889 31709 93975 31732
rect 94057 31709 94143 31732
rect 4409 31016 4495 31039
rect 4577 31016 4663 31039
rect 4409 30976 4434 31016
rect 4434 30976 4474 31016
rect 4474 30976 4495 31016
rect 4577 30976 4598 31016
rect 4598 30976 4638 31016
rect 4638 30976 4663 31016
rect 4409 30953 4495 30976
rect 4577 30953 4663 30976
rect 19529 31016 19615 31039
rect 19697 31016 19783 31039
rect 19529 30976 19554 31016
rect 19554 30976 19594 31016
rect 19594 30976 19615 31016
rect 19697 30976 19718 31016
rect 19718 30976 19758 31016
rect 19758 30976 19783 31016
rect 19529 30953 19615 30976
rect 19697 30953 19783 30976
rect 34649 31016 34735 31039
rect 34817 31016 34903 31039
rect 34649 30976 34674 31016
rect 34674 30976 34714 31016
rect 34714 30976 34735 31016
rect 34817 30976 34838 31016
rect 34838 30976 34878 31016
rect 34878 30976 34903 31016
rect 34649 30953 34735 30976
rect 34817 30953 34903 30976
rect 49769 31016 49855 31039
rect 49937 31016 50023 31039
rect 49769 30976 49794 31016
rect 49794 30976 49834 31016
rect 49834 30976 49855 31016
rect 49937 30976 49958 31016
rect 49958 30976 49998 31016
rect 49998 30976 50023 31016
rect 49769 30953 49855 30976
rect 49937 30953 50023 30976
rect 64889 31016 64975 31039
rect 65057 31016 65143 31039
rect 64889 30976 64914 31016
rect 64914 30976 64954 31016
rect 64954 30976 64975 31016
rect 65057 30976 65078 31016
rect 65078 30976 65118 31016
rect 65118 30976 65143 31016
rect 64889 30953 64975 30976
rect 65057 30953 65143 30976
rect 80009 31016 80095 31039
rect 80177 31016 80263 31039
rect 80009 30976 80034 31016
rect 80034 30976 80074 31016
rect 80074 30976 80095 31016
rect 80177 30976 80198 31016
rect 80198 30976 80238 31016
rect 80238 30976 80263 31016
rect 80009 30953 80095 30976
rect 80177 30953 80263 30976
rect 95129 31016 95215 31039
rect 95297 31016 95383 31039
rect 95129 30976 95154 31016
rect 95154 30976 95194 31016
rect 95194 30976 95215 31016
rect 95297 30976 95318 31016
rect 95318 30976 95358 31016
rect 95358 30976 95383 31016
rect 95129 30953 95215 30976
rect 95297 30953 95383 30976
rect 3169 30260 3255 30283
rect 3337 30260 3423 30283
rect 3169 30220 3194 30260
rect 3194 30220 3234 30260
rect 3234 30220 3255 30260
rect 3337 30220 3358 30260
rect 3358 30220 3398 30260
rect 3398 30220 3423 30260
rect 3169 30197 3255 30220
rect 3337 30197 3423 30220
rect 18289 30260 18375 30283
rect 18457 30260 18543 30283
rect 18289 30220 18314 30260
rect 18314 30220 18354 30260
rect 18354 30220 18375 30260
rect 18457 30220 18478 30260
rect 18478 30220 18518 30260
rect 18518 30220 18543 30260
rect 18289 30197 18375 30220
rect 18457 30197 18543 30220
rect 33409 30260 33495 30283
rect 33577 30260 33663 30283
rect 33409 30220 33434 30260
rect 33434 30220 33474 30260
rect 33474 30220 33495 30260
rect 33577 30220 33598 30260
rect 33598 30220 33638 30260
rect 33638 30220 33663 30260
rect 33409 30197 33495 30220
rect 33577 30197 33663 30220
rect 48529 30260 48615 30283
rect 48697 30260 48783 30283
rect 48529 30220 48554 30260
rect 48554 30220 48594 30260
rect 48594 30220 48615 30260
rect 48697 30220 48718 30260
rect 48718 30220 48758 30260
rect 48758 30220 48783 30260
rect 48529 30197 48615 30220
rect 48697 30197 48783 30220
rect 63649 30260 63735 30283
rect 63817 30260 63903 30283
rect 63649 30220 63674 30260
rect 63674 30220 63714 30260
rect 63714 30220 63735 30260
rect 63817 30220 63838 30260
rect 63838 30220 63878 30260
rect 63878 30220 63903 30260
rect 63649 30197 63735 30220
rect 63817 30197 63903 30220
rect 78769 30260 78855 30283
rect 78937 30260 79023 30283
rect 78769 30220 78794 30260
rect 78794 30220 78834 30260
rect 78834 30220 78855 30260
rect 78937 30220 78958 30260
rect 78958 30220 78998 30260
rect 78998 30220 79023 30260
rect 78769 30197 78855 30220
rect 78937 30197 79023 30220
rect 93889 30260 93975 30283
rect 94057 30260 94143 30283
rect 93889 30220 93914 30260
rect 93914 30220 93954 30260
rect 93954 30220 93975 30260
rect 94057 30220 94078 30260
rect 94078 30220 94118 30260
rect 94118 30220 94143 30260
rect 93889 30197 93975 30220
rect 94057 30197 94143 30220
rect 4409 29504 4495 29527
rect 4577 29504 4663 29527
rect 4409 29464 4434 29504
rect 4434 29464 4474 29504
rect 4474 29464 4495 29504
rect 4577 29464 4598 29504
rect 4598 29464 4638 29504
rect 4638 29464 4663 29504
rect 4409 29441 4495 29464
rect 4577 29441 4663 29464
rect 19529 29504 19615 29527
rect 19697 29504 19783 29527
rect 19529 29464 19554 29504
rect 19554 29464 19594 29504
rect 19594 29464 19615 29504
rect 19697 29464 19718 29504
rect 19718 29464 19758 29504
rect 19758 29464 19783 29504
rect 19529 29441 19615 29464
rect 19697 29441 19783 29464
rect 34649 29504 34735 29527
rect 34817 29504 34903 29527
rect 34649 29464 34674 29504
rect 34674 29464 34714 29504
rect 34714 29464 34735 29504
rect 34817 29464 34838 29504
rect 34838 29464 34878 29504
rect 34878 29464 34903 29504
rect 34649 29441 34735 29464
rect 34817 29441 34903 29464
rect 49769 29504 49855 29527
rect 49937 29504 50023 29527
rect 49769 29464 49794 29504
rect 49794 29464 49834 29504
rect 49834 29464 49855 29504
rect 49937 29464 49958 29504
rect 49958 29464 49998 29504
rect 49998 29464 50023 29504
rect 49769 29441 49855 29464
rect 49937 29441 50023 29464
rect 64889 29504 64975 29527
rect 65057 29504 65143 29527
rect 64889 29464 64914 29504
rect 64914 29464 64954 29504
rect 64954 29464 64975 29504
rect 65057 29464 65078 29504
rect 65078 29464 65118 29504
rect 65118 29464 65143 29504
rect 64889 29441 64975 29464
rect 65057 29441 65143 29464
rect 80009 29504 80095 29527
rect 80177 29504 80263 29527
rect 80009 29464 80034 29504
rect 80034 29464 80074 29504
rect 80074 29464 80095 29504
rect 80177 29464 80198 29504
rect 80198 29464 80238 29504
rect 80238 29464 80263 29504
rect 80009 29441 80095 29464
rect 80177 29441 80263 29464
rect 95129 29504 95215 29527
rect 95297 29504 95383 29527
rect 95129 29464 95154 29504
rect 95154 29464 95194 29504
rect 95194 29464 95215 29504
rect 95297 29464 95318 29504
rect 95318 29464 95358 29504
rect 95358 29464 95383 29504
rect 95129 29441 95215 29464
rect 95297 29441 95383 29464
rect 3169 28748 3255 28771
rect 3337 28748 3423 28771
rect 3169 28708 3194 28748
rect 3194 28708 3234 28748
rect 3234 28708 3255 28748
rect 3337 28708 3358 28748
rect 3358 28708 3398 28748
rect 3398 28708 3423 28748
rect 3169 28685 3255 28708
rect 3337 28685 3423 28708
rect 18289 28748 18375 28771
rect 18457 28748 18543 28771
rect 18289 28708 18314 28748
rect 18314 28708 18354 28748
rect 18354 28708 18375 28748
rect 18457 28708 18478 28748
rect 18478 28708 18518 28748
rect 18518 28708 18543 28748
rect 18289 28685 18375 28708
rect 18457 28685 18543 28708
rect 33409 28748 33495 28771
rect 33577 28748 33663 28771
rect 33409 28708 33434 28748
rect 33434 28708 33474 28748
rect 33474 28708 33495 28748
rect 33577 28708 33598 28748
rect 33598 28708 33638 28748
rect 33638 28708 33663 28748
rect 33409 28685 33495 28708
rect 33577 28685 33663 28708
rect 48529 28748 48615 28771
rect 48697 28748 48783 28771
rect 48529 28708 48554 28748
rect 48554 28708 48594 28748
rect 48594 28708 48615 28748
rect 48697 28708 48718 28748
rect 48718 28708 48758 28748
rect 48758 28708 48783 28748
rect 48529 28685 48615 28708
rect 48697 28685 48783 28708
rect 63649 28748 63735 28771
rect 63817 28748 63903 28771
rect 63649 28708 63674 28748
rect 63674 28708 63714 28748
rect 63714 28708 63735 28748
rect 63817 28708 63838 28748
rect 63838 28708 63878 28748
rect 63878 28708 63903 28748
rect 63649 28685 63735 28708
rect 63817 28685 63903 28708
rect 78769 28748 78855 28771
rect 78937 28748 79023 28771
rect 78769 28708 78794 28748
rect 78794 28708 78834 28748
rect 78834 28708 78855 28748
rect 78937 28708 78958 28748
rect 78958 28708 78998 28748
rect 78998 28708 79023 28748
rect 78769 28685 78855 28708
rect 78937 28685 79023 28708
rect 93889 28748 93975 28771
rect 94057 28748 94143 28771
rect 93889 28708 93914 28748
rect 93914 28708 93954 28748
rect 93954 28708 93975 28748
rect 94057 28708 94078 28748
rect 94078 28708 94118 28748
rect 94118 28708 94143 28748
rect 93889 28685 93975 28708
rect 94057 28685 94143 28708
rect 4409 27992 4495 28015
rect 4577 27992 4663 28015
rect 4409 27952 4434 27992
rect 4434 27952 4474 27992
rect 4474 27952 4495 27992
rect 4577 27952 4598 27992
rect 4598 27952 4638 27992
rect 4638 27952 4663 27992
rect 4409 27929 4495 27952
rect 4577 27929 4663 27952
rect 19529 27992 19615 28015
rect 19697 27992 19783 28015
rect 19529 27952 19554 27992
rect 19554 27952 19594 27992
rect 19594 27952 19615 27992
rect 19697 27952 19718 27992
rect 19718 27952 19758 27992
rect 19758 27952 19783 27992
rect 19529 27929 19615 27952
rect 19697 27929 19783 27952
rect 34649 27992 34735 28015
rect 34817 27992 34903 28015
rect 34649 27952 34674 27992
rect 34674 27952 34714 27992
rect 34714 27952 34735 27992
rect 34817 27952 34838 27992
rect 34838 27952 34878 27992
rect 34878 27952 34903 27992
rect 34649 27929 34735 27952
rect 34817 27929 34903 27952
rect 49769 27992 49855 28015
rect 49937 27992 50023 28015
rect 49769 27952 49794 27992
rect 49794 27952 49834 27992
rect 49834 27952 49855 27992
rect 49937 27952 49958 27992
rect 49958 27952 49998 27992
rect 49998 27952 50023 27992
rect 49769 27929 49855 27952
rect 49937 27929 50023 27952
rect 64889 27992 64975 28015
rect 65057 27992 65143 28015
rect 64889 27952 64914 27992
rect 64914 27952 64954 27992
rect 64954 27952 64975 27992
rect 65057 27952 65078 27992
rect 65078 27952 65118 27992
rect 65118 27952 65143 27992
rect 64889 27929 64975 27952
rect 65057 27929 65143 27952
rect 80009 27992 80095 28015
rect 80177 27992 80263 28015
rect 80009 27952 80034 27992
rect 80034 27952 80074 27992
rect 80074 27952 80095 27992
rect 80177 27952 80198 27992
rect 80198 27952 80238 27992
rect 80238 27952 80263 27992
rect 80009 27929 80095 27952
rect 80177 27929 80263 27952
rect 95129 27992 95215 28015
rect 95297 27992 95383 28015
rect 95129 27952 95154 27992
rect 95154 27952 95194 27992
rect 95194 27952 95215 27992
rect 95297 27952 95318 27992
rect 95318 27952 95358 27992
rect 95358 27952 95383 27992
rect 95129 27929 95215 27952
rect 95297 27929 95383 27952
rect 3169 27236 3255 27259
rect 3337 27236 3423 27259
rect 3169 27196 3194 27236
rect 3194 27196 3234 27236
rect 3234 27196 3255 27236
rect 3337 27196 3358 27236
rect 3358 27196 3398 27236
rect 3398 27196 3423 27236
rect 3169 27173 3255 27196
rect 3337 27173 3423 27196
rect 18289 27236 18375 27259
rect 18457 27236 18543 27259
rect 18289 27196 18314 27236
rect 18314 27196 18354 27236
rect 18354 27196 18375 27236
rect 18457 27196 18478 27236
rect 18478 27196 18518 27236
rect 18518 27196 18543 27236
rect 18289 27173 18375 27196
rect 18457 27173 18543 27196
rect 33409 27236 33495 27259
rect 33577 27236 33663 27259
rect 33409 27196 33434 27236
rect 33434 27196 33474 27236
rect 33474 27196 33495 27236
rect 33577 27196 33598 27236
rect 33598 27196 33638 27236
rect 33638 27196 33663 27236
rect 33409 27173 33495 27196
rect 33577 27173 33663 27196
rect 48529 27236 48615 27259
rect 48697 27236 48783 27259
rect 48529 27196 48554 27236
rect 48554 27196 48594 27236
rect 48594 27196 48615 27236
rect 48697 27196 48718 27236
rect 48718 27196 48758 27236
rect 48758 27196 48783 27236
rect 48529 27173 48615 27196
rect 48697 27173 48783 27196
rect 63649 27236 63735 27259
rect 63817 27236 63903 27259
rect 63649 27196 63674 27236
rect 63674 27196 63714 27236
rect 63714 27196 63735 27236
rect 63817 27196 63838 27236
rect 63838 27196 63878 27236
rect 63878 27196 63903 27236
rect 63649 27173 63735 27196
rect 63817 27173 63903 27196
rect 78769 27236 78855 27259
rect 78937 27236 79023 27259
rect 78769 27196 78794 27236
rect 78794 27196 78834 27236
rect 78834 27196 78855 27236
rect 78937 27196 78958 27236
rect 78958 27196 78998 27236
rect 78998 27196 79023 27236
rect 78769 27173 78855 27196
rect 78937 27173 79023 27196
rect 93889 27236 93975 27259
rect 94057 27236 94143 27259
rect 93889 27196 93914 27236
rect 93914 27196 93954 27236
rect 93954 27196 93975 27236
rect 94057 27196 94078 27236
rect 94078 27196 94118 27236
rect 94118 27196 94143 27236
rect 93889 27173 93975 27196
rect 94057 27173 94143 27196
rect 4409 26480 4495 26503
rect 4577 26480 4663 26503
rect 4409 26440 4434 26480
rect 4434 26440 4474 26480
rect 4474 26440 4495 26480
rect 4577 26440 4598 26480
rect 4598 26440 4638 26480
rect 4638 26440 4663 26480
rect 4409 26417 4495 26440
rect 4577 26417 4663 26440
rect 19529 26480 19615 26503
rect 19697 26480 19783 26503
rect 19529 26440 19554 26480
rect 19554 26440 19594 26480
rect 19594 26440 19615 26480
rect 19697 26440 19718 26480
rect 19718 26440 19758 26480
rect 19758 26440 19783 26480
rect 19529 26417 19615 26440
rect 19697 26417 19783 26440
rect 34649 26480 34735 26503
rect 34817 26480 34903 26503
rect 34649 26440 34674 26480
rect 34674 26440 34714 26480
rect 34714 26440 34735 26480
rect 34817 26440 34838 26480
rect 34838 26440 34878 26480
rect 34878 26440 34903 26480
rect 34649 26417 34735 26440
rect 34817 26417 34903 26440
rect 49769 26480 49855 26503
rect 49937 26480 50023 26503
rect 49769 26440 49794 26480
rect 49794 26440 49834 26480
rect 49834 26440 49855 26480
rect 49937 26440 49958 26480
rect 49958 26440 49998 26480
rect 49998 26440 50023 26480
rect 49769 26417 49855 26440
rect 49937 26417 50023 26440
rect 64889 26480 64975 26503
rect 65057 26480 65143 26503
rect 64889 26440 64914 26480
rect 64914 26440 64954 26480
rect 64954 26440 64975 26480
rect 65057 26440 65078 26480
rect 65078 26440 65118 26480
rect 65118 26440 65143 26480
rect 64889 26417 64975 26440
rect 65057 26417 65143 26440
rect 80009 26480 80095 26503
rect 80177 26480 80263 26503
rect 80009 26440 80034 26480
rect 80034 26440 80074 26480
rect 80074 26440 80095 26480
rect 80177 26440 80198 26480
rect 80198 26440 80238 26480
rect 80238 26440 80263 26480
rect 80009 26417 80095 26440
rect 80177 26417 80263 26440
rect 95129 26480 95215 26503
rect 95297 26480 95383 26503
rect 95129 26440 95154 26480
rect 95154 26440 95194 26480
rect 95194 26440 95215 26480
rect 95297 26440 95318 26480
rect 95318 26440 95358 26480
rect 95358 26440 95383 26480
rect 95129 26417 95215 26440
rect 95297 26417 95383 26440
rect 3169 25724 3255 25747
rect 3337 25724 3423 25747
rect 3169 25684 3194 25724
rect 3194 25684 3234 25724
rect 3234 25684 3255 25724
rect 3337 25684 3358 25724
rect 3358 25684 3398 25724
rect 3398 25684 3423 25724
rect 3169 25661 3255 25684
rect 3337 25661 3423 25684
rect 18289 25724 18375 25747
rect 18457 25724 18543 25747
rect 18289 25684 18314 25724
rect 18314 25684 18354 25724
rect 18354 25684 18375 25724
rect 18457 25684 18478 25724
rect 18478 25684 18518 25724
rect 18518 25684 18543 25724
rect 18289 25661 18375 25684
rect 18457 25661 18543 25684
rect 33409 25724 33495 25747
rect 33577 25724 33663 25747
rect 33409 25684 33434 25724
rect 33434 25684 33474 25724
rect 33474 25684 33495 25724
rect 33577 25684 33598 25724
rect 33598 25684 33638 25724
rect 33638 25684 33663 25724
rect 33409 25661 33495 25684
rect 33577 25661 33663 25684
rect 48529 25724 48615 25747
rect 48697 25724 48783 25747
rect 48529 25684 48554 25724
rect 48554 25684 48594 25724
rect 48594 25684 48615 25724
rect 48697 25684 48718 25724
rect 48718 25684 48758 25724
rect 48758 25684 48783 25724
rect 48529 25661 48615 25684
rect 48697 25661 48783 25684
rect 63649 25724 63735 25747
rect 63817 25724 63903 25747
rect 63649 25684 63674 25724
rect 63674 25684 63714 25724
rect 63714 25684 63735 25724
rect 63817 25684 63838 25724
rect 63838 25684 63878 25724
rect 63878 25684 63903 25724
rect 63649 25661 63735 25684
rect 63817 25661 63903 25684
rect 78769 25724 78855 25747
rect 78937 25724 79023 25747
rect 78769 25684 78794 25724
rect 78794 25684 78834 25724
rect 78834 25684 78855 25724
rect 78937 25684 78958 25724
rect 78958 25684 78998 25724
rect 78998 25684 79023 25724
rect 78769 25661 78855 25684
rect 78937 25661 79023 25684
rect 93889 25724 93975 25747
rect 94057 25724 94143 25747
rect 93889 25684 93914 25724
rect 93914 25684 93954 25724
rect 93954 25684 93975 25724
rect 94057 25684 94078 25724
rect 94078 25684 94118 25724
rect 94118 25684 94143 25724
rect 93889 25661 93975 25684
rect 94057 25661 94143 25684
rect 4409 24968 4495 24991
rect 4577 24968 4663 24991
rect 4409 24928 4434 24968
rect 4434 24928 4474 24968
rect 4474 24928 4495 24968
rect 4577 24928 4598 24968
rect 4598 24928 4638 24968
rect 4638 24928 4663 24968
rect 4409 24905 4495 24928
rect 4577 24905 4663 24928
rect 19529 24968 19615 24991
rect 19697 24968 19783 24991
rect 19529 24928 19554 24968
rect 19554 24928 19594 24968
rect 19594 24928 19615 24968
rect 19697 24928 19718 24968
rect 19718 24928 19758 24968
rect 19758 24928 19783 24968
rect 19529 24905 19615 24928
rect 19697 24905 19783 24928
rect 34649 24968 34735 24991
rect 34817 24968 34903 24991
rect 34649 24928 34674 24968
rect 34674 24928 34714 24968
rect 34714 24928 34735 24968
rect 34817 24928 34838 24968
rect 34838 24928 34878 24968
rect 34878 24928 34903 24968
rect 34649 24905 34735 24928
rect 34817 24905 34903 24928
rect 49769 24968 49855 24991
rect 49937 24968 50023 24991
rect 49769 24928 49794 24968
rect 49794 24928 49834 24968
rect 49834 24928 49855 24968
rect 49937 24928 49958 24968
rect 49958 24928 49998 24968
rect 49998 24928 50023 24968
rect 49769 24905 49855 24928
rect 49937 24905 50023 24928
rect 64889 24968 64975 24991
rect 65057 24968 65143 24991
rect 64889 24928 64914 24968
rect 64914 24928 64954 24968
rect 64954 24928 64975 24968
rect 65057 24928 65078 24968
rect 65078 24928 65118 24968
rect 65118 24928 65143 24968
rect 64889 24905 64975 24928
rect 65057 24905 65143 24928
rect 80009 24968 80095 24991
rect 80177 24968 80263 24991
rect 80009 24928 80034 24968
rect 80034 24928 80074 24968
rect 80074 24928 80095 24968
rect 80177 24928 80198 24968
rect 80198 24928 80238 24968
rect 80238 24928 80263 24968
rect 80009 24905 80095 24928
rect 80177 24905 80263 24928
rect 95129 24968 95215 24991
rect 95297 24968 95383 24991
rect 95129 24928 95154 24968
rect 95154 24928 95194 24968
rect 95194 24928 95215 24968
rect 95297 24928 95318 24968
rect 95318 24928 95358 24968
rect 95358 24928 95383 24968
rect 95129 24905 95215 24928
rect 95297 24905 95383 24928
rect 3169 24212 3255 24235
rect 3337 24212 3423 24235
rect 3169 24172 3194 24212
rect 3194 24172 3234 24212
rect 3234 24172 3255 24212
rect 3337 24172 3358 24212
rect 3358 24172 3398 24212
rect 3398 24172 3423 24212
rect 3169 24149 3255 24172
rect 3337 24149 3423 24172
rect 18289 24212 18375 24235
rect 18457 24212 18543 24235
rect 18289 24172 18314 24212
rect 18314 24172 18354 24212
rect 18354 24172 18375 24212
rect 18457 24172 18478 24212
rect 18478 24172 18518 24212
rect 18518 24172 18543 24212
rect 18289 24149 18375 24172
rect 18457 24149 18543 24172
rect 33409 24212 33495 24235
rect 33577 24212 33663 24235
rect 33409 24172 33434 24212
rect 33434 24172 33474 24212
rect 33474 24172 33495 24212
rect 33577 24172 33598 24212
rect 33598 24172 33638 24212
rect 33638 24172 33663 24212
rect 33409 24149 33495 24172
rect 33577 24149 33663 24172
rect 48529 24212 48615 24235
rect 48697 24212 48783 24235
rect 48529 24172 48554 24212
rect 48554 24172 48594 24212
rect 48594 24172 48615 24212
rect 48697 24172 48718 24212
rect 48718 24172 48758 24212
rect 48758 24172 48783 24212
rect 48529 24149 48615 24172
rect 48697 24149 48783 24172
rect 63649 24212 63735 24235
rect 63817 24212 63903 24235
rect 63649 24172 63674 24212
rect 63674 24172 63714 24212
rect 63714 24172 63735 24212
rect 63817 24172 63838 24212
rect 63838 24172 63878 24212
rect 63878 24172 63903 24212
rect 63649 24149 63735 24172
rect 63817 24149 63903 24172
rect 78769 24212 78855 24235
rect 78937 24212 79023 24235
rect 78769 24172 78794 24212
rect 78794 24172 78834 24212
rect 78834 24172 78855 24212
rect 78937 24172 78958 24212
rect 78958 24172 78998 24212
rect 78998 24172 79023 24212
rect 78769 24149 78855 24172
rect 78937 24149 79023 24172
rect 93889 24212 93975 24235
rect 94057 24212 94143 24235
rect 93889 24172 93914 24212
rect 93914 24172 93954 24212
rect 93954 24172 93975 24212
rect 94057 24172 94078 24212
rect 94078 24172 94118 24212
rect 94118 24172 94143 24212
rect 93889 24149 93975 24172
rect 94057 24149 94143 24172
rect 4409 23456 4495 23479
rect 4577 23456 4663 23479
rect 4409 23416 4434 23456
rect 4434 23416 4474 23456
rect 4474 23416 4495 23456
rect 4577 23416 4598 23456
rect 4598 23416 4638 23456
rect 4638 23416 4663 23456
rect 4409 23393 4495 23416
rect 4577 23393 4663 23416
rect 19529 23456 19615 23479
rect 19697 23456 19783 23479
rect 19529 23416 19554 23456
rect 19554 23416 19594 23456
rect 19594 23416 19615 23456
rect 19697 23416 19718 23456
rect 19718 23416 19758 23456
rect 19758 23416 19783 23456
rect 19529 23393 19615 23416
rect 19697 23393 19783 23416
rect 34649 23456 34735 23479
rect 34817 23456 34903 23479
rect 34649 23416 34674 23456
rect 34674 23416 34714 23456
rect 34714 23416 34735 23456
rect 34817 23416 34838 23456
rect 34838 23416 34878 23456
rect 34878 23416 34903 23456
rect 34649 23393 34735 23416
rect 34817 23393 34903 23416
rect 49769 23456 49855 23479
rect 49937 23456 50023 23479
rect 49769 23416 49794 23456
rect 49794 23416 49834 23456
rect 49834 23416 49855 23456
rect 49937 23416 49958 23456
rect 49958 23416 49998 23456
rect 49998 23416 50023 23456
rect 49769 23393 49855 23416
rect 49937 23393 50023 23416
rect 64889 23456 64975 23479
rect 65057 23456 65143 23479
rect 64889 23416 64914 23456
rect 64914 23416 64954 23456
rect 64954 23416 64975 23456
rect 65057 23416 65078 23456
rect 65078 23416 65118 23456
rect 65118 23416 65143 23456
rect 64889 23393 64975 23416
rect 65057 23393 65143 23416
rect 80009 23456 80095 23479
rect 80177 23456 80263 23479
rect 80009 23416 80034 23456
rect 80034 23416 80074 23456
rect 80074 23416 80095 23456
rect 80177 23416 80198 23456
rect 80198 23416 80238 23456
rect 80238 23416 80263 23456
rect 80009 23393 80095 23416
rect 80177 23393 80263 23416
rect 95129 23456 95215 23479
rect 95297 23456 95383 23479
rect 95129 23416 95154 23456
rect 95154 23416 95194 23456
rect 95194 23416 95215 23456
rect 95297 23416 95318 23456
rect 95318 23416 95358 23456
rect 95358 23416 95383 23456
rect 95129 23393 95215 23416
rect 95297 23393 95383 23416
rect 3169 22700 3255 22723
rect 3337 22700 3423 22723
rect 3169 22660 3194 22700
rect 3194 22660 3234 22700
rect 3234 22660 3255 22700
rect 3337 22660 3358 22700
rect 3358 22660 3398 22700
rect 3398 22660 3423 22700
rect 3169 22637 3255 22660
rect 3337 22637 3423 22660
rect 18289 22700 18375 22723
rect 18457 22700 18543 22723
rect 18289 22660 18314 22700
rect 18314 22660 18354 22700
rect 18354 22660 18375 22700
rect 18457 22660 18478 22700
rect 18478 22660 18518 22700
rect 18518 22660 18543 22700
rect 18289 22637 18375 22660
rect 18457 22637 18543 22660
rect 33409 22700 33495 22723
rect 33577 22700 33663 22723
rect 33409 22660 33434 22700
rect 33434 22660 33474 22700
rect 33474 22660 33495 22700
rect 33577 22660 33598 22700
rect 33598 22660 33638 22700
rect 33638 22660 33663 22700
rect 33409 22637 33495 22660
rect 33577 22637 33663 22660
rect 48529 22700 48615 22723
rect 48697 22700 48783 22723
rect 48529 22660 48554 22700
rect 48554 22660 48594 22700
rect 48594 22660 48615 22700
rect 48697 22660 48718 22700
rect 48718 22660 48758 22700
rect 48758 22660 48783 22700
rect 48529 22637 48615 22660
rect 48697 22637 48783 22660
rect 63649 22700 63735 22723
rect 63817 22700 63903 22723
rect 63649 22660 63674 22700
rect 63674 22660 63714 22700
rect 63714 22660 63735 22700
rect 63817 22660 63838 22700
rect 63838 22660 63878 22700
rect 63878 22660 63903 22700
rect 63649 22637 63735 22660
rect 63817 22637 63903 22660
rect 78769 22700 78855 22723
rect 78937 22700 79023 22723
rect 78769 22660 78794 22700
rect 78794 22660 78834 22700
rect 78834 22660 78855 22700
rect 78937 22660 78958 22700
rect 78958 22660 78998 22700
rect 78998 22660 79023 22700
rect 78769 22637 78855 22660
rect 78937 22637 79023 22660
rect 93889 22700 93975 22723
rect 94057 22700 94143 22723
rect 93889 22660 93914 22700
rect 93914 22660 93954 22700
rect 93954 22660 93975 22700
rect 94057 22660 94078 22700
rect 94078 22660 94118 22700
rect 94118 22660 94143 22700
rect 93889 22637 93975 22660
rect 94057 22637 94143 22660
rect 4409 21944 4495 21967
rect 4577 21944 4663 21967
rect 4409 21904 4434 21944
rect 4434 21904 4474 21944
rect 4474 21904 4495 21944
rect 4577 21904 4598 21944
rect 4598 21904 4638 21944
rect 4638 21904 4663 21944
rect 4409 21881 4495 21904
rect 4577 21881 4663 21904
rect 19529 21944 19615 21967
rect 19697 21944 19783 21967
rect 19529 21904 19554 21944
rect 19554 21904 19594 21944
rect 19594 21904 19615 21944
rect 19697 21904 19718 21944
rect 19718 21904 19758 21944
rect 19758 21904 19783 21944
rect 19529 21881 19615 21904
rect 19697 21881 19783 21904
rect 34649 21944 34735 21967
rect 34817 21944 34903 21967
rect 34649 21904 34674 21944
rect 34674 21904 34714 21944
rect 34714 21904 34735 21944
rect 34817 21904 34838 21944
rect 34838 21904 34878 21944
rect 34878 21904 34903 21944
rect 34649 21881 34735 21904
rect 34817 21881 34903 21904
rect 49769 21944 49855 21967
rect 49937 21944 50023 21967
rect 49769 21904 49794 21944
rect 49794 21904 49834 21944
rect 49834 21904 49855 21944
rect 49937 21904 49958 21944
rect 49958 21904 49998 21944
rect 49998 21904 50023 21944
rect 49769 21881 49855 21904
rect 49937 21881 50023 21904
rect 64889 21944 64975 21967
rect 65057 21944 65143 21967
rect 64889 21904 64914 21944
rect 64914 21904 64954 21944
rect 64954 21904 64975 21944
rect 65057 21904 65078 21944
rect 65078 21904 65118 21944
rect 65118 21904 65143 21944
rect 64889 21881 64975 21904
rect 65057 21881 65143 21904
rect 80009 21944 80095 21967
rect 80177 21944 80263 21967
rect 80009 21904 80034 21944
rect 80034 21904 80074 21944
rect 80074 21904 80095 21944
rect 80177 21904 80198 21944
rect 80198 21904 80238 21944
rect 80238 21904 80263 21944
rect 80009 21881 80095 21904
rect 80177 21881 80263 21904
rect 95129 21944 95215 21967
rect 95297 21944 95383 21967
rect 95129 21904 95154 21944
rect 95154 21904 95194 21944
rect 95194 21904 95215 21944
rect 95297 21904 95318 21944
rect 95318 21904 95358 21944
rect 95358 21904 95383 21944
rect 95129 21881 95215 21904
rect 95297 21881 95383 21904
rect 3169 21188 3255 21211
rect 3337 21188 3423 21211
rect 3169 21148 3194 21188
rect 3194 21148 3234 21188
rect 3234 21148 3255 21188
rect 3337 21148 3358 21188
rect 3358 21148 3398 21188
rect 3398 21148 3423 21188
rect 3169 21125 3255 21148
rect 3337 21125 3423 21148
rect 18289 21188 18375 21211
rect 18457 21188 18543 21211
rect 18289 21148 18314 21188
rect 18314 21148 18354 21188
rect 18354 21148 18375 21188
rect 18457 21148 18478 21188
rect 18478 21148 18518 21188
rect 18518 21148 18543 21188
rect 18289 21125 18375 21148
rect 18457 21125 18543 21148
rect 33409 21188 33495 21211
rect 33577 21188 33663 21211
rect 33409 21148 33434 21188
rect 33434 21148 33474 21188
rect 33474 21148 33495 21188
rect 33577 21148 33598 21188
rect 33598 21148 33638 21188
rect 33638 21148 33663 21188
rect 33409 21125 33495 21148
rect 33577 21125 33663 21148
rect 48529 21188 48615 21211
rect 48697 21188 48783 21211
rect 48529 21148 48554 21188
rect 48554 21148 48594 21188
rect 48594 21148 48615 21188
rect 48697 21148 48718 21188
rect 48718 21148 48758 21188
rect 48758 21148 48783 21188
rect 48529 21125 48615 21148
rect 48697 21125 48783 21148
rect 63649 21188 63735 21211
rect 63817 21188 63903 21211
rect 63649 21148 63674 21188
rect 63674 21148 63714 21188
rect 63714 21148 63735 21188
rect 63817 21148 63838 21188
rect 63838 21148 63878 21188
rect 63878 21148 63903 21188
rect 63649 21125 63735 21148
rect 63817 21125 63903 21148
rect 78769 21188 78855 21211
rect 78937 21188 79023 21211
rect 78769 21148 78794 21188
rect 78794 21148 78834 21188
rect 78834 21148 78855 21188
rect 78937 21148 78958 21188
rect 78958 21148 78998 21188
rect 78998 21148 79023 21188
rect 78769 21125 78855 21148
rect 78937 21125 79023 21148
rect 93889 21188 93975 21211
rect 94057 21188 94143 21211
rect 93889 21148 93914 21188
rect 93914 21148 93954 21188
rect 93954 21148 93975 21188
rect 94057 21148 94078 21188
rect 94078 21148 94118 21188
rect 94118 21148 94143 21188
rect 93889 21125 93975 21148
rect 94057 21125 94143 21148
rect 4409 20432 4495 20455
rect 4577 20432 4663 20455
rect 4409 20392 4434 20432
rect 4434 20392 4474 20432
rect 4474 20392 4495 20432
rect 4577 20392 4598 20432
rect 4598 20392 4638 20432
rect 4638 20392 4663 20432
rect 4409 20369 4495 20392
rect 4577 20369 4663 20392
rect 19529 20432 19615 20455
rect 19697 20432 19783 20455
rect 19529 20392 19554 20432
rect 19554 20392 19594 20432
rect 19594 20392 19615 20432
rect 19697 20392 19718 20432
rect 19718 20392 19758 20432
rect 19758 20392 19783 20432
rect 19529 20369 19615 20392
rect 19697 20369 19783 20392
rect 34649 20432 34735 20455
rect 34817 20432 34903 20455
rect 34649 20392 34674 20432
rect 34674 20392 34714 20432
rect 34714 20392 34735 20432
rect 34817 20392 34838 20432
rect 34838 20392 34878 20432
rect 34878 20392 34903 20432
rect 34649 20369 34735 20392
rect 34817 20369 34903 20392
rect 49769 20432 49855 20455
rect 49937 20432 50023 20455
rect 49769 20392 49794 20432
rect 49794 20392 49834 20432
rect 49834 20392 49855 20432
rect 49937 20392 49958 20432
rect 49958 20392 49998 20432
rect 49998 20392 50023 20432
rect 49769 20369 49855 20392
rect 49937 20369 50023 20392
rect 64889 20432 64975 20455
rect 65057 20432 65143 20455
rect 64889 20392 64914 20432
rect 64914 20392 64954 20432
rect 64954 20392 64975 20432
rect 65057 20392 65078 20432
rect 65078 20392 65118 20432
rect 65118 20392 65143 20432
rect 64889 20369 64975 20392
rect 65057 20369 65143 20392
rect 80009 20432 80095 20455
rect 80177 20432 80263 20455
rect 80009 20392 80034 20432
rect 80034 20392 80074 20432
rect 80074 20392 80095 20432
rect 80177 20392 80198 20432
rect 80198 20392 80238 20432
rect 80238 20392 80263 20432
rect 80009 20369 80095 20392
rect 80177 20369 80263 20392
rect 95129 20432 95215 20455
rect 95297 20432 95383 20455
rect 95129 20392 95154 20432
rect 95154 20392 95194 20432
rect 95194 20392 95215 20432
rect 95297 20392 95318 20432
rect 95318 20392 95358 20432
rect 95358 20392 95383 20432
rect 95129 20369 95215 20392
rect 95297 20369 95383 20392
rect 3169 19676 3255 19699
rect 3337 19676 3423 19699
rect 3169 19636 3194 19676
rect 3194 19636 3234 19676
rect 3234 19636 3255 19676
rect 3337 19636 3358 19676
rect 3358 19636 3398 19676
rect 3398 19636 3423 19676
rect 3169 19613 3255 19636
rect 3337 19613 3423 19636
rect 18289 19676 18375 19699
rect 18457 19676 18543 19699
rect 18289 19636 18314 19676
rect 18314 19636 18354 19676
rect 18354 19636 18375 19676
rect 18457 19636 18478 19676
rect 18478 19636 18518 19676
rect 18518 19636 18543 19676
rect 18289 19613 18375 19636
rect 18457 19613 18543 19636
rect 33409 19676 33495 19699
rect 33577 19676 33663 19699
rect 33409 19636 33434 19676
rect 33434 19636 33474 19676
rect 33474 19636 33495 19676
rect 33577 19636 33598 19676
rect 33598 19636 33638 19676
rect 33638 19636 33663 19676
rect 33409 19613 33495 19636
rect 33577 19613 33663 19636
rect 48529 19676 48615 19699
rect 48697 19676 48783 19699
rect 48529 19636 48554 19676
rect 48554 19636 48594 19676
rect 48594 19636 48615 19676
rect 48697 19636 48718 19676
rect 48718 19636 48758 19676
rect 48758 19636 48783 19676
rect 48529 19613 48615 19636
rect 48697 19613 48783 19636
rect 63649 19676 63735 19699
rect 63817 19676 63903 19699
rect 63649 19636 63674 19676
rect 63674 19636 63714 19676
rect 63714 19636 63735 19676
rect 63817 19636 63838 19676
rect 63838 19636 63878 19676
rect 63878 19636 63903 19676
rect 63649 19613 63735 19636
rect 63817 19613 63903 19636
rect 78769 19676 78855 19699
rect 78937 19676 79023 19699
rect 78769 19636 78794 19676
rect 78794 19636 78834 19676
rect 78834 19636 78855 19676
rect 78937 19636 78958 19676
rect 78958 19636 78998 19676
rect 78998 19636 79023 19676
rect 78769 19613 78855 19636
rect 78937 19613 79023 19636
rect 93889 19676 93975 19699
rect 94057 19676 94143 19699
rect 93889 19636 93914 19676
rect 93914 19636 93954 19676
rect 93954 19636 93975 19676
rect 94057 19636 94078 19676
rect 94078 19636 94118 19676
rect 94118 19636 94143 19676
rect 93889 19613 93975 19636
rect 94057 19613 94143 19636
rect 4409 18920 4495 18943
rect 4577 18920 4663 18943
rect 4409 18880 4434 18920
rect 4434 18880 4474 18920
rect 4474 18880 4495 18920
rect 4577 18880 4598 18920
rect 4598 18880 4638 18920
rect 4638 18880 4663 18920
rect 4409 18857 4495 18880
rect 4577 18857 4663 18880
rect 19529 18920 19615 18943
rect 19697 18920 19783 18943
rect 19529 18880 19554 18920
rect 19554 18880 19594 18920
rect 19594 18880 19615 18920
rect 19697 18880 19718 18920
rect 19718 18880 19758 18920
rect 19758 18880 19783 18920
rect 19529 18857 19615 18880
rect 19697 18857 19783 18880
rect 34649 18920 34735 18943
rect 34817 18920 34903 18943
rect 34649 18880 34674 18920
rect 34674 18880 34714 18920
rect 34714 18880 34735 18920
rect 34817 18880 34838 18920
rect 34838 18880 34878 18920
rect 34878 18880 34903 18920
rect 34649 18857 34735 18880
rect 34817 18857 34903 18880
rect 49769 18920 49855 18943
rect 49937 18920 50023 18943
rect 49769 18880 49794 18920
rect 49794 18880 49834 18920
rect 49834 18880 49855 18920
rect 49937 18880 49958 18920
rect 49958 18880 49998 18920
rect 49998 18880 50023 18920
rect 49769 18857 49855 18880
rect 49937 18857 50023 18880
rect 64889 18920 64975 18943
rect 65057 18920 65143 18943
rect 64889 18880 64914 18920
rect 64914 18880 64954 18920
rect 64954 18880 64975 18920
rect 65057 18880 65078 18920
rect 65078 18880 65118 18920
rect 65118 18880 65143 18920
rect 64889 18857 64975 18880
rect 65057 18857 65143 18880
rect 80009 18920 80095 18943
rect 80177 18920 80263 18943
rect 80009 18880 80034 18920
rect 80034 18880 80074 18920
rect 80074 18880 80095 18920
rect 80177 18880 80198 18920
rect 80198 18880 80238 18920
rect 80238 18880 80263 18920
rect 80009 18857 80095 18880
rect 80177 18857 80263 18880
rect 95129 18920 95215 18943
rect 95297 18920 95383 18943
rect 95129 18880 95154 18920
rect 95154 18880 95194 18920
rect 95194 18880 95215 18920
rect 95297 18880 95318 18920
rect 95318 18880 95358 18920
rect 95358 18880 95383 18920
rect 95129 18857 95215 18880
rect 95297 18857 95383 18880
rect 3169 18164 3255 18187
rect 3337 18164 3423 18187
rect 3169 18124 3194 18164
rect 3194 18124 3234 18164
rect 3234 18124 3255 18164
rect 3337 18124 3358 18164
rect 3358 18124 3398 18164
rect 3398 18124 3423 18164
rect 3169 18101 3255 18124
rect 3337 18101 3423 18124
rect 18289 18164 18375 18187
rect 18457 18164 18543 18187
rect 18289 18124 18314 18164
rect 18314 18124 18354 18164
rect 18354 18124 18375 18164
rect 18457 18124 18478 18164
rect 18478 18124 18518 18164
rect 18518 18124 18543 18164
rect 18289 18101 18375 18124
rect 18457 18101 18543 18124
rect 33409 18164 33495 18187
rect 33577 18164 33663 18187
rect 33409 18124 33434 18164
rect 33434 18124 33474 18164
rect 33474 18124 33495 18164
rect 33577 18124 33598 18164
rect 33598 18124 33638 18164
rect 33638 18124 33663 18164
rect 33409 18101 33495 18124
rect 33577 18101 33663 18124
rect 48529 18164 48615 18187
rect 48697 18164 48783 18187
rect 48529 18124 48554 18164
rect 48554 18124 48594 18164
rect 48594 18124 48615 18164
rect 48697 18124 48718 18164
rect 48718 18124 48758 18164
rect 48758 18124 48783 18164
rect 48529 18101 48615 18124
rect 48697 18101 48783 18124
rect 63649 18164 63735 18187
rect 63817 18164 63903 18187
rect 63649 18124 63674 18164
rect 63674 18124 63714 18164
rect 63714 18124 63735 18164
rect 63817 18124 63838 18164
rect 63838 18124 63878 18164
rect 63878 18124 63903 18164
rect 63649 18101 63735 18124
rect 63817 18101 63903 18124
rect 78769 18164 78855 18187
rect 78937 18164 79023 18187
rect 78769 18124 78794 18164
rect 78794 18124 78834 18164
rect 78834 18124 78855 18164
rect 78937 18124 78958 18164
rect 78958 18124 78998 18164
rect 78998 18124 79023 18164
rect 78769 18101 78855 18124
rect 78937 18101 79023 18124
rect 93889 18164 93975 18187
rect 94057 18164 94143 18187
rect 93889 18124 93914 18164
rect 93914 18124 93954 18164
rect 93954 18124 93975 18164
rect 94057 18124 94078 18164
rect 94078 18124 94118 18164
rect 94118 18124 94143 18164
rect 93889 18101 93975 18124
rect 94057 18101 94143 18124
rect 4409 17408 4495 17431
rect 4577 17408 4663 17431
rect 4409 17368 4434 17408
rect 4434 17368 4474 17408
rect 4474 17368 4495 17408
rect 4577 17368 4598 17408
rect 4598 17368 4638 17408
rect 4638 17368 4663 17408
rect 4409 17345 4495 17368
rect 4577 17345 4663 17368
rect 19529 17408 19615 17431
rect 19697 17408 19783 17431
rect 19529 17368 19554 17408
rect 19554 17368 19594 17408
rect 19594 17368 19615 17408
rect 19697 17368 19718 17408
rect 19718 17368 19758 17408
rect 19758 17368 19783 17408
rect 19529 17345 19615 17368
rect 19697 17345 19783 17368
rect 34649 17408 34735 17431
rect 34817 17408 34903 17431
rect 34649 17368 34674 17408
rect 34674 17368 34714 17408
rect 34714 17368 34735 17408
rect 34817 17368 34838 17408
rect 34838 17368 34878 17408
rect 34878 17368 34903 17408
rect 34649 17345 34735 17368
rect 34817 17345 34903 17368
rect 49769 17408 49855 17431
rect 49937 17408 50023 17431
rect 49769 17368 49794 17408
rect 49794 17368 49834 17408
rect 49834 17368 49855 17408
rect 49937 17368 49958 17408
rect 49958 17368 49998 17408
rect 49998 17368 50023 17408
rect 49769 17345 49855 17368
rect 49937 17345 50023 17368
rect 64889 17408 64975 17431
rect 65057 17408 65143 17431
rect 64889 17368 64914 17408
rect 64914 17368 64954 17408
rect 64954 17368 64975 17408
rect 65057 17368 65078 17408
rect 65078 17368 65118 17408
rect 65118 17368 65143 17408
rect 64889 17345 64975 17368
rect 65057 17345 65143 17368
rect 80009 17408 80095 17431
rect 80177 17408 80263 17431
rect 80009 17368 80034 17408
rect 80034 17368 80074 17408
rect 80074 17368 80095 17408
rect 80177 17368 80198 17408
rect 80198 17368 80238 17408
rect 80238 17368 80263 17408
rect 80009 17345 80095 17368
rect 80177 17345 80263 17368
rect 95129 17408 95215 17431
rect 95297 17408 95383 17431
rect 95129 17368 95154 17408
rect 95154 17368 95194 17408
rect 95194 17368 95215 17408
rect 95297 17368 95318 17408
rect 95318 17368 95358 17408
rect 95358 17368 95383 17408
rect 95129 17345 95215 17368
rect 95297 17345 95383 17368
rect 3169 16652 3255 16675
rect 3337 16652 3423 16675
rect 3169 16612 3194 16652
rect 3194 16612 3234 16652
rect 3234 16612 3255 16652
rect 3337 16612 3358 16652
rect 3358 16612 3398 16652
rect 3398 16612 3423 16652
rect 3169 16589 3255 16612
rect 3337 16589 3423 16612
rect 18289 16652 18375 16675
rect 18457 16652 18543 16675
rect 18289 16612 18314 16652
rect 18314 16612 18354 16652
rect 18354 16612 18375 16652
rect 18457 16612 18478 16652
rect 18478 16612 18518 16652
rect 18518 16612 18543 16652
rect 18289 16589 18375 16612
rect 18457 16589 18543 16612
rect 33409 16652 33495 16675
rect 33577 16652 33663 16675
rect 33409 16612 33434 16652
rect 33434 16612 33474 16652
rect 33474 16612 33495 16652
rect 33577 16612 33598 16652
rect 33598 16612 33638 16652
rect 33638 16612 33663 16652
rect 33409 16589 33495 16612
rect 33577 16589 33663 16612
rect 48529 16652 48615 16675
rect 48697 16652 48783 16675
rect 48529 16612 48554 16652
rect 48554 16612 48594 16652
rect 48594 16612 48615 16652
rect 48697 16612 48718 16652
rect 48718 16612 48758 16652
rect 48758 16612 48783 16652
rect 48529 16589 48615 16612
rect 48697 16589 48783 16612
rect 63649 16652 63735 16675
rect 63817 16652 63903 16675
rect 63649 16612 63674 16652
rect 63674 16612 63714 16652
rect 63714 16612 63735 16652
rect 63817 16612 63838 16652
rect 63838 16612 63878 16652
rect 63878 16612 63903 16652
rect 63649 16589 63735 16612
rect 63817 16589 63903 16612
rect 78769 16652 78855 16675
rect 78937 16652 79023 16675
rect 78769 16612 78794 16652
rect 78794 16612 78834 16652
rect 78834 16612 78855 16652
rect 78937 16612 78958 16652
rect 78958 16612 78998 16652
rect 78998 16612 79023 16652
rect 78769 16589 78855 16612
rect 78937 16589 79023 16612
rect 93889 16652 93975 16675
rect 94057 16652 94143 16675
rect 93889 16612 93914 16652
rect 93914 16612 93954 16652
rect 93954 16612 93975 16652
rect 94057 16612 94078 16652
rect 94078 16612 94118 16652
rect 94118 16612 94143 16652
rect 93889 16589 93975 16612
rect 94057 16589 94143 16612
rect 4409 15896 4495 15919
rect 4577 15896 4663 15919
rect 4409 15856 4434 15896
rect 4434 15856 4474 15896
rect 4474 15856 4495 15896
rect 4577 15856 4598 15896
rect 4598 15856 4638 15896
rect 4638 15856 4663 15896
rect 4409 15833 4495 15856
rect 4577 15833 4663 15856
rect 19529 15896 19615 15919
rect 19697 15896 19783 15919
rect 19529 15856 19554 15896
rect 19554 15856 19594 15896
rect 19594 15856 19615 15896
rect 19697 15856 19718 15896
rect 19718 15856 19758 15896
rect 19758 15856 19783 15896
rect 19529 15833 19615 15856
rect 19697 15833 19783 15856
rect 34649 15896 34735 15919
rect 34817 15896 34903 15919
rect 34649 15856 34674 15896
rect 34674 15856 34714 15896
rect 34714 15856 34735 15896
rect 34817 15856 34838 15896
rect 34838 15856 34878 15896
rect 34878 15856 34903 15896
rect 34649 15833 34735 15856
rect 34817 15833 34903 15856
rect 49769 15896 49855 15919
rect 49937 15896 50023 15919
rect 49769 15856 49794 15896
rect 49794 15856 49834 15896
rect 49834 15856 49855 15896
rect 49937 15856 49958 15896
rect 49958 15856 49998 15896
rect 49998 15856 50023 15896
rect 49769 15833 49855 15856
rect 49937 15833 50023 15856
rect 64889 15896 64975 15919
rect 65057 15896 65143 15919
rect 64889 15856 64914 15896
rect 64914 15856 64954 15896
rect 64954 15856 64975 15896
rect 65057 15856 65078 15896
rect 65078 15856 65118 15896
rect 65118 15856 65143 15896
rect 64889 15833 64975 15856
rect 65057 15833 65143 15856
rect 80009 15896 80095 15919
rect 80177 15896 80263 15919
rect 80009 15856 80034 15896
rect 80034 15856 80074 15896
rect 80074 15856 80095 15896
rect 80177 15856 80198 15896
rect 80198 15856 80238 15896
rect 80238 15856 80263 15896
rect 80009 15833 80095 15856
rect 80177 15833 80263 15856
rect 95129 15896 95215 15919
rect 95297 15896 95383 15919
rect 95129 15856 95154 15896
rect 95154 15856 95194 15896
rect 95194 15856 95215 15896
rect 95297 15856 95318 15896
rect 95318 15856 95358 15896
rect 95358 15856 95383 15896
rect 95129 15833 95215 15856
rect 95297 15833 95383 15856
rect 3169 15140 3255 15163
rect 3337 15140 3423 15163
rect 3169 15100 3194 15140
rect 3194 15100 3234 15140
rect 3234 15100 3255 15140
rect 3337 15100 3358 15140
rect 3358 15100 3398 15140
rect 3398 15100 3423 15140
rect 3169 15077 3255 15100
rect 3337 15077 3423 15100
rect 18289 15140 18375 15163
rect 18457 15140 18543 15163
rect 18289 15100 18314 15140
rect 18314 15100 18354 15140
rect 18354 15100 18375 15140
rect 18457 15100 18478 15140
rect 18478 15100 18518 15140
rect 18518 15100 18543 15140
rect 18289 15077 18375 15100
rect 18457 15077 18543 15100
rect 33409 15140 33495 15163
rect 33577 15140 33663 15163
rect 33409 15100 33434 15140
rect 33434 15100 33474 15140
rect 33474 15100 33495 15140
rect 33577 15100 33598 15140
rect 33598 15100 33638 15140
rect 33638 15100 33663 15140
rect 33409 15077 33495 15100
rect 33577 15077 33663 15100
rect 48529 15140 48615 15163
rect 48697 15140 48783 15163
rect 48529 15100 48554 15140
rect 48554 15100 48594 15140
rect 48594 15100 48615 15140
rect 48697 15100 48718 15140
rect 48718 15100 48758 15140
rect 48758 15100 48783 15140
rect 48529 15077 48615 15100
rect 48697 15077 48783 15100
rect 63649 15140 63735 15163
rect 63817 15140 63903 15163
rect 63649 15100 63674 15140
rect 63674 15100 63714 15140
rect 63714 15100 63735 15140
rect 63817 15100 63838 15140
rect 63838 15100 63878 15140
rect 63878 15100 63903 15140
rect 63649 15077 63735 15100
rect 63817 15077 63903 15100
rect 78769 15140 78855 15163
rect 78937 15140 79023 15163
rect 78769 15100 78794 15140
rect 78794 15100 78834 15140
rect 78834 15100 78855 15140
rect 78937 15100 78958 15140
rect 78958 15100 78998 15140
rect 78998 15100 79023 15140
rect 78769 15077 78855 15100
rect 78937 15077 79023 15100
rect 93889 15140 93975 15163
rect 94057 15140 94143 15163
rect 93889 15100 93914 15140
rect 93914 15100 93954 15140
rect 93954 15100 93975 15140
rect 94057 15100 94078 15140
rect 94078 15100 94118 15140
rect 94118 15100 94143 15140
rect 93889 15077 93975 15100
rect 94057 15077 94143 15100
rect 4409 14384 4495 14407
rect 4577 14384 4663 14407
rect 4409 14344 4434 14384
rect 4434 14344 4474 14384
rect 4474 14344 4495 14384
rect 4577 14344 4598 14384
rect 4598 14344 4638 14384
rect 4638 14344 4663 14384
rect 4409 14321 4495 14344
rect 4577 14321 4663 14344
rect 19529 14384 19615 14407
rect 19697 14384 19783 14407
rect 19529 14344 19554 14384
rect 19554 14344 19594 14384
rect 19594 14344 19615 14384
rect 19697 14344 19718 14384
rect 19718 14344 19758 14384
rect 19758 14344 19783 14384
rect 19529 14321 19615 14344
rect 19697 14321 19783 14344
rect 34649 14384 34735 14407
rect 34817 14384 34903 14407
rect 34649 14344 34674 14384
rect 34674 14344 34714 14384
rect 34714 14344 34735 14384
rect 34817 14344 34838 14384
rect 34838 14344 34878 14384
rect 34878 14344 34903 14384
rect 34649 14321 34735 14344
rect 34817 14321 34903 14344
rect 49769 14384 49855 14407
rect 49937 14384 50023 14407
rect 49769 14344 49794 14384
rect 49794 14344 49834 14384
rect 49834 14344 49855 14384
rect 49937 14344 49958 14384
rect 49958 14344 49998 14384
rect 49998 14344 50023 14384
rect 49769 14321 49855 14344
rect 49937 14321 50023 14344
rect 64889 14384 64975 14407
rect 65057 14384 65143 14407
rect 64889 14344 64914 14384
rect 64914 14344 64954 14384
rect 64954 14344 64975 14384
rect 65057 14344 65078 14384
rect 65078 14344 65118 14384
rect 65118 14344 65143 14384
rect 64889 14321 64975 14344
rect 65057 14321 65143 14344
rect 80009 14384 80095 14407
rect 80177 14384 80263 14407
rect 80009 14344 80034 14384
rect 80034 14344 80074 14384
rect 80074 14344 80095 14384
rect 80177 14344 80198 14384
rect 80198 14344 80238 14384
rect 80238 14344 80263 14384
rect 80009 14321 80095 14344
rect 80177 14321 80263 14344
rect 95129 14384 95215 14407
rect 95297 14384 95383 14407
rect 95129 14344 95154 14384
rect 95154 14344 95194 14384
rect 95194 14344 95215 14384
rect 95297 14344 95318 14384
rect 95318 14344 95358 14384
rect 95358 14344 95383 14384
rect 95129 14321 95215 14344
rect 95297 14321 95383 14344
rect 3169 13628 3255 13651
rect 3337 13628 3423 13651
rect 3169 13588 3194 13628
rect 3194 13588 3234 13628
rect 3234 13588 3255 13628
rect 3337 13588 3358 13628
rect 3358 13588 3398 13628
rect 3398 13588 3423 13628
rect 3169 13565 3255 13588
rect 3337 13565 3423 13588
rect 18289 13628 18375 13651
rect 18457 13628 18543 13651
rect 18289 13588 18314 13628
rect 18314 13588 18354 13628
rect 18354 13588 18375 13628
rect 18457 13588 18478 13628
rect 18478 13588 18518 13628
rect 18518 13588 18543 13628
rect 18289 13565 18375 13588
rect 18457 13565 18543 13588
rect 33409 13628 33495 13651
rect 33577 13628 33663 13651
rect 33409 13588 33434 13628
rect 33434 13588 33474 13628
rect 33474 13588 33495 13628
rect 33577 13588 33598 13628
rect 33598 13588 33638 13628
rect 33638 13588 33663 13628
rect 33409 13565 33495 13588
rect 33577 13565 33663 13588
rect 48529 13628 48615 13651
rect 48697 13628 48783 13651
rect 48529 13588 48554 13628
rect 48554 13588 48594 13628
rect 48594 13588 48615 13628
rect 48697 13588 48718 13628
rect 48718 13588 48758 13628
rect 48758 13588 48783 13628
rect 48529 13565 48615 13588
rect 48697 13565 48783 13588
rect 63649 13628 63735 13651
rect 63817 13628 63903 13651
rect 63649 13588 63674 13628
rect 63674 13588 63714 13628
rect 63714 13588 63735 13628
rect 63817 13588 63838 13628
rect 63838 13588 63878 13628
rect 63878 13588 63903 13628
rect 63649 13565 63735 13588
rect 63817 13565 63903 13588
rect 78769 13628 78855 13651
rect 78937 13628 79023 13651
rect 78769 13588 78794 13628
rect 78794 13588 78834 13628
rect 78834 13588 78855 13628
rect 78937 13588 78958 13628
rect 78958 13588 78998 13628
rect 78998 13588 79023 13628
rect 78769 13565 78855 13588
rect 78937 13565 79023 13588
rect 93889 13628 93975 13651
rect 94057 13628 94143 13651
rect 93889 13588 93914 13628
rect 93914 13588 93954 13628
rect 93954 13588 93975 13628
rect 94057 13588 94078 13628
rect 94078 13588 94118 13628
rect 94118 13588 94143 13628
rect 93889 13565 93975 13588
rect 94057 13565 94143 13588
rect 4409 12872 4495 12895
rect 4577 12872 4663 12895
rect 4409 12832 4434 12872
rect 4434 12832 4474 12872
rect 4474 12832 4495 12872
rect 4577 12832 4598 12872
rect 4598 12832 4638 12872
rect 4638 12832 4663 12872
rect 4409 12809 4495 12832
rect 4577 12809 4663 12832
rect 19529 12872 19615 12895
rect 19697 12872 19783 12895
rect 19529 12832 19554 12872
rect 19554 12832 19594 12872
rect 19594 12832 19615 12872
rect 19697 12832 19718 12872
rect 19718 12832 19758 12872
rect 19758 12832 19783 12872
rect 19529 12809 19615 12832
rect 19697 12809 19783 12832
rect 34649 12872 34735 12895
rect 34817 12872 34903 12895
rect 34649 12832 34674 12872
rect 34674 12832 34714 12872
rect 34714 12832 34735 12872
rect 34817 12832 34838 12872
rect 34838 12832 34878 12872
rect 34878 12832 34903 12872
rect 34649 12809 34735 12832
rect 34817 12809 34903 12832
rect 49769 12872 49855 12895
rect 49937 12872 50023 12895
rect 49769 12832 49794 12872
rect 49794 12832 49834 12872
rect 49834 12832 49855 12872
rect 49937 12832 49958 12872
rect 49958 12832 49998 12872
rect 49998 12832 50023 12872
rect 49769 12809 49855 12832
rect 49937 12809 50023 12832
rect 64889 12872 64975 12895
rect 65057 12872 65143 12895
rect 64889 12832 64914 12872
rect 64914 12832 64954 12872
rect 64954 12832 64975 12872
rect 65057 12832 65078 12872
rect 65078 12832 65118 12872
rect 65118 12832 65143 12872
rect 64889 12809 64975 12832
rect 65057 12809 65143 12832
rect 80009 12872 80095 12895
rect 80177 12872 80263 12895
rect 80009 12832 80034 12872
rect 80034 12832 80074 12872
rect 80074 12832 80095 12872
rect 80177 12832 80198 12872
rect 80198 12832 80238 12872
rect 80238 12832 80263 12872
rect 80009 12809 80095 12832
rect 80177 12809 80263 12832
rect 95129 12872 95215 12895
rect 95297 12872 95383 12895
rect 95129 12832 95154 12872
rect 95154 12832 95194 12872
rect 95194 12832 95215 12872
rect 95297 12832 95318 12872
rect 95318 12832 95358 12872
rect 95358 12832 95383 12872
rect 95129 12809 95215 12832
rect 95297 12809 95383 12832
rect 3169 12116 3255 12139
rect 3337 12116 3423 12139
rect 3169 12076 3194 12116
rect 3194 12076 3234 12116
rect 3234 12076 3255 12116
rect 3337 12076 3358 12116
rect 3358 12076 3398 12116
rect 3398 12076 3423 12116
rect 3169 12053 3255 12076
rect 3337 12053 3423 12076
rect 18289 12116 18375 12139
rect 18457 12116 18543 12139
rect 18289 12076 18314 12116
rect 18314 12076 18354 12116
rect 18354 12076 18375 12116
rect 18457 12076 18478 12116
rect 18478 12076 18518 12116
rect 18518 12076 18543 12116
rect 18289 12053 18375 12076
rect 18457 12053 18543 12076
rect 33409 12116 33495 12139
rect 33577 12116 33663 12139
rect 33409 12076 33434 12116
rect 33434 12076 33474 12116
rect 33474 12076 33495 12116
rect 33577 12076 33598 12116
rect 33598 12076 33638 12116
rect 33638 12076 33663 12116
rect 33409 12053 33495 12076
rect 33577 12053 33663 12076
rect 48529 12116 48615 12139
rect 48697 12116 48783 12139
rect 48529 12076 48554 12116
rect 48554 12076 48594 12116
rect 48594 12076 48615 12116
rect 48697 12076 48718 12116
rect 48718 12076 48758 12116
rect 48758 12076 48783 12116
rect 48529 12053 48615 12076
rect 48697 12053 48783 12076
rect 63649 12116 63735 12139
rect 63817 12116 63903 12139
rect 63649 12076 63674 12116
rect 63674 12076 63714 12116
rect 63714 12076 63735 12116
rect 63817 12076 63838 12116
rect 63838 12076 63878 12116
rect 63878 12076 63903 12116
rect 63649 12053 63735 12076
rect 63817 12053 63903 12076
rect 78769 12116 78855 12139
rect 78937 12116 79023 12139
rect 78769 12076 78794 12116
rect 78794 12076 78834 12116
rect 78834 12076 78855 12116
rect 78937 12076 78958 12116
rect 78958 12076 78998 12116
rect 78998 12076 79023 12116
rect 78769 12053 78855 12076
rect 78937 12053 79023 12076
rect 93889 12116 93975 12139
rect 94057 12116 94143 12139
rect 93889 12076 93914 12116
rect 93914 12076 93954 12116
rect 93954 12076 93975 12116
rect 94057 12076 94078 12116
rect 94078 12076 94118 12116
rect 94118 12076 94143 12116
rect 93889 12053 93975 12076
rect 94057 12053 94143 12076
rect 4409 11360 4495 11383
rect 4577 11360 4663 11383
rect 4409 11320 4434 11360
rect 4434 11320 4474 11360
rect 4474 11320 4495 11360
rect 4577 11320 4598 11360
rect 4598 11320 4638 11360
rect 4638 11320 4663 11360
rect 4409 11297 4495 11320
rect 4577 11297 4663 11320
rect 19529 11360 19615 11383
rect 19697 11360 19783 11383
rect 19529 11320 19554 11360
rect 19554 11320 19594 11360
rect 19594 11320 19615 11360
rect 19697 11320 19718 11360
rect 19718 11320 19758 11360
rect 19758 11320 19783 11360
rect 19529 11297 19615 11320
rect 19697 11297 19783 11320
rect 34649 11360 34735 11383
rect 34817 11360 34903 11383
rect 34649 11320 34674 11360
rect 34674 11320 34714 11360
rect 34714 11320 34735 11360
rect 34817 11320 34838 11360
rect 34838 11320 34878 11360
rect 34878 11320 34903 11360
rect 34649 11297 34735 11320
rect 34817 11297 34903 11320
rect 49769 11360 49855 11383
rect 49937 11360 50023 11383
rect 49769 11320 49794 11360
rect 49794 11320 49834 11360
rect 49834 11320 49855 11360
rect 49937 11320 49958 11360
rect 49958 11320 49998 11360
rect 49998 11320 50023 11360
rect 49769 11297 49855 11320
rect 49937 11297 50023 11320
rect 64889 11360 64975 11383
rect 65057 11360 65143 11383
rect 64889 11320 64914 11360
rect 64914 11320 64954 11360
rect 64954 11320 64975 11360
rect 65057 11320 65078 11360
rect 65078 11320 65118 11360
rect 65118 11320 65143 11360
rect 64889 11297 64975 11320
rect 65057 11297 65143 11320
rect 80009 11360 80095 11383
rect 80177 11360 80263 11383
rect 80009 11320 80034 11360
rect 80034 11320 80074 11360
rect 80074 11320 80095 11360
rect 80177 11320 80198 11360
rect 80198 11320 80238 11360
rect 80238 11320 80263 11360
rect 80009 11297 80095 11320
rect 80177 11297 80263 11320
rect 95129 11360 95215 11383
rect 95297 11360 95383 11383
rect 95129 11320 95154 11360
rect 95154 11320 95194 11360
rect 95194 11320 95215 11360
rect 95297 11320 95318 11360
rect 95318 11320 95358 11360
rect 95358 11320 95383 11360
rect 95129 11297 95215 11320
rect 95297 11297 95383 11320
rect 3169 10604 3255 10627
rect 3337 10604 3423 10627
rect 3169 10564 3194 10604
rect 3194 10564 3234 10604
rect 3234 10564 3255 10604
rect 3337 10564 3358 10604
rect 3358 10564 3398 10604
rect 3398 10564 3423 10604
rect 3169 10541 3255 10564
rect 3337 10541 3423 10564
rect 18289 10604 18375 10627
rect 18457 10604 18543 10627
rect 18289 10564 18314 10604
rect 18314 10564 18354 10604
rect 18354 10564 18375 10604
rect 18457 10564 18478 10604
rect 18478 10564 18518 10604
rect 18518 10564 18543 10604
rect 18289 10541 18375 10564
rect 18457 10541 18543 10564
rect 33409 10604 33495 10627
rect 33577 10604 33663 10627
rect 33409 10564 33434 10604
rect 33434 10564 33474 10604
rect 33474 10564 33495 10604
rect 33577 10564 33598 10604
rect 33598 10564 33638 10604
rect 33638 10564 33663 10604
rect 33409 10541 33495 10564
rect 33577 10541 33663 10564
rect 48529 10604 48615 10627
rect 48697 10604 48783 10627
rect 48529 10564 48554 10604
rect 48554 10564 48594 10604
rect 48594 10564 48615 10604
rect 48697 10564 48718 10604
rect 48718 10564 48758 10604
rect 48758 10564 48783 10604
rect 48529 10541 48615 10564
rect 48697 10541 48783 10564
rect 63649 10604 63735 10627
rect 63817 10604 63903 10627
rect 63649 10564 63674 10604
rect 63674 10564 63714 10604
rect 63714 10564 63735 10604
rect 63817 10564 63838 10604
rect 63838 10564 63878 10604
rect 63878 10564 63903 10604
rect 63649 10541 63735 10564
rect 63817 10541 63903 10564
rect 78769 10604 78855 10627
rect 78937 10604 79023 10627
rect 78769 10564 78794 10604
rect 78794 10564 78834 10604
rect 78834 10564 78855 10604
rect 78937 10564 78958 10604
rect 78958 10564 78998 10604
rect 78998 10564 79023 10604
rect 78769 10541 78855 10564
rect 78937 10541 79023 10564
rect 93889 10604 93975 10627
rect 94057 10604 94143 10627
rect 93889 10564 93914 10604
rect 93914 10564 93954 10604
rect 93954 10564 93975 10604
rect 94057 10564 94078 10604
rect 94078 10564 94118 10604
rect 94118 10564 94143 10604
rect 93889 10541 93975 10564
rect 94057 10541 94143 10564
rect 4409 9848 4495 9871
rect 4577 9848 4663 9871
rect 4409 9808 4434 9848
rect 4434 9808 4474 9848
rect 4474 9808 4495 9848
rect 4577 9808 4598 9848
rect 4598 9808 4638 9848
rect 4638 9808 4663 9848
rect 4409 9785 4495 9808
rect 4577 9785 4663 9808
rect 19529 9848 19615 9871
rect 19697 9848 19783 9871
rect 19529 9808 19554 9848
rect 19554 9808 19594 9848
rect 19594 9808 19615 9848
rect 19697 9808 19718 9848
rect 19718 9808 19758 9848
rect 19758 9808 19783 9848
rect 19529 9785 19615 9808
rect 19697 9785 19783 9808
rect 34649 9848 34735 9871
rect 34817 9848 34903 9871
rect 34649 9808 34674 9848
rect 34674 9808 34714 9848
rect 34714 9808 34735 9848
rect 34817 9808 34838 9848
rect 34838 9808 34878 9848
rect 34878 9808 34903 9848
rect 34649 9785 34735 9808
rect 34817 9785 34903 9808
rect 49769 9848 49855 9871
rect 49937 9848 50023 9871
rect 49769 9808 49794 9848
rect 49794 9808 49834 9848
rect 49834 9808 49855 9848
rect 49937 9808 49958 9848
rect 49958 9808 49998 9848
rect 49998 9808 50023 9848
rect 49769 9785 49855 9808
rect 49937 9785 50023 9808
rect 64889 9848 64975 9871
rect 65057 9848 65143 9871
rect 64889 9808 64914 9848
rect 64914 9808 64954 9848
rect 64954 9808 64975 9848
rect 65057 9808 65078 9848
rect 65078 9808 65118 9848
rect 65118 9808 65143 9848
rect 64889 9785 64975 9808
rect 65057 9785 65143 9808
rect 80009 9848 80095 9871
rect 80177 9848 80263 9871
rect 80009 9808 80034 9848
rect 80034 9808 80074 9848
rect 80074 9808 80095 9848
rect 80177 9808 80198 9848
rect 80198 9808 80238 9848
rect 80238 9808 80263 9848
rect 80009 9785 80095 9808
rect 80177 9785 80263 9808
rect 95129 9848 95215 9871
rect 95297 9848 95383 9871
rect 95129 9808 95154 9848
rect 95154 9808 95194 9848
rect 95194 9808 95215 9848
rect 95297 9808 95318 9848
rect 95318 9808 95358 9848
rect 95358 9808 95383 9848
rect 95129 9785 95215 9808
rect 95297 9785 95383 9808
rect 3169 9092 3255 9115
rect 3337 9092 3423 9115
rect 3169 9052 3194 9092
rect 3194 9052 3234 9092
rect 3234 9052 3255 9092
rect 3337 9052 3358 9092
rect 3358 9052 3398 9092
rect 3398 9052 3423 9092
rect 3169 9029 3255 9052
rect 3337 9029 3423 9052
rect 18289 9092 18375 9115
rect 18457 9092 18543 9115
rect 18289 9052 18314 9092
rect 18314 9052 18354 9092
rect 18354 9052 18375 9092
rect 18457 9052 18478 9092
rect 18478 9052 18518 9092
rect 18518 9052 18543 9092
rect 18289 9029 18375 9052
rect 18457 9029 18543 9052
rect 33409 9092 33495 9115
rect 33577 9092 33663 9115
rect 33409 9052 33434 9092
rect 33434 9052 33474 9092
rect 33474 9052 33495 9092
rect 33577 9052 33598 9092
rect 33598 9052 33638 9092
rect 33638 9052 33663 9092
rect 33409 9029 33495 9052
rect 33577 9029 33663 9052
rect 48529 9092 48615 9115
rect 48697 9092 48783 9115
rect 48529 9052 48554 9092
rect 48554 9052 48594 9092
rect 48594 9052 48615 9092
rect 48697 9052 48718 9092
rect 48718 9052 48758 9092
rect 48758 9052 48783 9092
rect 48529 9029 48615 9052
rect 48697 9029 48783 9052
rect 63649 9092 63735 9115
rect 63817 9092 63903 9115
rect 63649 9052 63674 9092
rect 63674 9052 63714 9092
rect 63714 9052 63735 9092
rect 63817 9052 63838 9092
rect 63838 9052 63878 9092
rect 63878 9052 63903 9092
rect 63649 9029 63735 9052
rect 63817 9029 63903 9052
rect 78769 9092 78855 9115
rect 78937 9092 79023 9115
rect 78769 9052 78794 9092
rect 78794 9052 78834 9092
rect 78834 9052 78855 9092
rect 78937 9052 78958 9092
rect 78958 9052 78998 9092
rect 78998 9052 79023 9092
rect 78769 9029 78855 9052
rect 78937 9029 79023 9052
rect 93889 9092 93975 9115
rect 94057 9092 94143 9115
rect 93889 9052 93914 9092
rect 93914 9052 93954 9092
rect 93954 9052 93975 9092
rect 94057 9052 94078 9092
rect 94078 9052 94118 9092
rect 94118 9052 94143 9092
rect 93889 9029 93975 9052
rect 94057 9029 94143 9052
rect 4409 8336 4495 8359
rect 4577 8336 4663 8359
rect 4409 8296 4434 8336
rect 4434 8296 4474 8336
rect 4474 8296 4495 8336
rect 4577 8296 4598 8336
rect 4598 8296 4638 8336
rect 4638 8296 4663 8336
rect 4409 8273 4495 8296
rect 4577 8273 4663 8296
rect 19529 8336 19615 8359
rect 19697 8336 19783 8359
rect 19529 8296 19554 8336
rect 19554 8296 19594 8336
rect 19594 8296 19615 8336
rect 19697 8296 19718 8336
rect 19718 8296 19758 8336
rect 19758 8296 19783 8336
rect 19529 8273 19615 8296
rect 19697 8273 19783 8296
rect 34649 8336 34735 8359
rect 34817 8336 34903 8359
rect 34649 8296 34674 8336
rect 34674 8296 34714 8336
rect 34714 8296 34735 8336
rect 34817 8296 34838 8336
rect 34838 8296 34878 8336
rect 34878 8296 34903 8336
rect 34649 8273 34735 8296
rect 34817 8273 34903 8296
rect 49769 8336 49855 8359
rect 49937 8336 50023 8359
rect 49769 8296 49794 8336
rect 49794 8296 49834 8336
rect 49834 8296 49855 8336
rect 49937 8296 49958 8336
rect 49958 8296 49998 8336
rect 49998 8296 50023 8336
rect 49769 8273 49855 8296
rect 49937 8273 50023 8296
rect 64889 8336 64975 8359
rect 65057 8336 65143 8359
rect 64889 8296 64914 8336
rect 64914 8296 64954 8336
rect 64954 8296 64975 8336
rect 65057 8296 65078 8336
rect 65078 8296 65118 8336
rect 65118 8296 65143 8336
rect 64889 8273 64975 8296
rect 65057 8273 65143 8296
rect 80009 8336 80095 8359
rect 80177 8336 80263 8359
rect 80009 8296 80034 8336
rect 80034 8296 80074 8336
rect 80074 8296 80095 8336
rect 80177 8296 80198 8336
rect 80198 8296 80238 8336
rect 80238 8296 80263 8336
rect 80009 8273 80095 8296
rect 80177 8273 80263 8296
rect 95129 8336 95215 8359
rect 95297 8336 95383 8359
rect 95129 8296 95154 8336
rect 95154 8296 95194 8336
rect 95194 8296 95215 8336
rect 95297 8296 95318 8336
rect 95318 8296 95358 8336
rect 95358 8296 95383 8336
rect 95129 8273 95215 8296
rect 95297 8273 95383 8296
rect 3169 7580 3255 7603
rect 3337 7580 3423 7603
rect 3169 7540 3194 7580
rect 3194 7540 3234 7580
rect 3234 7540 3255 7580
rect 3337 7540 3358 7580
rect 3358 7540 3398 7580
rect 3398 7540 3423 7580
rect 3169 7517 3255 7540
rect 3337 7517 3423 7540
rect 18289 7580 18375 7603
rect 18457 7580 18543 7603
rect 18289 7540 18314 7580
rect 18314 7540 18354 7580
rect 18354 7540 18375 7580
rect 18457 7540 18478 7580
rect 18478 7540 18518 7580
rect 18518 7540 18543 7580
rect 18289 7517 18375 7540
rect 18457 7517 18543 7540
rect 33409 7580 33495 7603
rect 33577 7580 33663 7603
rect 33409 7540 33434 7580
rect 33434 7540 33474 7580
rect 33474 7540 33495 7580
rect 33577 7540 33598 7580
rect 33598 7540 33638 7580
rect 33638 7540 33663 7580
rect 33409 7517 33495 7540
rect 33577 7517 33663 7540
rect 48529 7580 48615 7603
rect 48697 7580 48783 7603
rect 48529 7540 48554 7580
rect 48554 7540 48594 7580
rect 48594 7540 48615 7580
rect 48697 7540 48718 7580
rect 48718 7540 48758 7580
rect 48758 7540 48783 7580
rect 48529 7517 48615 7540
rect 48697 7517 48783 7540
rect 63649 7580 63735 7603
rect 63817 7580 63903 7603
rect 63649 7540 63674 7580
rect 63674 7540 63714 7580
rect 63714 7540 63735 7580
rect 63817 7540 63838 7580
rect 63838 7540 63878 7580
rect 63878 7540 63903 7580
rect 63649 7517 63735 7540
rect 63817 7517 63903 7540
rect 78769 7580 78855 7603
rect 78937 7580 79023 7603
rect 78769 7540 78794 7580
rect 78794 7540 78834 7580
rect 78834 7540 78855 7580
rect 78937 7540 78958 7580
rect 78958 7540 78998 7580
rect 78998 7540 79023 7580
rect 78769 7517 78855 7540
rect 78937 7517 79023 7540
rect 93889 7580 93975 7603
rect 94057 7580 94143 7603
rect 93889 7540 93914 7580
rect 93914 7540 93954 7580
rect 93954 7540 93975 7580
rect 94057 7540 94078 7580
rect 94078 7540 94118 7580
rect 94118 7540 94143 7580
rect 93889 7517 93975 7540
rect 94057 7517 94143 7540
rect 4409 6824 4495 6847
rect 4577 6824 4663 6847
rect 4409 6784 4434 6824
rect 4434 6784 4474 6824
rect 4474 6784 4495 6824
rect 4577 6784 4598 6824
rect 4598 6784 4638 6824
rect 4638 6784 4663 6824
rect 4409 6761 4495 6784
rect 4577 6761 4663 6784
rect 19529 6824 19615 6847
rect 19697 6824 19783 6847
rect 19529 6784 19554 6824
rect 19554 6784 19594 6824
rect 19594 6784 19615 6824
rect 19697 6784 19718 6824
rect 19718 6784 19758 6824
rect 19758 6784 19783 6824
rect 19529 6761 19615 6784
rect 19697 6761 19783 6784
rect 34649 6824 34735 6847
rect 34817 6824 34903 6847
rect 34649 6784 34674 6824
rect 34674 6784 34714 6824
rect 34714 6784 34735 6824
rect 34817 6784 34838 6824
rect 34838 6784 34878 6824
rect 34878 6784 34903 6824
rect 34649 6761 34735 6784
rect 34817 6761 34903 6784
rect 49769 6824 49855 6847
rect 49937 6824 50023 6847
rect 49769 6784 49794 6824
rect 49794 6784 49834 6824
rect 49834 6784 49855 6824
rect 49937 6784 49958 6824
rect 49958 6784 49998 6824
rect 49998 6784 50023 6824
rect 49769 6761 49855 6784
rect 49937 6761 50023 6784
rect 64889 6824 64975 6847
rect 65057 6824 65143 6847
rect 64889 6784 64914 6824
rect 64914 6784 64954 6824
rect 64954 6784 64975 6824
rect 65057 6784 65078 6824
rect 65078 6784 65118 6824
rect 65118 6784 65143 6824
rect 64889 6761 64975 6784
rect 65057 6761 65143 6784
rect 80009 6824 80095 6847
rect 80177 6824 80263 6847
rect 80009 6784 80034 6824
rect 80034 6784 80074 6824
rect 80074 6784 80095 6824
rect 80177 6784 80198 6824
rect 80198 6784 80238 6824
rect 80238 6784 80263 6824
rect 80009 6761 80095 6784
rect 80177 6761 80263 6784
rect 95129 6824 95215 6847
rect 95297 6824 95383 6847
rect 95129 6784 95154 6824
rect 95154 6784 95194 6824
rect 95194 6784 95215 6824
rect 95297 6784 95318 6824
rect 95318 6784 95358 6824
rect 95358 6784 95383 6824
rect 95129 6761 95215 6784
rect 95297 6761 95383 6784
rect 3169 6068 3255 6091
rect 3337 6068 3423 6091
rect 3169 6028 3194 6068
rect 3194 6028 3234 6068
rect 3234 6028 3255 6068
rect 3337 6028 3358 6068
rect 3358 6028 3398 6068
rect 3398 6028 3423 6068
rect 3169 6005 3255 6028
rect 3337 6005 3423 6028
rect 18289 6068 18375 6091
rect 18457 6068 18543 6091
rect 18289 6028 18314 6068
rect 18314 6028 18354 6068
rect 18354 6028 18375 6068
rect 18457 6028 18478 6068
rect 18478 6028 18518 6068
rect 18518 6028 18543 6068
rect 18289 6005 18375 6028
rect 18457 6005 18543 6028
rect 33409 6068 33495 6091
rect 33577 6068 33663 6091
rect 33409 6028 33434 6068
rect 33434 6028 33474 6068
rect 33474 6028 33495 6068
rect 33577 6028 33598 6068
rect 33598 6028 33638 6068
rect 33638 6028 33663 6068
rect 33409 6005 33495 6028
rect 33577 6005 33663 6028
rect 48529 6068 48615 6091
rect 48697 6068 48783 6091
rect 48529 6028 48554 6068
rect 48554 6028 48594 6068
rect 48594 6028 48615 6068
rect 48697 6028 48718 6068
rect 48718 6028 48758 6068
rect 48758 6028 48783 6068
rect 48529 6005 48615 6028
rect 48697 6005 48783 6028
rect 63649 6068 63735 6091
rect 63817 6068 63903 6091
rect 63649 6028 63674 6068
rect 63674 6028 63714 6068
rect 63714 6028 63735 6068
rect 63817 6028 63838 6068
rect 63838 6028 63878 6068
rect 63878 6028 63903 6068
rect 63649 6005 63735 6028
rect 63817 6005 63903 6028
rect 78769 6068 78855 6091
rect 78937 6068 79023 6091
rect 78769 6028 78794 6068
rect 78794 6028 78834 6068
rect 78834 6028 78855 6068
rect 78937 6028 78958 6068
rect 78958 6028 78998 6068
rect 78998 6028 79023 6068
rect 78769 6005 78855 6028
rect 78937 6005 79023 6028
rect 93889 6068 93975 6091
rect 94057 6068 94143 6091
rect 93889 6028 93914 6068
rect 93914 6028 93954 6068
rect 93954 6028 93975 6068
rect 94057 6028 94078 6068
rect 94078 6028 94118 6068
rect 94118 6028 94143 6068
rect 93889 6005 93975 6028
rect 94057 6005 94143 6028
rect 4409 5312 4495 5335
rect 4577 5312 4663 5335
rect 4409 5272 4434 5312
rect 4434 5272 4474 5312
rect 4474 5272 4495 5312
rect 4577 5272 4598 5312
rect 4598 5272 4638 5312
rect 4638 5272 4663 5312
rect 4409 5249 4495 5272
rect 4577 5249 4663 5272
rect 19529 5312 19615 5335
rect 19697 5312 19783 5335
rect 19529 5272 19554 5312
rect 19554 5272 19594 5312
rect 19594 5272 19615 5312
rect 19697 5272 19718 5312
rect 19718 5272 19758 5312
rect 19758 5272 19783 5312
rect 19529 5249 19615 5272
rect 19697 5249 19783 5272
rect 34649 5312 34735 5335
rect 34817 5312 34903 5335
rect 34649 5272 34674 5312
rect 34674 5272 34714 5312
rect 34714 5272 34735 5312
rect 34817 5272 34838 5312
rect 34838 5272 34878 5312
rect 34878 5272 34903 5312
rect 34649 5249 34735 5272
rect 34817 5249 34903 5272
rect 49769 5312 49855 5335
rect 49937 5312 50023 5335
rect 49769 5272 49794 5312
rect 49794 5272 49834 5312
rect 49834 5272 49855 5312
rect 49937 5272 49958 5312
rect 49958 5272 49998 5312
rect 49998 5272 50023 5312
rect 49769 5249 49855 5272
rect 49937 5249 50023 5272
rect 64889 5312 64975 5335
rect 65057 5312 65143 5335
rect 64889 5272 64914 5312
rect 64914 5272 64954 5312
rect 64954 5272 64975 5312
rect 65057 5272 65078 5312
rect 65078 5272 65118 5312
rect 65118 5272 65143 5312
rect 64889 5249 64975 5272
rect 65057 5249 65143 5272
rect 80009 5312 80095 5335
rect 80177 5312 80263 5335
rect 80009 5272 80034 5312
rect 80034 5272 80074 5312
rect 80074 5272 80095 5312
rect 80177 5272 80198 5312
rect 80198 5272 80238 5312
rect 80238 5272 80263 5312
rect 80009 5249 80095 5272
rect 80177 5249 80263 5272
rect 95129 5312 95215 5335
rect 95297 5312 95383 5335
rect 95129 5272 95154 5312
rect 95154 5272 95194 5312
rect 95194 5272 95215 5312
rect 95297 5272 95318 5312
rect 95318 5272 95358 5312
rect 95358 5272 95383 5312
rect 95129 5249 95215 5272
rect 95297 5249 95383 5272
rect 3169 4556 3255 4579
rect 3337 4556 3423 4579
rect 3169 4516 3194 4556
rect 3194 4516 3234 4556
rect 3234 4516 3255 4556
rect 3337 4516 3358 4556
rect 3358 4516 3398 4556
rect 3398 4516 3423 4556
rect 3169 4493 3255 4516
rect 3337 4493 3423 4516
rect 18289 4556 18375 4579
rect 18457 4556 18543 4579
rect 18289 4516 18314 4556
rect 18314 4516 18354 4556
rect 18354 4516 18375 4556
rect 18457 4516 18478 4556
rect 18478 4516 18518 4556
rect 18518 4516 18543 4556
rect 18289 4493 18375 4516
rect 18457 4493 18543 4516
rect 33409 4556 33495 4579
rect 33577 4556 33663 4579
rect 33409 4516 33434 4556
rect 33434 4516 33474 4556
rect 33474 4516 33495 4556
rect 33577 4516 33598 4556
rect 33598 4516 33638 4556
rect 33638 4516 33663 4556
rect 33409 4493 33495 4516
rect 33577 4493 33663 4516
rect 48529 4556 48615 4579
rect 48697 4556 48783 4579
rect 48529 4516 48554 4556
rect 48554 4516 48594 4556
rect 48594 4516 48615 4556
rect 48697 4516 48718 4556
rect 48718 4516 48758 4556
rect 48758 4516 48783 4556
rect 48529 4493 48615 4516
rect 48697 4493 48783 4516
rect 63649 4556 63735 4579
rect 63817 4556 63903 4579
rect 63649 4516 63674 4556
rect 63674 4516 63714 4556
rect 63714 4516 63735 4556
rect 63817 4516 63838 4556
rect 63838 4516 63878 4556
rect 63878 4516 63903 4556
rect 63649 4493 63735 4516
rect 63817 4493 63903 4516
rect 78769 4556 78855 4579
rect 78937 4556 79023 4579
rect 78769 4516 78794 4556
rect 78794 4516 78834 4556
rect 78834 4516 78855 4556
rect 78937 4516 78958 4556
rect 78958 4516 78998 4556
rect 78998 4516 79023 4556
rect 78769 4493 78855 4516
rect 78937 4493 79023 4516
rect 93889 4556 93975 4579
rect 94057 4556 94143 4579
rect 93889 4516 93914 4556
rect 93914 4516 93954 4556
rect 93954 4516 93975 4556
rect 94057 4516 94078 4556
rect 94078 4516 94118 4556
rect 94118 4516 94143 4556
rect 93889 4493 93975 4516
rect 94057 4493 94143 4516
rect 4409 3800 4495 3823
rect 4577 3800 4663 3823
rect 4409 3760 4434 3800
rect 4434 3760 4474 3800
rect 4474 3760 4495 3800
rect 4577 3760 4598 3800
rect 4598 3760 4638 3800
rect 4638 3760 4663 3800
rect 4409 3737 4495 3760
rect 4577 3737 4663 3760
rect 19529 3800 19615 3823
rect 19697 3800 19783 3823
rect 19529 3760 19554 3800
rect 19554 3760 19594 3800
rect 19594 3760 19615 3800
rect 19697 3760 19718 3800
rect 19718 3760 19758 3800
rect 19758 3760 19783 3800
rect 19529 3737 19615 3760
rect 19697 3737 19783 3760
rect 34649 3800 34735 3823
rect 34817 3800 34903 3823
rect 34649 3760 34674 3800
rect 34674 3760 34714 3800
rect 34714 3760 34735 3800
rect 34817 3760 34838 3800
rect 34838 3760 34878 3800
rect 34878 3760 34903 3800
rect 34649 3737 34735 3760
rect 34817 3737 34903 3760
rect 49769 3800 49855 3823
rect 49937 3800 50023 3823
rect 49769 3760 49794 3800
rect 49794 3760 49834 3800
rect 49834 3760 49855 3800
rect 49937 3760 49958 3800
rect 49958 3760 49998 3800
rect 49998 3760 50023 3800
rect 49769 3737 49855 3760
rect 49937 3737 50023 3760
rect 64889 3800 64975 3823
rect 65057 3800 65143 3823
rect 64889 3760 64914 3800
rect 64914 3760 64954 3800
rect 64954 3760 64975 3800
rect 65057 3760 65078 3800
rect 65078 3760 65118 3800
rect 65118 3760 65143 3800
rect 64889 3737 64975 3760
rect 65057 3737 65143 3760
rect 80009 3800 80095 3823
rect 80177 3800 80263 3823
rect 80009 3760 80034 3800
rect 80034 3760 80074 3800
rect 80074 3760 80095 3800
rect 80177 3760 80198 3800
rect 80198 3760 80238 3800
rect 80238 3760 80263 3800
rect 80009 3737 80095 3760
rect 80177 3737 80263 3760
rect 95129 3800 95215 3823
rect 95297 3800 95383 3823
rect 95129 3760 95154 3800
rect 95154 3760 95194 3800
rect 95194 3760 95215 3800
rect 95297 3760 95318 3800
rect 95318 3760 95358 3800
rect 95358 3760 95383 3800
rect 95129 3737 95215 3760
rect 95297 3737 95383 3760
rect 3169 3044 3255 3067
rect 3337 3044 3423 3067
rect 3169 3004 3194 3044
rect 3194 3004 3234 3044
rect 3234 3004 3255 3044
rect 3337 3004 3358 3044
rect 3358 3004 3398 3044
rect 3398 3004 3423 3044
rect 3169 2981 3255 3004
rect 3337 2981 3423 3004
rect 18289 3044 18375 3067
rect 18457 3044 18543 3067
rect 18289 3004 18314 3044
rect 18314 3004 18354 3044
rect 18354 3004 18375 3044
rect 18457 3004 18478 3044
rect 18478 3004 18518 3044
rect 18518 3004 18543 3044
rect 18289 2981 18375 3004
rect 18457 2981 18543 3004
rect 33409 3044 33495 3067
rect 33577 3044 33663 3067
rect 33409 3004 33434 3044
rect 33434 3004 33474 3044
rect 33474 3004 33495 3044
rect 33577 3004 33598 3044
rect 33598 3004 33638 3044
rect 33638 3004 33663 3044
rect 33409 2981 33495 3004
rect 33577 2981 33663 3004
rect 48529 3044 48615 3067
rect 48697 3044 48783 3067
rect 48529 3004 48554 3044
rect 48554 3004 48594 3044
rect 48594 3004 48615 3044
rect 48697 3004 48718 3044
rect 48718 3004 48758 3044
rect 48758 3004 48783 3044
rect 48529 2981 48615 3004
rect 48697 2981 48783 3004
rect 63649 3044 63735 3067
rect 63817 3044 63903 3067
rect 63649 3004 63674 3044
rect 63674 3004 63714 3044
rect 63714 3004 63735 3044
rect 63817 3004 63838 3044
rect 63838 3004 63878 3044
rect 63878 3004 63903 3044
rect 63649 2981 63735 3004
rect 63817 2981 63903 3004
rect 78769 3044 78855 3067
rect 78937 3044 79023 3067
rect 78769 3004 78794 3044
rect 78794 3004 78834 3044
rect 78834 3004 78855 3044
rect 78937 3004 78958 3044
rect 78958 3004 78998 3044
rect 78998 3004 79023 3044
rect 78769 2981 78855 3004
rect 78937 2981 79023 3004
rect 93889 3044 93975 3067
rect 94057 3044 94143 3067
rect 93889 3004 93914 3044
rect 93914 3004 93954 3044
rect 93954 3004 93975 3044
rect 94057 3004 94078 3044
rect 94078 3004 94118 3044
rect 94118 3004 94143 3044
rect 93889 2981 93975 3004
rect 94057 2981 94143 3004
rect 4409 2288 4495 2311
rect 4577 2288 4663 2311
rect 4409 2248 4434 2288
rect 4434 2248 4474 2288
rect 4474 2248 4495 2288
rect 4577 2248 4598 2288
rect 4598 2248 4638 2288
rect 4638 2248 4663 2288
rect 4409 2225 4495 2248
rect 4577 2225 4663 2248
rect 19529 2288 19615 2311
rect 19697 2288 19783 2311
rect 19529 2248 19554 2288
rect 19554 2248 19594 2288
rect 19594 2248 19615 2288
rect 19697 2248 19718 2288
rect 19718 2248 19758 2288
rect 19758 2248 19783 2288
rect 19529 2225 19615 2248
rect 19697 2225 19783 2248
rect 34649 2288 34735 2311
rect 34817 2288 34903 2311
rect 34649 2248 34674 2288
rect 34674 2248 34714 2288
rect 34714 2248 34735 2288
rect 34817 2248 34838 2288
rect 34838 2248 34878 2288
rect 34878 2248 34903 2288
rect 34649 2225 34735 2248
rect 34817 2225 34903 2248
rect 49769 2288 49855 2311
rect 49937 2288 50023 2311
rect 49769 2248 49794 2288
rect 49794 2248 49834 2288
rect 49834 2248 49855 2288
rect 49937 2248 49958 2288
rect 49958 2248 49998 2288
rect 49998 2248 50023 2288
rect 49769 2225 49855 2248
rect 49937 2225 50023 2248
rect 64889 2288 64975 2311
rect 65057 2288 65143 2311
rect 64889 2248 64914 2288
rect 64914 2248 64954 2288
rect 64954 2248 64975 2288
rect 65057 2248 65078 2288
rect 65078 2248 65118 2288
rect 65118 2248 65143 2288
rect 64889 2225 64975 2248
rect 65057 2225 65143 2248
rect 80009 2288 80095 2311
rect 80177 2288 80263 2311
rect 80009 2248 80034 2288
rect 80034 2248 80074 2288
rect 80074 2248 80095 2288
rect 80177 2248 80198 2288
rect 80198 2248 80238 2288
rect 80238 2248 80263 2288
rect 80009 2225 80095 2248
rect 80177 2225 80263 2248
rect 95129 2288 95215 2311
rect 95297 2288 95383 2311
rect 95129 2248 95154 2288
rect 95154 2248 95194 2288
rect 95194 2248 95215 2288
rect 95297 2248 95318 2288
rect 95318 2248 95358 2288
rect 95358 2248 95383 2288
rect 95129 2225 95215 2248
rect 95297 2225 95383 2248
rect 3169 1532 3255 1555
rect 3337 1532 3423 1555
rect 3169 1492 3194 1532
rect 3194 1492 3234 1532
rect 3234 1492 3255 1532
rect 3337 1492 3358 1532
rect 3358 1492 3398 1532
rect 3398 1492 3423 1532
rect 3169 1469 3255 1492
rect 3337 1469 3423 1492
rect 18289 1532 18375 1555
rect 18457 1532 18543 1555
rect 18289 1492 18314 1532
rect 18314 1492 18354 1532
rect 18354 1492 18375 1532
rect 18457 1492 18478 1532
rect 18478 1492 18518 1532
rect 18518 1492 18543 1532
rect 18289 1469 18375 1492
rect 18457 1469 18543 1492
rect 33409 1532 33495 1555
rect 33577 1532 33663 1555
rect 33409 1492 33434 1532
rect 33434 1492 33474 1532
rect 33474 1492 33495 1532
rect 33577 1492 33598 1532
rect 33598 1492 33638 1532
rect 33638 1492 33663 1532
rect 33409 1469 33495 1492
rect 33577 1469 33663 1492
rect 48529 1532 48615 1555
rect 48697 1532 48783 1555
rect 48529 1492 48554 1532
rect 48554 1492 48594 1532
rect 48594 1492 48615 1532
rect 48697 1492 48718 1532
rect 48718 1492 48758 1532
rect 48758 1492 48783 1532
rect 48529 1469 48615 1492
rect 48697 1469 48783 1492
rect 63649 1532 63735 1555
rect 63817 1532 63903 1555
rect 63649 1492 63674 1532
rect 63674 1492 63714 1532
rect 63714 1492 63735 1532
rect 63817 1492 63838 1532
rect 63838 1492 63878 1532
rect 63878 1492 63903 1532
rect 63649 1469 63735 1492
rect 63817 1469 63903 1492
rect 78769 1532 78855 1555
rect 78937 1532 79023 1555
rect 78769 1492 78794 1532
rect 78794 1492 78834 1532
rect 78834 1492 78855 1532
rect 78937 1492 78958 1532
rect 78958 1492 78998 1532
rect 78998 1492 79023 1532
rect 78769 1469 78855 1492
rect 78937 1469 79023 1492
rect 93889 1532 93975 1555
rect 94057 1532 94143 1555
rect 93889 1492 93914 1532
rect 93914 1492 93954 1532
rect 93954 1492 93975 1532
rect 94057 1492 94078 1532
rect 94078 1492 94118 1532
rect 94118 1492 94143 1532
rect 93889 1469 93975 1492
rect 94057 1469 94143 1492
rect 4409 776 4495 799
rect 4577 776 4663 799
rect 4409 736 4434 776
rect 4434 736 4474 776
rect 4474 736 4495 776
rect 4577 736 4598 776
rect 4598 736 4638 776
rect 4638 736 4663 776
rect 4409 713 4495 736
rect 4577 713 4663 736
rect 19529 776 19615 799
rect 19697 776 19783 799
rect 19529 736 19554 776
rect 19554 736 19594 776
rect 19594 736 19615 776
rect 19697 736 19718 776
rect 19718 736 19758 776
rect 19758 736 19783 776
rect 19529 713 19615 736
rect 19697 713 19783 736
rect 34649 776 34735 799
rect 34817 776 34903 799
rect 34649 736 34674 776
rect 34674 736 34714 776
rect 34714 736 34735 776
rect 34817 736 34838 776
rect 34838 736 34878 776
rect 34878 736 34903 776
rect 34649 713 34735 736
rect 34817 713 34903 736
rect 49769 776 49855 799
rect 49937 776 50023 799
rect 49769 736 49794 776
rect 49794 736 49834 776
rect 49834 736 49855 776
rect 49937 736 49958 776
rect 49958 736 49998 776
rect 49998 736 50023 776
rect 49769 713 49855 736
rect 49937 713 50023 736
rect 64889 776 64975 799
rect 65057 776 65143 799
rect 64889 736 64914 776
rect 64914 736 64954 776
rect 64954 736 64975 776
rect 65057 736 65078 776
rect 65078 736 65118 776
rect 65118 736 65143 776
rect 64889 713 64975 736
rect 65057 713 65143 736
rect 80009 776 80095 799
rect 80177 776 80263 799
rect 80009 736 80034 776
rect 80034 736 80074 776
rect 80074 736 80095 776
rect 80177 736 80198 776
rect 80198 736 80238 776
rect 80238 736 80263 776
rect 80009 713 80095 736
rect 80177 713 80263 736
rect 95129 776 95215 799
rect 95297 776 95383 799
rect 95129 736 95154 776
rect 95154 736 95194 776
rect 95194 736 95215 776
rect 95297 736 95318 776
rect 95318 736 95358 776
rect 95358 736 95383 776
rect 95129 713 95215 736
rect 95297 713 95383 736
<< metal6 >>
rect 3076 81691 3516 81774
rect 3076 81605 3169 81691
rect 3255 81605 3337 81691
rect 3423 81605 3516 81691
rect 3076 80179 3516 81605
rect 3076 80093 3169 80179
rect 3255 80093 3337 80179
rect 3423 80093 3516 80179
rect 3076 78667 3516 80093
rect 3076 78581 3169 78667
rect 3255 78581 3337 78667
rect 3423 78581 3516 78667
rect 3076 77155 3516 78581
rect 3076 77069 3169 77155
rect 3255 77069 3337 77155
rect 3423 77069 3516 77155
rect 3076 75643 3516 77069
rect 3076 75557 3169 75643
rect 3255 75557 3337 75643
rect 3423 75557 3516 75643
rect 3076 74131 3516 75557
rect 3076 74045 3169 74131
rect 3255 74045 3337 74131
rect 3423 74045 3516 74131
rect 3076 72619 3516 74045
rect 3076 72533 3169 72619
rect 3255 72533 3337 72619
rect 3423 72533 3516 72619
rect 3076 71107 3516 72533
rect 3076 71021 3169 71107
rect 3255 71021 3337 71107
rect 3423 71021 3516 71107
rect 3076 69595 3516 71021
rect 3076 69509 3169 69595
rect 3255 69509 3337 69595
rect 3423 69509 3516 69595
rect 3076 68083 3516 69509
rect 3076 67997 3169 68083
rect 3255 67997 3337 68083
rect 3423 67997 3516 68083
rect 3076 66571 3516 67997
rect 3076 66485 3169 66571
rect 3255 66485 3337 66571
rect 3423 66485 3516 66571
rect 3076 65059 3516 66485
rect 3076 64973 3169 65059
rect 3255 64973 3337 65059
rect 3423 64973 3516 65059
rect 3076 63547 3516 64973
rect 3076 63461 3169 63547
rect 3255 63461 3337 63547
rect 3423 63461 3516 63547
rect 3076 62035 3516 63461
rect 3076 61949 3169 62035
rect 3255 61949 3337 62035
rect 3423 61949 3516 62035
rect 3076 60523 3516 61949
rect 3076 60437 3169 60523
rect 3255 60437 3337 60523
rect 3423 60437 3516 60523
rect 3076 59011 3516 60437
rect 3076 58925 3169 59011
rect 3255 58925 3337 59011
rect 3423 58925 3516 59011
rect 3076 57499 3516 58925
rect 3076 57413 3169 57499
rect 3255 57413 3337 57499
rect 3423 57413 3516 57499
rect 3076 55987 3516 57413
rect 3076 55901 3169 55987
rect 3255 55901 3337 55987
rect 3423 55901 3516 55987
rect 3076 54475 3516 55901
rect 3076 54389 3169 54475
rect 3255 54389 3337 54475
rect 3423 54389 3516 54475
rect 3076 52963 3516 54389
rect 3076 52877 3169 52963
rect 3255 52877 3337 52963
rect 3423 52877 3516 52963
rect 3076 51451 3516 52877
rect 3076 51365 3169 51451
rect 3255 51365 3337 51451
rect 3423 51365 3516 51451
rect 3076 49939 3516 51365
rect 3076 49853 3169 49939
rect 3255 49853 3337 49939
rect 3423 49853 3516 49939
rect 3076 48427 3516 49853
rect 3076 48341 3169 48427
rect 3255 48341 3337 48427
rect 3423 48341 3516 48427
rect 3076 46915 3516 48341
rect 3076 46829 3169 46915
rect 3255 46829 3337 46915
rect 3423 46829 3516 46915
rect 3076 45403 3516 46829
rect 3076 45317 3169 45403
rect 3255 45317 3337 45403
rect 3423 45317 3516 45403
rect 3076 43891 3516 45317
rect 3076 43805 3169 43891
rect 3255 43805 3337 43891
rect 3423 43805 3516 43891
rect 3076 42379 3516 43805
rect 3076 42293 3169 42379
rect 3255 42293 3337 42379
rect 3423 42293 3516 42379
rect 3076 40867 3516 42293
rect 3076 40781 3169 40867
rect 3255 40781 3337 40867
rect 3423 40781 3516 40867
rect 3076 39355 3516 40781
rect 3076 39269 3169 39355
rect 3255 39269 3337 39355
rect 3423 39269 3516 39355
rect 3076 37843 3516 39269
rect 3076 37757 3169 37843
rect 3255 37757 3337 37843
rect 3423 37757 3516 37843
rect 3076 36331 3516 37757
rect 3076 36245 3169 36331
rect 3255 36245 3337 36331
rect 3423 36245 3516 36331
rect 3076 34819 3516 36245
rect 3076 34733 3169 34819
rect 3255 34733 3337 34819
rect 3423 34733 3516 34819
rect 3076 33307 3516 34733
rect 3076 33221 3169 33307
rect 3255 33221 3337 33307
rect 3423 33221 3516 33307
rect 3076 31795 3516 33221
rect 3076 31709 3169 31795
rect 3255 31709 3337 31795
rect 3423 31709 3516 31795
rect 3076 30283 3516 31709
rect 3076 30197 3169 30283
rect 3255 30197 3337 30283
rect 3423 30197 3516 30283
rect 3076 28771 3516 30197
rect 3076 28685 3169 28771
rect 3255 28685 3337 28771
rect 3423 28685 3516 28771
rect 3076 27259 3516 28685
rect 3076 27173 3169 27259
rect 3255 27173 3337 27259
rect 3423 27173 3516 27259
rect 3076 25747 3516 27173
rect 3076 25661 3169 25747
rect 3255 25661 3337 25747
rect 3423 25661 3516 25747
rect 3076 24235 3516 25661
rect 3076 24149 3169 24235
rect 3255 24149 3337 24235
rect 3423 24149 3516 24235
rect 3076 22723 3516 24149
rect 3076 22637 3169 22723
rect 3255 22637 3337 22723
rect 3423 22637 3516 22723
rect 3076 21211 3516 22637
rect 3076 21125 3169 21211
rect 3255 21125 3337 21211
rect 3423 21125 3516 21211
rect 3076 19699 3516 21125
rect 3076 19613 3169 19699
rect 3255 19613 3337 19699
rect 3423 19613 3516 19699
rect 3076 18187 3516 19613
rect 3076 18101 3169 18187
rect 3255 18101 3337 18187
rect 3423 18101 3516 18187
rect 3076 16675 3516 18101
rect 3076 16589 3169 16675
rect 3255 16589 3337 16675
rect 3423 16589 3516 16675
rect 3076 15163 3516 16589
rect 3076 15077 3169 15163
rect 3255 15077 3337 15163
rect 3423 15077 3516 15163
rect 3076 13651 3516 15077
rect 3076 13565 3169 13651
rect 3255 13565 3337 13651
rect 3423 13565 3516 13651
rect 3076 12139 3516 13565
rect 3076 12053 3169 12139
rect 3255 12053 3337 12139
rect 3423 12053 3516 12139
rect 3076 10627 3516 12053
rect 3076 10541 3169 10627
rect 3255 10541 3337 10627
rect 3423 10541 3516 10627
rect 3076 9115 3516 10541
rect 3076 9029 3169 9115
rect 3255 9029 3337 9115
rect 3423 9029 3516 9115
rect 3076 7603 3516 9029
rect 3076 7517 3169 7603
rect 3255 7517 3337 7603
rect 3423 7517 3516 7603
rect 3076 6091 3516 7517
rect 3076 6005 3169 6091
rect 3255 6005 3337 6091
rect 3423 6005 3516 6091
rect 3076 4579 3516 6005
rect 3076 4493 3169 4579
rect 3255 4493 3337 4579
rect 3423 4493 3516 4579
rect 3076 3067 3516 4493
rect 3076 2981 3169 3067
rect 3255 2981 3337 3067
rect 3423 2981 3516 3067
rect 3076 1555 3516 2981
rect 3076 1469 3169 1555
rect 3255 1469 3337 1555
rect 3423 1469 3516 1555
rect 3076 712 3516 1469
rect 4316 80935 4756 81692
rect 4316 80849 4409 80935
rect 4495 80849 4577 80935
rect 4663 80849 4756 80935
rect 4316 79423 4756 80849
rect 4316 79337 4409 79423
rect 4495 79337 4577 79423
rect 4663 79337 4756 79423
rect 4316 77911 4756 79337
rect 4316 77825 4409 77911
rect 4495 77825 4577 77911
rect 4663 77825 4756 77911
rect 4316 76399 4756 77825
rect 4316 76313 4409 76399
rect 4495 76313 4577 76399
rect 4663 76313 4756 76399
rect 4316 74887 4756 76313
rect 4316 74801 4409 74887
rect 4495 74801 4577 74887
rect 4663 74801 4756 74887
rect 4316 73375 4756 74801
rect 4316 73289 4409 73375
rect 4495 73289 4577 73375
rect 4663 73289 4756 73375
rect 4316 71863 4756 73289
rect 4316 71777 4409 71863
rect 4495 71777 4577 71863
rect 4663 71777 4756 71863
rect 4316 70351 4756 71777
rect 4316 70265 4409 70351
rect 4495 70265 4577 70351
rect 4663 70265 4756 70351
rect 4316 68839 4756 70265
rect 4316 68753 4409 68839
rect 4495 68753 4577 68839
rect 4663 68753 4756 68839
rect 4316 67327 4756 68753
rect 4316 67241 4409 67327
rect 4495 67241 4577 67327
rect 4663 67241 4756 67327
rect 4316 65815 4756 67241
rect 4316 65729 4409 65815
rect 4495 65729 4577 65815
rect 4663 65729 4756 65815
rect 4316 64303 4756 65729
rect 4316 64217 4409 64303
rect 4495 64217 4577 64303
rect 4663 64217 4756 64303
rect 4316 62791 4756 64217
rect 4316 62705 4409 62791
rect 4495 62705 4577 62791
rect 4663 62705 4756 62791
rect 4316 61279 4756 62705
rect 4316 61193 4409 61279
rect 4495 61193 4577 61279
rect 4663 61193 4756 61279
rect 4316 59767 4756 61193
rect 4316 59681 4409 59767
rect 4495 59681 4577 59767
rect 4663 59681 4756 59767
rect 4316 58255 4756 59681
rect 4316 58169 4409 58255
rect 4495 58169 4577 58255
rect 4663 58169 4756 58255
rect 4316 56743 4756 58169
rect 4316 56657 4409 56743
rect 4495 56657 4577 56743
rect 4663 56657 4756 56743
rect 4316 55231 4756 56657
rect 4316 55145 4409 55231
rect 4495 55145 4577 55231
rect 4663 55145 4756 55231
rect 4316 53719 4756 55145
rect 4316 53633 4409 53719
rect 4495 53633 4577 53719
rect 4663 53633 4756 53719
rect 4316 52207 4756 53633
rect 4316 52121 4409 52207
rect 4495 52121 4577 52207
rect 4663 52121 4756 52207
rect 4316 50695 4756 52121
rect 4316 50609 4409 50695
rect 4495 50609 4577 50695
rect 4663 50609 4756 50695
rect 4316 49183 4756 50609
rect 4316 49097 4409 49183
rect 4495 49097 4577 49183
rect 4663 49097 4756 49183
rect 4316 47671 4756 49097
rect 4316 47585 4409 47671
rect 4495 47585 4577 47671
rect 4663 47585 4756 47671
rect 4316 46159 4756 47585
rect 4316 46073 4409 46159
rect 4495 46073 4577 46159
rect 4663 46073 4756 46159
rect 4316 44647 4756 46073
rect 4316 44561 4409 44647
rect 4495 44561 4577 44647
rect 4663 44561 4756 44647
rect 4316 43135 4756 44561
rect 4316 43049 4409 43135
rect 4495 43049 4577 43135
rect 4663 43049 4756 43135
rect 4316 41623 4756 43049
rect 4316 41537 4409 41623
rect 4495 41537 4577 41623
rect 4663 41537 4756 41623
rect 4316 40111 4756 41537
rect 4316 40025 4409 40111
rect 4495 40025 4577 40111
rect 4663 40025 4756 40111
rect 4316 38599 4756 40025
rect 4316 38513 4409 38599
rect 4495 38513 4577 38599
rect 4663 38513 4756 38599
rect 4316 37087 4756 38513
rect 4316 37001 4409 37087
rect 4495 37001 4577 37087
rect 4663 37001 4756 37087
rect 4316 35575 4756 37001
rect 4316 35489 4409 35575
rect 4495 35489 4577 35575
rect 4663 35489 4756 35575
rect 4316 34063 4756 35489
rect 4316 33977 4409 34063
rect 4495 33977 4577 34063
rect 4663 33977 4756 34063
rect 4316 32551 4756 33977
rect 4316 32465 4409 32551
rect 4495 32465 4577 32551
rect 4663 32465 4756 32551
rect 4316 31039 4756 32465
rect 4316 30953 4409 31039
rect 4495 30953 4577 31039
rect 4663 30953 4756 31039
rect 4316 29527 4756 30953
rect 4316 29441 4409 29527
rect 4495 29441 4577 29527
rect 4663 29441 4756 29527
rect 4316 28015 4756 29441
rect 4316 27929 4409 28015
rect 4495 27929 4577 28015
rect 4663 27929 4756 28015
rect 4316 26503 4756 27929
rect 4316 26417 4409 26503
rect 4495 26417 4577 26503
rect 4663 26417 4756 26503
rect 4316 24991 4756 26417
rect 4316 24905 4409 24991
rect 4495 24905 4577 24991
rect 4663 24905 4756 24991
rect 4316 23479 4756 24905
rect 4316 23393 4409 23479
rect 4495 23393 4577 23479
rect 4663 23393 4756 23479
rect 4316 21967 4756 23393
rect 4316 21881 4409 21967
rect 4495 21881 4577 21967
rect 4663 21881 4756 21967
rect 4316 20455 4756 21881
rect 4316 20369 4409 20455
rect 4495 20369 4577 20455
rect 4663 20369 4756 20455
rect 4316 18943 4756 20369
rect 4316 18857 4409 18943
rect 4495 18857 4577 18943
rect 4663 18857 4756 18943
rect 4316 17431 4756 18857
rect 4316 17345 4409 17431
rect 4495 17345 4577 17431
rect 4663 17345 4756 17431
rect 4316 15919 4756 17345
rect 4316 15833 4409 15919
rect 4495 15833 4577 15919
rect 4663 15833 4756 15919
rect 4316 14407 4756 15833
rect 4316 14321 4409 14407
rect 4495 14321 4577 14407
rect 4663 14321 4756 14407
rect 4316 12895 4756 14321
rect 4316 12809 4409 12895
rect 4495 12809 4577 12895
rect 4663 12809 4756 12895
rect 4316 11383 4756 12809
rect 4316 11297 4409 11383
rect 4495 11297 4577 11383
rect 4663 11297 4756 11383
rect 4316 9871 4756 11297
rect 4316 9785 4409 9871
rect 4495 9785 4577 9871
rect 4663 9785 4756 9871
rect 4316 8359 4756 9785
rect 4316 8273 4409 8359
rect 4495 8273 4577 8359
rect 4663 8273 4756 8359
rect 4316 6847 4756 8273
rect 4316 6761 4409 6847
rect 4495 6761 4577 6847
rect 4663 6761 4756 6847
rect 4316 5335 4756 6761
rect 4316 5249 4409 5335
rect 4495 5249 4577 5335
rect 4663 5249 4756 5335
rect 4316 3823 4756 5249
rect 4316 3737 4409 3823
rect 4495 3737 4577 3823
rect 4663 3737 4756 3823
rect 4316 2311 4756 3737
rect 4316 2225 4409 2311
rect 4495 2225 4577 2311
rect 4663 2225 4756 2311
rect 4316 799 4756 2225
rect 4316 713 4409 799
rect 4495 713 4577 799
rect 4663 713 4756 799
rect 4316 630 4756 713
rect 18196 81691 18636 81774
rect 18196 81605 18289 81691
rect 18375 81605 18457 81691
rect 18543 81605 18636 81691
rect 18196 80179 18636 81605
rect 18196 80093 18289 80179
rect 18375 80093 18457 80179
rect 18543 80093 18636 80179
rect 18196 78667 18636 80093
rect 18196 78581 18289 78667
rect 18375 78581 18457 78667
rect 18543 78581 18636 78667
rect 18196 77155 18636 78581
rect 18196 77069 18289 77155
rect 18375 77069 18457 77155
rect 18543 77069 18636 77155
rect 18196 75643 18636 77069
rect 18196 75557 18289 75643
rect 18375 75557 18457 75643
rect 18543 75557 18636 75643
rect 18196 74131 18636 75557
rect 18196 74045 18289 74131
rect 18375 74045 18457 74131
rect 18543 74045 18636 74131
rect 18196 72619 18636 74045
rect 18196 72533 18289 72619
rect 18375 72533 18457 72619
rect 18543 72533 18636 72619
rect 18196 71107 18636 72533
rect 18196 71021 18289 71107
rect 18375 71021 18457 71107
rect 18543 71021 18636 71107
rect 18196 69595 18636 71021
rect 18196 69509 18289 69595
rect 18375 69509 18457 69595
rect 18543 69509 18636 69595
rect 18196 68083 18636 69509
rect 18196 67997 18289 68083
rect 18375 67997 18457 68083
rect 18543 67997 18636 68083
rect 18196 66571 18636 67997
rect 18196 66485 18289 66571
rect 18375 66485 18457 66571
rect 18543 66485 18636 66571
rect 18196 65059 18636 66485
rect 18196 64973 18289 65059
rect 18375 64973 18457 65059
rect 18543 64973 18636 65059
rect 18196 63547 18636 64973
rect 18196 63461 18289 63547
rect 18375 63461 18457 63547
rect 18543 63461 18636 63547
rect 18196 62035 18636 63461
rect 18196 61949 18289 62035
rect 18375 61949 18457 62035
rect 18543 61949 18636 62035
rect 18196 60523 18636 61949
rect 18196 60437 18289 60523
rect 18375 60437 18457 60523
rect 18543 60437 18636 60523
rect 18196 59011 18636 60437
rect 18196 58925 18289 59011
rect 18375 58925 18457 59011
rect 18543 58925 18636 59011
rect 18196 57499 18636 58925
rect 18196 57413 18289 57499
rect 18375 57413 18457 57499
rect 18543 57413 18636 57499
rect 18196 55987 18636 57413
rect 18196 55901 18289 55987
rect 18375 55901 18457 55987
rect 18543 55901 18636 55987
rect 18196 54475 18636 55901
rect 18196 54389 18289 54475
rect 18375 54389 18457 54475
rect 18543 54389 18636 54475
rect 18196 52963 18636 54389
rect 18196 52877 18289 52963
rect 18375 52877 18457 52963
rect 18543 52877 18636 52963
rect 18196 51451 18636 52877
rect 18196 51365 18289 51451
rect 18375 51365 18457 51451
rect 18543 51365 18636 51451
rect 18196 49939 18636 51365
rect 18196 49853 18289 49939
rect 18375 49853 18457 49939
rect 18543 49853 18636 49939
rect 18196 48427 18636 49853
rect 18196 48341 18289 48427
rect 18375 48341 18457 48427
rect 18543 48341 18636 48427
rect 18196 46915 18636 48341
rect 18196 46829 18289 46915
rect 18375 46829 18457 46915
rect 18543 46829 18636 46915
rect 18196 45403 18636 46829
rect 18196 45317 18289 45403
rect 18375 45317 18457 45403
rect 18543 45317 18636 45403
rect 18196 43891 18636 45317
rect 18196 43805 18289 43891
rect 18375 43805 18457 43891
rect 18543 43805 18636 43891
rect 18196 42379 18636 43805
rect 18196 42293 18289 42379
rect 18375 42293 18457 42379
rect 18543 42293 18636 42379
rect 18196 40867 18636 42293
rect 18196 40781 18289 40867
rect 18375 40781 18457 40867
rect 18543 40781 18636 40867
rect 18196 39355 18636 40781
rect 18196 39269 18289 39355
rect 18375 39269 18457 39355
rect 18543 39269 18636 39355
rect 18196 37843 18636 39269
rect 18196 37757 18289 37843
rect 18375 37757 18457 37843
rect 18543 37757 18636 37843
rect 18196 36331 18636 37757
rect 18196 36245 18289 36331
rect 18375 36245 18457 36331
rect 18543 36245 18636 36331
rect 18196 34819 18636 36245
rect 18196 34733 18289 34819
rect 18375 34733 18457 34819
rect 18543 34733 18636 34819
rect 18196 33307 18636 34733
rect 18196 33221 18289 33307
rect 18375 33221 18457 33307
rect 18543 33221 18636 33307
rect 18196 31795 18636 33221
rect 18196 31709 18289 31795
rect 18375 31709 18457 31795
rect 18543 31709 18636 31795
rect 18196 30283 18636 31709
rect 18196 30197 18289 30283
rect 18375 30197 18457 30283
rect 18543 30197 18636 30283
rect 18196 28771 18636 30197
rect 18196 28685 18289 28771
rect 18375 28685 18457 28771
rect 18543 28685 18636 28771
rect 18196 27259 18636 28685
rect 18196 27173 18289 27259
rect 18375 27173 18457 27259
rect 18543 27173 18636 27259
rect 18196 25747 18636 27173
rect 18196 25661 18289 25747
rect 18375 25661 18457 25747
rect 18543 25661 18636 25747
rect 18196 24235 18636 25661
rect 18196 24149 18289 24235
rect 18375 24149 18457 24235
rect 18543 24149 18636 24235
rect 18196 22723 18636 24149
rect 18196 22637 18289 22723
rect 18375 22637 18457 22723
rect 18543 22637 18636 22723
rect 18196 21211 18636 22637
rect 18196 21125 18289 21211
rect 18375 21125 18457 21211
rect 18543 21125 18636 21211
rect 18196 19699 18636 21125
rect 18196 19613 18289 19699
rect 18375 19613 18457 19699
rect 18543 19613 18636 19699
rect 18196 18187 18636 19613
rect 18196 18101 18289 18187
rect 18375 18101 18457 18187
rect 18543 18101 18636 18187
rect 18196 16675 18636 18101
rect 18196 16589 18289 16675
rect 18375 16589 18457 16675
rect 18543 16589 18636 16675
rect 18196 15163 18636 16589
rect 18196 15077 18289 15163
rect 18375 15077 18457 15163
rect 18543 15077 18636 15163
rect 18196 13651 18636 15077
rect 18196 13565 18289 13651
rect 18375 13565 18457 13651
rect 18543 13565 18636 13651
rect 18196 12139 18636 13565
rect 18196 12053 18289 12139
rect 18375 12053 18457 12139
rect 18543 12053 18636 12139
rect 18196 10627 18636 12053
rect 18196 10541 18289 10627
rect 18375 10541 18457 10627
rect 18543 10541 18636 10627
rect 18196 9115 18636 10541
rect 18196 9029 18289 9115
rect 18375 9029 18457 9115
rect 18543 9029 18636 9115
rect 18196 7603 18636 9029
rect 18196 7517 18289 7603
rect 18375 7517 18457 7603
rect 18543 7517 18636 7603
rect 18196 6091 18636 7517
rect 18196 6005 18289 6091
rect 18375 6005 18457 6091
rect 18543 6005 18636 6091
rect 18196 4579 18636 6005
rect 18196 4493 18289 4579
rect 18375 4493 18457 4579
rect 18543 4493 18636 4579
rect 18196 3067 18636 4493
rect 18196 2981 18289 3067
rect 18375 2981 18457 3067
rect 18543 2981 18636 3067
rect 18196 1555 18636 2981
rect 18196 1469 18289 1555
rect 18375 1469 18457 1555
rect 18543 1469 18636 1555
rect 18196 712 18636 1469
rect 19436 80935 19876 81692
rect 19436 80849 19529 80935
rect 19615 80849 19697 80935
rect 19783 80849 19876 80935
rect 19436 79423 19876 80849
rect 19436 79337 19529 79423
rect 19615 79337 19697 79423
rect 19783 79337 19876 79423
rect 19436 77911 19876 79337
rect 19436 77825 19529 77911
rect 19615 77825 19697 77911
rect 19783 77825 19876 77911
rect 19436 76399 19876 77825
rect 19436 76313 19529 76399
rect 19615 76313 19697 76399
rect 19783 76313 19876 76399
rect 19436 74887 19876 76313
rect 19436 74801 19529 74887
rect 19615 74801 19697 74887
rect 19783 74801 19876 74887
rect 19436 73375 19876 74801
rect 19436 73289 19529 73375
rect 19615 73289 19697 73375
rect 19783 73289 19876 73375
rect 19436 71863 19876 73289
rect 19436 71777 19529 71863
rect 19615 71777 19697 71863
rect 19783 71777 19876 71863
rect 19436 70351 19876 71777
rect 19436 70265 19529 70351
rect 19615 70265 19697 70351
rect 19783 70265 19876 70351
rect 19436 68839 19876 70265
rect 19436 68753 19529 68839
rect 19615 68753 19697 68839
rect 19783 68753 19876 68839
rect 19436 67327 19876 68753
rect 19436 67241 19529 67327
rect 19615 67241 19697 67327
rect 19783 67241 19876 67327
rect 19436 65815 19876 67241
rect 19436 65729 19529 65815
rect 19615 65729 19697 65815
rect 19783 65729 19876 65815
rect 19436 64303 19876 65729
rect 19436 64217 19529 64303
rect 19615 64217 19697 64303
rect 19783 64217 19876 64303
rect 19436 62791 19876 64217
rect 19436 62705 19529 62791
rect 19615 62705 19697 62791
rect 19783 62705 19876 62791
rect 19436 61279 19876 62705
rect 19436 61193 19529 61279
rect 19615 61193 19697 61279
rect 19783 61193 19876 61279
rect 19436 59767 19876 61193
rect 19436 59681 19529 59767
rect 19615 59681 19697 59767
rect 19783 59681 19876 59767
rect 19436 58255 19876 59681
rect 19436 58169 19529 58255
rect 19615 58169 19697 58255
rect 19783 58169 19876 58255
rect 19436 56743 19876 58169
rect 19436 56657 19529 56743
rect 19615 56657 19697 56743
rect 19783 56657 19876 56743
rect 19436 55231 19876 56657
rect 19436 55145 19529 55231
rect 19615 55145 19697 55231
rect 19783 55145 19876 55231
rect 19436 53719 19876 55145
rect 19436 53633 19529 53719
rect 19615 53633 19697 53719
rect 19783 53633 19876 53719
rect 19436 52207 19876 53633
rect 19436 52121 19529 52207
rect 19615 52121 19697 52207
rect 19783 52121 19876 52207
rect 19436 50695 19876 52121
rect 19436 50609 19529 50695
rect 19615 50609 19697 50695
rect 19783 50609 19876 50695
rect 19436 49183 19876 50609
rect 19436 49097 19529 49183
rect 19615 49097 19697 49183
rect 19783 49097 19876 49183
rect 19436 47671 19876 49097
rect 19436 47585 19529 47671
rect 19615 47585 19697 47671
rect 19783 47585 19876 47671
rect 19436 46159 19876 47585
rect 19436 46073 19529 46159
rect 19615 46073 19697 46159
rect 19783 46073 19876 46159
rect 19436 44647 19876 46073
rect 19436 44561 19529 44647
rect 19615 44561 19697 44647
rect 19783 44561 19876 44647
rect 19436 43135 19876 44561
rect 19436 43049 19529 43135
rect 19615 43049 19697 43135
rect 19783 43049 19876 43135
rect 19436 41623 19876 43049
rect 19436 41537 19529 41623
rect 19615 41537 19697 41623
rect 19783 41537 19876 41623
rect 19436 40111 19876 41537
rect 19436 40025 19529 40111
rect 19615 40025 19697 40111
rect 19783 40025 19876 40111
rect 19436 38599 19876 40025
rect 19436 38513 19529 38599
rect 19615 38513 19697 38599
rect 19783 38513 19876 38599
rect 19436 37087 19876 38513
rect 19436 37001 19529 37087
rect 19615 37001 19697 37087
rect 19783 37001 19876 37087
rect 19436 35575 19876 37001
rect 19436 35489 19529 35575
rect 19615 35489 19697 35575
rect 19783 35489 19876 35575
rect 19436 34063 19876 35489
rect 19436 33977 19529 34063
rect 19615 33977 19697 34063
rect 19783 33977 19876 34063
rect 19436 32551 19876 33977
rect 19436 32465 19529 32551
rect 19615 32465 19697 32551
rect 19783 32465 19876 32551
rect 19436 31039 19876 32465
rect 19436 30953 19529 31039
rect 19615 30953 19697 31039
rect 19783 30953 19876 31039
rect 19436 29527 19876 30953
rect 19436 29441 19529 29527
rect 19615 29441 19697 29527
rect 19783 29441 19876 29527
rect 19436 28015 19876 29441
rect 19436 27929 19529 28015
rect 19615 27929 19697 28015
rect 19783 27929 19876 28015
rect 19436 26503 19876 27929
rect 19436 26417 19529 26503
rect 19615 26417 19697 26503
rect 19783 26417 19876 26503
rect 19436 24991 19876 26417
rect 19436 24905 19529 24991
rect 19615 24905 19697 24991
rect 19783 24905 19876 24991
rect 19436 23479 19876 24905
rect 19436 23393 19529 23479
rect 19615 23393 19697 23479
rect 19783 23393 19876 23479
rect 19436 21967 19876 23393
rect 19436 21881 19529 21967
rect 19615 21881 19697 21967
rect 19783 21881 19876 21967
rect 19436 20455 19876 21881
rect 19436 20369 19529 20455
rect 19615 20369 19697 20455
rect 19783 20369 19876 20455
rect 19436 18943 19876 20369
rect 19436 18857 19529 18943
rect 19615 18857 19697 18943
rect 19783 18857 19876 18943
rect 19436 17431 19876 18857
rect 19436 17345 19529 17431
rect 19615 17345 19697 17431
rect 19783 17345 19876 17431
rect 19436 15919 19876 17345
rect 19436 15833 19529 15919
rect 19615 15833 19697 15919
rect 19783 15833 19876 15919
rect 19436 14407 19876 15833
rect 19436 14321 19529 14407
rect 19615 14321 19697 14407
rect 19783 14321 19876 14407
rect 19436 12895 19876 14321
rect 19436 12809 19529 12895
rect 19615 12809 19697 12895
rect 19783 12809 19876 12895
rect 19436 11383 19876 12809
rect 19436 11297 19529 11383
rect 19615 11297 19697 11383
rect 19783 11297 19876 11383
rect 19436 9871 19876 11297
rect 19436 9785 19529 9871
rect 19615 9785 19697 9871
rect 19783 9785 19876 9871
rect 19436 8359 19876 9785
rect 19436 8273 19529 8359
rect 19615 8273 19697 8359
rect 19783 8273 19876 8359
rect 19436 6847 19876 8273
rect 19436 6761 19529 6847
rect 19615 6761 19697 6847
rect 19783 6761 19876 6847
rect 19436 5335 19876 6761
rect 19436 5249 19529 5335
rect 19615 5249 19697 5335
rect 19783 5249 19876 5335
rect 19436 3823 19876 5249
rect 19436 3737 19529 3823
rect 19615 3737 19697 3823
rect 19783 3737 19876 3823
rect 19436 2311 19876 3737
rect 19436 2225 19529 2311
rect 19615 2225 19697 2311
rect 19783 2225 19876 2311
rect 19436 799 19876 2225
rect 19436 713 19529 799
rect 19615 713 19697 799
rect 19783 713 19876 799
rect 19436 630 19876 713
rect 33316 81691 33756 81774
rect 33316 81605 33409 81691
rect 33495 81605 33577 81691
rect 33663 81605 33756 81691
rect 33316 80179 33756 81605
rect 33316 80093 33409 80179
rect 33495 80093 33577 80179
rect 33663 80093 33756 80179
rect 33316 78667 33756 80093
rect 33316 78581 33409 78667
rect 33495 78581 33577 78667
rect 33663 78581 33756 78667
rect 33316 77155 33756 78581
rect 33316 77069 33409 77155
rect 33495 77069 33577 77155
rect 33663 77069 33756 77155
rect 33316 75643 33756 77069
rect 33316 75557 33409 75643
rect 33495 75557 33577 75643
rect 33663 75557 33756 75643
rect 33316 74131 33756 75557
rect 33316 74045 33409 74131
rect 33495 74045 33577 74131
rect 33663 74045 33756 74131
rect 33316 72619 33756 74045
rect 33316 72533 33409 72619
rect 33495 72533 33577 72619
rect 33663 72533 33756 72619
rect 33316 71107 33756 72533
rect 33316 71021 33409 71107
rect 33495 71021 33577 71107
rect 33663 71021 33756 71107
rect 33316 69595 33756 71021
rect 33316 69509 33409 69595
rect 33495 69509 33577 69595
rect 33663 69509 33756 69595
rect 33316 68083 33756 69509
rect 33316 67997 33409 68083
rect 33495 67997 33577 68083
rect 33663 67997 33756 68083
rect 33316 66571 33756 67997
rect 33316 66485 33409 66571
rect 33495 66485 33577 66571
rect 33663 66485 33756 66571
rect 33316 65059 33756 66485
rect 33316 64973 33409 65059
rect 33495 64973 33577 65059
rect 33663 64973 33756 65059
rect 33316 63547 33756 64973
rect 33316 63461 33409 63547
rect 33495 63461 33577 63547
rect 33663 63461 33756 63547
rect 33316 62035 33756 63461
rect 33316 61949 33409 62035
rect 33495 61949 33577 62035
rect 33663 61949 33756 62035
rect 33316 60523 33756 61949
rect 33316 60437 33409 60523
rect 33495 60437 33577 60523
rect 33663 60437 33756 60523
rect 33316 59011 33756 60437
rect 33316 58925 33409 59011
rect 33495 58925 33577 59011
rect 33663 58925 33756 59011
rect 33316 57499 33756 58925
rect 33316 57413 33409 57499
rect 33495 57413 33577 57499
rect 33663 57413 33756 57499
rect 33316 55987 33756 57413
rect 33316 55901 33409 55987
rect 33495 55901 33577 55987
rect 33663 55901 33756 55987
rect 33316 54475 33756 55901
rect 33316 54389 33409 54475
rect 33495 54389 33577 54475
rect 33663 54389 33756 54475
rect 33316 52963 33756 54389
rect 33316 52877 33409 52963
rect 33495 52877 33577 52963
rect 33663 52877 33756 52963
rect 33316 51451 33756 52877
rect 33316 51365 33409 51451
rect 33495 51365 33577 51451
rect 33663 51365 33756 51451
rect 33316 49939 33756 51365
rect 33316 49853 33409 49939
rect 33495 49853 33577 49939
rect 33663 49853 33756 49939
rect 33316 48427 33756 49853
rect 33316 48341 33409 48427
rect 33495 48341 33577 48427
rect 33663 48341 33756 48427
rect 33316 46915 33756 48341
rect 33316 46829 33409 46915
rect 33495 46829 33577 46915
rect 33663 46829 33756 46915
rect 33316 45403 33756 46829
rect 33316 45317 33409 45403
rect 33495 45317 33577 45403
rect 33663 45317 33756 45403
rect 33316 43891 33756 45317
rect 33316 43805 33409 43891
rect 33495 43805 33577 43891
rect 33663 43805 33756 43891
rect 33316 42379 33756 43805
rect 33316 42293 33409 42379
rect 33495 42293 33577 42379
rect 33663 42293 33756 42379
rect 33316 40867 33756 42293
rect 33316 40781 33409 40867
rect 33495 40781 33577 40867
rect 33663 40781 33756 40867
rect 33316 39355 33756 40781
rect 33316 39269 33409 39355
rect 33495 39269 33577 39355
rect 33663 39269 33756 39355
rect 33316 37843 33756 39269
rect 33316 37757 33409 37843
rect 33495 37757 33577 37843
rect 33663 37757 33756 37843
rect 33316 36331 33756 37757
rect 33316 36245 33409 36331
rect 33495 36245 33577 36331
rect 33663 36245 33756 36331
rect 33316 34819 33756 36245
rect 33316 34733 33409 34819
rect 33495 34733 33577 34819
rect 33663 34733 33756 34819
rect 33316 33307 33756 34733
rect 33316 33221 33409 33307
rect 33495 33221 33577 33307
rect 33663 33221 33756 33307
rect 33316 31795 33756 33221
rect 33316 31709 33409 31795
rect 33495 31709 33577 31795
rect 33663 31709 33756 31795
rect 33316 30283 33756 31709
rect 33316 30197 33409 30283
rect 33495 30197 33577 30283
rect 33663 30197 33756 30283
rect 33316 28771 33756 30197
rect 33316 28685 33409 28771
rect 33495 28685 33577 28771
rect 33663 28685 33756 28771
rect 33316 27259 33756 28685
rect 33316 27173 33409 27259
rect 33495 27173 33577 27259
rect 33663 27173 33756 27259
rect 33316 25747 33756 27173
rect 33316 25661 33409 25747
rect 33495 25661 33577 25747
rect 33663 25661 33756 25747
rect 33316 24235 33756 25661
rect 33316 24149 33409 24235
rect 33495 24149 33577 24235
rect 33663 24149 33756 24235
rect 33316 22723 33756 24149
rect 33316 22637 33409 22723
rect 33495 22637 33577 22723
rect 33663 22637 33756 22723
rect 33316 21211 33756 22637
rect 33316 21125 33409 21211
rect 33495 21125 33577 21211
rect 33663 21125 33756 21211
rect 33316 19699 33756 21125
rect 33316 19613 33409 19699
rect 33495 19613 33577 19699
rect 33663 19613 33756 19699
rect 33316 18187 33756 19613
rect 33316 18101 33409 18187
rect 33495 18101 33577 18187
rect 33663 18101 33756 18187
rect 33316 16675 33756 18101
rect 33316 16589 33409 16675
rect 33495 16589 33577 16675
rect 33663 16589 33756 16675
rect 33316 15163 33756 16589
rect 33316 15077 33409 15163
rect 33495 15077 33577 15163
rect 33663 15077 33756 15163
rect 33316 13651 33756 15077
rect 33316 13565 33409 13651
rect 33495 13565 33577 13651
rect 33663 13565 33756 13651
rect 33316 12139 33756 13565
rect 33316 12053 33409 12139
rect 33495 12053 33577 12139
rect 33663 12053 33756 12139
rect 33316 10627 33756 12053
rect 33316 10541 33409 10627
rect 33495 10541 33577 10627
rect 33663 10541 33756 10627
rect 33316 9115 33756 10541
rect 33316 9029 33409 9115
rect 33495 9029 33577 9115
rect 33663 9029 33756 9115
rect 33316 7603 33756 9029
rect 33316 7517 33409 7603
rect 33495 7517 33577 7603
rect 33663 7517 33756 7603
rect 33316 6091 33756 7517
rect 33316 6005 33409 6091
rect 33495 6005 33577 6091
rect 33663 6005 33756 6091
rect 33316 4579 33756 6005
rect 33316 4493 33409 4579
rect 33495 4493 33577 4579
rect 33663 4493 33756 4579
rect 33316 3067 33756 4493
rect 33316 2981 33409 3067
rect 33495 2981 33577 3067
rect 33663 2981 33756 3067
rect 33316 1555 33756 2981
rect 33316 1469 33409 1555
rect 33495 1469 33577 1555
rect 33663 1469 33756 1555
rect 33316 712 33756 1469
rect 34556 80935 34996 81692
rect 34556 80849 34649 80935
rect 34735 80849 34817 80935
rect 34903 80849 34996 80935
rect 34556 79423 34996 80849
rect 34556 79337 34649 79423
rect 34735 79337 34817 79423
rect 34903 79337 34996 79423
rect 34556 77911 34996 79337
rect 34556 77825 34649 77911
rect 34735 77825 34817 77911
rect 34903 77825 34996 77911
rect 34556 76399 34996 77825
rect 34556 76313 34649 76399
rect 34735 76313 34817 76399
rect 34903 76313 34996 76399
rect 34556 74887 34996 76313
rect 34556 74801 34649 74887
rect 34735 74801 34817 74887
rect 34903 74801 34996 74887
rect 34556 73375 34996 74801
rect 34556 73289 34649 73375
rect 34735 73289 34817 73375
rect 34903 73289 34996 73375
rect 34556 71863 34996 73289
rect 34556 71777 34649 71863
rect 34735 71777 34817 71863
rect 34903 71777 34996 71863
rect 34556 70351 34996 71777
rect 34556 70265 34649 70351
rect 34735 70265 34817 70351
rect 34903 70265 34996 70351
rect 34556 68839 34996 70265
rect 34556 68753 34649 68839
rect 34735 68753 34817 68839
rect 34903 68753 34996 68839
rect 34556 67327 34996 68753
rect 34556 67241 34649 67327
rect 34735 67241 34817 67327
rect 34903 67241 34996 67327
rect 34556 65815 34996 67241
rect 34556 65729 34649 65815
rect 34735 65729 34817 65815
rect 34903 65729 34996 65815
rect 34556 64303 34996 65729
rect 34556 64217 34649 64303
rect 34735 64217 34817 64303
rect 34903 64217 34996 64303
rect 34556 62791 34996 64217
rect 34556 62705 34649 62791
rect 34735 62705 34817 62791
rect 34903 62705 34996 62791
rect 34556 61279 34996 62705
rect 34556 61193 34649 61279
rect 34735 61193 34817 61279
rect 34903 61193 34996 61279
rect 34556 59767 34996 61193
rect 34556 59681 34649 59767
rect 34735 59681 34817 59767
rect 34903 59681 34996 59767
rect 34556 58255 34996 59681
rect 34556 58169 34649 58255
rect 34735 58169 34817 58255
rect 34903 58169 34996 58255
rect 34556 56743 34996 58169
rect 34556 56657 34649 56743
rect 34735 56657 34817 56743
rect 34903 56657 34996 56743
rect 34556 55231 34996 56657
rect 34556 55145 34649 55231
rect 34735 55145 34817 55231
rect 34903 55145 34996 55231
rect 34556 53719 34996 55145
rect 34556 53633 34649 53719
rect 34735 53633 34817 53719
rect 34903 53633 34996 53719
rect 34556 52207 34996 53633
rect 34556 52121 34649 52207
rect 34735 52121 34817 52207
rect 34903 52121 34996 52207
rect 34556 50695 34996 52121
rect 34556 50609 34649 50695
rect 34735 50609 34817 50695
rect 34903 50609 34996 50695
rect 34556 49183 34996 50609
rect 34556 49097 34649 49183
rect 34735 49097 34817 49183
rect 34903 49097 34996 49183
rect 34556 47671 34996 49097
rect 34556 47585 34649 47671
rect 34735 47585 34817 47671
rect 34903 47585 34996 47671
rect 34556 46159 34996 47585
rect 34556 46073 34649 46159
rect 34735 46073 34817 46159
rect 34903 46073 34996 46159
rect 34556 44647 34996 46073
rect 34556 44561 34649 44647
rect 34735 44561 34817 44647
rect 34903 44561 34996 44647
rect 34556 43135 34996 44561
rect 34556 43049 34649 43135
rect 34735 43049 34817 43135
rect 34903 43049 34996 43135
rect 34556 41623 34996 43049
rect 34556 41537 34649 41623
rect 34735 41537 34817 41623
rect 34903 41537 34996 41623
rect 34556 40111 34996 41537
rect 34556 40025 34649 40111
rect 34735 40025 34817 40111
rect 34903 40025 34996 40111
rect 34556 38599 34996 40025
rect 34556 38513 34649 38599
rect 34735 38513 34817 38599
rect 34903 38513 34996 38599
rect 34556 37087 34996 38513
rect 34556 37001 34649 37087
rect 34735 37001 34817 37087
rect 34903 37001 34996 37087
rect 34556 35575 34996 37001
rect 34556 35489 34649 35575
rect 34735 35489 34817 35575
rect 34903 35489 34996 35575
rect 34556 34063 34996 35489
rect 34556 33977 34649 34063
rect 34735 33977 34817 34063
rect 34903 33977 34996 34063
rect 34556 32551 34996 33977
rect 34556 32465 34649 32551
rect 34735 32465 34817 32551
rect 34903 32465 34996 32551
rect 34556 31039 34996 32465
rect 34556 30953 34649 31039
rect 34735 30953 34817 31039
rect 34903 30953 34996 31039
rect 34556 29527 34996 30953
rect 34556 29441 34649 29527
rect 34735 29441 34817 29527
rect 34903 29441 34996 29527
rect 34556 28015 34996 29441
rect 34556 27929 34649 28015
rect 34735 27929 34817 28015
rect 34903 27929 34996 28015
rect 34556 26503 34996 27929
rect 34556 26417 34649 26503
rect 34735 26417 34817 26503
rect 34903 26417 34996 26503
rect 34556 24991 34996 26417
rect 34556 24905 34649 24991
rect 34735 24905 34817 24991
rect 34903 24905 34996 24991
rect 34556 23479 34996 24905
rect 34556 23393 34649 23479
rect 34735 23393 34817 23479
rect 34903 23393 34996 23479
rect 34556 21967 34996 23393
rect 34556 21881 34649 21967
rect 34735 21881 34817 21967
rect 34903 21881 34996 21967
rect 34556 20455 34996 21881
rect 34556 20369 34649 20455
rect 34735 20369 34817 20455
rect 34903 20369 34996 20455
rect 34556 18943 34996 20369
rect 34556 18857 34649 18943
rect 34735 18857 34817 18943
rect 34903 18857 34996 18943
rect 34556 17431 34996 18857
rect 34556 17345 34649 17431
rect 34735 17345 34817 17431
rect 34903 17345 34996 17431
rect 34556 15919 34996 17345
rect 34556 15833 34649 15919
rect 34735 15833 34817 15919
rect 34903 15833 34996 15919
rect 34556 14407 34996 15833
rect 34556 14321 34649 14407
rect 34735 14321 34817 14407
rect 34903 14321 34996 14407
rect 34556 12895 34996 14321
rect 34556 12809 34649 12895
rect 34735 12809 34817 12895
rect 34903 12809 34996 12895
rect 34556 11383 34996 12809
rect 34556 11297 34649 11383
rect 34735 11297 34817 11383
rect 34903 11297 34996 11383
rect 34556 9871 34996 11297
rect 34556 9785 34649 9871
rect 34735 9785 34817 9871
rect 34903 9785 34996 9871
rect 34556 8359 34996 9785
rect 34556 8273 34649 8359
rect 34735 8273 34817 8359
rect 34903 8273 34996 8359
rect 34556 6847 34996 8273
rect 34556 6761 34649 6847
rect 34735 6761 34817 6847
rect 34903 6761 34996 6847
rect 34556 5335 34996 6761
rect 34556 5249 34649 5335
rect 34735 5249 34817 5335
rect 34903 5249 34996 5335
rect 34556 3823 34996 5249
rect 34556 3737 34649 3823
rect 34735 3737 34817 3823
rect 34903 3737 34996 3823
rect 34556 2311 34996 3737
rect 34556 2225 34649 2311
rect 34735 2225 34817 2311
rect 34903 2225 34996 2311
rect 34556 799 34996 2225
rect 34556 713 34649 799
rect 34735 713 34817 799
rect 34903 713 34996 799
rect 34556 630 34996 713
rect 48436 81691 48876 81774
rect 48436 81605 48529 81691
rect 48615 81605 48697 81691
rect 48783 81605 48876 81691
rect 48436 80179 48876 81605
rect 48436 80093 48529 80179
rect 48615 80093 48697 80179
rect 48783 80093 48876 80179
rect 48436 78667 48876 80093
rect 48436 78581 48529 78667
rect 48615 78581 48697 78667
rect 48783 78581 48876 78667
rect 48436 77155 48876 78581
rect 48436 77069 48529 77155
rect 48615 77069 48697 77155
rect 48783 77069 48876 77155
rect 48436 75643 48876 77069
rect 48436 75557 48529 75643
rect 48615 75557 48697 75643
rect 48783 75557 48876 75643
rect 48436 74131 48876 75557
rect 48436 74045 48529 74131
rect 48615 74045 48697 74131
rect 48783 74045 48876 74131
rect 48436 72619 48876 74045
rect 48436 72533 48529 72619
rect 48615 72533 48697 72619
rect 48783 72533 48876 72619
rect 48436 71107 48876 72533
rect 48436 71021 48529 71107
rect 48615 71021 48697 71107
rect 48783 71021 48876 71107
rect 48436 69595 48876 71021
rect 48436 69509 48529 69595
rect 48615 69509 48697 69595
rect 48783 69509 48876 69595
rect 48436 68083 48876 69509
rect 48436 67997 48529 68083
rect 48615 67997 48697 68083
rect 48783 67997 48876 68083
rect 48436 66571 48876 67997
rect 48436 66485 48529 66571
rect 48615 66485 48697 66571
rect 48783 66485 48876 66571
rect 48436 65059 48876 66485
rect 48436 64973 48529 65059
rect 48615 64973 48697 65059
rect 48783 64973 48876 65059
rect 48436 63547 48876 64973
rect 48436 63461 48529 63547
rect 48615 63461 48697 63547
rect 48783 63461 48876 63547
rect 48436 62035 48876 63461
rect 48436 61949 48529 62035
rect 48615 61949 48697 62035
rect 48783 61949 48876 62035
rect 48436 60523 48876 61949
rect 48436 60437 48529 60523
rect 48615 60437 48697 60523
rect 48783 60437 48876 60523
rect 48436 59011 48876 60437
rect 48436 58925 48529 59011
rect 48615 58925 48697 59011
rect 48783 58925 48876 59011
rect 48436 57499 48876 58925
rect 48436 57413 48529 57499
rect 48615 57413 48697 57499
rect 48783 57413 48876 57499
rect 48436 55987 48876 57413
rect 48436 55901 48529 55987
rect 48615 55901 48697 55987
rect 48783 55901 48876 55987
rect 48436 54475 48876 55901
rect 48436 54389 48529 54475
rect 48615 54389 48697 54475
rect 48783 54389 48876 54475
rect 48436 52963 48876 54389
rect 48436 52877 48529 52963
rect 48615 52877 48697 52963
rect 48783 52877 48876 52963
rect 48436 51451 48876 52877
rect 48436 51365 48529 51451
rect 48615 51365 48697 51451
rect 48783 51365 48876 51451
rect 48436 49939 48876 51365
rect 48436 49853 48529 49939
rect 48615 49853 48697 49939
rect 48783 49853 48876 49939
rect 48436 48427 48876 49853
rect 48436 48341 48529 48427
rect 48615 48341 48697 48427
rect 48783 48341 48876 48427
rect 48436 46915 48876 48341
rect 48436 46829 48529 46915
rect 48615 46829 48697 46915
rect 48783 46829 48876 46915
rect 48436 45403 48876 46829
rect 48436 45317 48529 45403
rect 48615 45317 48697 45403
rect 48783 45317 48876 45403
rect 48436 43891 48876 45317
rect 48436 43805 48529 43891
rect 48615 43805 48697 43891
rect 48783 43805 48876 43891
rect 48436 42379 48876 43805
rect 48436 42293 48529 42379
rect 48615 42293 48697 42379
rect 48783 42293 48876 42379
rect 48436 40867 48876 42293
rect 48436 40781 48529 40867
rect 48615 40781 48697 40867
rect 48783 40781 48876 40867
rect 48436 39355 48876 40781
rect 48436 39269 48529 39355
rect 48615 39269 48697 39355
rect 48783 39269 48876 39355
rect 48436 37843 48876 39269
rect 48436 37757 48529 37843
rect 48615 37757 48697 37843
rect 48783 37757 48876 37843
rect 48436 36331 48876 37757
rect 48436 36245 48529 36331
rect 48615 36245 48697 36331
rect 48783 36245 48876 36331
rect 48436 34819 48876 36245
rect 48436 34733 48529 34819
rect 48615 34733 48697 34819
rect 48783 34733 48876 34819
rect 48436 33307 48876 34733
rect 48436 33221 48529 33307
rect 48615 33221 48697 33307
rect 48783 33221 48876 33307
rect 48436 31795 48876 33221
rect 48436 31709 48529 31795
rect 48615 31709 48697 31795
rect 48783 31709 48876 31795
rect 48436 30283 48876 31709
rect 48436 30197 48529 30283
rect 48615 30197 48697 30283
rect 48783 30197 48876 30283
rect 48436 28771 48876 30197
rect 48436 28685 48529 28771
rect 48615 28685 48697 28771
rect 48783 28685 48876 28771
rect 48436 27259 48876 28685
rect 48436 27173 48529 27259
rect 48615 27173 48697 27259
rect 48783 27173 48876 27259
rect 48436 25747 48876 27173
rect 48436 25661 48529 25747
rect 48615 25661 48697 25747
rect 48783 25661 48876 25747
rect 48436 24235 48876 25661
rect 48436 24149 48529 24235
rect 48615 24149 48697 24235
rect 48783 24149 48876 24235
rect 48436 22723 48876 24149
rect 48436 22637 48529 22723
rect 48615 22637 48697 22723
rect 48783 22637 48876 22723
rect 48436 21211 48876 22637
rect 48436 21125 48529 21211
rect 48615 21125 48697 21211
rect 48783 21125 48876 21211
rect 48436 19699 48876 21125
rect 48436 19613 48529 19699
rect 48615 19613 48697 19699
rect 48783 19613 48876 19699
rect 48436 18187 48876 19613
rect 48436 18101 48529 18187
rect 48615 18101 48697 18187
rect 48783 18101 48876 18187
rect 48436 16675 48876 18101
rect 48436 16589 48529 16675
rect 48615 16589 48697 16675
rect 48783 16589 48876 16675
rect 48436 15163 48876 16589
rect 48436 15077 48529 15163
rect 48615 15077 48697 15163
rect 48783 15077 48876 15163
rect 48436 13651 48876 15077
rect 48436 13565 48529 13651
rect 48615 13565 48697 13651
rect 48783 13565 48876 13651
rect 48436 12139 48876 13565
rect 48436 12053 48529 12139
rect 48615 12053 48697 12139
rect 48783 12053 48876 12139
rect 48436 10627 48876 12053
rect 48436 10541 48529 10627
rect 48615 10541 48697 10627
rect 48783 10541 48876 10627
rect 48436 9115 48876 10541
rect 48436 9029 48529 9115
rect 48615 9029 48697 9115
rect 48783 9029 48876 9115
rect 48436 7603 48876 9029
rect 48436 7517 48529 7603
rect 48615 7517 48697 7603
rect 48783 7517 48876 7603
rect 48436 6091 48876 7517
rect 48436 6005 48529 6091
rect 48615 6005 48697 6091
rect 48783 6005 48876 6091
rect 48436 4579 48876 6005
rect 48436 4493 48529 4579
rect 48615 4493 48697 4579
rect 48783 4493 48876 4579
rect 48436 3067 48876 4493
rect 48436 2981 48529 3067
rect 48615 2981 48697 3067
rect 48783 2981 48876 3067
rect 48436 1555 48876 2981
rect 48436 1469 48529 1555
rect 48615 1469 48697 1555
rect 48783 1469 48876 1555
rect 48436 712 48876 1469
rect 49676 80935 50116 81692
rect 49676 80849 49769 80935
rect 49855 80849 49937 80935
rect 50023 80849 50116 80935
rect 49676 79423 50116 80849
rect 49676 79337 49769 79423
rect 49855 79337 49937 79423
rect 50023 79337 50116 79423
rect 49676 77911 50116 79337
rect 49676 77825 49769 77911
rect 49855 77825 49937 77911
rect 50023 77825 50116 77911
rect 49676 76399 50116 77825
rect 49676 76313 49769 76399
rect 49855 76313 49937 76399
rect 50023 76313 50116 76399
rect 49676 74887 50116 76313
rect 49676 74801 49769 74887
rect 49855 74801 49937 74887
rect 50023 74801 50116 74887
rect 49676 73375 50116 74801
rect 49676 73289 49769 73375
rect 49855 73289 49937 73375
rect 50023 73289 50116 73375
rect 49676 71863 50116 73289
rect 49676 71777 49769 71863
rect 49855 71777 49937 71863
rect 50023 71777 50116 71863
rect 49676 70351 50116 71777
rect 49676 70265 49769 70351
rect 49855 70265 49937 70351
rect 50023 70265 50116 70351
rect 49676 68839 50116 70265
rect 49676 68753 49769 68839
rect 49855 68753 49937 68839
rect 50023 68753 50116 68839
rect 49676 67327 50116 68753
rect 49676 67241 49769 67327
rect 49855 67241 49937 67327
rect 50023 67241 50116 67327
rect 49676 65815 50116 67241
rect 49676 65729 49769 65815
rect 49855 65729 49937 65815
rect 50023 65729 50116 65815
rect 49676 64303 50116 65729
rect 49676 64217 49769 64303
rect 49855 64217 49937 64303
rect 50023 64217 50116 64303
rect 49676 62791 50116 64217
rect 49676 62705 49769 62791
rect 49855 62705 49937 62791
rect 50023 62705 50116 62791
rect 49676 61279 50116 62705
rect 49676 61193 49769 61279
rect 49855 61193 49937 61279
rect 50023 61193 50116 61279
rect 49676 59767 50116 61193
rect 49676 59681 49769 59767
rect 49855 59681 49937 59767
rect 50023 59681 50116 59767
rect 49676 58255 50116 59681
rect 49676 58169 49769 58255
rect 49855 58169 49937 58255
rect 50023 58169 50116 58255
rect 49676 56743 50116 58169
rect 49676 56657 49769 56743
rect 49855 56657 49937 56743
rect 50023 56657 50116 56743
rect 49676 55231 50116 56657
rect 49676 55145 49769 55231
rect 49855 55145 49937 55231
rect 50023 55145 50116 55231
rect 49676 53719 50116 55145
rect 49676 53633 49769 53719
rect 49855 53633 49937 53719
rect 50023 53633 50116 53719
rect 49676 52207 50116 53633
rect 49676 52121 49769 52207
rect 49855 52121 49937 52207
rect 50023 52121 50116 52207
rect 49676 50695 50116 52121
rect 49676 50609 49769 50695
rect 49855 50609 49937 50695
rect 50023 50609 50116 50695
rect 49676 49183 50116 50609
rect 49676 49097 49769 49183
rect 49855 49097 49937 49183
rect 50023 49097 50116 49183
rect 49676 47671 50116 49097
rect 49676 47585 49769 47671
rect 49855 47585 49937 47671
rect 50023 47585 50116 47671
rect 49676 46159 50116 47585
rect 49676 46073 49769 46159
rect 49855 46073 49937 46159
rect 50023 46073 50116 46159
rect 49676 44647 50116 46073
rect 49676 44561 49769 44647
rect 49855 44561 49937 44647
rect 50023 44561 50116 44647
rect 49676 43135 50116 44561
rect 49676 43049 49769 43135
rect 49855 43049 49937 43135
rect 50023 43049 50116 43135
rect 49676 41623 50116 43049
rect 49676 41537 49769 41623
rect 49855 41537 49937 41623
rect 50023 41537 50116 41623
rect 49676 40111 50116 41537
rect 49676 40025 49769 40111
rect 49855 40025 49937 40111
rect 50023 40025 50116 40111
rect 49676 38599 50116 40025
rect 49676 38513 49769 38599
rect 49855 38513 49937 38599
rect 50023 38513 50116 38599
rect 49676 37087 50116 38513
rect 49676 37001 49769 37087
rect 49855 37001 49937 37087
rect 50023 37001 50116 37087
rect 49676 35575 50116 37001
rect 49676 35489 49769 35575
rect 49855 35489 49937 35575
rect 50023 35489 50116 35575
rect 49676 34063 50116 35489
rect 49676 33977 49769 34063
rect 49855 33977 49937 34063
rect 50023 33977 50116 34063
rect 49676 32551 50116 33977
rect 49676 32465 49769 32551
rect 49855 32465 49937 32551
rect 50023 32465 50116 32551
rect 49676 31039 50116 32465
rect 49676 30953 49769 31039
rect 49855 30953 49937 31039
rect 50023 30953 50116 31039
rect 49676 29527 50116 30953
rect 49676 29441 49769 29527
rect 49855 29441 49937 29527
rect 50023 29441 50116 29527
rect 49676 28015 50116 29441
rect 49676 27929 49769 28015
rect 49855 27929 49937 28015
rect 50023 27929 50116 28015
rect 49676 26503 50116 27929
rect 49676 26417 49769 26503
rect 49855 26417 49937 26503
rect 50023 26417 50116 26503
rect 49676 24991 50116 26417
rect 49676 24905 49769 24991
rect 49855 24905 49937 24991
rect 50023 24905 50116 24991
rect 49676 23479 50116 24905
rect 49676 23393 49769 23479
rect 49855 23393 49937 23479
rect 50023 23393 50116 23479
rect 49676 21967 50116 23393
rect 49676 21881 49769 21967
rect 49855 21881 49937 21967
rect 50023 21881 50116 21967
rect 49676 20455 50116 21881
rect 49676 20369 49769 20455
rect 49855 20369 49937 20455
rect 50023 20369 50116 20455
rect 49676 18943 50116 20369
rect 49676 18857 49769 18943
rect 49855 18857 49937 18943
rect 50023 18857 50116 18943
rect 49676 17431 50116 18857
rect 49676 17345 49769 17431
rect 49855 17345 49937 17431
rect 50023 17345 50116 17431
rect 49676 15919 50116 17345
rect 49676 15833 49769 15919
rect 49855 15833 49937 15919
rect 50023 15833 50116 15919
rect 49676 14407 50116 15833
rect 49676 14321 49769 14407
rect 49855 14321 49937 14407
rect 50023 14321 50116 14407
rect 49676 12895 50116 14321
rect 49676 12809 49769 12895
rect 49855 12809 49937 12895
rect 50023 12809 50116 12895
rect 49676 11383 50116 12809
rect 49676 11297 49769 11383
rect 49855 11297 49937 11383
rect 50023 11297 50116 11383
rect 49676 9871 50116 11297
rect 49676 9785 49769 9871
rect 49855 9785 49937 9871
rect 50023 9785 50116 9871
rect 49676 8359 50116 9785
rect 49676 8273 49769 8359
rect 49855 8273 49937 8359
rect 50023 8273 50116 8359
rect 49676 6847 50116 8273
rect 49676 6761 49769 6847
rect 49855 6761 49937 6847
rect 50023 6761 50116 6847
rect 49676 5335 50116 6761
rect 49676 5249 49769 5335
rect 49855 5249 49937 5335
rect 50023 5249 50116 5335
rect 49676 3823 50116 5249
rect 49676 3737 49769 3823
rect 49855 3737 49937 3823
rect 50023 3737 50116 3823
rect 49676 2311 50116 3737
rect 49676 2225 49769 2311
rect 49855 2225 49937 2311
rect 50023 2225 50116 2311
rect 49676 799 50116 2225
rect 49676 713 49769 799
rect 49855 713 49937 799
rect 50023 713 50116 799
rect 49676 630 50116 713
rect 63556 81691 63996 81774
rect 63556 81605 63649 81691
rect 63735 81605 63817 81691
rect 63903 81605 63996 81691
rect 63556 80179 63996 81605
rect 63556 80093 63649 80179
rect 63735 80093 63817 80179
rect 63903 80093 63996 80179
rect 63556 78667 63996 80093
rect 63556 78581 63649 78667
rect 63735 78581 63817 78667
rect 63903 78581 63996 78667
rect 63556 77155 63996 78581
rect 63556 77069 63649 77155
rect 63735 77069 63817 77155
rect 63903 77069 63996 77155
rect 63556 75643 63996 77069
rect 63556 75557 63649 75643
rect 63735 75557 63817 75643
rect 63903 75557 63996 75643
rect 63556 74131 63996 75557
rect 63556 74045 63649 74131
rect 63735 74045 63817 74131
rect 63903 74045 63996 74131
rect 63556 72619 63996 74045
rect 63556 72533 63649 72619
rect 63735 72533 63817 72619
rect 63903 72533 63996 72619
rect 63556 71107 63996 72533
rect 63556 71021 63649 71107
rect 63735 71021 63817 71107
rect 63903 71021 63996 71107
rect 63556 69595 63996 71021
rect 63556 69509 63649 69595
rect 63735 69509 63817 69595
rect 63903 69509 63996 69595
rect 63556 68083 63996 69509
rect 63556 67997 63649 68083
rect 63735 67997 63817 68083
rect 63903 67997 63996 68083
rect 63556 66571 63996 67997
rect 63556 66485 63649 66571
rect 63735 66485 63817 66571
rect 63903 66485 63996 66571
rect 63556 65059 63996 66485
rect 63556 64973 63649 65059
rect 63735 64973 63817 65059
rect 63903 64973 63996 65059
rect 63556 63547 63996 64973
rect 63556 63461 63649 63547
rect 63735 63461 63817 63547
rect 63903 63461 63996 63547
rect 63556 62035 63996 63461
rect 63556 61949 63649 62035
rect 63735 61949 63817 62035
rect 63903 61949 63996 62035
rect 63556 60523 63996 61949
rect 63556 60437 63649 60523
rect 63735 60437 63817 60523
rect 63903 60437 63996 60523
rect 63556 59011 63996 60437
rect 63556 58925 63649 59011
rect 63735 58925 63817 59011
rect 63903 58925 63996 59011
rect 63556 57499 63996 58925
rect 63556 57413 63649 57499
rect 63735 57413 63817 57499
rect 63903 57413 63996 57499
rect 63556 55987 63996 57413
rect 63556 55901 63649 55987
rect 63735 55901 63817 55987
rect 63903 55901 63996 55987
rect 63556 54475 63996 55901
rect 63556 54389 63649 54475
rect 63735 54389 63817 54475
rect 63903 54389 63996 54475
rect 63556 52963 63996 54389
rect 63556 52877 63649 52963
rect 63735 52877 63817 52963
rect 63903 52877 63996 52963
rect 63556 51451 63996 52877
rect 63556 51365 63649 51451
rect 63735 51365 63817 51451
rect 63903 51365 63996 51451
rect 63556 49939 63996 51365
rect 63556 49853 63649 49939
rect 63735 49853 63817 49939
rect 63903 49853 63996 49939
rect 63556 48427 63996 49853
rect 63556 48341 63649 48427
rect 63735 48341 63817 48427
rect 63903 48341 63996 48427
rect 63556 46915 63996 48341
rect 63556 46829 63649 46915
rect 63735 46829 63817 46915
rect 63903 46829 63996 46915
rect 63556 45403 63996 46829
rect 63556 45317 63649 45403
rect 63735 45317 63817 45403
rect 63903 45317 63996 45403
rect 63556 43891 63996 45317
rect 63556 43805 63649 43891
rect 63735 43805 63817 43891
rect 63903 43805 63996 43891
rect 63556 42379 63996 43805
rect 63556 42293 63649 42379
rect 63735 42293 63817 42379
rect 63903 42293 63996 42379
rect 63556 40867 63996 42293
rect 63556 40781 63649 40867
rect 63735 40781 63817 40867
rect 63903 40781 63996 40867
rect 63556 39355 63996 40781
rect 63556 39269 63649 39355
rect 63735 39269 63817 39355
rect 63903 39269 63996 39355
rect 63556 37843 63996 39269
rect 63556 37757 63649 37843
rect 63735 37757 63817 37843
rect 63903 37757 63996 37843
rect 63556 36331 63996 37757
rect 63556 36245 63649 36331
rect 63735 36245 63817 36331
rect 63903 36245 63996 36331
rect 63556 34819 63996 36245
rect 63556 34733 63649 34819
rect 63735 34733 63817 34819
rect 63903 34733 63996 34819
rect 63556 33307 63996 34733
rect 63556 33221 63649 33307
rect 63735 33221 63817 33307
rect 63903 33221 63996 33307
rect 63556 31795 63996 33221
rect 63556 31709 63649 31795
rect 63735 31709 63817 31795
rect 63903 31709 63996 31795
rect 63556 30283 63996 31709
rect 63556 30197 63649 30283
rect 63735 30197 63817 30283
rect 63903 30197 63996 30283
rect 63556 28771 63996 30197
rect 63556 28685 63649 28771
rect 63735 28685 63817 28771
rect 63903 28685 63996 28771
rect 63556 27259 63996 28685
rect 63556 27173 63649 27259
rect 63735 27173 63817 27259
rect 63903 27173 63996 27259
rect 63556 25747 63996 27173
rect 63556 25661 63649 25747
rect 63735 25661 63817 25747
rect 63903 25661 63996 25747
rect 63556 24235 63996 25661
rect 63556 24149 63649 24235
rect 63735 24149 63817 24235
rect 63903 24149 63996 24235
rect 63556 22723 63996 24149
rect 63556 22637 63649 22723
rect 63735 22637 63817 22723
rect 63903 22637 63996 22723
rect 63556 21211 63996 22637
rect 63556 21125 63649 21211
rect 63735 21125 63817 21211
rect 63903 21125 63996 21211
rect 63556 19699 63996 21125
rect 63556 19613 63649 19699
rect 63735 19613 63817 19699
rect 63903 19613 63996 19699
rect 63556 18187 63996 19613
rect 63556 18101 63649 18187
rect 63735 18101 63817 18187
rect 63903 18101 63996 18187
rect 63556 16675 63996 18101
rect 63556 16589 63649 16675
rect 63735 16589 63817 16675
rect 63903 16589 63996 16675
rect 63556 15163 63996 16589
rect 63556 15077 63649 15163
rect 63735 15077 63817 15163
rect 63903 15077 63996 15163
rect 63556 13651 63996 15077
rect 63556 13565 63649 13651
rect 63735 13565 63817 13651
rect 63903 13565 63996 13651
rect 63556 12139 63996 13565
rect 63556 12053 63649 12139
rect 63735 12053 63817 12139
rect 63903 12053 63996 12139
rect 63556 10627 63996 12053
rect 63556 10541 63649 10627
rect 63735 10541 63817 10627
rect 63903 10541 63996 10627
rect 63556 9115 63996 10541
rect 63556 9029 63649 9115
rect 63735 9029 63817 9115
rect 63903 9029 63996 9115
rect 63556 7603 63996 9029
rect 63556 7517 63649 7603
rect 63735 7517 63817 7603
rect 63903 7517 63996 7603
rect 63556 6091 63996 7517
rect 63556 6005 63649 6091
rect 63735 6005 63817 6091
rect 63903 6005 63996 6091
rect 63556 4579 63996 6005
rect 63556 4493 63649 4579
rect 63735 4493 63817 4579
rect 63903 4493 63996 4579
rect 63556 3067 63996 4493
rect 63556 2981 63649 3067
rect 63735 2981 63817 3067
rect 63903 2981 63996 3067
rect 63556 1555 63996 2981
rect 63556 1469 63649 1555
rect 63735 1469 63817 1555
rect 63903 1469 63996 1555
rect 63556 712 63996 1469
rect 64796 80935 65236 81692
rect 64796 80849 64889 80935
rect 64975 80849 65057 80935
rect 65143 80849 65236 80935
rect 64796 79423 65236 80849
rect 64796 79337 64889 79423
rect 64975 79337 65057 79423
rect 65143 79337 65236 79423
rect 64796 77911 65236 79337
rect 64796 77825 64889 77911
rect 64975 77825 65057 77911
rect 65143 77825 65236 77911
rect 64796 76399 65236 77825
rect 64796 76313 64889 76399
rect 64975 76313 65057 76399
rect 65143 76313 65236 76399
rect 64796 74887 65236 76313
rect 64796 74801 64889 74887
rect 64975 74801 65057 74887
rect 65143 74801 65236 74887
rect 64796 73375 65236 74801
rect 64796 73289 64889 73375
rect 64975 73289 65057 73375
rect 65143 73289 65236 73375
rect 64796 71863 65236 73289
rect 64796 71777 64889 71863
rect 64975 71777 65057 71863
rect 65143 71777 65236 71863
rect 64796 70351 65236 71777
rect 64796 70265 64889 70351
rect 64975 70265 65057 70351
rect 65143 70265 65236 70351
rect 64796 68839 65236 70265
rect 64796 68753 64889 68839
rect 64975 68753 65057 68839
rect 65143 68753 65236 68839
rect 64796 67327 65236 68753
rect 64796 67241 64889 67327
rect 64975 67241 65057 67327
rect 65143 67241 65236 67327
rect 64796 65815 65236 67241
rect 64796 65729 64889 65815
rect 64975 65729 65057 65815
rect 65143 65729 65236 65815
rect 64796 64303 65236 65729
rect 64796 64217 64889 64303
rect 64975 64217 65057 64303
rect 65143 64217 65236 64303
rect 64796 62791 65236 64217
rect 64796 62705 64889 62791
rect 64975 62705 65057 62791
rect 65143 62705 65236 62791
rect 64796 61279 65236 62705
rect 64796 61193 64889 61279
rect 64975 61193 65057 61279
rect 65143 61193 65236 61279
rect 64796 59767 65236 61193
rect 64796 59681 64889 59767
rect 64975 59681 65057 59767
rect 65143 59681 65236 59767
rect 64796 58255 65236 59681
rect 64796 58169 64889 58255
rect 64975 58169 65057 58255
rect 65143 58169 65236 58255
rect 64796 56743 65236 58169
rect 64796 56657 64889 56743
rect 64975 56657 65057 56743
rect 65143 56657 65236 56743
rect 64796 55231 65236 56657
rect 64796 55145 64889 55231
rect 64975 55145 65057 55231
rect 65143 55145 65236 55231
rect 64796 53719 65236 55145
rect 64796 53633 64889 53719
rect 64975 53633 65057 53719
rect 65143 53633 65236 53719
rect 64796 52207 65236 53633
rect 64796 52121 64889 52207
rect 64975 52121 65057 52207
rect 65143 52121 65236 52207
rect 64796 50695 65236 52121
rect 64796 50609 64889 50695
rect 64975 50609 65057 50695
rect 65143 50609 65236 50695
rect 64796 49183 65236 50609
rect 64796 49097 64889 49183
rect 64975 49097 65057 49183
rect 65143 49097 65236 49183
rect 64796 47671 65236 49097
rect 64796 47585 64889 47671
rect 64975 47585 65057 47671
rect 65143 47585 65236 47671
rect 64796 46159 65236 47585
rect 64796 46073 64889 46159
rect 64975 46073 65057 46159
rect 65143 46073 65236 46159
rect 64796 44647 65236 46073
rect 64796 44561 64889 44647
rect 64975 44561 65057 44647
rect 65143 44561 65236 44647
rect 64796 43135 65236 44561
rect 64796 43049 64889 43135
rect 64975 43049 65057 43135
rect 65143 43049 65236 43135
rect 64796 41623 65236 43049
rect 64796 41537 64889 41623
rect 64975 41537 65057 41623
rect 65143 41537 65236 41623
rect 64796 40111 65236 41537
rect 64796 40025 64889 40111
rect 64975 40025 65057 40111
rect 65143 40025 65236 40111
rect 64796 38599 65236 40025
rect 64796 38513 64889 38599
rect 64975 38513 65057 38599
rect 65143 38513 65236 38599
rect 64796 37087 65236 38513
rect 64796 37001 64889 37087
rect 64975 37001 65057 37087
rect 65143 37001 65236 37087
rect 64796 35575 65236 37001
rect 64796 35489 64889 35575
rect 64975 35489 65057 35575
rect 65143 35489 65236 35575
rect 64796 34063 65236 35489
rect 64796 33977 64889 34063
rect 64975 33977 65057 34063
rect 65143 33977 65236 34063
rect 64796 32551 65236 33977
rect 64796 32465 64889 32551
rect 64975 32465 65057 32551
rect 65143 32465 65236 32551
rect 64796 31039 65236 32465
rect 64796 30953 64889 31039
rect 64975 30953 65057 31039
rect 65143 30953 65236 31039
rect 64796 29527 65236 30953
rect 64796 29441 64889 29527
rect 64975 29441 65057 29527
rect 65143 29441 65236 29527
rect 64796 28015 65236 29441
rect 64796 27929 64889 28015
rect 64975 27929 65057 28015
rect 65143 27929 65236 28015
rect 64796 26503 65236 27929
rect 64796 26417 64889 26503
rect 64975 26417 65057 26503
rect 65143 26417 65236 26503
rect 64796 24991 65236 26417
rect 64796 24905 64889 24991
rect 64975 24905 65057 24991
rect 65143 24905 65236 24991
rect 64796 23479 65236 24905
rect 64796 23393 64889 23479
rect 64975 23393 65057 23479
rect 65143 23393 65236 23479
rect 64796 21967 65236 23393
rect 64796 21881 64889 21967
rect 64975 21881 65057 21967
rect 65143 21881 65236 21967
rect 64796 20455 65236 21881
rect 64796 20369 64889 20455
rect 64975 20369 65057 20455
rect 65143 20369 65236 20455
rect 64796 18943 65236 20369
rect 64796 18857 64889 18943
rect 64975 18857 65057 18943
rect 65143 18857 65236 18943
rect 64796 17431 65236 18857
rect 64796 17345 64889 17431
rect 64975 17345 65057 17431
rect 65143 17345 65236 17431
rect 64796 15919 65236 17345
rect 64796 15833 64889 15919
rect 64975 15833 65057 15919
rect 65143 15833 65236 15919
rect 64796 14407 65236 15833
rect 64796 14321 64889 14407
rect 64975 14321 65057 14407
rect 65143 14321 65236 14407
rect 64796 12895 65236 14321
rect 64796 12809 64889 12895
rect 64975 12809 65057 12895
rect 65143 12809 65236 12895
rect 64796 11383 65236 12809
rect 64796 11297 64889 11383
rect 64975 11297 65057 11383
rect 65143 11297 65236 11383
rect 64796 9871 65236 11297
rect 64796 9785 64889 9871
rect 64975 9785 65057 9871
rect 65143 9785 65236 9871
rect 64796 8359 65236 9785
rect 64796 8273 64889 8359
rect 64975 8273 65057 8359
rect 65143 8273 65236 8359
rect 64796 6847 65236 8273
rect 64796 6761 64889 6847
rect 64975 6761 65057 6847
rect 65143 6761 65236 6847
rect 64796 5335 65236 6761
rect 64796 5249 64889 5335
rect 64975 5249 65057 5335
rect 65143 5249 65236 5335
rect 64796 3823 65236 5249
rect 64796 3737 64889 3823
rect 64975 3737 65057 3823
rect 65143 3737 65236 3823
rect 64796 2311 65236 3737
rect 64796 2225 64889 2311
rect 64975 2225 65057 2311
rect 65143 2225 65236 2311
rect 64796 799 65236 2225
rect 64796 713 64889 799
rect 64975 713 65057 799
rect 65143 713 65236 799
rect 64796 630 65236 713
rect 78676 81691 79116 81774
rect 78676 81605 78769 81691
rect 78855 81605 78937 81691
rect 79023 81605 79116 81691
rect 78676 80179 79116 81605
rect 78676 80093 78769 80179
rect 78855 80093 78937 80179
rect 79023 80093 79116 80179
rect 78676 78667 79116 80093
rect 78676 78581 78769 78667
rect 78855 78581 78937 78667
rect 79023 78581 79116 78667
rect 78676 77155 79116 78581
rect 78676 77069 78769 77155
rect 78855 77069 78937 77155
rect 79023 77069 79116 77155
rect 78676 75643 79116 77069
rect 78676 75557 78769 75643
rect 78855 75557 78937 75643
rect 79023 75557 79116 75643
rect 78676 74131 79116 75557
rect 78676 74045 78769 74131
rect 78855 74045 78937 74131
rect 79023 74045 79116 74131
rect 78676 72619 79116 74045
rect 78676 72533 78769 72619
rect 78855 72533 78937 72619
rect 79023 72533 79116 72619
rect 78676 71107 79116 72533
rect 78676 71021 78769 71107
rect 78855 71021 78937 71107
rect 79023 71021 79116 71107
rect 78676 69595 79116 71021
rect 78676 69509 78769 69595
rect 78855 69509 78937 69595
rect 79023 69509 79116 69595
rect 78676 68083 79116 69509
rect 78676 67997 78769 68083
rect 78855 67997 78937 68083
rect 79023 67997 79116 68083
rect 78676 66571 79116 67997
rect 78676 66485 78769 66571
rect 78855 66485 78937 66571
rect 79023 66485 79116 66571
rect 78676 65059 79116 66485
rect 78676 64973 78769 65059
rect 78855 64973 78937 65059
rect 79023 64973 79116 65059
rect 78676 63547 79116 64973
rect 78676 63461 78769 63547
rect 78855 63461 78937 63547
rect 79023 63461 79116 63547
rect 78676 62035 79116 63461
rect 78676 61949 78769 62035
rect 78855 61949 78937 62035
rect 79023 61949 79116 62035
rect 78676 60523 79116 61949
rect 78676 60437 78769 60523
rect 78855 60437 78937 60523
rect 79023 60437 79116 60523
rect 78676 59011 79116 60437
rect 78676 58925 78769 59011
rect 78855 58925 78937 59011
rect 79023 58925 79116 59011
rect 78676 57499 79116 58925
rect 78676 57413 78769 57499
rect 78855 57413 78937 57499
rect 79023 57413 79116 57499
rect 78676 55987 79116 57413
rect 78676 55901 78769 55987
rect 78855 55901 78937 55987
rect 79023 55901 79116 55987
rect 78676 54475 79116 55901
rect 78676 54389 78769 54475
rect 78855 54389 78937 54475
rect 79023 54389 79116 54475
rect 78676 52963 79116 54389
rect 78676 52877 78769 52963
rect 78855 52877 78937 52963
rect 79023 52877 79116 52963
rect 78676 51451 79116 52877
rect 78676 51365 78769 51451
rect 78855 51365 78937 51451
rect 79023 51365 79116 51451
rect 78676 49939 79116 51365
rect 78676 49853 78769 49939
rect 78855 49853 78937 49939
rect 79023 49853 79116 49939
rect 78676 48427 79116 49853
rect 78676 48341 78769 48427
rect 78855 48341 78937 48427
rect 79023 48341 79116 48427
rect 78676 46915 79116 48341
rect 78676 46829 78769 46915
rect 78855 46829 78937 46915
rect 79023 46829 79116 46915
rect 78676 45403 79116 46829
rect 78676 45317 78769 45403
rect 78855 45317 78937 45403
rect 79023 45317 79116 45403
rect 78676 43891 79116 45317
rect 78676 43805 78769 43891
rect 78855 43805 78937 43891
rect 79023 43805 79116 43891
rect 78676 42379 79116 43805
rect 78676 42293 78769 42379
rect 78855 42293 78937 42379
rect 79023 42293 79116 42379
rect 78676 40867 79116 42293
rect 78676 40781 78769 40867
rect 78855 40781 78937 40867
rect 79023 40781 79116 40867
rect 78676 39355 79116 40781
rect 78676 39269 78769 39355
rect 78855 39269 78937 39355
rect 79023 39269 79116 39355
rect 78676 37843 79116 39269
rect 78676 37757 78769 37843
rect 78855 37757 78937 37843
rect 79023 37757 79116 37843
rect 78676 36331 79116 37757
rect 78676 36245 78769 36331
rect 78855 36245 78937 36331
rect 79023 36245 79116 36331
rect 78676 34819 79116 36245
rect 78676 34733 78769 34819
rect 78855 34733 78937 34819
rect 79023 34733 79116 34819
rect 78676 33307 79116 34733
rect 78676 33221 78769 33307
rect 78855 33221 78937 33307
rect 79023 33221 79116 33307
rect 78676 31795 79116 33221
rect 78676 31709 78769 31795
rect 78855 31709 78937 31795
rect 79023 31709 79116 31795
rect 78676 30283 79116 31709
rect 78676 30197 78769 30283
rect 78855 30197 78937 30283
rect 79023 30197 79116 30283
rect 78676 28771 79116 30197
rect 78676 28685 78769 28771
rect 78855 28685 78937 28771
rect 79023 28685 79116 28771
rect 78676 27259 79116 28685
rect 78676 27173 78769 27259
rect 78855 27173 78937 27259
rect 79023 27173 79116 27259
rect 78676 25747 79116 27173
rect 78676 25661 78769 25747
rect 78855 25661 78937 25747
rect 79023 25661 79116 25747
rect 78676 24235 79116 25661
rect 78676 24149 78769 24235
rect 78855 24149 78937 24235
rect 79023 24149 79116 24235
rect 78676 22723 79116 24149
rect 78676 22637 78769 22723
rect 78855 22637 78937 22723
rect 79023 22637 79116 22723
rect 78676 21211 79116 22637
rect 78676 21125 78769 21211
rect 78855 21125 78937 21211
rect 79023 21125 79116 21211
rect 78676 19699 79116 21125
rect 78676 19613 78769 19699
rect 78855 19613 78937 19699
rect 79023 19613 79116 19699
rect 78676 18187 79116 19613
rect 78676 18101 78769 18187
rect 78855 18101 78937 18187
rect 79023 18101 79116 18187
rect 78676 16675 79116 18101
rect 78676 16589 78769 16675
rect 78855 16589 78937 16675
rect 79023 16589 79116 16675
rect 78676 15163 79116 16589
rect 78676 15077 78769 15163
rect 78855 15077 78937 15163
rect 79023 15077 79116 15163
rect 78676 13651 79116 15077
rect 78676 13565 78769 13651
rect 78855 13565 78937 13651
rect 79023 13565 79116 13651
rect 78676 12139 79116 13565
rect 78676 12053 78769 12139
rect 78855 12053 78937 12139
rect 79023 12053 79116 12139
rect 78676 10627 79116 12053
rect 78676 10541 78769 10627
rect 78855 10541 78937 10627
rect 79023 10541 79116 10627
rect 78676 9115 79116 10541
rect 78676 9029 78769 9115
rect 78855 9029 78937 9115
rect 79023 9029 79116 9115
rect 78676 7603 79116 9029
rect 78676 7517 78769 7603
rect 78855 7517 78937 7603
rect 79023 7517 79116 7603
rect 78676 6091 79116 7517
rect 78676 6005 78769 6091
rect 78855 6005 78937 6091
rect 79023 6005 79116 6091
rect 78676 4579 79116 6005
rect 78676 4493 78769 4579
rect 78855 4493 78937 4579
rect 79023 4493 79116 4579
rect 78676 3067 79116 4493
rect 78676 2981 78769 3067
rect 78855 2981 78937 3067
rect 79023 2981 79116 3067
rect 78676 1555 79116 2981
rect 78676 1469 78769 1555
rect 78855 1469 78937 1555
rect 79023 1469 79116 1555
rect 78676 712 79116 1469
rect 79916 80935 80356 81692
rect 79916 80849 80009 80935
rect 80095 80849 80177 80935
rect 80263 80849 80356 80935
rect 79916 79423 80356 80849
rect 79916 79337 80009 79423
rect 80095 79337 80177 79423
rect 80263 79337 80356 79423
rect 79916 77911 80356 79337
rect 79916 77825 80009 77911
rect 80095 77825 80177 77911
rect 80263 77825 80356 77911
rect 79916 76399 80356 77825
rect 79916 76313 80009 76399
rect 80095 76313 80177 76399
rect 80263 76313 80356 76399
rect 79916 74887 80356 76313
rect 79916 74801 80009 74887
rect 80095 74801 80177 74887
rect 80263 74801 80356 74887
rect 79916 73375 80356 74801
rect 79916 73289 80009 73375
rect 80095 73289 80177 73375
rect 80263 73289 80356 73375
rect 79916 71863 80356 73289
rect 79916 71777 80009 71863
rect 80095 71777 80177 71863
rect 80263 71777 80356 71863
rect 79916 70351 80356 71777
rect 79916 70265 80009 70351
rect 80095 70265 80177 70351
rect 80263 70265 80356 70351
rect 79916 68839 80356 70265
rect 79916 68753 80009 68839
rect 80095 68753 80177 68839
rect 80263 68753 80356 68839
rect 79916 67327 80356 68753
rect 79916 67241 80009 67327
rect 80095 67241 80177 67327
rect 80263 67241 80356 67327
rect 79916 65815 80356 67241
rect 79916 65729 80009 65815
rect 80095 65729 80177 65815
rect 80263 65729 80356 65815
rect 79916 64303 80356 65729
rect 79916 64217 80009 64303
rect 80095 64217 80177 64303
rect 80263 64217 80356 64303
rect 79916 62791 80356 64217
rect 79916 62705 80009 62791
rect 80095 62705 80177 62791
rect 80263 62705 80356 62791
rect 79916 61279 80356 62705
rect 79916 61193 80009 61279
rect 80095 61193 80177 61279
rect 80263 61193 80356 61279
rect 79916 59767 80356 61193
rect 79916 59681 80009 59767
rect 80095 59681 80177 59767
rect 80263 59681 80356 59767
rect 79916 58255 80356 59681
rect 79916 58169 80009 58255
rect 80095 58169 80177 58255
rect 80263 58169 80356 58255
rect 79916 56743 80356 58169
rect 79916 56657 80009 56743
rect 80095 56657 80177 56743
rect 80263 56657 80356 56743
rect 79916 55231 80356 56657
rect 79916 55145 80009 55231
rect 80095 55145 80177 55231
rect 80263 55145 80356 55231
rect 79916 53719 80356 55145
rect 79916 53633 80009 53719
rect 80095 53633 80177 53719
rect 80263 53633 80356 53719
rect 79916 52207 80356 53633
rect 79916 52121 80009 52207
rect 80095 52121 80177 52207
rect 80263 52121 80356 52207
rect 79916 50695 80356 52121
rect 79916 50609 80009 50695
rect 80095 50609 80177 50695
rect 80263 50609 80356 50695
rect 79916 49183 80356 50609
rect 79916 49097 80009 49183
rect 80095 49097 80177 49183
rect 80263 49097 80356 49183
rect 79916 47671 80356 49097
rect 79916 47585 80009 47671
rect 80095 47585 80177 47671
rect 80263 47585 80356 47671
rect 79916 46159 80356 47585
rect 79916 46073 80009 46159
rect 80095 46073 80177 46159
rect 80263 46073 80356 46159
rect 79916 44647 80356 46073
rect 79916 44561 80009 44647
rect 80095 44561 80177 44647
rect 80263 44561 80356 44647
rect 79916 43135 80356 44561
rect 79916 43049 80009 43135
rect 80095 43049 80177 43135
rect 80263 43049 80356 43135
rect 79916 41623 80356 43049
rect 79916 41537 80009 41623
rect 80095 41537 80177 41623
rect 80263 41537 80356 41623
rect 79916 40111 80356 41537
rect 79916 40025 80009 40111
rect 80095 40025 80177 40111
rect 80263 40025 80356 40111
rect 79916 38599 80356 40025
rect 79916 38513 80009 38599
rect 80095 38513 80177 38599
rect 80263 38513 80356 38599
rect 79916 37087 80356 38513
rect 79916 37001 80009 37087
rect 80095 37001 80177 37087
rect 80263 37001 80356 37087
rect 79916 35575 80356 37001
rect 79916 35489 80009 35575
rect 80095 35489 80177 35575
rect 80263 35489 80356 35575
rect 79916 34063 80356 35489
rect 79916 33977 80009 34063
rect 80095 33977 80177 34063
rect 80263 33977 80356 34063
rect 79916 32551 80356 33977
rect 79916 32465 80009 32551
rect 80095 32465 80177 32551
rect 80263 32465 80356 32551
rect 79916 31039 80356 32465
rect 79916 30953 80009 31039
rect 80095 30953 80177 31039
rect 80263 30953 80356 31039
rect 79916 29527 80356 30953
rect 79916 29441 80009 29527
rect 80095 29441 80177 29527
rect 80263 29441 80356 29527
rect 79916 28015 80356 29441
rect 79916 27929 80009 28015
rect 80095 27929 80177 28015
rect 80263 27929 80356 28015
rect 79916 26503 80356 27929
rect 79916 26417 80009 26503
rect 80095 26417 80177 26503
rect 80263 26417 80356 26503
rect 79916 24991 80356 26417
rect 79916 24905 80009 24991
rect 80095 24905 80177 24991
rect 80263 24905 80356 24991
rect 79916 23479 80356 24905
rect 79916 23393 80009 23479
rect 80095 23393 80177 23479
rect 80263 23393 80356 23479
rect 79916 21967 80356 23393
rect 79916 21881 80009 21967
rect 80095 21881 80177 21967
rect 80263 21881 80356 21967
rect 79916 20455 80356 21881
rect 79916 20369 80009 20455
rect 80095 20369 80177 20455
rect 80263 20369 80356 20455
rect 79916 18943 80356 20369
rect 79916 18857 80009 18943
rect 80095 18857 80177 18943
rect 80263 18857 80356 18943
rect 79916 17431 80356 18857
rect 79916 17345 80009 17431
rect 80095 17345 80177 17431
rect 80263 17345 80356 17431
rect 79916 15919 80356 17345
rect 79916 15833 80009 15919
rect 80095 15833 80177 15919
rect 80263 15833 80356 15919
rect 79916 14407 80356 15833
rect 79916 14321 80009 14407
rect 80095 14321 80177 14407
rect 80263 14321 80356 14407
rect 79916 12895 80356 14321
rect 79916 12809 80009 12895
rect 80095 12809 80177 12895
rect 80263 12809 80356 12895
rect 79916 11383 80356 12809
rect 79916 11297 80009 11383
rect 80095 11297 80177 11383
rect 80263 11297 80356 11383
rect 79916 9871 80356 11297
rect 79916 9785 80009 9871
rect 80095 9785 80177 9871
rect 80263 9785 80356 9871
rect 79916 8359 80356 9785
rect 79916 8273 80009 8359
rect 80095 8273 80177 8359
rect 80263 8273 80356 8359
rect 79916 6847 80356 8273
rect 79916 6761 80009 6847
rect 80095 6761 80177 6847
rect 80263 6761 80356 6847
rect 79916 5335 80356 6761
rect 79916 5249 80009 5335
rect 80095 5249 80177 5335
rect 80263 5249 80356 5335
rect 79916 3823 80356 5249
rect 79916 3737 80009 3823
rect 80095 3737 80177 3823
rect 80263 3737 80356 3823
rect 79916 2311 80356 3737
rect 79916 2225 80009 2311
rect 80095 2225 80177 2311
rect 80263 2225 80356 2311
rect 79916 799 80356 2225
rect 79916 713 80009 799
rect 80095 713 80177 799
rect 80263 713 80356 799
rect 79916 630 80356 713
rect 93796 81691 94236 81774
rect 93796 81605 93889 81691
rect 93975 81605 94057 81691
rect 94143 81605 94236 81691
rect 93796 80179 94236 81605
rect 93796 80093 93889 80179
rect 93975 80093 94057 80179
rect 94143 80093 94236 80179
rect 93796 78667 94236 80093
rect 93796 78581 93889 78667
rect 93975 78581 94057 78667
rect 94143 78581 94236 78667
rect 93796 77155 94236 78581
rect 93796 77069 93889 77155
rect 93975 77069 94057 77155
rect 94143 77069 94236 77155
rect 93796 75643 94236 77069
rect 93796 75557 93889 75643
rect 93975 75557 94057 75643
rect 94143 75557 94236 75643
rect 93796 74131 94236 75557
rect 93796 74045 93889 74131
rect 93975 74045 94057 74131
rect 94143 74045 94236 74131
rect 93796 72619 94236 74045
rect 93796 72533 93889 72619
rect 93975 72533 94057 72619
rect 94143 72533 94236 72619
rect 93796 71107 94236 72533
rect 93796 71021 93889 71107
rect 93975 71021 94057 71107
rect 94143 71021 94236 71107
rect 93796 69595 94236 71021
rect 93796 69509 93889 69595
rect 93975 69509 94057 69595
rect 94143 69509 94236 69595
rect 93796 68083 94236 69509
rect 93796 67997 93889 68083
rect 93975 67997 94057 68083
rect 94143 67997 94236 68083
rect 93796 66571 94236 67997
rect 93796 66485 93889 66571
rect 93975 66485 94057 66571
rect 94143 66485 94236 66571
rect 93796 65059 94236 66485
rect 93796 64973 93889 65059
rect 93975 64973 94057 65059
rect 94143 64973 94236 65059
rect 93796 63547 94236 64973
rect 93796 63461 93889 63547
rect 93975 63461 94057 63547
rect 94143 63461 94236 63547
rect 93796 62035 94236 63461
rect 93796 61949 93889 62035
rect 93975 61949 94057 62035
rect 94143 61949 94236 62035
rect 93796 60523 94236 61949
rect 93796 60437 93889 60523
rect 93975 60437 94057 60523
rect 94143 60437 94236 60523
rect 93796 59011 94236 60437
rect 93796 58925 93889 59011
rect 93975 58925 94057 59011
rect 94143 58925 94236 59011
rect 93796 57499 94236 58925
rect 93796 57413 93889 57499
rect 93975 57413 94057 57499
rect 94143 57413 94236 57499
rect 93796 55987 94236 57413
rect 93796 55901 93889 55987
rect 93975 55901 94057 55987
rect 94143 55901 94236 55987
rect 93796 54475 94236 55901
rect 93796 54389 93889 54475
rect 93975 54389 94057 54475
rect 94143 54389 94236 54475
rect 93796 52963 94236 54389
rect 93796 52877 93889 52963
rect 93975 52877 94057 52963
rect 94143 52877 94236 52963
rect 93796 51451 94236 52877
rect 93796 51365 93889 51451
rect 93975 51365 94057 51451
rect 94143 51365 94236 51451
rect 93796 49939 94236 51365
rect 93796 49853 93889 49939
rect 93975 49853 94057 49939
rect 94143 49853 94236 49939
rect 93796 48427 94236 49853
rect 93796 48341 93889 48427
rect 93975 48341 94057 48427
rect 94143 48341 94236 48427
rect 93796 46915 94236 48341
rect 93796 46829 93889 46915
rect 93975 46829 94057 46915
rect 94143 46829 94236 46915
rect 93796 45403 94236 46829
rect 93796 45317 93889 45403
rect 93975 45317 94057 45403
rect 94143 45317 94236 45403
rect 93796 43891 94236 45317
rect 93796 43805 93889 43891
rect 93975 43805 94057 43891
rect 94143 43805 94236 43891
rect 93796 42379 94236 43805
rect 93796 42293 93889 42379
rect 93975 42293 94057 42379
rect 94143 42293 94236 42379
rect 93796 40867 94236 42293
rect 93796 40781 93889 40867
rect 93975 40781 94057 40867
rect 94143 40781 94236 40867
rect 93796 39355 94236 40781
rect 93796 39269 93889 39355
rect 93975 39269 94057 39355
rect 94143 39269 94236 39355
rect 93796 37843 94236 39269
rect 93796 37757 93889 37843
rect 93975 37757 94057 37843
rect 94143 37757 94236 37843
rect 93796 36331 94236 37757
rect 93796 36245 93889 36331
rect 93975 36245 94057 36331
rect 94143 36245 94236 36331
rect 93796 34819 94236 36245
rect 93796 34733 93889 34819
rect 93975 34733 94057 34819
rect 94143 34733 94236 34819
rect 93796 33307 94236 34733
rect 93796 33221 93889 33307
rect 93975 33221 94057 33307
rect 94143 33221 94236 33307
rect 93796 31795 94236 33221
rect 93796 31709 93889 31795
rect 93975 31709 94057 31795
rect 94143 31709 94236 31795
rect 93796 30283 94236 31709
rect 93796 30197 93889 30283
rect 93975 30197 94057 30283
rect 94143 30197 94236 30283
rect 93796 28771 94236 30197
rect 93796 28685 93889 28771
rect 93975 28685 94057 28771
rect 94143 28685 94236 28771
rect 93796 27259 94236 28685
rect 93796 27173 93889 27259
rect 93975 27173 94057 27259
rect 94143 27173 94236 27259
rect 93796 25747 94236 27173
rect 93796 25661 93889 25747
rect 93975 25661 94057 25747
rect 94143 25661 94236 25747
rect 93796 24235 94236 25661
rect 93796 24149 93889 24235
rect 93975 24149 94057 24235
rect 94143 24149 94236 24235
rect 93796 22723 94236 24149
rect 93796 22637 93889 22723
rect 93975 22637 94057 22723
rect 94143 22637 94236 22723
rect 93796 21211 94236 22637
rect 93796 21125 93889 21211
rect 93975 21125 94057 21211
rect 94143 21125 94236 21211
rect 93796 19699 94236 21125
rect 93796 19613 93889 19699
rect 93975 19613 94057 19699
rect 94143 19613 94236 19699
rect 93796 18187 94236 19613
rect 93796 18101 93889 18187
rect 93975 18101 94057 18187
rect 94143 18101 94236 18187
rect 93796 16675 94236 18101
rect 93796 16589 93889 16675
rect 93975 16589 94057 16675
rect 94143 16589 94236 16675
rect 93796 15163 94236 16589
rect 93796 15077 93889 15163
rect 93975 15077 94057 15163
rect 94143 15077 94236 15163
rect 93796 13651 94236 15077
rect 93796 13565 93889 13651
rect 93975 13565 94057 13651
rect 94143 13565 94236 13651
rect 93796 12139 94236 13565
rect 93796 12053 93889 12139
rect 93975 12053 94057 12139
rect 94143 12053 94236 12139
rect 93796 10627 94236 12053
rect 93796 10541 93889 10627
rect 93975 10541 94057 10627
rect 94143 10541 94236 10627
rect 93796 9115 94236 10541
rect 93796 9029 93889 9115
rect 93975 9029 94057 9115
rect 94143 9029 94236 9115
rect 93796 7603 94236 9029
rect 93796 7517 93889 7603
rect 93975 7517 94057 7603
rect 94143 7517 94236 7603
rect 93796 6091 94236 7517
rect 93796 6005 93889 6091
rect 93975 6005 94057 6091
rect 94143 6005 94236 6091
rect 93796 4579 94236 6005
rect 93796 4493 93889 4579
rect 93975 4493 94057 4579
rect 94143 4493 94236 4579
rect 93796 3067 94236 4493
rect 93796 2981 93889 3067
rect 93975 2981 94057 3067
rect 94143 2981 94236 3067
rect 93796 1555 94236 2981
rect 93796 1469 93889 1555
rect 93975 1469 94057 1555
rect 94143 1469 94236 1555
rect 93796 712 94236 1469
rect 95036 80935 95476 81692
rect 95036 80849 95129 80935
rect 95215 80849 95297 80935
rect 95383 80849 95476 80935
rect 95036 79423 95476 80849
rect 95036 79337 95129 79423
rect 95215 79337 95297 79423
rect 95383 79337 95476 79423
rect 95036 77911 95476 79337
rect 95036 77825 95129 77911
rect 95215 77825 95297 77911
rect 95383 77825 95476 77911
rect 95036 76399 95476 77825
rect 95036 76313 95129 76399
rect 95215 76313 95297 76399
rect 95383 76313 95476 76399
rect 95036 74887 95476 76313
rect 95036 74801 95129 74887
rect 95215 74801 95297 74887
rect 95383 74801 95476 74887
rect 95036 73375 95476 74801
rect 95036 73289 95129 73375
rect 95215 73289 95297 73375
rect 95383 73289 95476 73375
rect 95036 71863 95476 73289
rect 95036 71777 95129 71863
rect 95215 71777 95297 71863
rect 95383 71777 95476 71863
rect 95036 70351 95476 71777
rect 95036 70265 95129 70351
rect 95215 70265 95297 70351
rect 95383 70265 95476 70351
rect 95036 68839 95476 70265
rect 95036 68753 95129 68839
rect 95215 68753 95297 68839
rect 95383 68753 95476 68839
rect 95036 67327 95476 68753
rect 95036 67241 95129 67327
rect 95215 67241 95297 67327
rect 95383 67241 95476 67327
rect 95036 65815 95476 67241
rect 95036 65729 95129 65815
rect 95215 65729 95297 65815
rect 95383 65729 95476 65815
rect 95036 64303 95476 65729
rect 95036 64217 95129 64303
rect 95215 64217 95297 64303
rect 95383 64217 95476 64303
rect 95036 62791 95476 64217
rect 95036 62705 95129 62791
rect 95215 62705 95297 62791
rect 95383 62705 95476 62791
rect 95036 61279 95476 62705
rect 95036 61193 95129 61279
rect 95215 61193 95297 61279
rect 95383 61193 95476 61279
rect 95036 59767 95476 61193
rect 95036 59681 95129 59767
rect 95215 59681 95297 59767
rect 95383 59681 95476 59767
rect 95036 58255 95476 59681
rect 95036 58169 95129 58255
rect 95215 58169 95297 58255
rect 95383 58169 95476 58255
rect 95036 56743 95476 58169
rect 95036 56657 95129 56743
rect 95215 56657 95297 56743
rect 95383 56657 95476 56743
rect 95036 55231 95476 56657
rect 95036 55145 95129 55231
rect 95215 55145 95297 55231
rect 95383 55145 95476 55231
rect 95036 53719 95476 55145
rect 95036 53633 95129 53719
rect 95215 53633 95297 53719
rect 95383 53633 95476 53719
rect 95036 52207 95476 53633
rect 95036 52121 95129 52207
rect 95215 52121 95297 52207
rect 95383 52121 95476 52207
rect 95036 50695 95476 52121
rect 95036 50609 95129 50695
rect 95215 50609 95297 50695
rect 95383 50609 95476 50695
rect 95036 49183 95476 50609
rect 95036 49097 95129 49183
rect 95215 49097 95297 49183
rect 95383 49097 95476 49183
rect 95036 47671 95476 49097
rect 95036 47585 95129 47671
rect 95215 47585 95297 47671
rect 95383 47585 95476 47671
rect 95036 46159 95476 47585
rect 95036 46073 95129 46159
rect 95215 46073 95297 46159
rect 95383 46073 95476 46159
rect 95036 44647 95476 46073
rect 95036 44561 95129 44647
rect 95215 44561 95297 44647
rect 95383 44561 95476 44647
rect 95036 43135 95476 44561
rect 95036 43049 95129 43135
rect 95215 43049 95297 43135
rect 95383 43049 95476 43135
rect 95036 41623 95476 43049
rect 95036 41537 95129 41623
rect 95215 41537 95297 41623
rect 95383 41537 95476 41623
rect 95036 40111 95476 41537
rect 95036 40025 95129 40111
rect 95215 40025 95297 40111
rect 95383 40025 95476 40111
rect 95036 38599 95476 40025
rect 95036 38513 95129 38599
rect 95215 38513 95297 38599
rect 95383 38513 95476 38599
rect 95036 37087 95476 38513
rect 95036 37001 95129 37087
rect 95215 37001 95297 37087
rect 95383 37001 95476 37087
rect 95036 35575 95476 37001
rect 95036 35489 95129 35575
rect 95215 35489 95297 35575
rect 95383 35489 95476 35575
rect 95036 34063 95476 35489
rect 95036 33977 95129 34063
rect 95215 33977 95297 34063
rect 95383 33977 95476 34063
rect 95036 32551 95476 33977
rect 95036 32465 95129 32551
rect 95215 32465 95297 32551
rect 95383 32465 95476 32551
rect 95036 31039 95476 32465
rect 95036 30953 95129 31039
rect 95215 30953 95297 31039
rect 95383 30953 95476 31039
rect 95036 29527 95476 30953
rect 95036 29441 95129 29527
rect 95215 29441 95297 29527
rect 95383 29441 95476 29527
rect 95036 28015 95476 29441
rect 95036 27929 95129 28015
rect 95215 27929 95297 28015
rect 95383 27929 95476 28015
rect 95036 26503 95476 27929
rect 95036 26417 95129 26503
rect 95215 26417 95297 26503
rect 95383 26417 95476 26503
rect 95036 24991 95476 26417
rect 95036 24905 95129 24991
rect 95215 24905 95297 24991
rect 95383 24905 95476 24991
rect 95036 23479 95476 24905
rect 95036 23393 95129 23479
rect 95215 23393 95297 23479
rect 95383 23393 95476 23479
rect 95036 21967 95476 23393
rect 95036 21881 95129 21967
rect 95215 21881 95297 21967
rect 95383 21881 95476 21967
rect 95036 20455 95476 21881
rect 95036 20369 95129 20455
rect 95215 20369 95297 20455
rect 95383 20369 95476 20455
rect 95036 18943 95476 20369
rect 95036 18857 95129 18943
rect 95215 18857 95297 18943
rect 95383 18857 95476 18943
rect 95036 17431 95476 18857
rect 95036 17345 95129 17431
rect 95215 17345 95297 17431
rect 95383 17345 95476 17431
rect 95036 15919 95476 17345
rect 95036 15833 95129 15919
rect 95215 15833 95297 15919
rect 95383 15833 95476 15919
rect 95036 14407 95476 15833
rect 95036 14321 95129 14407
rect 95215 14321 95297 14407
rect 95383 14321 95476 14407
rect 95036 12895 95476 14321
rect 95036 12809 95129 12895
rect 95215 12809 95297 12895
rect 95383 12809 95476 12895
rect 95036 11383 95476 12809
rect 95036 11297 95129 11383
rect 95215 11297 95297 11383
rect 95383 11297 95476 11383
rect 95036 9871 95476 11297
rect 95036 9785 95129 9871
rect 95215 9785 95297 9871
rect 95383 9785 95476 9871
rect 95036 8359 95476 9785
rect 95036 8273 95129 8359
rect 95215 8273 95297 8359
rect 95383 8273 95476 8359
rect 95036 6847 95476 8273
rect 95036 6761 95129 6847
rect 95215 6761 95297 6847
rect 95383 6761 95476 6847
rect 95036 5335 95476 6761
rect 95036 5249 95129 5335
rect 95215 5249 95297 5335
rect 95383 5249 95476 5335
rect 95036 3823 95476 5249
rect 95036 3737 95129 3823
rect 95215 3737 95297 3823
rect 95383 3737 95476 3823
rect 95036 2311 95476 3737
rect 95036 2225 95129 2311
rect 95215 2225 95297 2311
rect 95383 2225 95476 2311
rect 95036 799 95476 2225
rect 95036 713 95129 799
rect 95215 713 95297 799
rect 95383 713 95476 799
rect 95036 630 95476 713
use sg13g2_and2_1  _29_
timestamp 1676901763
transform 1 0 14016 0 -1 46116
box -48 -56 528 834
use sg13g2_and2_1  _30_
timestamp 1676901763
transform 1 0 13056 0 -1 47628
box -48 -56 528 834
use sg13g2_xor2_1  _31_
timestamp 1677577977
transform 1 0 13536 0 -1 47628
box -48 -56 816 834
use sg13g2_xor2_1  _32_
timestamp 1677577977
transform -1 0 15072 0 -1 47628
box -48 -56 816 834
use sg13g2_a21oi_2  _33_
timestamp 1685174172
transform -1 0 14400 0 1 46116
box -48 -56 816 834
use sg13g2_and2_1  _34_
timestamp 1676901763
transform -1 0 7968 0 -1 46116
box -48 -56 528 834
use sg13g2_xnor2_1  _35_
timestamp 1677516600
transform -1 0 8736 0 -1 46116
box -48 -56 816 834
use sg13g2_nor2_1  _36_
timestamp 1676627187
transform -1 0 7680 0 -1 47628
box -48 -56 432 834
use sg13g2_xor2_1  _37_
timestamp 1677577977
transform -1 0 9984 0 1 47628
box -48 -56 816 834
use sg13g2_or2_1  _38_
timestamp 1684236171
transform 1 0 2496 0 1 46116
box -48 -56 528 834
use sg13g2_and2_1  _39_
timestamp 1676901763
transform 1 0 1920 0 -1 47628
box -48 -56 528 834
use sg13g2_xor2_1  _40_
timestamp 1677577977
transform 1 0 2400 0 -1 47628
box -48 -56 816 834
use sg13g2_nor2_1  _41_
timestamp 1676627187
transform 1 0 6720 0 -1 47628
box -48 -56 432 834
use sg13g2_xnor2_1  _42_
timestamp 1677516600
transform -1 0 6240 0 -1 47628
box -48 -56 816 834
use sg13g2_nand2b_1  _43_
timestamp 1676567195
transform -1 0 6720 0 -1 47628
box -48 -56 528 834
use sg13g2_a21oi_1  _44_
timestamp 1683973020
transform -1 0 4128 0 -1 47628
box -48 -56 528 834
use sg13g2_o21ai_1  _45_
timestamp 1685175443
transform -1 0 6528 0 1 47628
box -48 -56 538 834
use sg13g2_nand2_1  _46_
timestamp 1676557249
transform 1 0 2016 0 -1 52164
box -48 -56 432 834
use sg13g2_xor2_1  _47_
timestamp 1677577977
transform 1 0 2400 0 -1 52164
box -48 -56 816 834
use sg13g2_inv_1  _48_
timestamp 1676382929
transform 1 0 5184 0 -1 52164
box -48 -56 336 834
use sg13g2_nand2_1  _49_
timestamp 1676557249
transform 1 0 3840 0 -1 52164
box -48 -56 432 834
use sg13g2_xnor2_1  _50_
timestamp 1677516600
transform -1 0 7296 0 -1 52164
box -48 -56 816 834
use sg13g2_nor2_1  _51_
timestamp 1676627187
transform -1 0 6720 0 -1 53676
box -48 -56 432 834
use sg13g2_xnor2_1  _52_
timestamp 1677516600
transform -1 0 7104 0 1 52164
box -48 -56 816 834
use sg13g2_nand2_1  _53_
timestamp 1676557249
transform -1 0 3552 0 -1 52164
box -48 -56 432 834
use sg13g2_xnor2_1  _54_
timestamp 1677516600
transform -1 0 3168 0 1 50652
box -48 -56 816 834
use sg13g2_nor2_1  _55_
timestamp 1676627187
transform -1 0 6528 0 -1 52164
box -48 -56 432 834
use sg13g2_nor2_1  _56_
timestamp 1676627187
transform 1 0 5472 0 -1 52164
box -48 -56 432 834
use sg13g2_a221oi_1  _57_
timestamp 1685197497
transform 1 0 5568 0 1 52164
box -48 -56 816 834
use sg13g2_nand2_1  _58_
timestamp 1676557249
transform 1 0 5760 0 1 56700
box -48 -56 432 834
use sg13g2_nor2_1  _59_
timestamp 1676627187
transform 1 0 6240 0 -1 58212
box -48 -56 432 834
use sg13g2_xor2_1  _60_
timestamp 1677577977
transform 1 0 6144 0 1 56700
box -48 -56 816 834
use sg13g2_xnor2_1  _61_
timestamp 1677516600
transform -1 0 7008 0 -1 56700
box -48 -56 816 834
use sg13g2_o21ai_1  _62_
timestamp 1685175443
transform 1 0 6912 0 1 56700
box -48 -56 538 834
use sg13g2_xnor2_1  _63_
timestamp 1677516600
transform 1 0 6240 0 -1 61236
box -48 -56 816 834
use sg13g2_xnor2_1  _64_
timestamp 1677516600
transform -1 0 7200 0 1 59724
box -48 -56 816 834
use sg13g2_xor2_1  _65_
timestamp 1677577977
transform -1 0 14688 0 1 44604
box -48 -56 816 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1679581782
transform 1 0 576 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1679581782
transform 1 0 1248 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1679581782
transform 1 0 1920 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_21
timestamp 1679581782
transform 1 0 2592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_28
timestamp 1679581782
transform 1 0 3264 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_35
timestamp 1679581782
transform 1 0 3936 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_42
timestamp 1679581782
transform 1 0 4608 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_49
timestamp 1679581782
transform 1 0 5280 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_56
timestamp 1679581782
transform 1 0 5952 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_63
timestamp 1679581782
transform 1 0 6624 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_70
timestamp 1679581782
transform 1 0 7296 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_77
timestamp 1679581782
transform 1 0 7968 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_84
timestamp 1679581782
transform 1 0 8640 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_91
timestamp 1679581782
transform 1 0 9312 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_98
timestamp 1679581782
transform 1 0 9984 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_105
timestamp 1679581782
transform 1 0 10656 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_112
timestamp 1679581782
transform 1 0 11328 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_119
timestamp 1679581782
transform 1 0 12000 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_126
timestamp 1679581782
transform 1 0 12672 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_133
timestamp 1679581782
transform 1 0 13344 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_140
timestamp 1679581782
transform 1 0 14016 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_147
timestamp 1679581782
transform 1 0 14688 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_154
timestamp 1679581782
transform 1 0 15360 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_161
timestamp 1679581782
transform 1 0 16032 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_168
timestamp 1679581782
transform 1 0 16704 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_175
timestamp 1679581782
transform 1 0 17376 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_182
timestamp 1679581782
transform 1 0 18048 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_189
timestamp 1679581782
transform 1 0 18720 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_196
timestamp 1679581782
transform 1 0 19392 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_203
timestamp 1679581782
transform 1 0 20064 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_210
timestamp 1679581782
transform 1 0 20736 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_217
timestamp 1679581782
transform 1 0 21408 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_224
timestamp 1679581782
transform 1 0 22080 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_231
timestamp 1679581782
transform 1 0 22752 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_238
timestamp 1679581782
transform 1 0 23424 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_245
timestamp 1679581782
transform 1 0 24096 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_252
timestamp 1679581782
transform 1 0 24768 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_259
timestamp 1679581782
transform 1 0 25440 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_266
timestamp 1679581782
transform 1 0 26112 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_273
timestamp 1679581782
transform 1 0 26784 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_280
timestamp 1679581782
transform 1 0 27456 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_287
timestamp 1679581782
transform 1 0 28128 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_294
timestamp 1679581782
transform 1 0 28800 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_301
timestamp 1679581782
transform 1 0 29472 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_308
timestamp 1679581782
transform 1 0 30144 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_315
timestamp 1679581782
transform 1 0 30816 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_322
timestamp 1679581782
transform 1 0 31488 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_329
timestamp 1679581782
transform 1 0 32160 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_336
timestamp 1679581782
transform 1 0 32832 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_343
timestamp 1679581782
transform 1 0 33504 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_350
timestamp 1679581782
transform 1 0 34176 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_357
timestamp 1679581782
transform 1 0 34848 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_364
timestamp 1679581782
transform 1 0 35520 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_371
timestamp 1679581782
transform 1 0 36192 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_378
timestamp 1679581782
transform 1 0 36864 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_385
timestamp 1679581782
transform 1 0 37536 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_392
timestamp 1679581782
transform 1 0 38208 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_399
timestamp 1679581782
transform 1 0 38880 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_406
timestamp 1679581782
transform 1 0 39552 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_413
timestamp 1679581782
transform 1 0 40224 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_420
timestamp 1679581782
transform 1 0 40896 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_427
timestamp 1679581782
transform 1 0 41568 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_434
timestamp 1679581782
transform 1 0 42240 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_441
timestamp 1679581782
transform 1 0 42912 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_448
timestamp 1679581782
transform 1 0 43584 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_455
timestamp 1679581782
transform 1 0 44256 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_462
timestamp 1679581782
transform 1 0 44928 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_469
timestamp 1679581782
transform 1 0 45600 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_476
timestamp 1679581782
transform 1 0 46272 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_483
timestamp 1679581782
transform 1 0 46944 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_490
timestamp 1679581782
transform 1 0 47616 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_497
timestamp 1679581782
transform 1 0 48288 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_504
timestamp 1679581782
transform 1 0 48960 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_511
timestamp 1679581782
transform 1 0 49632 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_518
timestamp 1679581782
transform 1 0 50304 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_525
timestamp 1679581782
transform 1 0 50976 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_532
timestamp 1679581782
transform 1 0 51648 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_539
timestamp 1679581782
transform 1 0 52320 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_546
timestamp 1679581782
transform 1 0 52992 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_553
timestamp 1679581782
transform 1 0 53664 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_560
timestamp 1679581782
transform 1 0 54336 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_567
timestamp 1679581782
transform 1 0 55008 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_574
timestamp 1679581782
transform 1 0 55680 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_581
timestamp 1679581782
transform 1 0 56352 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_588
timestamp 1679581782
transform 1 0 57024 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_595
timestamp 1679581782
transform 1 0 57696 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_602
timestamp 1679581782
transform 1 0 58368 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_609
timestamp 1679581782
transform 1 0 59040 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_616
timestamp 1679581782
transform 1 0 59712 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_623
timestamp 1679581782
transform 1 0 60384 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_630
timestamp 1679581782
transform 1 0 61056 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_637
timestamp 1679581782
transform 1 0 61728 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_644
timestamp 1679581782
transform 1 0 62400 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_651
timestamp 1679581782
transform 1 0 63072 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_658
timestamp 1679581782
transform 1 0 63744 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_665
timestamp 1679581782
transform 1 0 64416 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_672
timestamp 1679581782
transform 1 0 65088 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_679
timestamp 1679581782
transform 1 0 65760 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_686
timestamp 1679581782
transform 1 0 66432 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_693
timestamp 1679581782
transform 1 0 67104 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_700
timestamp 1679581782
transform 1 0 67776 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_707
timestamp 1679581782
transform 1 0 68448 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_714
timestamp 1679581782
transform 1 0 69120 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_721
timestamp 1679581782
transform 1 0 69792 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_728
timestamp 1679581782
transform 1 0 70464 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_735
timestamp 1679581782
transform 1 0 71136 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_742
timestamp 1679581782
transform 1 0 71808 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_749
timestamp 1679581782
transform 1 0 72480 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_756
timestamp 1679581782
transform 1 0 73152 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_763
timestamp 1679581782
transform 1 0 73824 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_770
timestamp 1679581782
transform 1 0 74496 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_777
timestamp 1679581782
transform 1 0 75168 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_784
timestamp 1679581782
transform 1 0 75840 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_791
timestamp 1679581782
transform 1 0 76512 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_798
timestamp 1679581782
transform 1 0 77184 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_805
timestamp 1679581782
transform 1 0 77856 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_812
timestamp 1679581782
transform 1 0 78528 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_819
timestamp 1679581782
transform 1 0 79200 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_826
timestamp 1679581782
transform 1 0 79872 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_833
timestamp 1679581782
transform 1 0 80544 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_840
timestamp 1679581782
transform 1 0 81216 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_847
timestamp 1679581782
transform 1 0 81888 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_854
timestamp 1679581782
transform 1 0 82560 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_861
timestamp 1679581782
transform 1 0 83232 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_868
timestamp 1679581782
transform 1 0 83904 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_875
timestamp 1679581782
transform 1 0 84576 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_882
timestamp 1679581782
transform 1 0 85248 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_889
timestamp 1679581782
transform 1 0 85920 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_896
timestamp 1679581782
transform 1 0 86592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_903
timestamp 1679581782
transform 1 0 87264 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_910
timestamp 1679581782
transform 1 0 87936 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_917
timestamp 1679581782
transform 1 0 88608 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_924
timestamp 1679581782
transform 1 0 89280 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_931
timestamp 1679581782
transform 1 0 89952 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_938
timestamp 1679581782
transform 1 0 90624 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_945
timestamp 1679581782
transform 1 0 91296 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_952
timestamp 1679581782
transform 1 0 91968 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_959
timestamp 1679581782
transform 1 0 92640 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_966
timestamp 1679581782
transform 1 0 93312 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_973
timestamp 1679581782
transform 1 0 93984 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_980
timestamp 1679581782
transform 1 0 94656 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_987
timestamp 1679581782
transform 1 0 95328 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_994
timestamp 1679581782
transform 1 0 96000 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_1001
timestamp 1679581782
transform 1 0 96672 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_1008
timestamp 1679581782
transform 1 0 97344 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_1015
timestamp 1679581782
transform 1 0 98016 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_1022
timestamp 1679581782
transform 1 0 98688 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679581782
transform 1 0 576 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_7
timestamp 1679581782
transform 1 0 1248 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_14
timestamp 1679581782
transform 1 0 1920 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_21
timestamp 1679581782
transform 1 0 2592 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_28
timestamp 1679581782
transform 1 0 3264 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_35
timestamp 1679581782
transform 1 0 3936 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_42
timestamp 1679581782
transform 1 0 4608 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_49
timestamp 1679581782
transform 1 0 5280 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_56
timestamp 1679581782
transform 1 0 5952 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_63
timestamp 1679581782
transform 1 0 6624 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_70
timestamp 1679581782
transform 1 0 7296 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_77
timestamp 1679581782
transform 1 0 7968 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_84
timestamp 1679581782
transform 1 0 8640 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_91
timestamp 1679581782
transform 1 0 9312 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_98
timestamp 1679581782
transform 1 0 9984 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_105
timestamp 1679581782
transform 1 0 10656 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_112
timestamp 1679581782
transform 1 0 11328 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_119
timestamp 1679581782
transform 1 0 12000 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_126
timestamp 1679581782
transform 1 0 12672 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_133
timestamp 1679581782
transform 1 0 13344 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_140
timestamp 1679581782
transform 1 0 14016 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_147
timestamp 1679581782
transform 1 0 14688 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_154
timestamp 1679581782
transform 1 0 15360 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_161
timestamp 1679581782
transform 1 0 16032 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_168
timestamp 1679581782
transform 1 0 16704 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_175
timestamp 1679581782
transform 1 0 17376 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_182
timestamp 1679581782
transform 1 0 18048 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_189
timestamp 1679581782
transform 1 0 18720 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_196
timestamp 1679581782
transform 1 0 19392 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_203
timestamp 1679581782
transform 1 0 20064 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_210
timestamp 1679581782
transform 1 0 20736 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_217
timestamp 1679581782
transform 1 0 21408 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_224
timestamp 1679581782
transform 1 0 22080 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_231
timestamp 1679581782
transform 1 0 22752 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_238
timestamp 1679581782
transform 1 0 23424 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_245
timestamp 1679581782
transform 1 0 24096 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_252
timestamp 1679581782
transform 1 0 24768 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_259
timestamp 1679581782
transform 1 0 25440 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_266
timestamp 1679581782
transform 1 0 26112 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_273
timestamp 1679581782
transform 1 0 26784 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_280
timestamp 1679581782
transform 1 0 27456 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_287
timestamp 1679581782
transform 1 0 28128 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_294
timestamp 1679581782
transform 1 0 28800 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_301
timestamp 1679581782
transform 1 0 29472 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_308
timestamp 1679581782
transform 1 0 30144 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_315
timestamp 1679581782
transform 1 0 30816 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_322
timestamp 1679581782
transform 1 0 31488 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_329
timestamp 1679581782
transform 1 0 32160 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_336
timestamp 1679581782
transform 1 0 32832 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_343
timestamp 1679581782
transform 1 0 33504 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_350
timestamp 1679581782
transform 1 0 34176 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_357
timestamp 1679581782
transform 1 0 34848 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_364
timestamp 1679581782
transform 1 0 35520 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_371
timestamp 1679581782
transform 1 0 36192 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_378
timestamp 1679581782
transform 1 0 36864 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_385
timestamp 1679581782
transform 1 0 37536 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_392
timestamp 1679581782
transform 1 0 38208 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_399
timestamp 1679581782
transform 1 0 38880 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_406
timestamp 1679581782
transform 1 0 39552 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_413
timestamp 1679581782
transform 1 0 40224 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_420
timestamp 1679581782
transform 1 0 40896 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_427
timestamp 1679581782
transform 1 0 41568 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_434
timestamp 1679581782
transform 1 0 42240 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_441
timestamp 1679581782
transform 1 0 42912 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_448
timestamp 1679581782
transform 1 0 43584 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_455
timestamp 1679581782
transform 1 0 44256 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_462
timestamp 1679581782
transform 1 0 44928 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_469
timestamp 1679581782
transform 1 0 45600 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_476
timestamp 1679581782
transform 1 0 46272 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_483
timestamp 1679581782
transform 1 0 46944 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_490
timestamp 1679581782
transform 1 0 47616 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_497
timestamp 1679581782
transform 1 0 48288 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_504
timestamp 1679581782
transform 1 0 48960 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_511
timestamp 1679581782
transform 1 0 49632 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_518
timestamp 1679581782
transform 1 0 50304 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_525
timestamp 1679581782
transform 1 0 50976 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_532
timestamp 1679581782
transform 1 0 51648 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_539
timestamp 1679581782
transform 1 0 52320 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_546
timestamp 1679581782
transform 1 0 52992 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_553
timestamp 1679581782
transform 1 0 53664 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_560
timestamp 1679581782
transform 1 0 54336 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_567
timestamp 1679581782
transform 1 0 55008 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_574
timestamp 1679581782
transform 1 0 55680 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_581
timestamp 1679581782
transform 1 0 56352 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_588
timestamp 1679581782
transform 1 0 57024 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_595
timestamp 1679581782
transform 1 0 57696 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_602
timestamp 1679581782
transform 1 0 58368 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_609
timestamp 1679581782
transform 1 0 59040 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_616
timestamp 1679581782
transform 1 0 59712 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_623
timestamp 1679581782
transform 1 0 60384 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_630
timestamp 1679581782
transform 1 0 61056 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_637
timestamp 1679581782
transform 1 0 61728 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_644
timestamp 1679581782
transform 1 0 62400 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_651
timestamp 1679581782
transform 1 0 63072 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_658
timestamp 1679581782
transform 1 0 63744 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_665
timestamp 1679581782
transform 1 0 64416 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_672
timestamp 1679581782
transform 1 0 65088 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_679
timestamp 1679581782
transform 1 0 65760 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_686
timestamp 1679581782
transform 1 0 66432 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_693
timestamp 1679581782
transform 1 0 67104 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_700
timestamp 1679581782
transform 1 0 67776 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_707
timestamp 1679581782
transform 1 0 68448 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_714
timestamp 1679581782
transform 1 0 69120 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_721
timestamp 1679581782
transform 1 0 69792 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_728
timestamp 1679581782
transform 1 0 70464 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_735
timestamp 1679581782
transform 1 0 71136 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_742
timestamp 1679581782
transform 1 0 71808 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_749
timestamp 1679581782
transform 1 0 72480 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_756
timestamp 1679581782
transform 1 0 73152 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_763
timestamp 1679581782
transform 1 0 73824 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_770
timestamp 1679581782
transform 1 0 74496 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_777
timestamp 1679581782
transform 1 0 75168 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_784
timestamp 1679581782
transform 1 0 75840 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_791
timestamp 1679581782
transform 1 0 76512 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_798
timestamp 1679581782
transform 1 0 77184 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_805
timestamp 1679581782
transform 1 0 77856 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_812
timestamp 1679581782
transform 1 0 78528 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_819
timestamp 1679581782
transform 1 0 79200 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_826
timestamp 1679581782
transform 1 0 79872 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_833
timestamp 1679581782
transform 1 0 80544 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_840
timestamp 1679581782
transform 1 0 81216 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_847
timestamp 1679581782
transform 1 0 81888 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_854
timestamp 1679581782
transform 1 0 82560 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_861
timestamp 1679581782
transform 1 0 83232 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_868
timestamp 1679581782
transform 1 0 83904 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_875
timestamp 1679581782
transform 1 0 84576 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_882
timestamp 1679581782
transform 1 0 85248 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_889
timestamp 1679581782
transform 1 0 85920 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_896
timestamp 1679581782
transform 1 0 86592 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_903
timestamp 1679581782
transform 1 0 87264 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_910
timestamp 1679581782
transform 1 0 87936 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_917
timestamp 1679581782
transform 1 0 88608 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_924
timestamp 1679581782
transform 1 0 89280 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_931
timestamp 1679581782
transform 1 0 89952 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_938
timestamp 1679581782
transform 1 0 90624 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_945
timestamp 1679581782
transform 1 0 91296 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_952
timestamp 1679581782
transform 1 0 91968 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_959
timestamp 1679581782
transform 1 0 92640 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_966
timestamp 1679581782
transform 1 0 93312 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_973
timestamp 1679581782
transform 1 0 93984 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_980
timestamp 1679581782
transform 1 0 94656 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_987
timestamp 1679581782
transform 1 0 95328 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_994
timestamp 1679581782
transform 1 0 96000 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_1001
timestamp 1679581782
transform 1 0 96672 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_1008
timestamp 1679581782
transform 1 0 97344 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_1015
timestamp 1679581782
transform 1 0 98016 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_1022
timestamp 1679581782
transform 1 0 98688 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_4
timestamp 1679581782
transform 1 0 960 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_11
timestamp 1679581782
transform 1 0 1632 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_18
timestamp 1679581782
transform 1 0 2304 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_25
timestamp 1679581782
transform 1 0 2976 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_32
timestamp 1679581782
transform 1 0 3648 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_39
timestamp 1679581782
transform 1 0 4320 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_46
timestamp 1679581782
transform 1 0 4992 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_53
timestamp 1679581782
transform 1 0 5664 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_60
timestamp 1679581782
transform 1 0 6336 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_67
timestamp 1679581782
transform 1 0 7008 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_74
timestamp 1679581782
transform 1 0 7680 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_81
timestamp 1679581782
transform 1 0 8352 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_88
timestamp 1679581782
transform 1 0 9024 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_95
timestamp 1679581782
transform 1 0 9696 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_102
timestamp 1679581782
transform 1 0 10368 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_109
timestamp 1679581782
transform 1 0 11040 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_116
timestamp 1679581782
transform 1 0 11712 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_123
timestamp 1679581782
transform 1 0 12384 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_130
timestamp 1679581782
transform 1 0 13056 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_137
timestamp 1679581782
transform 1 0 13728 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_144
timestamp 1679581782
transform 1 0 14400 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_151
timestamp 1679581782
transform 1 0 15072 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_158
timestamp 1679581782
transform 1 0 15744 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_165
timestamp 1679581782
transform 1 0 16416 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_172
timestamp 1679581782
transform 1 0 17088 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_179
timestamp 1679581782
transform 1 0 17760 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_186
timestamp 1679581782
transform 1 0 18432 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_193
timestamp 1679581782
transform 1 0 19104 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_200
timestamp 1679581782
transform 1 0 19776 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_207
timestamp 1679581782
transform 1 0 20448 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_214
timestamp 1679581782
transform 1 0 21120 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_221
timestamp 1679581782
transform 1 0 21792 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_228
timestamp 1679581782
transform 1 0 22464 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_235
timestamp 1679581782
transform 1 0 23136 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_242
timestamp 1679581782
transform 1 0 23808 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_249
timestamp 1679581782
transform 1 0 24480 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_256
timestamp 1679581782
transform 1 0 25152 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_263
timestamp 1679581782
transform 1 0 25824 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_270
timestamp 1679581782
transform 1 0 26496 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_277
timestamp 1679581782
transform 1 0 27168 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_284
timestamp 1679581782
transform 1 0 27840 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_291
timestamp 1679581782
transform 1 0 28512 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_298
timestamp 1679581782
transform 1 0 29184 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_305
timestamp 1679581782
transform 1 0 29856 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_312
timestamp 1679581782
transform 1 0 30528 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_319
timestamp 1679581782
transform 1 0 31200 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_326
timestamp 1679581782
transform 1 0 31872 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_333
timestamp 1679581782
transform 1 0 32544 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_340
timestamp 1679581782
transform 1 0 33216 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_347
timestamp 1679581782
transform 1 0 33888 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_354
timestamp 1679581782
transform 1 0 34560 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_361
timestamp 1679581782
transform 1 0 35232 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_368
timestamp 1679581782
transform 1 0 35904 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_375
timestamp 1679581782
transform 1 0 36576 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_382
timestamp 1679581782
transform 1 0 37248 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_389
timestamp 1679581782
transform 1 0 37920 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_396
timestamp 1679581782
transform 1 0 38592 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_403
timestamp 1679581782
transform 1 0 39264 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_410
timestamp 1679581782
transform 1 0 39936 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_417
timestamp 1679581782
transform 1 0 40608 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_424
timestamp 1679581782
transform 1 0 41280 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_431
timestamp 1679581782
transform 1 0 41952 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_438
timestamp 1679581782
transform 1 0 42624 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_445
timestamp 1679581782
transform 1 0 43296 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_452
timestamp 1679581782
transform 1 0 43968 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_459
timestamp 1679581782
transform 1 0 44640 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_466
timestamp 1679581782
transform 1 0 45312 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_473
timestamp 1679581782
transform 1 0 45984 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_480
timestamp 1679581782
transform 1 0 46656 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_487
timestamp 1679581782
transform 1 0 47328 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_494
timestamp 1679581782
transform 1 0 48000 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_501
timestamp 1679581782
transform 1 0 48672 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_508
timestamp 1679581782
transform 1 0 49344 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_515
timestamp 1679581782
transform 1 0 50016 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_522
timestamp 1679581782
transform 1 0 50688 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_529
timestamp 1679581782
transform 1 0 51360 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_536
timestamp 1679581782
transform 1 0 52032 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_543
timestamp 1679581782
transform 1 0 52704 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_550
timestamp 1679581782
transform 1 0 53376 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_557
timestamp 1679581782
transform 1 0 54048 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_564
timestamp 1679581782
transform 1 0 54720 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_571
timestamp 1679581782
transform 1 0 55392 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_578
timestamp 1679581782
transform 1 0 56064 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_585
timestamp 1679581782
transform 1 0 56736 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_592
timestamp 1679581782
transform 1 0 57408 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_599
timestamp 1679581782
transform 1 0 58080 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_606
timestamp 1679581782
transform 1 0 58752 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_613
timestamp 1679581782
transform 1 0 59424 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_620
timestamp 1679581782
transform 1 0 60096 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_627
timestamp 1679581782
transform 1 0 60768 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_634
timestamp 1679581782
transform 1 0 61440 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_641
timestamp 1679581782
transform 1 0 62112 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_648
timestamp 1679581782
transform 1 0 62784 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_655
timestamp 1679581782
transform 1 0 63456 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_662
timestamp 1679581782
transform 1 0 64128 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_669
timestamp 1679581782
transform 1 0 64800 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_676
timestamp 1679581782
transform 1 0 65472 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_683
timestamp 1679581782
transform 1 0 66144 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_690
timestamp 1679581782
transform 1 0 66816 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_697
timestamp 1679581782
transform 1 0 67488 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_704
timestamp 1679581782
transform 1 0 68160 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_711
timestamp 1679581782
transform 1 0 68832 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_718
timestamp 1679581782
transform 1 0 69504 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_725
timestamp 1679581782
transform 1 0 70176 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_732
timestamp 1679581782
transform 1 0 70848 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_739
timestamp 1679581782
transform 1 0 71520 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_746
timestamp 1679581782
transform 1 0 72192 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_753
timestamp 1679581782
transform 1 0 72864 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_760
timestamp 1679581782
transform 1 0 73536 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_767
timestamp 1679581782
transform 1 0 74208 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_774
timestamp 1679581782
transform 1 0 74880 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_781
timestamp 1679581782
transform 1 0 75552 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_788
timestamp 1679581782
transform 1 0 76224 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_795
timestamp 1679581782
transform 1 0 76896 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_802
timestamp 1679581782
transform 1 0 77568 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_809
timestamp 1679581782
transform 1 0 78240 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_816
timestamp 1679581782
transform 1 0 78912 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_823
timestamp 1679581782
transform 1 0 79584 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_830
timestamp 1679581782
transform 1 0 80256 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_837
timestamp 1679581782
transform 1 0 80928 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_844
timestamp 1679581782
transform 1 0 81600 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_851
timestamp 1679581782
transform 1 0 82272 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_858
timestamp 1679581782
transform 1 0 82944 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_865
timestamp 1679581782
transform 1 0 83616 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_872
timestamp 1679581782
transform 1 0 84288 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_879
timestamp 1679581782
transform 1 0 84960 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_886
timestamp 1679581782
transform 1 0 85632 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_893
timestamp 1679581782
transform 1 0 86304 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_900
timestamp 1679581782
transform 1 0 86976 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_907
timestamp 1679581782
transform 1 0 87648 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_914
timestamp 1679581782
transform 1 0 88320 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_921
timestamp 1679581782
transform 1 0 88992 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_928
timestamp 1679581782
transform 1 0 89664 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_935
timestamp 1679581782
transform 1 0 90336 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_942
timestamp 1679581782
transform 1 0 91008 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_949
timestamp 1679581782
transform 1 0 91680 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_956
timestamp 1679581782
transform 1 0 92352 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_963
timestamp 1679581782
transform 1 0 93024 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_970
timestamp 1679581782
transform 1 0 93696 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_977
timestamp 1679581782
transform 1 0 94368 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_984
timestamp 1679581782
transform 1 0 95040 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_991
timestamp 1679581782
transform 1 0 95712 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_998
timestamp 1679581782
transform 1 0 96384 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_1005
timestamp 1679581782
transform 1 0 97056 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_1012
timestamp 1679581782
transform 1 0 97728 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_1019
timestamp 1679581782
transform 1 0 98400 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_1026
timestamp 1677580104
transform 1 0 99072 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_1028
timestamp 1677579658
transform 1 0 99264 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_0
timestamp 1679581782
transform 1 0 576 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_7
timestamp 1679581782
transform 1 0 1248 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_14
timestamp 1679581782
transform 1 0 1920 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_21
timestamp 1679581782
transform 1 0 2592 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_28
timestamp 1679581782
transform 1 0 3264 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_35
timestamp 1679581782
transform 1 0 3936 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_42
timestamp 1679581782
transform 1 0 4608 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_49
timestamp 1679581782
transform 1 0 5280 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_56
timestamp 1679581782
transform 1 0 5952 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_63
timestamp 1679581782
transform 1 0 6624 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_70
timestamp 1679581782
transform 1 0 7296 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_77
timestamp 1679581782
transform 1 0 7968 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_84
timestamp 1679581782
transform 1 0 8640 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_91
timestamp 1679581782
transform 1 0 9312 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_98
timestamp 1679581782
transform 1 0 9984 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_105
timestamp 1679581782
transform 1 0 10656 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_112
timestamp 1679581782
transform 1 0 11328 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_119
timestamp 1679581782
transform 1 0 12000 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_126
timestamp 1679581782
transform 1 0 12672 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_133
timestamp 1679581782
transform 1 0 13344 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_140
timestamp 1679581782
transform 1 0 14016 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_147
timestamp 1679581782
transform 1 0 14688 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_154
timestamp 1679581782
transform 1 0 15360 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_161
timestamp 1679581782
transform 1 0 16032 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_168
timestamp 1679581782
transform 1 0 16704 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_175
timestamp 1679581782
transform 1 0 17376 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_182
timestamp 1679581782
transform 1 0 18048 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_189
timestamp 1679581782
transform 1 0 18720 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_196
timestamp 1679581782
transform 1 0 19392 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_203
timestamp 1679581782
transform 1 0 20064 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_210
timestamp 1679581782
transform 1 0 20736 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_217
timestamp 1679581782
transform 1 0 21408 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_224
timestamp 1679581782
transform 1 0 22080 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_231
timestamp 1679581782
transform 1 0 22752 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_238
timestamp 1679581782
transform 1 0 23424 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_245
timestamp 1679581782
transform 1 0 24096 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_252
timestamp 1679581782
transform 1 0 24768 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_259
timestamp 1679581782
transform 1 0 25440 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_266
timestamp 1679581782
transform 1 0 26112 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_273
timestamp 1679581782
transform 1 0 26784 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_280
timestamp 1679581782
transform 1 0 27456 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_287
timestamp 1679581782
transform 1 0 28128 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_294
timestamp 1679581782
transform 1 0 28800 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_301
timestamp 1679581782
transform 1 0 29472 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_308
timestamp 1679581782
transform 1 0 30144 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_315
timestamp 1679581782
transform 1 0 30816 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_322
timestamp 1679581782
transform 1 0 31488 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_329
timestamp 1679581782
transform 1 0 32160 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_336
timestamp 1679581782
transform 1 0 32832 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_343
timestamp 1679581782
transform 1 0 33504 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_350
timestamp 1679581782
transform 1 0 34176 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_357
timestamp 1679581782
transform 1 0 34848 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_364
timestamp 1679581782
transform 1 0 35520 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_371
timestamp 1679581782
transform 1 0 36192 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_378
timestamp 1679581782
transform 1 0 36864 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_385
timestamp 1679581782
transform 1 0 37536 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_392
timestamp 1679581782
transform 1 0 38208 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_399
timestamp 1679581782
transform 1 0 38880 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_406
timestamp 1679581782
transform 1 0 39552 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_413
timestamp 1679581782
transform 1 0 40224 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_420
timestamp 1679581782
transform 1 0 40896 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_427
timestamp 1679581782
transform 1 0 41568 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_434
timestamp 1679581782
transform 1 0 42240 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_441
timestamp 1679581782
transform 1 0 42912 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_448
timestamp 1679581782
transform 1 0 43584 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_455
timestamp 1679581782
transform 1 0 44256 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_462
timestamp 1679581782
transform 1 0 44928 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_469
timestamp 1679581782
transform 1 0 45600 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_476
timestamp 1679581782
transform 1 0 46272 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_483
timestamp 1679581782
transform 1 0 46944 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_490
timestamp 1679581782
transform 1 0 47616 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_497
timestamp 1679581782
transform 1 0 48288 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_504
timestamp 1679581782
transform 1 0 48960 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_511
timestamp 1679581782
transform 1 0 49632 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_518
timestamp 1679581782
transform 1 0 50304 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_525
timestamp 1679581782
transform 1 0 50976 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_532
timestamp 1679581782
transform 1 0 51648 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_539
timestamp 1679581782
transform 1 0 52320 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_546
timestamp 1679581782
transform 1 0 52992 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_553
timestamp 1679581782
transform 1 0 53664 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_560
timestamp 1679581782
transform 1 0 54336 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_567
timestamp 1679581782
transform 1 0 55008 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_574
timestamp 1679581782
transform 1 0 55680 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_581
timestamp 1679581782
transform 1 0 56352 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_588
timestamp 1679581782
transform 1 0 57024 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_595
timestamp 1679581782
transform 1 0 57696 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_602
timestamp 1679581782
transform 1 0 58368 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_609
timestamp 1679581782
transform 1 0 59040 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_616
timestamp 1679581782
transform 1 0 59712 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_623
timestamp 1679581782
transform 1 0 60384 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_630
timestamp 1679581782
transform 1 0 61056 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_637
timestamp 1679581782
transform 1 0 61728 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_644
timestamp 1679581782
transform 1 0 62400 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_651
timestamp 1679581782
transform 1 0 63072 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_658
timestamp 1679581782
transform 1 0 63744 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_665
timestamp 1679581782
transform 1 0 64416 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_672
timestamp 1679581782
transform 1 0 65088 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_679
timestamp 1679581782
transform 1 0 65760 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_686
timestamp 1679581782
transform 1 0 66432 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_693
timestamp 1679581782
transform 1 0 67104 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_700
timestamp 1679581782
transform 1 0 67776 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_707
timestamp 1679581782
transform 1 0 68448 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_714
timestamp 1679581782
transform 1 0 69120 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_721
timestamp 1679581782
transform 1 0 69792 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_728
timestamp 1679581782
transform 1 0 70464 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_735
timestamp 1679581782
transform 1 0 71136 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_742
timestamp 1679581782
transform 1 0 71808 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_749
timestamp 1679581782
transform 1 0 72480 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_756
timestamp 1679581782
transform 1 0 73152 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_763
timestamp 1679581782
transform 1 0 73824 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_770
timestamp 1679581782
transform 1 0 74496 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_777
timestamp 1679581782
transform 1 0 75168 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_784
timestamp 1679581782
transform 1 0 75840 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_791
timestamp 1679581782
transform 1 0 76512 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_798
timestamp 1679581782
transform 1 0 77184 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_805
timestamp 1679581782
transform 1 0 77856 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_812
timestamp 1679581782
transform 1 0 78528 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_819
timestamp 1679581782
transform 1 0 79200 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_826
timestamp 1679581782
transform 1 0 79872 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_833
timestamp 1679581782
transform 1 0 80544 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_840
timestamp 1679581782
transform 1 0 81216 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_847
timestamp 1679581782
transform 1 0 81888 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_854
timestamp 1679581782
transform 1 0 82560 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_861
timestamp 1679581782
transform 1 0 83232 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_868
timestamp 1679581782
transform 1 0 83904 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_875
timestamp 1679581782
transform 1 0 84576 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_882
timestamp 1679581782
transform 1 0 85248 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_889
timestamp 1679581782
transform 1 0 85920 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_896
timestamp 1679581782
transform 1 0 86592 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_903
timestamp 1679581782
transform 1 0 87264 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_910
timestamp 1679581782
transform 1 0 87936 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_917
timestamp 1679581782
transform 1 0 88608 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_924
timestamp 1679581782
transform 1 0 89280 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_931
timestamp 1679581782
transform 1 0 89952 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_938
timestamp 1679581782
transform 1 0 90624 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_945
timestamp 1679581782
transform 1 0 91296 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_952
timestamp 1679581782
transform 1 0 91968 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_959
timestamp 1679581782
transform 1 0 92640 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_966
timestamp 1679581782
transform 1 0 93312 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_973
timestamp 1679581782
transform 1 0 93984 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_980
timestamp 1679581782
transform 1 0 94656 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_987
timestamp 1679581782
transform 1 0 95328 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_994
timestamp 1679581782
transform 1 0 96000 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_1001
timestamp 1679581782
transform 1 0 96672 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_1008
timestamp 1679581782
transform 1 0 97344 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_1015
timestamp 1679581782
transform 1 0 98016 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_1022
timestamp 1679581782
transform 1 0 98688 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_0
timestamp 1679581782
transform 1 0 576 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_7
timestamp 1679581782
transform 1 0 1248 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_14
timestamp 1679581782
transform 1 0 1920 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_21
timestamp 1679581782
transform 1 0 2592 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_28
timestamp 1679581782
transform 1 0 3264 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_35
timestamp 1679581782
transform 1 0 3936 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_42
timestamp 1679581782
transform 1 0 4608 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_49
timestamp 1679581782
transform 1 0 5280 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_56
timestamp 1679581782
transform 1 0 5952 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_63
timestamp 1679581782
transform 1 0 6624 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_70
timestamp 1679581782
transform 1 0 7296 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_77
timestamp 1679581782
transform 1 0 7968 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_84
timestamp 1679581782
transform 1 0 8640 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_91
timestamp 1679581782
transform 1 0 9312 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_98
timestamp 1679581782
transform 1 0 9984 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_105
timestamp 1679581782
transform 1 0 10656 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_112
timestamp 1679581782
transform 1 0 11328 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_119
timestamp 1679581782
transform 1 0 12000 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_126
timestamp 1679581782
transform 1 0 12672 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_133
timestamp 1679581782
transform 1 0 13344 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_140
timestamp 1679581782
transform 1 0 14016 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_147
timestamp 1679581782
transform 1 0 14688 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_154
timestamp 1679581782
transform 1 0 15360 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_161
timestamp 1679581782
transform 1 0 16032 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_168
timestamp 1679581782
transform 1 0 16704 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_175
timestamp 1679581782
transform 1 0 17376 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_182
timestamp 1679581782
transform 1 0 18048 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_189
timestamp 1679581782
transform 1 0 18720 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_196
timestamp 1679581782
transform 1 0 19392 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_203
timestamp 1679581782
transform 1 0 20064 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_210
timestamp 1679581782
transform 1 0 20736 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_217
timestamp 1679581782
transform 1 0 21408 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_224
timestamp 1679581782
transform 1 0 22080 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_231
timestamp 1679581782
transform 1 0 22752 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_238
timestamp 1679581782
transform 1 0 23424 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_245
timestamp 1679581782
transform 1 0 24096 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_252
timestamp 1679581782
transform 1 0 24768 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_259
timestamp 1679581782
transform 1 0 25440 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_266
timestamp 1679581782
transform 1 0 26112 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_273
timestamp 1679581782
transform 1 0 26784 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_280
timestamp 1679581782
transform 1 0 27456 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_287
timestamp 1679581782
transform 1 0 28128 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_294
timestamp 1679581782
transform 1 0 28800 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_301
timestamp 1679581782
transform 1 0 29472 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_308
timestamp 1679581782
transform 1 0 30144 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_315
timestamp 1679581782
transform 1 0 30816 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_322
timestamp 1679581782
transform 1 0 31488 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_329
timestamp 1679581782
transform 1 0 32160 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_336
timestamp 1679581782
transform 1 0 32832 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_343
timestamp 1679581782
transform 1 0 33504 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_350
timestamp 1679581782
transform 1 0 34176 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_357
timestamp 1679581782
transform 1 0 34848 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_364
timestamp 1679581782
transform 1 0 35520 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_371
timestamp 1679581782
transform 1 0 36192 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_378
timestamp 1679581782
transform 1 0 36864 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_385
timestamp 1679581782
transform 1 0 37536 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_392
timestamp 1679581782
transform 1 0 38208 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_399
timestamp 1679581782
transform 1 0 38880 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_406
timestamp 1679581782
transform 1 0 39552 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_413
timestamp 1679581782
transform 1 0 40224 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_420
timestamp 1679581782
transform 1 0 40896 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_427
timestamp 1679581782
transform 1 0 41568 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_434
timestamp 1679581782
transform 1 0 42240 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_441
timestamp 1679581782
transform 1 0 42912 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_448
timestamp 1679581782
transform 1 0 43584 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_455
timestamp 1679581782
transform 1 0 44256 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_462
timestamp 1679581782
transform 1 0 44928 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_469
timestamp 1679581782
transform 1 0 45600 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_476
timestamp 1679581782
transform 1 0 46272 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_483
timestamp 1679581782
transform 1 0 46944 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_490
timestamp 1679581782
transform 1 0 47616 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_497
timestamp 1679581782
transform 1 0 48288 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_504
timestamp 1679581782
transform 1 0 48960 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_511
timestamp 1679581782
transform 1 0 49632 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_518
timestamp 1679581782
transform 1 0 50304 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_525
timestamp 1679581782
transform 1 0 50976 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_532
timestamp 1679581782
transform 1 0 51648 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_539
timestamp 1679581782
transform 1 0 52320 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_546
timestamp 1679581782
transform 1 0 52992 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_553
timestamp 1679581782
transform 1 0 53664 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_560
timestamp 1679581782
transform 1 0 54336 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_567
timestamp 1679581782
transform 1 0 55008 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_574
timestamp 1679581782
transform 1 0 55680 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_581
timestamp 1679581782
transform 1 0 56352 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_588
timestamp 1679581782
transform 1 0 57024 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_595
timestamp 1679581782
transform 1 0 57696 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_602
timestamp 1679581782
transform 1 0 58368 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_609
timestamp 1679581782
transform 1 0 59040 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_616
timestamp 1679581782
transform 1 0 59712 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_623
timestamp 1679581782
transform 1 0 60384 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_630
timestamp 1679581782
transform 1 0 61056 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_637
timestamp 1679581782
transform 1 0 61728 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_644
timestamp 1679581782
transform 1 0 62400 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_651
timestamp 1679581782
transform 1 0 63072 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_658
timestamp 1679581782
transform 1 0 63744 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_665
timestamp 1679581782
transform 1 0 64416 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_672
timestamp 1679581782
transform 1 0 65088 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_679
timestamp 1679581782
transform 1 0 65760 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_686
timestamp 1679581782
transform 1 0 66432 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_693
timestamp 1679581782
transform 1 0 67104 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_700
timestamp 1679581782
transform 1 0 67776 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_707
timestamp 1679581782
transform 1 0 68448 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_714
timestamp 1679581782
transform 1 0 69120 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_721
timestamp 1679581782
transform 1 0 69792 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_728
timestamp 1679581782
transform 1 0 70464 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_735
timestamp 1679581782
transform 1 0 71136 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_742
timestamp 1679581782
transform 1 0 71808 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_749
timestamp 1679581782
transform 1 0 72480 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_756
timestamp 1679581782
transform 1 0 73152 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_763
timestamp 1679581782
transform 1 0 73824 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_770
timestamp 1679581782
transform 1 0 74496 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_777
timestamp 1679581782
transform 1 0 75168 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_784
timestamp 1679581782
transform 1 0 75840 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_791
timestamp 1679581782
transform 1 0 76512 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_798
timestamp 1679581782
transform 1 0 77184 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_805
timestamp 1679581782
transform 1 0 77856 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_812
timestamp 1679581782
transform 1 0 78528 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_819
timestamp 1679581782
transform 1 0 79200 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_826
timestamp 1679581782
transform 1 0 79872 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_833
timestamp 1679581782
transform 1 0 80544 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_840
timestamp 1679581782
transform 1 0 81216 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_847
timestamp 1679581782
transform 1 0 81888 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_854
timestamp 1679581782
transform 1 0 82560 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_861
timestamp 1679581782
transform 1 0 83232 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_868
timestamp 1679581782
transform 1 0 83904 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_875
timestamp 1679581782
transform 1 0 84576 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_882
timestamp 1679581782
transform 1 0 85248 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_889
timestamp 1679581782
transform 1 0 85920 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_896
timestamp 1679581782
transform 1 0 86592 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_903
timestamp 1679581782
transform 1 0 87264 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_910
timestamp 1679581782
transform 1 0 87936 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_917
timestamp 1679581782
transform 1 0 88608 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_924
timestamp 1679581782
transform 1 0 89280 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_931
timestamp 1679581782
transform 1 0 89952 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_938
timestamp 1679581782
transform 1 0 90624 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_945
timestamp 1679581782
transform 1 0 91296 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_952
timestamp 1679581782
transform 1 0 91968 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_959
timestamp 1679581782
transform 1 0 92640 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_966
timestamp 1679581782
transform 1 0 93312 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_973
timestamp 1679581782
transform 1 0 93984 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_980
timestamp 1679581782
transform 1 0 94656 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_987
timestamp 1679581782
transform 1 0 95328 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_994
timestamp 1679581782
transform 1 0 96000 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_1001
timestamp 1679581782
transform 1 0 96672 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_1008
timestamp 1679581782
transform 1 0 97344 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_1015
timestamp 1679581782
transform 1 0 98016 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_1022
timestamp 1679581782
transform 1 0 98688 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_4
timestamp 1679581782
transform 1 0 960 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_11
timestamp 1679581782
transform 1 0 1632 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_18
timestamp 1679581782
transform 1 0 2304 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_25
timestamp 1679581782
transform 1 0 2976 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_32
timestamp 1679581782
transform 1 0 3648 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_39
timestamp 1679581782
transform 1 0 4320 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_46
timestamp 1679581782
transform 1 0 4992 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_53
timestamp 1679581782
transform 1 0 5664 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_60
timestamp 1679581782
transform 1 0 6336 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_67
timestamp 1679581782
transform 1 0 7008 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_74
timestamp 1679581782
transform 1 0 7680 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_81
timestamp 1679581782
transform 1 0 8352 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_88
timestamp 1679581782
transform 1 0 9024 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_95
timestamp 1679581782
transform 1 0 9696 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_102
timestamp 1679581782
transform 1 0 10368 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_109
timestamp 1679581782
transform 1 0 11040 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_116
timestamp 1679581782
transform 1 0 11712 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_123
timestamp 1679581782
transform 1 0 12384 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_130
timestamp 1679581782
transform 1 0 13056 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_137
timestamp 1679581782
transform 1 0 13728 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_144
timestamp 1679581782
transform 1 0 14400 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_151
timestamp 1679581782
transform 1 0 15072 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_158
timestamp 1679581782
transform 1 0 15744 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_165
timestamp 1679581782
transform 1 0 16416 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_172
timestamp 1679581782
transform 1 0 17088 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_179
timestamp 1679581782
transform 1 0 17760 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_186
timestamp 1679581782
transform 1 0 18432 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_193
timestamp 1679581782
transform 1 0 19104 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_200
timestamp 1679581782
transform 1 0 19776 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_207
timestamp 1679581782
transform 1 0 20448 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_214
timestamp 1679581782
transform 1 0 21120 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_221
timestamp 1679581782
transform 1 0 21792 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_228
timestamp 1679581782
transform 1 0 22464 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_235
timestamp 1679581782
transform 1 0 23136 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_242
timestamp 1679581782
transform 1 0 23808 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_249
timestamp 1679581782
transform 1 0 24480 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_256
timestamp 1679581782
transform 1 0 25152 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_263
timestamp 1679581782
transform 1 0 25824 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_270
timestamp 1679581782
transform 1 0 26496 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_277
timestamp 1679581782
transform 1 0 27168 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_284
timestamp 1679581782
transform 1 0 27840 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_291
timestamp 1679581782
transform 1 0 28512 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_298
timestamp 1679581782
transform 1 0 29184 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_305
timestamp 1679581782
transform 1 0 29856 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_312
timestamp 1679581782
transform 1 0 30528 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_319
timestamp 1679581782
transform 1 0 31200 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_326
timestamp 1679581782
transform 1 0 31872 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_333
timestamp 1679581782
transform 1 0 32544 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_340
timestamp 1679581782
transform 1 0 33216 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_347
timestamp 1679581782
transform 1 0 33888 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_354
timestamp 1679581782
transform 1 0 34560 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_361
timestamp 1679581782
transform 1 0 35232 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_368
timestamp 1679581782
transform 1 0 35904 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_375
timestamp 1679581782
transform 1 0 36576 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_382
timestamp 1679581782
transform 1 0 37248 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_389
timestamp 1679581782
transform 1 0 37920 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_396
timestamp 1679581782
transform 1 0 38592 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_403
timestamp 1679581782
transform 1 0 39264 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_410
timestamp 1679581782
transform 1 0 39936 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_417
timestamp 1679581782
transform 1 0 40608 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_424
timestamp 1679581782
transform 1 0 41280 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_431
timestamp 1679581782
transform 1 0 41952 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_438
timestamp 1679581782
transform 1 0 42624 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_445
timestamp 1679581782
transform 1 0 43296 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_452
timestamp 1679581782
transform 1 0 43968 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_459
timestamp 1679581782
transform 1 0 44640 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_466
timestamp 1679581782
transform 1 0 45312 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_473
timestamp 1679581782
transform 1 0 45984 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_480
timestamp 1679581782
transform 1 0 46656 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_487
timestamp 1679581782
transform 1 0 47328 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_494
timestamp 1679581782
transform 1 0 48000 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_501
timestamp 1679581782
transform 1 0 48672 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_508
timestamp 1679581782
transform 1 0 49344 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_515
timestamp 1679581782
transform 1 0 50016 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_522
timestamp 1679581782
transform 1 0 50688 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_529
timestamp 1679581782
transform 1 0 51360 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_536
timestamp 1679581782
transform 1 0 52032 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_543
timestamp 1679581782
transform 1 0 52704 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_550
timestamp 1679581782
transform 1 0 53376 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_557
timestamp 1679581782
transform 1 0 54048 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_564
timestamp 1679581782
transform 1 0 54720 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_571
timestamp 1679581782
transform 1 0 55392 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_578
timestamp 1679581782
transform 1 0 56064 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_585
timestamp 1679581782
transform 1 0 56736 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_592
timestamp 1679581782
transform 1 0 57408 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_599
timestamp 1679581782
transform 1 0 58080 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_606
timestamp 1679581782
transform 1 0 58752 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_613
timestamp 1679581782
transform 1 0 59424 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_620
timestamp 1679581782
transform 1 0 60096 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_627
timestamp 1679581782
transform 1 0 60768 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_634
timestamp 1679581782
transform 1 0 61440 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_641
timestamp 1679581782
transform 1 0 62112 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_648
timestamp 1679581782
transform 1 0 62784 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_655
timestamp 1679581782
transform 1 0 63456 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_662
timestamp 1679581782
transform 1 0 64128 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_669
timestamp 1679581782
transform 1 0 64800 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_676
timestamp 1679581782
transform 1 0 65472 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_683
timestamp 1679581782
transform 1 0 66144 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_690
timestamp 1679581782
transform 1 0 66816 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_697
timestamp 1679581782
transform 1 0 67488 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_704
timestamp 1679581782
transform 1 0 68160 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_711
timestamp 1679581782
transform 1 0 68832 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_718
timestamp 1679581782
transform 1 0 69504 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_725
timestamp 1679581782
transform 1 0 70176 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_732
timestamp 1679581782
transform 1 0 70848 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_739
timestamp 1679581782
transform 1 0 71520 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_746
timestamp 1679581782
transform 1 0 72192 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_753
timestamp 1679581782
transform 1 0 72864 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_760
timestamp 1679581782
transform 1 0 73536 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_767
timestamp 1679581782
transform 1 0 74208 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_774
timestamp 1679581782
transform 1 0 74880 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_781
timestamp 1679581782
transform 1 0 75552 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_788
timestamp 1679581782
transform 1 0 76224 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_795
timestamp 1679581782
transform 1 0 76896 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_802
timestamp 1679581782
transform 1 0 77568 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_809
timestamp 1679581782
transform 1 0 78240 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_816
timestamp 1679581782
transform 1 0 78912 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_823
timestamp 1679581782
transform 1 0 79584 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_830
timestamp 1679581782
transform 1 0 80256 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_837
timestamp 1679581782
transform 1 0 80928 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_844
timestamp 1679581782
transform 1 0 81600 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_851
timestamp 1679581782
transform 1 0 82272 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_858
timestamp 1679581782
transform 1 0 82944 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_865
timestamp 1679581782
transform 1 0 83616 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_872
timestamp 1679581782
transform 1 0 84288 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_879
timestamp 1679581782
transform 1 0 84960 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_886
timestamp 1679581782
transform 1 0 85632 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_893
timestamp 1679581782
transform 1 0 86304 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_900
timestamp 1679581782
transform 1 0 86976 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_907
timestamp 1679581782
transform 1 0 87648 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_914
timestamp 1679581782
transform 1 0 88320 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_921
timestamp 1679581782
transform 1 0 88992 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_928
timestamp 1679581782
transform 1 0 89664 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_935
timestamp 1679581782
transform 1 0 90336 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_942
timestamp 1679581782
transform 1 0 91008 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_949
timestamp 1679581782
transform 1 0 91680 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_956
timestamp 1679581782
transform 1 0 92352 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_963
timestamp 1679581782
transform 1 0 93024 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_970
timestamp 1679581782
transform 1 0 93696 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_977
timestamp 1679581782
transform 1 0 94368 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_984
timestamp 1679581782
transform 1 0 95040 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_991
timestamp 1679581782
transform 1 0 95712 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_998
timestamp 1679581782
transform 1 0 96384 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_1005
timestamp 1679581782
transform 1 0 97056 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_1012
timestamp 1679581782
transform 1 0 97728 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_1019
timestamp 1679581782
transform 1 0 98400 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_1026
timestamp 1677580104
transform 1 0 99072 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_1028
timestamp 1677579658
transform 1 0 99264 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_0
timestamp 1679581782
transform 1 0 576 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_7
timestamp 1679581782
transform 1 0 1248 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_14
timestamp 1679581782
transform 1 0 1920 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_21
timestamp 1679581782
transform 1 0 2592 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_28
timestamp 1679581782
transform 1 0 3264 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_35
timestamp 1679581782
transform 1 0 3936 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_42
timestamp 1679581782
transform 1 0 4608 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_49
timestamp 1679581782
transform 1 0 5280 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_56
timestamp 1679581782
transform 1 0 5952 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_63
timestamp 1679581782
transform 1 0 6624 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_70
timestamp 1679581782
transform 1 0 7296 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_77
timestamp 1679581782
transform 1 0 7968 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_84
timestamp 1679581782
transform 1 0 8640 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_91
timestamp 1679581782
transform 1 0 9312 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_98
timestamp 1679581782
transform 1 0 9984 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_105
timestamp 1679581782
transform 1 0 10656 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_112
timestamp 1679581782
transform 1 0 11328 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_119
timestamp 1679581782
transform 1 0 12000 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_126
timestamp 1679581782
transform 1 0 12672 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_133
timestamp 1679581782
transform 1 0 13344 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_140
timestamp 1679581782
transform 1 0 14016 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_147
timestamp 1679581782
transform 1 0 14688 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_154
timestamp 1679581782
transform 1 0 15360 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_161
timestamp 1679581782
transform 1 0 16032 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_168
timestamp 1679581782
transform 1 0 16704 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_175
timestamp 1679581782
transform 1 0 17376 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_182
timestamp 1679581782
transform 1 0 18048 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_189
timestamp 1679581782
transform 1 0 18720 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_196
timestamp 1679581782
transform 1 0 19392 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_203
timestamp 1679581782
transform 1 0 20064 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_210
timestamp 1679581782
transform 1 0 20736 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_217
timestamp 1679581782
transform 1 0 21408 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_224
timestamp 1679581782
transform 1 0 22080 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_231
timestamp 1679581782
transform 1 0 22752 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_238
timestamp 1679581782
transform 1 0 23424 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_245
timestamp 1679581782
transform 1 0 24096 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_252
timestamp 1679581782
transform 1 0 24768 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_259
timestamp 1679581782
transform 1 0 25440 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_266
timestamp 1679581782
transform 1 0 26112 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_273
timestamp 1679581782
transform 1 0 26784 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_280
timestamp 1679581782
transform 1 0 27456 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_287
timestamp 1679581782
transform 1 0 28128 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_294
timestamp 1679581782
transform 1 0 28800 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_301
timestamp 1679581782
transform 1 0 29472 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_308
timestamp 1679581782
transform 1 0 30144 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_315
timestamp 1679581782
transform 1 0 30816 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_322
timestamp 1679581782
transform 1 0 31488 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_329
timestamp 1679581782
transform 1 0 32160 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_336
timestamp 1679581782
transform 1 0 32832 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_343
timestamp 1679581782
transform 1 0 33504 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_350
timestamp 1679581782
transform 1 0 34176 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_357
timestamp 1679581782
transform 1 0 34848 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_364
timestamp 1679581782
transform 1 0 35520 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_371
timestamp 1679581782
transform 1 0 36192 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_378
timestamp 1679581782
transform 1 0 36864 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_385
timestamp 1679581782
transform 1 0 37536 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_392
timestamp 1679581782
transform 1 0 38208 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_399
timestamp 1679581782
transform 1 0 38880 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_406
timestamp 1679581782
transform 1 0 39552 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_413
timestamp 1679581782
transform 1 0 40224 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_420
timestamp 1679581782
transform 1 0 40896 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_427
timestamp 1679581782
transform 1 0 41568 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_434
timestamp 1679581782
transform 1 0 42240 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_441
timestamp 1679581782
transform 1 0 42912 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_448
timestamp 1679581782
transform 1 0 43584 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_455
timestamp 1679581782
transform 1 0 44256 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_462
timestamp 1679581782
transform 1 0 44928 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_469
timestamp 1679581782
transform 1 0 45600 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_476
timestamp 1679581782
transform 1 0 46272 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_483
timestamp 1679581782
transform 1 0 46944 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_490
timestamp 1679581782
transform 1 0 47616 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_497
timestamp 1679581782
transform 1 0 48288 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_504
timestamp 1679581782
transform 1 0 48960 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_511
timestamp 1679581782
transform 1 0 49632 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_518
timestamp 1679581782
transform 1 0 50304 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_525
timestamp 1679581782
transform 1 0 50976 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_532
timestamp 1679581782
transform 1 0 51648 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_539
timestamp 1679581782
transform 1 0 52320 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_546
timestamp 1679581782
transform 1 0 52992 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_553
timestamp 1679581782
transform 1 0 53664 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_560
timestamp 1679581782
transform 1 0 54336 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_567
timestamp 1679581782
transform 1 0 55008 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_574
timestamp 1679581782
transform 1 0 55680 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_581
timestamp 1679581782
transform 1 0 56352 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_588
timestamp 1679581782
transform 1 0 57024 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_595
timestamp 1679581782
transform 1 0 57696 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_602
timestamp 1679581782
transform 1 0 58368 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_609
timestamp 1679581782
transform 1 0 59040 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_616
timestamp 1679581782
transform 1 0 59712 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_623
timestamp 1679581782
transform 1 0 60384 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_630
timestamp 1679581782
transform 1 0 61056 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_637
timestamp 1679581782
transform 1 0 61728 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_644
timestamp 1679581782
transform 1 0 62400 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_651
timestamp 1679581782
transform 1 0 63072 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_658
timestamp 1679581782
transform 1 0 63744 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_665
timestamp 1679581782
transform 1 0 64416 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_672
timestamp 1679581782
transform 1 0 65088 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_679
timestamp 1679581782
transform 1 0 65760 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_686
timestamp 1679581782
transform 1 0 66432 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_693
timestamp 1679581782
transform 1 0 67104 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_700
timestamp 1679581782
transform 1 0 67776 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_707
timestamp 1679581782
transform 1 0 68448 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_714
timestamp 1679581782
transform 1 0 69120 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_721
timestamp 1679581782
transform 1 0 69792 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_728
timestamp 1679581782
transform 1 0 70464 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_735
timestamp 1679581782
transform 1 0 71136 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_742
timestamp 1679581782
transform 1 0 71808 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_749
timestamp 1679581782
transform 1 0 72480 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_756
timestamp 1679581782
transform 1 0 73152 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_763
timestamp 1679581782
transform 1 0 73824 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_770
timestamp 1679581782
transform 1 0 74496 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_777
timestamp 1679581782
transform 1 0 75168 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_784
timestamp 1679581782
transform 1 0 75840 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_791
timestamp 1679581782
transform 1 0 76512 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_798
timestamp 1679581782
transform 1 0 77184 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_805
timestamp 1679581782
transform 1 0 77856 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_812
timestamp 1679581782
transform 1 0 78528 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_819
timestamp 1679581782
transform 1 0 79200 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_826
timestamp 1679581782
transform 1 0 79872 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_833
timestamp 1679581782
transform 1 0 80544 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_840
timestamp 1679581782
transform 1 0 81216 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_847
timestamp 1679581782
transform 1 0 81888 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_854
timestamp 1679581782
transform 1 0 82560 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_861
timestamp 1679581782
transform 1 0 83232 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_868
timestamp 1679581782
transform 1 0 83904 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_875
timestamp 1679581782
transform 1 0 84576 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_882
timestamp 1679581782
transform 1 0 85248 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_889
timestamp 1679581782
transform 1 0 85920 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_896
timestamp 1679581782
transform 1 0 86592 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_903
timestamp 1679581782
transform 1 0 87264 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_910
timestamp 1679581782
transform 1 0 87936 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_917
timestamp 1679581782
transform 1 0 88608 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_924
timestamp 1679581782
transform 1 0 89280 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_931
timestamp 1679581782
transform 1 0 89952 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_938
timestamp 1679581782
transform 1 0 90624 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_945
timestamp 1679581782
transform 1 0 91296 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_952
timestamp 1679581782
transform 1 0 91968 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_959
timestamp 1679581782
transform 1 0 92640 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_966
timestamp 1679581782
transform 1 0 93312 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_973
timestamp 1679581782
transform 1 0 93984 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_980
timestamp 1679581782
transform 1 0 94656 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_987
timestamp 1679581782
transform 1 0 95328 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_994
timestamp 1679581782
transform 1 0 96000 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_1001
timestamp 1679581782
transform 1 0 96672 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_1008
timestamp 1679581782
transform 1 0 97344 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_1015
timestamp 1679581782
transform 1 0 98016 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_1022
timestamp 1679581782
transform 1 0 98688 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_4
timestamp 1679581782
transform 1 0 960 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_11
timestamp 1679581782
transform 1 0 1632 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_18
timestamp 1679581782
transform 1 0 2304 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_25
timestamp 1679581782
transform 1 0 2976 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_32
timestamp 1679581782
transform 1 0 3648 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_39
timestamp 1679581782
transform 1 0 4320 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_46
timestamp 1679581782
transform 1 0 4992 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_53
timestamp 1679581782
transform 1 0 5664 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_60
timestamp 1679581782
transform 1 0 6336 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_67
timestamp 1679581782
transform 1 0 7008 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_74
timestamp 1679581782
transform 1 0 7680 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_81
timestamp 1679581782
transform 1 0 8352 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_88
timestamp 1679581782
transform 1 0 9024 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_95
timestamp 1679581782
transform 1 0 9696 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_102
timestamp 1679581782
transform 1 0 10368 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_109
timestamp 1679581782
transform 1 0 11040 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_116
timestamp 1679581782
transform 1 0 11712 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_123
timestamp 1679581782
transform 1 0 12384 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_130
timestamp 1679581782
transform 1 0 13056 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_137
timestamp 1679581782
transform 1 0 13728 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_144
timestamp 1679581782
transform 1 0 14400 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_151
timestamp 1679581782
transform 1 0 15072 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_158
timestamp 1679581782
transform 1 0 15744 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_165
timestamp 1679581782
transform 1 0 16416 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_172
timestamp 1679581782
transform 1 0 17088 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_179
timestamp 1679581782
transform 1 0 17760 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_186
timestamp 1679581782
transform 1 0 18432 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_193
timestamp 1679581782
transform 1 0 19104 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_200
timestamp 1679581782
transform 1 0 19776 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_207
timestamp 1679581782
transform 1 0 20448 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_214
timestamp 1679581782
transform 1 0 21120 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_221
timestamp 1679581782
transform 1 0 21792 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_228
timestamp 1679581782
transform 1 0 22464 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_235
timestamp 1679581782
transform 1 0 23136 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_242
timestamp 1679581782
transform 1 0 23808 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_249
timestamp 1679581782
transform 1 0 24480 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_256
timestamp 1679581782
transform 1 0 25152 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_263
timestamp 1679581782
transform 1 0 25824 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_270
timestamp 1679581782
transform 1 0 26496 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_277
timestamp 1679581782
transform 1 0 27168 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_284
timestamp 1679581782
transform 1 0 27840 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_291
timestamp 1679581782
transform 1 0 28512 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_298
timestamp 1679581782
transform 1 0 29184 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_305
timestamp 1679581782
transform 1 0 29856 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_312
timestamp 1679581782
transform 1 0 30528 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_319
timestamp 1679581782
transform 1 0 31200 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_326
timestamp 1679581782
transform 1 0 31872 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_333
timestamp 1679581782
transform 1 0 32544 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_340
timestamp 1679581782
transform 1 0 33216 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_347
timestamp 1679581782
transform 1 0 33888 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_354
timestamp 1679581782
transform 1 0 34560 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_361
timestamp 1679581782
transform 1 0 35232 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_368
timestamp 1679581782
transform 1 0 35904 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_375
timestamp 1679581782
transform 1 0 36576 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_382
timestamp 1679581782
transform 1 0 37248 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_389
timestamp 1679581782
transform 1 0 37920 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_396
timestamp 1679581782
transform 1 0 38592 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_403
timestamp 1679581782
transform 1 0 39264 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_410
timestamp 1679581782
transform 1 0 39936 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_417
timestamp 1679581782
transform 1 0 40608 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_424
timestamp 1679581782
transform 1 0 41280 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_431
timestamp 1679581782
transform 1 0 41952 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_438
timestamp 1679581782
transform 1 0 42624 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_445
timestamp 1679581782
transform 1 0 43296 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_452
timestamp 1679581782
transform 1 0 43968 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_459
timestamp 1679581782
transform 1 0 44640 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_466
timestamp 1679581782
transform 1 0 45312 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_473
timestamp 1679581782
transform 1 0 45984 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_480
timestamp 1679581782
transform 1 0 46656 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_487
timestamp 1679581782
transform 1 0 47328 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_494
timestamp 1679581782
transform 1 0 48000 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_501
timestamp 1679581782
transform 1 0 48672 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_508
timestamp 1679581782
transform 1 0 49344 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_515
timestamp 1679581782
transform 1 0 50016 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_522
timestamp 1679581782
transform 1 0 50688 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_529
timestamp 1679581782
transform 1 0 51360 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_536
timestamp 1679581782
transform 1 0 52032 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_543
timestamp 1679581782
transform 1 0 52704 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_550
timestamp 1679581782
transform 1 0 53376 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_557
timestamp 1679581782
transform 1 0 54048 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_564
timestamp 1679581782
transform 1 0 54720 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_571
timestamp 1679581782
transform 1 0 55392 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_578
timestamp 1679581782
transform 1 0 56064 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_585
timestamp 1679581782
transform 1 0 56736 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_592
timestamp 1679581782
transform 1 0 57408 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_599
timestamp 1679581782
transform 1 0 58080 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_606
timestamp 1679581782
transform 1 0 58752 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_613
timestamp 1679581782
transform 1 0 59424 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_620
timestamp 1679581782
transform 1 0 60096 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_627
timestamp 1679581782
transform 1 0 60768 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_634
timestamp 1679581782
transform 1 0 61440 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_641
timestamp 1679581782
transform 1 0 62112 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_648
timestamp 1679581782
transform 1 0 62784 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_655
timestamp 1679581782
transform 1 0 63456 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_662
timestamp 1679581782
transform 1 0 64128 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_669
timestamp 1679581782
transform 1 0 64800 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_676
timestamp 1679581782
transform 1 0 65472 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_683
timestamp 1679581782
transform 1 0 66144 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_690
timestamp 1679581782
transform 1 0 66816 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_697
timestamp 1679581782
transform 1 0 67488 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_704
timestamp 1679581782
transform 1 0 68160 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_711
timestamp 1679581782
transform 1 0 68832 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_718
timestamp 1679581782
transform 1 0 69504 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_725
timestamp 1679581782
transform 1 0 70176 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_732
timestamp 1679581782
transform 1 0 70848 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_739
timestamp 1679581782
transform 1 0 71520 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_746
timestamp 1679581782
transform 1 0 72192 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_753
timestamp 1679581782
transform 1 0 72864 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_760
timestamp 1679581782
transform 1 0 73536 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_767
timestamp 1679581782
transform 1 0 74208 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_774
timestamp 1679581782
transform 1 0 74880 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_781
timestamp 1679581782
transform 1 0 75552 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_788
timestamp 1679581782
transform 1 0 76224 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_795
timestamp 1679581782
transform 1 0 76896 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_802
timestamp 1679581782
transform 1 0 77568 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_809
timestamp 1679581782
transform 1 0 78240 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_816
timestamp 1679581782
transform 1 0 78912 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_823
timestamp 1679581782
transform 1 0 79584 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_830
timestamp 1679581782
transform 1 0 80256 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_837
timestamp 1679581782
transform 1 0 80928 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_844
timestamp 1679581782
transform 1 0 81600 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_851
timestamp 1679581782
transform 1 0 82272 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_858
timestamp 1679581782
transform 1 0 82944 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_865
timestamp 1679581782
transform 1 0 83616 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_872
timestamp 1679581782
transform 1 0 84288 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_879
timestamp 1679581782
transform 1 0 84960 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_886
timestamp 1679581782
transform 1 0 85632 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_893
timestamp 1679581782
transform 1 0 86304 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_900
timestamp 1679581782
transform 1 0 86976 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_907
timestamp 1679581782
transform 1 0 87648 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_914
timestamp 1679581782
transform 1 0 88320 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_921
timestamp 1679581782
transform 1 0 88992 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_928
timestamp 1679581782
transform 1 0 89664 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_935
timestamp 1679581782
transform 1 0 90336 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_942
timestamp 1679581782
transform 1 0 91008 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_949
timestamp 1679581782
transform 1 0 91680 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_956
timestamp 1679581782
transform 1 0 92352 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_963
timestamp 1679581782
transform 1 0 93024 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_970
timestamp 1679581782
transform 1 0 93696 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_977
timestamp 1679581782
transform 1 0 94368 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_984
timestamp 1679581782
transform 1 0 95040 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_991
timestamp 1679581782
transform 1 0 95712 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_998
timestamp 1679581782
transform 1 0 96384 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_1005
timestamp 1679581782
transform 1 0 97056 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_1012
timestamp 1679581782
transform 1 0 97728 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_1019
timestamp 1679581782
transform 1 0 98400 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_1026
timestamp 1677580104
transform 1 0 99072 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_1028
timestamp 1677579658
transform 1 0 99264 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_0
timestamp 1679581782
transform 1 0 576 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_7
timestamp 1679581782
transform 1 0 1248 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_14
timestamp 1679581782
transform 1 0 1920 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_21
timestamp 1679581782
transform 1 0 2592 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_28
timestamp 1679581782
transform 1 0 3264 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_35
timestamp 1679581782
transform 1 0 3936 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_42
timestamp 1679581782
transform 1 0 4608 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_49
timestamp 1679581782
transform 1 0 5280 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_56
timestamp 1679581782
transform 1 0 5952 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_63
timestamp 1679581782
transform 1 0 6624 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_70
timestamp 1679581782
transform 1 0 7296 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_77
timestamp 1679581782
transform 1 0 7968 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_84
timestamp 1679581782
transform 1 0 8640 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_91
timestamp 1679581782
transform 1 0 9312 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_98
timestamp 1679581782
transform 1 0 9984 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_105
timestamp 1679581782
transform 1 0 10656 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_112
timestamp 1679581782
transform 1 0 11328 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_119
timestamp 1679581782
transform 1 0 12000 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_126
timestamp 1679581782
transform 1 0 12672 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_133
timestamp 1679581782
transform 1 0 13344 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_140
timestamp 1679581782
transform 1 0 14016 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_147
timestamp 1679581782
transform 1 0 14688 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_154
timestamp 1679581782
transform 1 0 15360 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_161
timestamp 1679581782
transform 1 0 16032 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_168
timestamp 1679581782
transform 1 0 16704 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_175
timestamp 1679581782
transform 1 0 17376 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_182
timestamp 1679581782
transform 1 0 18048 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_189
timestamp 1679581782
transform 1 0 18720 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_196
timestamp 1679581782
transform 1 0 19392 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_203
timestamp 1679581782
transform 1 0 20064 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_210
timestamp 1679581782
transform 1 0 20736 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_217
timestamp 1679581782
transform 1 0 21408 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_224
timestamp 1679581782
transform 1 0 22080 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_231
timestamp 1679581782
transform 1 0 22752 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_238
timestamp 1679581782
transform 1 0 23424 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_245
timestamp 1679581782
transform 1 0 24096 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_252
timestamp 1679581782
transform 1 0 24768 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_259
timestamp 1679581782
transform 1 0 25440 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_266
timestamp 1679581782
transform 1 0 26112 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_273
timestamp 1679581782
transform 1 0 26784 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_280
timestamp 1679581782
transform 1 0 27456 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_287
timestamp 1679581782
transform 1 0 28128 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_294
timestamp 1679581782
transform 1 0 28800 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_301
timestamp 1679581782
transform 1 0 29472 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_308
timestamp 1679581782
transform 1 0 30144 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_315
timestamp 1679581782
transform 1 0 30816 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_322
timestamp 1679581782
transform 1 0 31488 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_329
timestamp 1679581782
transform 1 0 32160 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_336
timestamp 1679581782
transform 1 0 32832 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_343
timestamp 1679581782
transform 1 0 33504 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_350
timestamp 1679581782
transform 1 0 34176 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_357
timestamp 1679581782
transform 1 0 34848 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_364
timestamp 1679581782
transform 1 0 35520 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_371
timestamp 1679581782
transform 1 0 36192 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_378
timestamp 1679581782
transform 1 0 36864 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_385
timestamp 1679581782
transform 1 0 37536 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_392
timestamp 1679581782
transform 1 0 38208 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_399
timestamp 1679581782
transform 1 0 38880 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_406
timestamp 1679581782
transform 1 0 39552 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_413
timestamp 1679581782
transform 1 0 40224 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_420
timestamp 1679581782
transform 1 0 40896 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_427
timestamp 1679581782
transform 1 0 41568 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_434
timestamp 1679581782
transform 1 0 42240 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_441
timestamp 1679581782
transform 1 0 42912 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_448
timestamp 1679581782
transform 1 0 43584 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_455
timestamp 1679581782
transform 1 0 44256 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_462
timestamp 1679581782
transform 1 0 44928 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_469
timestamp 1679581782
transform 1 0 45600 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_476
timestamp 1679581782
transform 1 0 46272 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_483
timestamp 1679581782
transform 1 0 46944 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_490
timestamp 1679581782
transform 1 0 47616 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_497
timestamp 1679581782
transform 1 0 48288 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_504
timestamp 1679581782
transform 1 0 48960 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_511
timestamp 1679581782
transform 1 0 49632 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_518
timestamp 1679581782
transform 1 0 50304 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_525
timestamp 1679581782
transform 1 0 50976 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_532
timestamp 1679581782
transform 1 0 51648 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_539
timestamp 1679581782
transform 1 0 52320 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_546
timestamp 1679581782
transform 1 0 52992 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_553
timestamp 1679581782
transform 1 0 53664 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_560
timestamp 1679581782
transform 1 0 54336 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_567
timestamp 1679581782
transform 1 0 55008 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_574
timestamp 1679581782
transform 1 0 55680 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_581
timestamp 1679581782
transform 1 0 56352 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_588
timestamp 1679581782
transform 1 0 57024 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_595
timestamp 1679581782
transform 1 0 57696 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_602
timestamp 1679581782
transform 1 0 58368 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_609
timestamp 1679581782
transform 1 0 59040 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_616
timestamp 1679581782
transform 1 0 59712 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_623
timestamp 1679581782
transform 1 0 60384 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_630
timestamp 1679581782
transform 1 0 61056 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_637
timestamp 1679581782
transform 1 0 61728 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_644
timestamp 1679581782
transform 1 0 62400 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_651
timestamp 1679581782
transform 1 0 63072 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_658
timestamp 1679581782
transform 1 0 63744 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_665
timestamp 1679581782
transform 1 0 64416 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_672
timestamp 1679581782
transform 1 0 65088 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_679
timestamp 1679581782
transform 1 0 65760 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_686
timestamp 1679581782
transform 1 0 66432 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_693
timestamp 1679581782
transform 1 0 67104 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_700
timestamp 1679581782
transform 1 0 67776 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_707
timestamp 1679581782
transform 1 0 68448 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_714
timestamp 1679581782
transform 1 0 69120 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_721
timestamp 1679581782
transform 1 0 69792 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_728
timestamp 1679581782
transform 1 0 70464 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_735
timestamp 1679581782
transform 1 0 71136 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_742
timestamp 1679581782
transform 1 0 71808 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_749
timestamp 1679581782
transform 1 0 72480 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_756
timestamp 1679581782
transform 1 0 73152 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_763
timestamp 1679581782
transform 1 0 73824 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_770
timestamp 1679581782
transform 1 0 74496 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_777
timestamp 1679581782
transform 1 0 75168 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_784
timestamp 1679581782
transform 1 0 75840 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_791
timestamp 1679581782
transform 1 0 76512 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_798
timestamp 1679581782
transform 1 0 77184 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_805
timestamp 1679581782
transform 1 0 77856 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_812
timestamp 1679581782
transform 1 0 78528 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_819
timestamp 1679581782
transform 1 0 79200 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_826
timestamp 1679581782
transform 1 0 79872 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_833
timestamp 1679581782
transform 1 0 80544 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_840
timestamp 1679581782
transform 1 0 81216 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_847
timestamp 1679581782
transform 1 0 81888 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_854
timestamp 1679581782
transform 1 0 82560 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_861
timestamp 1679581782
transform 1 0 83232 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_868
timestamp 1679581782
transform 1 0 83904 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_875
timestamp 1679581782
transform 1 0 84576 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_882
timestamp 1679581782
transform 1 0 85248 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_889
timestamp 1679581782
transform 1 0 85920 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_896
timestamp 1679581782
transform 1 0 86592 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_903
timestamp 1679581782
transform 1 0 87264 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_910
timestamp 1679581782
transform 1 0 87936 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_917
timestamp 1679581782
transform 1 0 88608 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_924
timestamp 1679581782
transform 1 0 89280 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_931
timestamp 1679581782
transform 1 0 89952 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_938
timestamp 1679581782
transform 1 0 90624 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_945
timestamp 1679581782
transform 1 0 91296 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_952
timestamp 1679581782
transform 1 0 91968 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_959
timestamp 1679581782
transform 1 0 92640 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_966
timestamp 1679581782
transform 1 0 93312 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_973
timestamp 1679581782
transform 1 0 93984 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_980
timestamp 1679581782
transform 1 0 94656 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_987
timestamp 1679581782
transform 1 0 95328 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_994
timestamp 1679581782
transform 1 0 96000 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_1001
timestamp 1679581782
transform 1 0 96672 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_1008
timestamp 1679581782
transform 1 0 97344 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_1015
timestamp 1679581782
transform 1 0 98016 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_1022
timestamp 1679581782
transform 1 0 98688 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_0
timestamp 1679581782
transform 1 0 576 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_7
timestamp 1679581782
transform 1 0 1248 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_14
timestamp 1679581782
transform 1 0 1920 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_21
timestamp 1679581782
transform 1 0 2592 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_28
timestamp 1679581782
transform 1 0 3264 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_35
timestamp 1679581782
transform 1 0 3936 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_42
timestamp 1679581782
transform 1 0 4608 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_49
timestamp 1679581782
transform 1 0 5280 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_56
timestamp 1679581782
transform 1 0 5952 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_63
timestamp 1679581782
transform 1 0 6624 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_70
timestamp 1679581782
transform 1 0 7296 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_77
timestamp 1679581782
transform 1 0 7968 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_84
timestamp 1679581782
transform 1 0 8640 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_91
timestamp 1679581782
transform 1 0 9312 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_98
timestamp 1679581782
transform 1 0 9984 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_105
timestamp 1679581782
transform 1 0 10656 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_112
timestamp 1679581782
transform 1 0 11328 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_119
timestamp 1679581782
transform 1 0 12000 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_126
timestamp 1679581782
transform 1 0 12672 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_133
timestamp 1679581782
transform 1 0 13344 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_140
timestamp 1679581782
transform 1 0 14016 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_147
timestamp 1679581782
transform 1 0 14688 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_154
timestamp 1679581782
transform 1 0 15360 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_161
timestamp 1679581782
transform 1 0 16032 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_168
timestamp 1679581782
transform 1 0 16704 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_175
timestamp 1679581782
transform 1 0 17376 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_182
timestamp 1679581782
transform 1 0 18048 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_189
timestamp 1679581782
transform 1 0 18720 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_196
timestamp 1679581782
transform 1 0 19392 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_203
timestamp 1679581782
transform 1 0 20064 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_210
timestamp 1679581782
transform 1 0 20736 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_217
timestamp 1679581782
transform 1 0 21408 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_224
timestamp 1679581782
transform 1 0 22080 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_231
timestamp 1679581782
transform 1 0 22752 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_238
timestamp 1679581782
transform 1 0 23424 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_245
timestamp 1679581782
transform 1 0 24096 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_252
timestamp 1679581782
transform 1 0 24768 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_259
timestamp 1679581782
transform 1 0 25440 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_266
timestamp 1679581782
transform 1 0 26112 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_273
timestamp 1679581782
transform 1 0 26784 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_280
timestamp 1679581782
transform 1 0 27456 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_287
timestamp 1679581782
transform 1 0 28128 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_294
timestamp 1679581782
transform 1 0 28800 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_301
timestamp 1679581782
transform 1 0 29472 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_308
timestamp 1679581782
transform 1 0 30144 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_315
timestamp 1679581782
transform 1 0 30816 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_322
timestamp 1679581782
transform 1 0 31488 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_329
timestamp 1679581782
transform 1 0 32160 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_336
timestamp 1679581782
transform 1 0 32832 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_343
timestamp 1679581782
transform 1 0 33504 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_350
timestamp 1679581782
transform 1 0 34176 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_357
timestamp 1679581782
transform 1 0 34848 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_364
timestamp 1679581782
transform 1 0 35520 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_371
timestamp 1679581782
transform 1 0 36192 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_378
timestamp 1679581782
transform 1 0 36864 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_385
timestamp 1679581782
transform 1 0 37536 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_392
timestamp 1679581782
transform 1 0 38208 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_399
timestamp 1679581782
transform 1 0 38880 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_406
timestamp 1679581782
transform 1 0 39552 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_413
timestamp 1679581782
transform 1 0 40224 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_420
timestamp 1679581782
transform 1 0 40896 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_427
timestamp 1679581782
transform 1 0 41568 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_434
timestamp 1679581782
transform 1 0 42240 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_441
timestamp 1679581782
transform 1 0 42912 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_448
timestamp 1679581782
transform 1 0 43584 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_455
timestamp 1679581782
transform 1 0 44256 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_462
timestamp 1679581782
transform 1 0 44928 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_469
timestamp 1679581782
transform 1 0 45600 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_476
timestamp 1679581782
transform 1 0 46272 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_483
timestamp 1679581782
transform 1 0 46944 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_490
timestamp 1679581782
transform 1 0 47616 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_497
timestamp 1679581782
transform 1 0 48288 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_504
timestamp 1679581782
transform 1 0 48960 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_511
timestamp 1679581782
transform 1 0 49632 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_518
timestamp 1679581782
transform 1 0 50304 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_525
timestamp 1679581782
transform 1 0 50976 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_532
timestamp 1679581782
transform 1 0 51648 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_539
timestamp 1679581782
transform 1 0 52320 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_546
timestamp 1679581782
transform 1 0 52992 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_553
timestamp 1679581782
transform 1 0 53664 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_560
timestamp 1679581782
transform 1 0 54336 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_567
timestamp 1679581782
transform 1 0 55008 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_574
timestamp 1679581782
transform 1 0 55680 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_581
timestamp 1679581782
transform 1 0 56352 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_588
timestamp 1679581782
transform 1 0 57024 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_595
timestamp 1679581782
transform 1 0 57696 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_602
timestamp 1679581782
transform 1 0 58368 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_609
timestamp 1679581782
transform 1 0 59040 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_616
timestamp 1679581782
transform 1 0 59712 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_623
timestamp 1679581782
transform 1 0 60384 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_630
timestamp 1679581782
transform 1 0 61056 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_637
timestamp 1679581782
transform 1 0 61728 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_644
timestamp 1679581782
transform 1 0 62400 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_651
timestamp 1679581782
transform 1 0 63072 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_658
timestamp 1679581782
transform 1 0 63744 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_665
timestamp 1679581782
transform 1 0 64416 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_672
timestamp 1679581782
transform 1 0 65088 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_679
timestamp 1679581782
transform 1 0 65760 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_686
timestamp 1679581782
transform 1 0 66432 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_693
timestamp 1679581782
transform 1 0 67104 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_700
timestamp 1679581782
transform 1 0 67776 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_707
timestamp 1679581782
transform 1 0 68448 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_714
timestamp 1679581782
transform 1 0 69120 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_721
timestamp 1679581782
transform 1 0 69792 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_728
timestamp 1679581782
transform 1 0 70464 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_735
timestamp 1679581782
transform 1 0 71136 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_742
timestamp 1679581782
transform 1 0 71808 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_749
timestamp 1679581782
transform 1 0 72480 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_756
timestamp 1679581782
transform 1 0 73152 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_763
timestamp 1679581782
transform 1 0 73824 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_770
timestamp 1679581782
transform 1 0 74496 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_777
timestamp 1679581782
transform 1 0 75168 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_784
timestamp 1679581782
transform 1 0 75840 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_791
timestamp 1679581782
transform 1 0 76512 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_798
timestamp 1679581782
transform 1 0 77184 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_805
timestamp 1679581782
transform 1 0 77856 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_812
timestamp 1679581782
transform 1 0 78528 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_819
timestamp 1679581782
transform 1 0 79200 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_826
timestamp 1679581782
transform 1 0 79872 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_833
timestamp 1679581782
transform 1 0 80544 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_840
timestamp 1679581782
transform 1 0 81216 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_847
timestamp 1679581782
transform 1 0 81888 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_854
timestamp 1679581782
transform 1 0 82560 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_861
timestamp 1679581782
transform 1 0 83232 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_868
timestamp 1679581782
transform 1 0 83904 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_875
timestamp 1679581782
transform 1 0 84576 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_882
timestamp 1679581782
transform 1 0 85248 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_889
timestamp 1679581782
transform 1 0 85920 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_896
timestamp 1679581782
transform 1 0 86592 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_903
timestamp 1679581782
transform 1 0 87264 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_910
timestamp 1679581782
transform 1 0 87936 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_917
timestamp 1679581782
transform 1 0 88608 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_924
timestamp 1679581782
transform 1 0 89280 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_931
timestamp 1679581782
transform 1 0 89952 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_938
timestamp 1679581782
transform 1 0 90624 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_945
timestamp 1679581782
transform 1 0 91296 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_952
timestamp 1679581782
transform 1 0 91968 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_959
timestamp 1679581782
transform 1 0 92640 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_966
timestamp 1679581782
transform 1 0 93312 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_973
timestamp 1679581782
transform 1 0 93984 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_980
timestamp 1679581782
transform 1 0 94656 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_987
timestamp 1679581782
transform 1 0 95328 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_994
timestamp 1679581782
transform 1 0 96000 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_1001
timestamp 1679581782
transform 1 0 96672 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_1008
timestamp 1679581782
transform 1 0 97344 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_1015
timestamp 1679581782
transform 1 0 98016 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_1022
timestamp 1679581782
transform 1 0 98688 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_4
timestamp 1679581782
transform 1 0 960 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_11
timestamp 1679581782
transform 1 0 1632 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_18
timestamp 1679581782
transform 1 0 2304 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_25
timestamp 1679581782
transform 1 0 2976 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_32
timestamp 1679581782
transform 1 0 3648 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_39
timestamp 1679581782
transform 1 0 4320 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_46
timestamp 1679581782
transform 1 0 4992 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_53
timestamp 1679581782
transform 1 0 5664 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_60
timestamp 1679581782
transform 1 0 6336 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_67
timestamp 1679581782
transform 1 0 7008 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_74
timestamp 1679581782
transform 1 0 7680 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_81
timestamp 1679581782
transform 1 0 8352 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_88
timestamp 1679581782
transform 1 0 9024 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_95
timestamp 1679581782
transform 1 0 9696 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_102
timestamp 1679581782
transform 1 0 10368 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_109
timestamp 1679581782
transform 1 0 11040 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_116
timestamp 1679581782
transform 1 0 11712 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_123
timestamp 1679581782
transform 1 0 12384 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_130
timestamp 1679581782
transform 1 0 13056 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_137
timestamp 1679581782
transform 1 0 13728 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_144
timestamp 1679581782
transform 1 0 14400 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_151
timestamp 1679581782
transform 1 0 15072 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_158
timestamp 1679581782
transform 1 0 15744 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_165
timestamp 1679581782
transform 1 0 16416 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_172
timestamp 1679581782
transform 1 0 17088 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_179
timestamp 1679581782
transform 1 0 17760 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_186
timestamp 1679581782
transform 1 0 18432 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_193
timestamp 1679581782
transform 1 0 19104 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_200
timestamp 1679581782
transform 1 0 19776 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_207
timestamp 1679581782
transform 1 0 20448 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_214
timestamp 1679581782
transform 1 0 21120 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_221
timestamp 1679581782
transform 1 0 21792 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_228
timestamp 1679581782
transform 1 0 22464 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_235
timestamp 1679581782
transform 1 0 23136 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_242
timestamp 1679581782
transform 1 0 23808 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_249
timestamp 1679581782
transform 1 0 24480 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_256
timestamp 1679581782
transform 1 0 25152 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_263
timestamp 1679581782
transform 1 0 25824 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_270
timestamp 1679581782
transform 1 0 26496 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_277
timestamp 1679581782
transform 1 0 27168 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_284
timestamp 1679581782
transform 1 0 27840 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_291
timestamp 1679581782
transform 1 0 28512 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_298
timestamp 1679581782
transform 1 0 29184 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_305
timestamp 1679581782
transform 1 0 29856 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_312
timestamp 1679581782
transform 1 0 30528 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_319
timestamp 1679581782
transform 1 0 31200 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_326
timestamp 1679581782
transform 1 0 31872 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_333
timestamp 1679581782
transform 1 0 32544 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_340
timestamp 1679581782
transform 1 0 33216 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_347
timestamp 1679581782
transform 1 0 33888 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_354
timestamp 1679581782
transform 1 0 34560 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_361
timestamp 1679581782
transform 1 0 35232 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_368
timestamp 1679581782
transform 1 0 35904 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_375
timestamp 1679581782
transform 1 0 36576 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_382
timestamp 1679581782
transform 1 0 37248 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_389
timestamp 1679581782
transform 1 0 37920 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_396
timestamp 1679581782
transform 1 0 38592 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_403
timestamp 1679581782
transform 1 0 39264 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_410
timestamp 1679581782
transform 1 0 39936 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_417
timestamp 1679581782
transform 1 0 40608 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_424
timestamp 1679581782
transform 1 0 41280 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_431
timestamp 1679581782
transform 1 0 41952 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_438
timestamp 1679581782
transform 1 0 42624 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_445
timestamp 1679581782
transform 1 0 43296 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_452
timestamp 1679581782
transform 1 0 43968 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_459
timestamp 1679581782
transform 1 0 44640 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_466
timestamp 1679581782
transform 1 0 45312 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_473
timestamp 1679581782
transform 1 0 45984 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_480
timestamp 1679581782
transform 1 0 46656 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_487
timestamp 1679581782
transform 1 0 47328 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_494
timestamp 1679581782
transform 1 0 48000 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_501
timestamp 1679581782
transform 1 0 48672 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_508
timestamp 1679581782
transform 1 0 49344 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_515
timestamp 1679581782
transform 1 0 50016 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_522
timestamp 1679581782
transform 1 0 50688 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_529
timestamp 1679581782
transform 1 0 51360 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_536
timestamp 1679581782
transform 1 0 52032 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_543
timestamp 1679581782
transform 1 0 52704 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_550
timestamp 1679581782
transform 1 0 53376 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_557
timestamp 1679581782
transform 1 0 54048 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_564
timestamp 1679581782
transform 1 0 54720 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_571
timestamp 1679581782
transform 1 0 55392 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_578
timestamp 1679581782
transform 1 0 56064 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_585
timestamp 1679581782
transform 1 0 56736 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_592
timestamp 1679581782
transform 1 0 57408 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_599
timestamp 1679581782
transform 1 0 58080 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_606
timestamp 1679581782
transform 1 0 58752 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_613
timestamp 1679581782
transform 1 0 59424 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_620
timestamp 1679581782
transform 1 0 60096 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_627
timestamp 1679581782
transform 1 0 60768 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_634
timestamp 1679581782
transform 1 0 61440 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_641
timestamp 1679581782
transform 1 0 62112 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_648
timestamp 1679581782
transform 1 0 62784 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_655
timestamp 1679581782
transform 1 0 63456 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_662
timestamp 1679581782
transform 1 0 64128 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_669
timestamp 1679581782
transform 1 0 64800 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_676
timestamp 1679581782
transform 1 0 65472 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_683
timestamp 1679581782
transform 1 0 66144 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_690
timestamp 1679581782
transform 1 0 66816 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_697
timestamp 1679581782
transform 1 0 67488 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_704
timestamp 1679581782
transform 1 0 68160 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_711
timestamp 1679581782
transform 1 0 68832 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_718
timestamp 1679581782
transform 1 0 69504 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_725
timestamp 1679581782
transform 1 0 70176 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_732
timestamp 1679581782
transform 1 0 70848 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_739
timestamp 1679581782
transform 1 0 71520 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_746
timestamp 1679581782
transform 1 0 72192 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_753
timestamp 1679581782
transform 1 0 72864 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_760
timestamp 1679581782
transform 1 0 73536 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_767
timestamp 1679581782
transform 1 0 74208 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_774
timestamp 1679581782
transform 1 0 74880 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_781
timestamp 1679581782
transform 1 0 75552 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_788
timestamp 1679581782
transform 1 0 76224 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_795
timestamp 1679581782
transform 1 0 76896 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_802
timestamp 1679581782
transform 1 0 77568 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_809
timestamp 1679581782
transform 1 0 78240 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_816
timestamp 1679581782
transform 1 0 78912 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_823
timestamp 1679581782
transform 1 0 79584 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_830
timestamp 1679581782
transform 1 0 80256 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_837
timestamp 1679581782
transform 1 0 80928 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_844
timestamp 1679581782
transform 1 0 81600 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_851
timestamp 1679581782
transform 1 0 82272 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_858
timestamp 1679581782
transform 1 0 82944 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_865
timestamp 1679581782
transform 1 0 83616 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_872
timestamp 1679581782
transform 1 0 84288 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_879
timestamp 1679581782
transform 1 0 84960 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_886
timestamp 1679581782
transform 1 0 85632 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_893
timestamp 1679581782
transform 1 0 86304 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_900
timestamp 1679581782
transform 1 0 86976 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_907
timestamp 1679581782
transform 1 0 87648 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_914
timestamp 1679581782
transform 1 0 88320 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_921
timestamp 1679581782
transform 1 0 88992 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_928
timestamp 1679581782
transform 1 0 89664 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_935
timestamp 1679581782
transform 1 0 90336 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_942
timestamp 1679581782
transform 1 0 91008 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_949
timestamp 1679581782
transform 1 0 91680 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_956
timestamp 1679581782
transform 1 0 92352 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_963
timestamp 1679581782
transform 1 0 93024 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_970
timestamp 1679581782
transform 1 0 93696 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_977
timestamp 1679581782
transform 1 0 94368 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_984
timestamp 1679581782
transform 1 0 95040 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_991
timestamp 1679581782
transform 1 0 95712 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_998
timestamp 1679581782
transform 1 0 96384 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_1005
timestamp 1679581782
transform 1 0 97056 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_1012
timestamp 1679581782
transform 1 0 97728 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_1019
timestamp 1679581782
transform 1 0 98400 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_1026
timestamp 1677580104
transform 1 0 99072 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_1028
timestamp 1677579658
transform 1 0 99264 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_0
timestamp 1679581782
transform 1 0 576 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_7
timestamp 1679581782
transform 1 0 1248 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_14
timestamp 1679581782
transform 1 0 1920 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_21
timestamp 1679581782
transform 1 0 2592 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_28
timestamp 1679581782
transform 1 0 3264 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_35
timestamp 1679581782
transform 1 0 3936 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_42
timestamp 1679581782
transform 1 0 4608 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_49
timestamp 1679581782
transform 1 0 5280 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_56
timestamp 1679581782
transform 1 0 5952 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_63
timestamp 1679581782
transform 1 0 6624 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_70
timestamp 1679581782
transform 1 0 7296 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_77
timestamp 1679581782
transform 1 0 7968 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_84
timestamp 1679581782
transform 1 0 8640 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_91
timestamp 1679581782
transform 1 0 9312 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_98
timestamp 1679581782
transform 1 0 9984 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_105
timestamp 1679581782
transform 1 0 10656 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_112
timestamp 1679581782
transform 1 0 11328 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_119
timestamp 1679581782
transform 1 0 12000 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_126
timestamp 1679581782
transform 1 0 12672 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_133
timestamp 1679581782
transform 1 0 13344 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_140
timestamp 1679581782
transform 1 0 14016 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_147
timestamp 1679581782
transform 1 0 14688 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_154
timestamp 1679581782
transform 1 0 15360 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_161
timestamp 1679581782
transform 1 0 16032 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_168
timestamp 1679581782
transform 1 0 16704 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_175
timestamp 1679581782
transform 1 0 17376 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_182
timestamp 1679581782
transform 1 0 18048 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_189
timestamp 1679581782
transform 1 0 18720 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_196
timestamp 1679581782
transform 1 0 19392 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_203
timestamp 1679581782
transform 1 0 20064 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_210
timestamp 1679581782
transform 1 0 20736 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_217
timestamp 1679581782
transform 1 0 21408 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_224
timestamp 1679581782
transform 1 0 22080 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_231
timestamp 1679581782
transform 1 0 22752 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_238
timestamp 1679581782
transform 1 0 23424 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_245
timestamp 1679581782
transform 1 0 24096 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_252
timestamp 1679581782
transform 1 0 24768 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_259
timestamp 1679581782
transform 1 0 25440 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_266
timestamp 1679581782
transform 1 0 26112 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_273
timestamp 1679581782
transform 1 0 26784 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_280
timestamp 1679581782
transform 1 0 27456 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_287
timestamp 1679581782
transform 1 0 28128 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_294
timestamp 1679581782
transform 1 0 28800 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_301
timestamp 1679581782
transform 1 0 29472 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_308
timestamp 1679581782
transform 1 0 30144 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_315
timestamp 1679581782
transform 1 0 30816 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_322
timestamp 1679581782
transform 1 0 31488 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_329
timestamp 1679581782
transform 1 0 32160 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_336
timestamp 1679581782
transform 1 0 32832 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_343
timestamp 1679581782
transform 1 0 33504 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_350
timestamp 1679581782
transform 1 0 34176 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_357
timestamp 1679581782
transform 1 0 34848 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_364
timestamp 1679581782
transform 1 0 35520 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_371
timestamp 1679581782
transform 1 0 36192 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_378
timestamp 1679581782
transform 1 0 36864 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_385
timestamp 1679581782
transform 1 0 37536 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_392
timestamp 1679581782
transform 1 0 38208 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_399
timestamp 1679581782
transform 1 0 38880 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_406
timestamp 1679581782
transform 1 0 39552 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_413
timestamp 1679581782
transform 1 0 40224 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_420
timestamp 1679581782
transform 1 0 40896 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_427
timestamp 1679581782
transform 1 0 41568 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_434
timestamp 1679581782
transform 1 0 42240 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_441
timestamp 1679581782
transform 1 0 42912 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_448
timestamp 1679581782
transform 1 0 43584 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_455
timestamp 1679581782
transform 1 0 44256 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_462
timestamp 1679581782
transform 1 0 44928 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_469
timestamp 1679581782
transform 1 0 45600 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_476
timestamp 1679581782
transform 1 0 46272 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_483
timestamp 1679581782
transform 1 0 46944 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_490
timestamp 1679581782
transform 1 0 47616 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_497
timestamp 1679581782
transform 1 0 48288 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_504
timestamp 1679581782
transform 1 0 48960 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_511
timestamp 1679581782
transform 1 0 49632 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_518
timestamp 1679581782
transform 1 0 50304 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_525
timestamp 1679581782
transform 1 0 50976 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_532
timestamp 1679581782
transform 1 0 51648 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_539
timestamp 1679581782
transform 1 0 52320 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_546
timestamp 1679581782
transform 1 0 52992 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_553
timestamp 1679581782
transform 1 0 53664 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_560
timestamp 1679581782
transform 1 0 54336 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_567
timestamp 1679581782
transform 1 0 55008 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_574
timestamp 1679581782
transform 1 0 55680 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_581
timestamp 1679581782
transform 1 0 56352 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_588
timestamp 1679581782
transform 1 0 57024 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_595
timestamp 1679581782
transform 1 0 57696 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_602
timestamp 1679581782
transform 1 0 58368 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_609
timestamp 1679581782
transform 1 0 59040 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_616
timestamp 1679581782
transform 1 0 59712 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_623
timestamp 1679581782
transform 1 0 60384 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_630
timestamp 1679581782
transform 1 0 61056 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_637
timestamp 1679581782
transform 1 0 61728 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_644
timestamp 1679581782
transform 1 0 62400 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_651
timestamp 1679581782
transform 1 0 63072 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_658
timestamp 1679581782
transform 1 0 63744 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_665
timestamp 1679581782
transform 1 0 64416 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_672
timestamp 1679581782
transform 1 0 65088 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_679
timestamp 1679581782
transform 1 0 65760 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_686
timestamp 1679581782
transform 1 0 66432 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_693
timestamp 1679581782
transform 1 0 67104 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_700
timestamp 1679581782
transform 1 0 67776 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_707
timestamp 1679581782
transform 1 0 68448 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_714
timestamp 1679581782
transform 1 0 69120 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_721
timestamp 1679581782
transform 1 0 69792 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_728
timestamp 1679581782
transform 1 0 70464 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_735
timestamp 1679581782
transform 1 0 71136 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_742
timestamp 1679581782
transform 1 0 71808 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_749
timestamp 1679581782
transform 1 0 72480 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_756
timestamp 1679581782
transform 1 0 73152 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_763
timestamp 1679581782
transform 1 0 73824 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_770
timestamp 1679581782
transform 1 0 74496 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_777
timestamp 1679581782
transform 1 0 75168 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_784
timestamp 1679581782
transform 1 0 75840 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_791
timestamp 1679581782
transform 1 0 76512 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_798
timestamp 1679581782
transform 1 0 77184 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_805
timestamp 1679581782
transform 1 0 77856 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_812
timestamp 1679581782
transform 1 0 78528 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_819
timestamp 1679581782
transform 1 0 79200 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_826
timestamp 1679581782
transform 1 0 79872 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_833
timestamp 1679581782
transform 1 0 80544 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_840
timestamp 1679581782
transform 1 0 81216 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_847
timestamp 1679581782
transform 1 0 81888 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_854
timestamp 1679581782
transform 1 0 82560 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_861
timestamp 1679581782
transform 1 0 83232 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_868
timestamp 1679581782
transform 1 0 83904 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_875
timestamp 1679581782
transform 1 0 84576 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_882
timestamp 1679581782
transform 1 0 85248 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_889
timestamp 1679581782
transform 1 0 85920 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_896
timestamp 1679581782
transform 1 0 86592 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_903
timestamp 1679581782
transform 1 0 87264 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_910
timestamp 1679581782
transform 1 0 87936 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_917
timestamp 1679581782
transform 1 0 88608 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_924
timestamp 1679581782
transform 1 0 89280 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_931
timestamp 1679581782
transform 1 0 89952 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_938
timestamp 1679581782
transform 1 0 90624 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_945
timestamp 1679581782
transform 1 0 91296 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_952
timestamp 1679581782
transform 1 0 91968 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_959
timestamp 1679581782
transform 1 0 92640 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_966
timestamp 1679581782
transform 1 0 93312 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_973
timestamp 1679581782
transform 1 0 93984 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_980
timestamp 1679581782
transform 1 0 94656 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_987
timestamp 1679581782
transform 1 0 95328 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_994
timestamp 1679581782
transform 1 0 96000 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_1001
timestamp 1679581782
transform 1 0 96672 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_1008
timestamp 1679581782
transform 1 0 97344 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_1015
timestamp 1679581782
transform 1 0 98016 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_1022
timestamp 1679581782
transform 1 0 98688 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_4
timestamp 1679581782
transform 1 0 960 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_11
timestamp 1679581782
transform 1 0 1632 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_18
timestamp 1679581782
transform 1 0 2304 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_25
timestamp 1679581782
transform 1 0 2976 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_32
timestamp 1679581782
transform 1 0 3648 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_39
timestamp 1679581782
transform 1 0 4320 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_46
timestamp 1679581782
transform 1 0 4992 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_53
timestamp 1679581782
transform 1 0 5664 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_60
timestamp 1679581782
transform 1 0 6336 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_67
timestamp 1679581782
transform 1 0 7008 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_74
timestamp 1679581782
transform 1 0 7680 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_81
timestamp 1679581782
transform 1 0 8352 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_88
timestamp 1679581782
transform 1 0 9024 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_95
timestamp 1679581782
transform 1 0 9696 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_102
timestamp 1679581782
transform 1 0 10368 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_109
timestamp 1679581782
transform 1 0 11040 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_116
timestamp 1679581782
transform 1 0 11712 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_123
timestamp 1679581782
transform 1 0 12384 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_130
timestamp 1679581782
transform 1 0 13056 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_137
timestamp 1679581782
transform 1 0 13728 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_144
timestamp 1679581782
transform 1 0 14400 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_151
timestamp 1679581782
transform 1 0 15072 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_158
timestamp 1679581782
transform 1 0 15744 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_165
timestamp 1679581782
transform 1 0 16416 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_172
timestamp 1679581782
transform 1 0 17088 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_179
timestamp 1679581782
transform 1 0 17760 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_186
timestamp 1679581782
transform 1 0 18432 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_193
timestamp 1679581782
transform 1 0 19104 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_200
timestamp 1679581782
transform 1 0 19776 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_207
timestamp 1679581782
transform 1 0 20448 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_214
timestamp 1679581782
transform 1 0 21120 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_221
timestamp 1679581782
transform 1 0 21792 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_228
timestamp 1679581782
transform 1 0 22464 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_235
timestamp 1679581782
transform 1 0 23136 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_242
timestamp 1679581782
transform 1 0 23808 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_249
timestamp 1679581782
transform 1 0 24480 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_256
timestamp 1679581782
transform 1 0 25152 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_263
timestamp 1679581782
transform 1 0 25824 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_270
timestamp 1679581782
transform 1 0 26496 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_277
timestamp 1679581782
transform 1 0 27168 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_284
timestamp 1679581782
transform 1 0 27840 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_291
timestamp 1679581782
transform 1 0 28512 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_298
timestamp 1679581782
transform 1 0 29184 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_305
timestamp 1679581782
transform 1 0 29856 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_312
timestamp 1679581782
transform 1 0 30528 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_319
timestamp 1679581782
transform 1 0 31200 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_326
timestamp 1679581782
transform 1 0 31872 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_333
timestamp 1679581782
transform 1 0 32544 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_340
timestamp 1679581782
transform 1 0 33216 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_347
timestamp 1679581782
transform 1 0 33888 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_354
timestamp 1679581782
transform 1 0 34560 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_361
timestamp 1679581782
transform 1 0 35232 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_368
timestamp 1679581782
transform 1 0 35904 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_375
timestamp 1679581782
transform 1 0 36576 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_382
timestamp 1679581782
transform 1 0 37248 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_389
timestamp 1679581782
transform 1 0 37920 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_396
timestamp 1679581782
transform 1 0 38592 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_403
timestamp 1679581782
transform 1 0 39264 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_410
timestamp 1679581782
transform 1 0 39936 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_417
timestamp 1679581782
transform 1 0 40608 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_424
timestamp 1679581782
transform 1 0 41280 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_431
timestamp 1679581782
transform 1 0 41952 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_438
timestamp 1679581782
transform 1 0 42624 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_445
timestamp 1679581782
transform 1 0 43296 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_452
timestamp 1679581782
transform 1 0 43968 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_459
timestamp 1679581782
transform 1 0 44640 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_466
timestamp 1679581782
transform 1 0 45312 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_473
timestamp 1679581782
transform 1 0 45984 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_480
timestamp 1679581782
transform 1 0 46656 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_487
timestamp 1679581782
transform 1 0 47328 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_494
timestamp 1679581782
transform 1 0 48000 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_501
timestamp 1679581782
transform 1 0 48672 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_508
timestamp 1679581782
transform 1 0 49344 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_515
timestamp 1679581782
transform 1 0 50016 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_522
timestamp 1679581782
transform 1 0 50688 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_529
timestamp 1679581782
transform 1 0 51360 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_536
timestamp 1679581782
transform 1 0 52032 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_543
timestamp 1679581782
transform 1 0 52704 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_550
timestamp 1679581782
transform 1 0 53376 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_557
timestamp 1679581782
transform 1 0 54048 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_564
timestamp 1679581782
transform 1 0 54720 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_571
timestamp 1679581782
transform 1 0 55392 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_578
timestamp 1679581782
transform 1 0 56064 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_585
timestamp 1679581782
transform 1 0 56736 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_592
timestamp 1679581782
transform 1 0 57408 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_599
timestamp 1679581782
transform 1 0 58080 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_606
timestamp 1679581782
transform 1 0 58752 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_613
timestamp 1679581782
transform 1 0 59424 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_620
timestamp 1679581782
transform 1 0 60096 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_627
timestamp 1679581782
transform 1 0 60768 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_634
timestamp 1679581782
transform 1 0 61440 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_641
timestamp 1679581782
transform 1 0 62112 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_648
timestamp 1679581782
transform 1 0 62784 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_655
timestamp 1679581782
transform 1 0 63456 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_662
timestamp 1679581782
transform 1 0 64128 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_669
timestamp 1679581782
transform 1 0 64800 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_676
timestamp 1679581782
transform 1 0 65472 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_683
timestamp 1679581782
transform 1 0 66144 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_690
timestamp 1679581782
transform 1 0 66816 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_697
timestamp 1679581782
transform 1 0 67488 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_704
timestamp 1679581782
transform 1 0 68160 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_711
timestamp 1679581782
transform 1 0 68832 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_718
timestamp 1679581782
transform 1 0 69504 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_725
timestamp 1679581782
transform 1 0 70176 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_732
timestamp 1679581782
transform 1 0 70848 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_739
timestamp 1679581782
transform 1 0 71520 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_746
timestamp 1679581782
transform 1 0 72192 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_753
timestamp 1679581782
transform 1 0 72864 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_760
timestamp 1679581782
transform 1 0 73536 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_767
timestamp 1679581782
transform 1 0 74208 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_774
timestamp 1679581782
transform 1 0 74880 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_781
timestamp 1679581782
transform 1 0 75552 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_788
timestamp 1679581782
transform 1 0 76224 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_795
timestamp 1679581782
transform 1 0 76896 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_802
timestamp 1679581782
transform 1 0 77568 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_809
timestamp 1679581782
transform 1 0 78240 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_816
timestamp 1679581782
transform 1 0 78912 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_823
timestamp 1679581782
transform 1 0 79584 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_830
timestamp 1679581782
transform 1 0 80256 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_837
timestamp 1679581782
transform 1 0 80928 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_844
timestamp 1679581782
transform 1 0 81600 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_851
timestamp 1679581782
transform 1 0 82272 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_858
timestamp 1679581782
transform 1 0 82944 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_865
timestamp 1679581782
transform 1 0 83616 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_872
timestamp 1679581782
transform 1 0 84288 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_879
timestamp 1679581782
transform 1 0 84960 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_886
timestamp 1679581782
transform 1 0 85632 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_893
timestamp 1679581782
transform 1 0 86304 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_900
timestamp 1679581782
transform 1 0 86976 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_907
timestamp 1679581782
transform 1 0 87648 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_914
timestamp 1679581782
transform 1 0 88320 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_921
timestamp 1679581782
transform 1 0 88992 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_928
timestamp 1679581782
transform 1 0 89664 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_935
timestamp 1679581782
transform 1 0 90336 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_942
timestamp 1679581782
transform 1 0 91008 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_949
timestamp 1679581782
transform 1 0 91680 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_956
timestamp 1679581782
transform 1 0 92352 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_963
timestamp 1679581782
transform 1 0 93024 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_970
timestamp 1679581782
transform 1 0 93696 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_977
timestamp 1679581782
transform 1 0 94368 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_984
timestamp 1679581782
transform 1 0 95040 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_991
timestamp 1679581782
transform 1 0 95712 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_998
timestamp 1679581782
transform 1 0 96384 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_1005
timestamp 1679581782
transform 1 0 97056 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_1012
timestamp 1679581782
transform 1 0 97728 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_1019
timestamp 1679581782
transform 1 0 98400 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_1026
timestamp 1677580104
transform 1 0 99072 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_1028
timestamp 1677579658
transform 1 0 99264 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_0
timestamp 1679581782
transform 1 0 576 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_7
timestamp 1679581782
transform 1 0 1248 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_14
timestamp 1679581782
transform 1 0 1920 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_21
timestamp 1679581782
transform 1 0 2592 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_28
timestamp 1679581782
transform 1 0 3264 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_35
timestamp 1679581782
transform 1 0 3936 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_42
timestamp 1679581782
transform 1 0 4608 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_49
timestamp 1679581782
transform 1 0 5280 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_56
timestamp 1679581782
transform 1 0 5952 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_63
timestamp 1679581782
transform 1 0 6624 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_70
timestamp 1679581782
transform 1 0 7296 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_77
timestamp 1679581782
transform 1 0 7968 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_84
timestamp 1679581782
transform 1 0 8640 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_91
timestamp 1679581782
transform 1 0 9312 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_98
timestamp 1679581782
transform 1 0 9984 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_105
timestamp 1679581782
transform 1 0 10656 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_112
timestamp 1679581782
transform 1 0 11328 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_119
timestamp 1679581782
transform 1 0 12000 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_126
timestamp 1679581782
transform 1 0 12672 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_133
timestamp 1679581782
transform 1 0 13344 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_140
timestamp 1679581782
transform 1 0 14016 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_147
timestamp 1679581782
transform 1 0 14688 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_154
timestamp 1679581782
transform 1 0 15360 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_161
timestamp 1679581782
transform 1 0 16032 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_168
timestamp 1679581782
transform 1 0 16704 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_175
timestamp 1679581782
transform 1 0 17376 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_182
timestamp 1679581782
transform 1 0 18048 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_189
timestamp 1679581782
transform 1 0 18720 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_196
timestamp 1679581782
transform 1 0 19392 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_203
timestamp 1679581782
transform 1 0 20064 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_210
timestamp 1679581782
transform 1 0 20736 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_217
timestamp 1679581782
transform 1 0 21408 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_224
timestamp 1679581782
transform 1 0 22080 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_231
timestamp 1679581782
transform 1 0 22752 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_238
timestamp 1679581782
transform 1 0 23424 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_245
timestamp 1679581782
transform 1 0 24096 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_252
timestamp 1679581782
transform 1 0 24768 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_259
timestamp 1679581782
transform 1 0 25440 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_266
timestamp 1679581782
transform 1 0 26112 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_273
timestamp 1679581782
transform 1 0 26784 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_280
timestamp 1679581782
transform 1 0 27456 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_287
timestamp 1679581782
transform 1 0 28128 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_294
timestamp 1679581782
transform 1 0 28800 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_301
timestamp 1679581782
transform 1 0 29472 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_308
timestamp 1679581782
transform 1 0 30144 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_315
timestamp 1679581782
transform 1 0 30816 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_322
timestamp 1679581782
transform 1 0 31488 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_329
timestamp 1679581782
transform 1 0 32160 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_336
timestamp 1679581782
transform 1 0 32832 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_343
timestamp 1679581782
transform 1 0 33504 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_350
timestamp 1679581782
transform 1 0 34176 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_357
timestamp 1679581782
transform 1 0 34848 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_364
timestamp 1679581782
transform 1 0 35520 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_371
timestamp 1679581782
transform 1 0 36192 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_378
timestamp 1679581782
transform 1 0 36864 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_385
timestamp 1679581782
transform 1 0 37536 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_392
timestamp 1679581782
transform 1 0 38208 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_399
timestamp 1679581782
transform 1 0 38880 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_406
timestamp 1679581782
transform 1 0 39552 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_413
timestamp 1679581782
transform 1 0 40224 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_420
timestamp 1679581782
transform 1 0 40896 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_427
timestamp 1679581782
transform 1 0 41568 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_434
timestamp 1679581782
transform 1 0 42240 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_441
timestamp 1679581782
transform 1 0 42912 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_448
timestamp 1679581782
transform 1 0 43584 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_455
timestamp 1679581782
transform 1 0 44256 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_462
timestamp 1679581782
transform 1 0 44928 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_469
timestamp 1679581782
transform 1 0 45600 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_476
timestamp 1679581782
transform 1 0 46272 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_483
timestamp 1679581782
transform 1 0 46944 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_490
timestamp 1679581782
transform 1 0 47616 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_497
timestamp 1679581782
transform 1 0 48288 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_504
timestamp 1679581782
transform 1 0 48960 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_511
timestamp 1679581782
transform 1 0 49632 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_518
timestamp 1679581782
transform 1 0 50304 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_525
timestamp 1679581782
transform 1 0 50976 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_532
timestamp 1679581782
transform 1 0 51648 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_539
timestamp 1679581782
transform 1 0 52320 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_546
timestamp 1679581782
transform 1 0 52992 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_553
timestamp 1679581782
transform 1 0 53664 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_560
timestamp 1679581782
transform 1 0 54336 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_567
timestamp 1679581782
transform 1 0 55008 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_574
timestamp 1679581782
transform 1 0 55680 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_581
timestamp 1679581782
transform 1 0 56352 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_588
timestamp 1679581782
transform 1 0 57024 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_595
timestamp 1679581782
transform 1 0 57696 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_602
timestamp 1679581782
transform 1 0 58368 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_609
timestamp 1679581782
transform 1 0 59040 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_616
timestamp 1679581782
transform 1 0 59712 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_623
timestamp 1679581782
transform 1 0 60384 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_630
timestamp 1679581782
transform 1 0 61056 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_637
timestamp 1679581782
transform 1 0 61728 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_644
timestamp 1679581782
transform 1 0 62400 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_651
timestamp 1679581782
transform 1 0 63072 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_658
timestamp 1679581782
transform 1 0 63744 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_665
timestamp 1679581782
transform 1 0 64416 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_672
timestamp 1679581782
transform 1 0 65088 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_679
timestamp 1679581782
transform 1 0 65760 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_686
timestamp 1679581782
transform 1 0 66432 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_693
timestamp 1679581782
transform 1 0 67104 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_700
timestamp 1679581782
transform 1 0 67776 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_707
timestamp 1679581782
transform 1 0 68448 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_714
timestamp 1679581782
transform 1 0 69120 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_721
timestamp 1679581782
transform 1 0 69792 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_728
timestamp 1679581782
transform 1 0 70464 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_735
timestamp 1679581782
transform 1 0 71136 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_742
timestamp 1679581782
transform 1 0 71808 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_749
timestamp 1679581782
transform 1 0 72480 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_756
timestamp 1679581782
transform 1 0 73152 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_763
timestamp 1679581782
transform 1 0 73824 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_770
timestamp 1679581782
transform 1 0 74496 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_777
timestamp 1679581782
transform 1 0 75168 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_784
timestamp 1679581782
transform 1 0 75840 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_791
timestamp 1679581782
transform 1 0 76512 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_798
timestamp 1679581782
transform 1 0 77184 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_805
timestamp 1679581782
transform 1 0 77856 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_812
timestamp 1679581782
transform 1 0 78528 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_819
timestamp 1679581782
transform 1 0 79200 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_826
timestamp 1679581782
transform 1 0 79872 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_833
timestamp 1679581782
transform 1 0 80544 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_840
timestamp 1679581782
transform 1 0 81216 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_847
timestamp 1679581782
transform 1 0 81888 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_854
timestamp 1679581782
transform 1 0 82560 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_861
timestamp 1679581782
transform 1 0 83232 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_868
timestamp 1679581782
transform 1 0 83904 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_875
timestamp 1679581782
transform 1 0 84576 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_882
timestamp 1679581782
transform 1 0 85248 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_889
timestamp 1679581782
transform 1 0 85920 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_896
timestamp 1679581782
transform 1 0 86592 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_903
timestamp 1679581782
transform 1 0 87264 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_910
timestamp 1679581782
transform 1 0 87936 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_917
timestamp 1679581782
transform 1 0 88608 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_924
timestamp 1679581782
transform 1 0 89280 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_931
timestamp 1679581782
transform 1 0 89952 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_938
timestamp 1679581782
transform 1 0 90624 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_945
timestamp 1679581782
transform 1 0 91296 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_952
timestamp 1679581782
transform 1 0 91968 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_959
timestamp 1679581782
transform 1 0 92640 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_966
timestamp 1679581782
transform 1 0 93312 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_973
timestamp 1679581782
transform 1 0 93984 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_980
timestamp 1679581782
transform 1 0 94656 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_987
timestamp 1679581782
transform 1 0 95328 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_994
timestamp 1679581782
transform 1 0 96000 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_1001
timestamp 1679581782
transform 1 0 96672 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_1008
timestamp 1679581782
transform 1 0 97344 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_1015
timestamp 1679581782
transform 1 0 98016 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_1022
timestamp 1679581782
transform 1 0 98688 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_0
timestamp 1679581782
transform 1 0 576 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_7
timestamp 1679581782
transform 1 0 1248 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_14
timestamp 1679581782
transform 1 0 1920 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_21
timestamp 1679581782
transform 1 0 2592 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_28
timestamp 1679581782
transform 1 0 3264 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_35
timestamp 1679581782
transform 1 0 3936 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_42
timestamp 1679581782
transform 1 0 4608 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_49
timestamp 1679581782
transform 1 0 5280 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_56
timestamp 1679581782
transform 1 0 5952 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_63
timestamp 1679581782
transform 1 0 6624 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_70
timestamp 1679581782
transform 1 0 7296 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_77
timestamp 1679581782
transform 1 0 7968 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_84
timestamp 1679581782
transform 1 0 8640 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_91
timestamp 1679581782
transform 1 0 9312 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_98
timestamp 1679581782
transform 1 0 9984 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_105
timestamp 1679581782
transform 1 0 10656 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_112
timestamp 1679581782
transform 1 0 11328 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_119
timestamp 1679581782
transform 1 0 12000 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_126
timestamp 1679581782
transform 1 0 12672 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_133
timestamp 1679581782
transform 1 0 13344 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_140
timestamp 1679581782
transform 1 0 14016 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_147
timestamp 1679581782
transform 1 0 14688 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_154
timestamp 1679581782
transform 1 0 15360 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_161
timestamp 1679581782
transform 1 0 16032 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_168
timestamp 1679581782
transform 1 0 16704 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_175
timestamp 1679581782
transform 1 0 17376 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_182
timestamp 1679581782
transform 1 0 18048 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_189
timestamp 1679581782
transform 1 0 18720 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_196
timestamp 1679581782
transform 1 0 19392 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_203
timestamp 1679581782
transform 1 0 20064 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_210
timestamp 1679581782
transform 1 0 20736 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_217
timestamp 1679581782
transform 1 0 21408 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_224
timestamp 1679581782
transform 1 0 22080 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_231
timestamp 1679581782
transform 1 0 22752 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_238
timestamp 1679581782
transform 1 0 23424 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_245
timestamp 1679581782
transform 1 0 24096 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_252
timestamp 1679581782
transform 1 0 24768 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_259
timestamp 1679581782
transform 1 0 25440 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_266
timestamp 1679581782
transform 1 0 26112 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_273
timestamp 1679581782
transform 1 0 26784 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_280
timestamp 1679581782
transform 1 0 27456 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_287
timestamp 1679581782
transform 1 0 28128 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_294
timestamp 1679581782
transform 1 0 28800 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_301
timestamp 1679581782
transform 1 0 29472 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_308
timestamp 1679581782
transform 1 0 30144 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_315
timestamp 1679581782
transform 1 0 30816 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_322
timestamp 1679581782
transform 1 0 31488 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_329
timestamp 1679581782
transform 1 0 32160 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_336
timestamp 1679581782
transform 1 0 32832 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_343
timestamp 1679581782
transform 1 0 33504 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_350
timestamp 1679581782
transform 1 0 34176 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_357
timestamp 1679581782
transform 1 0 34848 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_364
timestamp 1679581782
transform 1 0 35520 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_371
timestamp 1679581782
transform 1 0 36192 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_378
timestamp 1679581782
transform 1 0 36864 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_385
timestamp 1679581782
transform 1 0 37536 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_392
timestamp 1679581782
transform 1 0 38208 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_399
timestamp 1679581782
transform 1 0 38880 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_406
timestamp 1679581782
transform 1 0 39552 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_413
timestamp 1679581782
transform 1 0 40224 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_420
timestamp 1679581782
transform 1 0 40896 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_427
timestamp 1679581782
transform 1 0 41568 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_434
timestamp 1679581782
transform 1 0 42240 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_441
timestamp 1679581782
transform 1 0 42912 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_448
timestamp 1679581782
transform 1 0 43584 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_455
timestamp 1679581782
transform 1 0 44256 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_462
timestamp 1679581782
transform 1 0 44928 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_469
timestamp 1679581782
transform 1 0 45600 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_476
timestamp 1679581782
transform 1 0 46272 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_483
timestamp 1679581782
transform 1 0 46944 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_490
timestamp 1679581782
transform 1 0 47616 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_497
timestamp 1679581782
transform 1 0 48288 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_504
timestamp 1679581782
transform 1 0 48960 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_511
timestamp 1679581782
transform 1 0 49632 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_518
timestamp 1679581782
transform 1 0 50304 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_525
timestamp 1679581782
transform 1 0 50976 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_532
timestamp 1679581782
transform 1 0 51648 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_539
timestamp 1679581782
transform 1 0 52320 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_546
timestamp 1679581782
transform 1 0 52992 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_553
timestamp 1679581782
transform 1 0 53664 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_560
timestamp 1679581782
transform 1 0 54336 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_567
timestamp 1679581782
transform 1 0 55008 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_574
timestamp 1679581782
transform 1 0 55680 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_581
timestamp 1679581782
transform 1 0 56352 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_588
timestamp 1679581782
transform 1 0 57024 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_595
timestamp 1679581782
transform 1 0 57696 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_602
timestamp 1679581782
transform 1 0 58368 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_609
timestamp 1679581782
transform 1 0 59040 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_616
timestamp 1679581782
transform 1 0 59712 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_623
timestamp 1679581782
transform 1 0 60384 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_630
timestamp 1679581782
transform 1 0 61056 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_637
timestamp 1679581782
transform 1 0 61728 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_644
timestamp 1679581782
transform 1 0 62400 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_651
timestamp 1679581782
transform 1 0 63072 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_658
timestamp 1679581782
transform 1 0 63744 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_665
timestamp 1679581782
transform 1 0 64416 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_672
timestamp 1679581782
transform 1 0 65088 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_679
timestamp 1679581782
transform 1 0 65760 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_686
timestamp 1679581782
transform 1 0 66432 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_693
timestamp 1679581782
transform 1 0 67104 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_700
timestamp 1679581782
transform 1 0 67776 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_707
timestamp 1679581782
transform 1 0 68448 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_714
timestamp 1679581782
transform 1 0 69120 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_721
timestamp 1679581782
transform 1 0 69792 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_728
timestamp 1679581782
transform 1 0 70464 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_735
timestamp 1679581782
transform 1 0 71136 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_742
timestamp 1679581782
transform 1 0 71808 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_749
timestamp 1679581782
transform 1 0 72480 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_756
timestamp 1679581782
transform 1 0 73152 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_763
timestamp 1679581782
transform 1 0 73824 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_770
timestamp 1679581782
transform 1 0 74496 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_777
timestamp 1679581782
transform 1 0 75168 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_784
timestamp 1679581782
transform 1 0 75840 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_791
timestamp 1679581782
transform 1 0 76512 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_798
timestamp 1679581782
transform 1 0 77184 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_805
timestamp 1679581782
transform 1 0 77856 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_812
timestamp 1679581782
transform 1 0 78528 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_819
timestamp 1679581782
transform 1 0 79200 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_826
timestamp 1679581782
transform 1 0 79872 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_833
timestamp 1679581782
transform 1 0 80544 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_840
timestamp 1679581782
transform 1 0 81216 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_847
timestamp 1679581782
transform 1 0 81888 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_854
timestamp 1679581782
transform 1 0 82560 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_861
timestamp 1679581782
transform 1 0 83232 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_868
timestamp 1679581782
transform 1 0 83904 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_875
timestamp 1679581782
transform 1 0 84576 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_882
timestamp 1679581782
transform 1 0 85248 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_889
timestamp 1679581782
transform 1 0 85920 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_896
timestamp 1679581782
transform 1 0 86592 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_903
timestamp 1679581782
transform 1 0 87264 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_910
timestamp 1679581782
transform 1 0 87936 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_917
timestamp 1679581782
transform 1 0 88608 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_924
timestamp 1679581782
transform 1 0 89280 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_931
timestamp 1679581782
transform 1 0 89952 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_938
timestamp 1679581782
transform 1 0 90624 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_945
timestamp 1679581782
transform 1 0 91296 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_952
timestamp 1679581782
transform 1 0 91968 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_959
timestamp 1679581782
transform 1 0 92640 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_966
timestamp 1679581782
transform 1 0 93312 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_973
timestamp 1679581782
transform 1 0 93984 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_980
timestamp 1679581782
transform 1 0 94656 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_987
timestamp 1679581782
transform 1 0 95328 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_994
timestamp 1679581782
transform 1 0 96000 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_1001
timestamp 1679581782
transform 1 0 96672 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_1008
timestamp 1679581782
transform 1 0 97344 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_1015
timestamp 1679581782
transform 1 0 98016 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_1022
timestamp 1679581782
transform 1 0 98688 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_4
timestamp 1679581782
transform 1 0 960 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_11
timestamp 1679581782
transform 1 0 1632 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_18
timestamp 1679581782
transform 1 0 2304 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_25
timestamp 1679581782
transform 1 0 2976 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_32
timestamp 1679581782
transform 1 0 3648 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_39
timestamp 1679581782
transform 1 0 4320 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_46
timestamp 1679581782
transform 1 0 4992 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_53
timestamp 1679581782
transform 1 0 5664 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_60
timestamp 1679581782
transform 1 0 6336 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_67
timestamp 1679581782
transform 1 0 7008 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_74
timestamp 1679581782
transform 1 0 7680 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_81
timestamp 1679581782
transform 1 0 8352 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_88
timestamp 1679581782
transform 1 0 9024 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_95
timestamp 1679581782
transform 1 0 9696 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_102
timestamp 1679581782
transform 1 0 10368 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_109
timestamp 1679581782
transform 1 0 11040 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_116
timestamp 1679581782
transform 1 0 11712 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_123
timestamp 1679581782
transform 1 0 12384 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_130
timestamp 1679581782
transform 1 0 13056 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_137
timestamp 1679581782
transform 1 0 13728 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_144
timestamp 1679581782
transform 1 0 14400 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_151
timestamp 1679581782
transform 1 0 15072 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_158
timestamp 1679581782
transform 1 0 15744 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_165
timestamp 1679581782
transform 1 0 16416 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_172
timestamp 1679581782
transform 1 0 17088 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_179
timestamp 1679581782
transform 1 0 17760 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_186
timestamp 1679581782
transform 1 0 18432 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_193
timestamp 1679581782
transform 1 0 19104 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_200
timestamp 1679581782
transform 1 0 19776 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_207
timestamp 1679581782
transform 1 0 20448 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_214
timestamp 1679581782
transform 1 0 21120 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_221
timestamp 1679581782
transform 1 0 21792 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_228
timestamp 1679581782
transform 1 0 22464 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_235
timestamp 1679581782
transform 1 0 23136 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_242
timestamp 1679581782
transform 1 0 23808 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_249
timestamp 1679581782
transform 1 0 24480 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_256
timestamp 1679581782
transform 1 0 25152 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_263
timestamp 1679581782
transform 1 0 25824 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_270
timestamp 1679581782
transform 1 0 26496 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_277
timestamp 1679581782
transform 1 0 27168 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_284
timestamp 1679581782
transform 1 0 27840 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_291
timestamp 1679581782
transform 1 0 28512 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_298
timestamp 1679581782
transform 1 0 29184 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_305
timestamp 1679581782
transform 1 0 29856 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_312
timestamp 1679581782
transform 1 0 30528 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_319
timestamp 1679581782
transform 1 0 31200 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_326
timestamp 1679581782
transform 1 0 31872 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_333
timestamp 1679581782
transform 1 0 32544 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_340
timestamp 1679581782
transform 1 0 33216 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_347
timestamp 1679581782
transform 1 0 33888 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_354
timestamp 1679581782
transform 1 0 34560 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_361
timestamp 1679581782
transform 1 0 35232 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_368
timestamp 1679581782
transform 1 0 35904 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_375
timestamp 1679581782
transform 1 0 36576 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_382
timestamp 1679581782
transform 1 0 37248 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_389
timestamp 1679581782
transform 1 0 37920 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_396
timestamp 1679581782
transform 1 0 38592 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_403
timestamp 1679581782
transform 1 0 39264 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_410
timestamp 1679581782
transform 1 0 39936 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_417
timestamp 1679581782
transform 1 0 40608 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_424
timestamp 1679581782
transform 1 0 41280 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_431
timestamp 1679581782
transform 1 0 41952 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_438
timestamp 1679581782
transform 1 0 42624 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_445
timestamp 1679581782
transform 1 0 43296 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_452
timestamp 1679581782
transform 1 0 43968 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_459
timestamp 1679581782
transform 1 0 44640 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_466
timestamp 1679581782
transform 1 0 45312 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_473
timestamp 1679581782
transform 1 0 45984 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_480
timestamp 1679581782
transform 1 0 46656 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_487
timestamp 1679581782
transform 1 0 47328 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_494
timestamp 1679581782
transform 1 0 48000 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_501
timestamp 1679581782
transform 1 0 48672 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_508
timestamp 1679581782
transform 1 0 49344 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_515
timestamp 1679581782
transform 1 0 50016 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_522
timestamp 1679581782
transform 1 0 50688 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_529
timestamp 1679581782
transform 1 0 51360 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_536
timestamp 1679581782
transform 1 0 52032 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_543
timestamp 1679581782
transform 1 0 52704 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_550
timestamp 1679581782
transform 1 0 53376 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_557
timestamp 1679581782
transform 1 0 54048 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_564
timestamp 1679581782
transform 1 0 54720 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_571
timestamp 1679581782
transform 1 0 55392 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_578
timestamp 1679581782
transform 1 0 56064 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_585
timestamp 1679581782
transform 1 0 56736 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_592
timestamp 1679581782
transform 1 0 57408 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_599
timestamp 1679581782
transform 1 0 58080 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_606
timestamp 1679581782
transform 1 0 58752 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_613
timestamp 1679581782
transform 1 0 59424 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_620
timestamp 1679581782
transform 1 0 60096 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_627
timestamp 1679581782
transform 1 0 60768 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_634
timestamp 1679581782
transform 1 0 61440 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_641
timestamp 1679581782
transform 1 0 62112 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_648
timestamp 1679581782
transform 1 0 62784 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_655
timestamp 1679581782
transform 1 0 63456 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_662
timestamp 1679581782
transform 1 0 64128 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_669
timestamp 1679581782
transform 1 0 64800 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_676
timestamp 1679581782
transform 1 0 65472 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_683
timestamp 1679581782
transform 1 0 66144 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_690
timestamp 1679581782
transform 1 0 66816 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_697
timestamp 1679581782
transform 1 0 67488 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_704
timestamp 1679581782
transform 1 0 68160 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_711
timestamp 1679581782
transform 1 0 68832 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_718
timestamp 1679581782
transform 1 0 69504 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_725
timestamp 1679581782
transform 1 0 70176 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_732
timestamp 1679581782
transform 1 0 70848 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_739
timestamp 1679581782
transform 1 0 71520 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_746
timestamp 1679581782
transform 1 0 72192 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_753
timestamp 1679581782
transform 1 0 72864 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_760
timestamp 1679581782
transform 1 0 73536 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_767
timestamp 1679581782
transform 1 0 74208 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_774
timestamp 1679581782
transform 1 0 74880 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_781
timestamp 1679581782
transform 1 0 75552 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_788
timestamp 1679581782
transform 1 0 76224 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_795
timestamp 1679581782
transform 1 0 76896 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_802
timestamp 1679581782
transform 1 0 77568 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_809
timestamp 1679581782
transform 1 0 78240 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_816
timestamp 1679581782
transform 1 0 78912 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_823
timestamp 1679581782
transform 1 0 79584 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_830
timestamp 1679581782
transform 1 0 80256 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_837
timestamp 1679581782
transform 1 0 80928 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_844
timestamp 1679581782
transform 1 0 81600 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_851
timestamp 1679581782
transform 1 0 82272 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_858
timestamp 1679581782
transform 1 0 82944 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_865
timestamp 1679581782
transform 1 0 83616 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_872
timestamp 1679581782
transform 1 0 84288 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_879
timestamp 1679581782
transform 1 0 84960 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_886
timestamp 1679581782
transform 1 0 85632 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_893
timestamp 1679581782
transform 1 0 86304 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_900
timestamp 1679581782
transform 1 0 86976 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_907
timestamp 1679581782
transform 1 0 87648 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_914
timestamp 1679581782
transform 1 0 88320 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_921
timestamp 1679581782
transform 1 0 88992 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_928
timestamp 1679581782
transform 1 0 89664 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_935
timestamp 1679581782
transform 1 0 90336 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_942
timestamp 1679581782
transform 1 0 91008 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_949
timestamp 1679581782
transform 1 0 91680 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_956
timestamp 1679581782
transform 1 0 92352 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_963
timestamp 1679581782
transform 1 0 93024 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_970
timestamp 1679581782
transform 1 0 93696 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_977
timestamp 1679581782
transform 1 0 94368 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_984
timestamp 1679581782
transform 1 0 95040 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_991
timestamp 1679581782
transform 1 0 95712 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_998
timestamp 1679581782
transform 1 0 96384 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_1005
timestamp 1679581782
transform 1 0 97056 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_1012
timestamp 1679581782
transform 1 0 97728 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_1019
timestamp 1679581782
transform 1 0 98400 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_15_1026
timestamp 1677580104
transform 1 0 99072 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_1028
timestamp 1677579658
transform 1 0 99264 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_0
timestamp 1679581782
transform 1 0 576 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_7
timestamp 1679581782
transform 1 0 1248 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_14
timestamp 1679581782
transform 1 0 1920 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_21
timestamp 1679581782
transform 1 0 2592 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_28
timestamp 1679581782
transform 1 0 3264 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_35
timestamp 1679581782
transform 1 0 3936 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_42
timestamp 1679581782
transform 1 0 4608 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_49
timestamp 1679581782
transform 1 0 5280 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_56
timestamp 1679581782
transform 1 0 5952 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_63
timestamp 1679581782
transform 1 0 6624 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_70
timestamp 1679581782
transform 1 0 7296 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_77
timestamp 1679581782
transform 1 0 7968 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_84
timestamp 1679581782
transform 1 0 8640 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_91
timestamp 1679581782
transform 1 0 9312 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_98
timestamp 1679581782
transform 1 0 9984 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_105
timestamp 1679581782
transform 1 0 10656 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_112
timestamp 1679581782
transform 1 0 11328 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_119
timestamp 1679581782
transform 1 0 12000 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_126
timestamp 1679581782
transform 1 0 12672 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_133
timestamp 1679581782
transform 1 0 13344 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_140
timestamp 1679581782
transform 1 0 14016 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_147
timestamp 1679581782
transform 1 0 14688 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_154
timestamp 1679581782
transform 1 0 15360 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_161
timestamp 1679581782
transform 1 0 16032 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_168
timestamp 1679581782
transform 1 0 16704 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_175
timestamp 1679581782
transform 1 0 17376 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_182
timestamp 1679581782
transform 1 0 18048 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_189
timestamp 1679581782
transform 1 0 18720 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_196
timestamp 1679581782
transform 1 0 19392 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_203
timestamp 1679581782
transform 1 0 20064 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_210
timestamp 1679581782
transform 1 0 20736 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_217
timestamp 1679581782
transform 1 0 21408 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_224
timestamp 1679581782
transform 1 0 22080 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_231
timestamp 1679581782
transform 1 0 22752 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_238
timestamp 1679581782
transform 1 0 23424 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_245
timestamp 1679581782
transform 1 0 24096 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_252
timestamp 1679581782
transform 1 0 24768 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_259
timestamp 1679581782
transform 1 0 25440 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_266
timestamp 1679581782
transform 1 0 26112 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_273
timestamp 1679581782
transform 1 0 26784 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_280
timestamp 1679581782
transform 1 0 27456 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_287
timestamp 1679581782
transform 1 0 28128 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_294
timestamp 1679581782
transform 1 0 28800 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_301
timestamp 1679581782
transform 1 0 29472 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_308
timestamp 1679581782
transform 1 0 30144 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_315
timestamp 1679581782
transform 1 0 30816 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_322
timestamp 1679581782
transform 1 0 31488 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_329
timestamp 1679581782
transform 1 0 32160 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_336
timestamp 1679581782
transform 1 0 32832 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_343
timestamp 1679581782
transform 1 0 33504 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_350
timestamp 1679581782
transform 1 0 34176 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_357
timestamp 1679581782
transform 1 0 34848 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_364
timestamp 1679581782
transform 1 0 35520 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_371
timestamp 1679581782
transform 1 0 36192 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_378
timestamp 1679581782
transform 1 0 36864 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_385
timestamp 1679581782
transform 1 0 37536 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_392
timestamp 1679581782
transform 1 0 38208 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_399
timestamp 1679581782
transform 1 0 38880 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_406
timestamp 1679581782
transform 1 0 39552 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_413
timestamp 1679581782
transform 1 0 40224 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_420
timestamp 1679581782
transform 1 0 40896 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_427
timestamp 1679581782
transform 1 0 41568 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_434
timestamp 1679581782
transform 1 0 42240 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_441
timestamp 1679581782
transform 1 0 42912 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_448
timestamp 1679581782
transform 1 0 43584 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_455
timestamp 1679581782
transform 1 0 44256 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_462
timestamp 1679581782
transform 1 0 44928 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_469
timestamp 1679581782
transform 1 0 45600 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_476
timestamp 1679581782
transform 1 0 46272 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_483
timestamp 1679581782
transform 1 0 46944 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_490
timestamp 1679581782
transform 1 0 47616 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_497
timestamp 1679581782
transform 1 0 48288 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_504
timestamp 1679581782
transform 1 0 48960 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_511
timestamp 1679581782
transform 1 0 49632 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_518
timestamp 1679581782
transform 1 0 50304 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_525
timestamp 1679581782
transform 1 0 50976 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_532
timestamp 1679581782
transform 1 0 51648 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_539
timestamp 1679581782
transform 1 0 52320 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_546
timestamp 1679581782
transform 1 0 52992 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_553
timestamp 1679581782
transform 1 0 53664 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_560
timestamp 1679581782
transform 1 0 54336 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_567
timestamp 1679581782
transform 1 0 55008 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_574
timestamp 1679581782
transform 1 0 55680 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_581
timestamp 1679581782
transform 1 0 56352 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_588
timestamp 1679581782
transform 1 0 57024 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_595
timestamp 1679581782
transform 1 0 57696 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_602
timestamp 1679581782
transform 1 0 58368 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_609
timestamp 1679581782
transform 1 0 59040 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_616
timestamp 1679581782
transform 1 0 59712 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_623
timestamp 1679581782
transform 1 0 60384 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_630
timestamp 1679581782
transform 1 0 61056 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_637
timestamp 1679581782
transform 1 0 61728 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_644
timestamp 1679581782
transform 1 0 62400 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_651
timestamp 1679581782
transform 1 0 63072 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_658
timestamp 1679581782
transform 1 0 63744 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_665
timestamp 1679581782
transform 1 0 64416 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_672
timestamp 1679581782
transform 1 0 65088 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_679
timestamp 1679581782
transform 1 0 65760 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_686
timestamp 1679581782
transform 1 0 66432 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_693
timestamp 1679581782
transform 1 0 67104 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_700
timestamp 1679581782
transform 1 0 67776 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_707
timestamp 1679581782
transform 1 0 68448 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_714
timestamp 1679581782
transform 1 0 69120 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_721
timestamp 1679581782
transform 1 0 69792 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_728
timestamp 1679581782
transform 1 0 70464 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_735
timestamp 1679581782
transform 1 0 71136 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_742
timestamp 1679581782
transform 1 0 71808 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_749
timestamp 1679581782
transform 1 0 72480 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_756
timestamp 1679581782
transform 1 0 73152 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_763
timestamp 1679581782
transform 1 0 73824 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_770
timestamp 1679581782
transform 1 0 74496 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_777
timestamp 1679581782
transform 1 0 75168 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_784
timestamp 1679581782
transform 1 0 75840 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_791
timestamp 1679581782
transform 1 0 76512 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_798
timestamp 1679581782
transform 1 0 77184 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_805
timestamp 1679581782
transform 1 0 77856 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_812
timestamp 1679581782
transform 1 0 78528 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_819
timestamp 1679581782
transform 1 0 79200 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_826
timestamp 1679581782
transform 1 0 79872 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_833
timestamp 1679581782
transform 1 0 80544 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_840
timestamp 1679581782
transform 1 0 81216 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_847
timestamp 1679581782
transform 1 0 81888 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_854
timestamp 1679581782
transform 1 0 82560 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_861
timestamp 1679581782
transform 1 0 83232 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_868
timestamp 1679581782
transform 1 0 83904 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_875
timestamp 1679581782
transform 1 0 84576 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_882
timestamp 1679581782
transform 1 0 85248 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_889
timestamp 1679581782
transform 1 0 85920 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_896
timestamp 1679581782
transform 1 0 86592 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_903
timestamp 1679581782
transform 1 0 87264 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_910
timestamp 1679581782
transform 1 0 87936 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_917
timestamp 1679581782
transform 1 0 88608 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_924
timestamp 1679581782
transform 1 0 89280 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_931
timestamp 1679581782
transform 1 0 89952 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_938
timestamp 1679581782
transform 1 0 90624 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_945
timestamp 1679581782
transform 1 0 91296 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_952
timestamp 1679581782
transform 1 0 91968 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_959
timestamp 1679581782
transform 1 0 92640 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_966
timestamp 1679581782
transform 1 0 93312 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_973
timestamp 1679581782
transform 1 0 93984 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_980
timestamp 1679581782
transform 1 0 94656 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_987
timestamp 1679581782
transform 1 0 95328 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_994
timestamp 1679581782
transform 1 0 96000 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_1001
timestamp 1679581782
transform 1 0 96672 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_1008
timestamp 1679581782
transform 1 0 97344 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_1015
timestamp 1679581782
transform 1 0 98016 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_1022
timestamp 1679581782
transform 1 0 98688 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_4
timestamp 1679581782
transform 1 0 960 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_11
timestamp 1679581782
transform 1 0 1632 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_18
timestamp 1679581782
transform 1 0 2304 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_25
timestamp 1679581782
transform 1 0 2976 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_32
timestamp 1679581782
transform 1 0 3648 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_39
timestamp 1679581782
transform 1 0 4320 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_46
timestamp 1679581782
transform 1 0 4992 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_53
timestamp 1679581782
transform 1 0 5664 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_60
timestamp 1679581782
transform 1 0 6336 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_67
timestamp 1679581782
transform 1 0 7008 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_74
timestamp 1679581782
transform 1 0 7680 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_81
timestamp 1679581782
transform 1 0 8352 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_88
timestamp 1679581782
transform 1 0 9024 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_95
timestamp 1679581782
transform 1 0 9696 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_102
timestamp 1679581782
transform 1 0 10368 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_109
timestamp 1679581782
transform 1 0 11040 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_116
timestamp 1679581782
transform 1 0 11712 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_123
timestamp 1679581782
transform 1 0 12384 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_130
timestamp 1679581782
transform 1 0 13056 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_137
timestamp 1679581782
transform 1 0 13728 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_144
timestamp 1679581782
transform 1 0 14400 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_151
timestamp 1679581782
transform 1 0 15072 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_158
timestamp 1679581782
transform 1 0 15744 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_165
timestamp 1679581782
transform 1 0 16416 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_172
timestamp 1679581782
transform 1 0 17088 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_179
timestamp 1679581782
transform 1 0 17760 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_186
timestamp 1679581782
transform 1 0 18432 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_193
timestamp 1679581782
transform 1 0 19104 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_200
timestamp 1679581782
transform 1 0 19776 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_207
timestamp 1679581782
transform 1 0 20448 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_214
timestamp 1679581782
transform 1 0 21120 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_221
timestamp 1679581782
transform 1 0 21792 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_228
timestamp 1679581782
transform 1 0 22464 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_235
timestamp 1679581782
transform 1 0 23136 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_242
timestamp 1679581782
transform 1 0 23808 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_249
timestamp 1679581782
transform 1 0 24480 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_256
timestamp 1679581782
transform 1 0 25152 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_263
timestamp 1679581782
transform 1 0 25824 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_270
timestamp 1679581782
transform 1 0 26496 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_277
timestamp 1679581782
transform 1 0 27168 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_284
timestamp 1679581782
transform 1 0 27840 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_291
timestamp 1679581782
transform 1 0 28512 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_298
timestamp 1679581782
transform 1 0 29184 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_305
timestamp 1679581782
transform 1 0 29856 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_312
timestamp 1679581782
transform 1 0 30528 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_319
timestamp 1679581782
transform 1 0 31200 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_326
timestamp 1679581782
transform 1 0 31872 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_333
timestamp 1679581782
transform 1 0 32544 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_340
timestamp 1679581782
transform 1 0 33216 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_347
timestamp 1679581782
transform 1 0 33888 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_354
timestamp 1679581782
transform 1 0 34560 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_361
timestamp 1679581782
transform 1 0 35232 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_368
timestamp 1679581782
transform 1 0 35904 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_375
timestamp 1679581782
transform 1 0 36576 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_382
timestamp 1679581782
transform 1 0 37248 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_389
timestamp 1679581782
transform 1 0 37920 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_396
timestamp 1679581782
transform 1 0 38592 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_403
timestamp 1679581782
transform 1 0 39264 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_410
timestamp 1679581782
transform 1 0 39936 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_417
timestamp 1679581782
transform 1 0 40608 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_424
timestamp 1679581782
transform 1 0 41280 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_431
timestamp 1679581782
transform 1 0 41952 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_438
timestamp 1679581782
transform 1 0 42624 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_445
timestamp 1679581782
transform 1 0 43296 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_452
timestamp 1679581782
transform 1 0 43968 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_459
timestamp 1679581782
transform 1 0 44640 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_466
timestamp 1679581782
transform 1 0 45312 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_473
timestamp 1679581782
transform 1 0 45984 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_480
timestamp 1679581782
transform 1 0 46656 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_487
timestamp 1679581782
transform 1 0 47328 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_494
timestamp 1679581782
transform 1 0 48000 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_501
timestamp 1679581782
transform 1 0 48672 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_508
timestamp 1679581782
transform 1 0 49344 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_515
timestamp 1679581782
transform 1 0 50016 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_522
timestamp 1679581782
transform 1 0 50688 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_529
timestamp 1679581782
transform 1 0 51360 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_536
timestamp 1679581782
transform 1 0 52032 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_543
timestamp 1679581782
transform 1 0 52704 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_550
timestamp 1679581782
transform 1 0 53376 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_557
timestamp 1679581782
transform 1 0 54048 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_564
timestamp 1679581782
transform 1 0 54720 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_571
timestamp 1679581782
transform 1 0 55392 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_578
timestamp 1679581782
transform 1 0 56064 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_585
timestamp 1679581782
transform 1 0 56736 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_592
timestamp 1679581782
transform 1 0 57408 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_599
timestamp 1679581782
transform 1 0 58080 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_606
timestamp 1679581782
transform 1 0 58752 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_613
timestamp 1679581782
transform 1 0 59424 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_620
timestamp 1679581782
transform 1 0 60096 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_627
timestamp 1679581782
transform 1 0 60768 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_634
timestamp 1679581782
transform 1 0 61440 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_641
timestamp 1679581782
transform 1 0 62112 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_648
timestamp 1679581782
transform 1 0 62784 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_655
timestamp 1679581782
transform 1 0 63456 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_662
timestamp 1679581782
transform 1 0 64128 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_669
timestamp 1679581782
transform 1 0 64800 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_676
timestamp 1679581782
transform 1 0 65472 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_683
timestamp 1679581782
transform 1 0 66144 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_690
timestamp 1679581782
transform 1 0 66816 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_697
timestamp 1679581782
transform 1 0 67488 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_704
timestamp 1679581782
transform 1 0 68160 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_711
timestamp 1679581782
transform 1 0 68832 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_718
timestamp 1679581782
transform 1 0 69504 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_725
timestamp 1679581782
transform 1 0 70176 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_732
timestamp 1679581782
transform 1 0 70848 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_739
timestamp 1679581782
transform 1 0 71520 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_746
timestamp 1679581782
transform 1 0 72192 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_753
timestamp 1679581782
transform 1 0 72864 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_760
timestamp 1679581782
transform 1 0 73536 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_767
timestamp 1679581782
transform 1 0 74208 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_774
timestamp 1679581782
transform 1 0 74880 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_781
timestamp 1679581782
transform 1 0 75552 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_788
timestamp 1679581782
transform 1 0 76224 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_795
timestamp 1679581782
transform 1 0 76896 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_802
timestamp 1679581782
transform 1 0 77568 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_809
timestamp 1679581782
transform 1 0 78240 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_816
timestamp 1679581782
transform 1 0 78912 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_823
timestamp 1679581782
transform 1 0 79584 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_830
timestamp 1679581782
transform 1 0 80256 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_837
timestamp 1679581782
transform 1 0 80928 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_844
timestamp 1679581782
transform 1 0 81600 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_851
timestamp 1679581782
transform 1 0 82272 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_858
timestamp 1679581782
transform 1 0 82944 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_865
timestamp 1679581782
transform 1 0 83616 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_872
timestamp 1679581782
transform 1 0 84288 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_879
timestamp 1679581782
transform 1 0 84960 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_886
timestamp 1679581782
transform 1 0 85632 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_893
timestamp 1679581782
transform 1 0 86304 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_900
timestamp 1679581782
transform 1 0 86976 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_907
timestamp 1679581782
transform 1 0 87648 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_914
timestamp 1679581782
transform 1 0 88320 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_921
timestamp 1679581782
transform 1 0 88992 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_928
timestamp 1679581782
transform 1 0 89664 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_935
timestamp 1679581782
transform 1 0 90336 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_942
timestamp 1679581782
transform 1 0 91008 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_949
timestamp 1679581782
transform 1 0 91680 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_956
timestamp 1679581782
transform 1 0 92352 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_963
timestamp 1679581782
transform 1 0 93024 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_970
timestamp 1679581782
transform 1 0 93696 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_977
timestamp 1679581782
transform 1 0 94368 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_984
timestamp 1679581782
transform 1 0 95040 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_991
timestamp 1679581782
transform 1 0 95712 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_998
timestamp 1679581782
transform 1 0 96384 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_1005
timestamp 1679581782
transform 1 0 97056 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_1012
timestamp 1679581782
transform 1 0 97728 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_1019
timestamp 1679581782
transform 1 0 98400 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_1026
timestamp 1677580104
transform 1 0 99072 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_1028
timestamp 1677579658
transform 1 0 99264 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_0
timestamp 1679581782
transform 1 0 576 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_7
timestamp 1679581782
transform 1 0 1248 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_14
timestamp 1679581782
transform 1 0 1920 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_21
timestamp 1679581782
transform 1 0 2592 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_28
timestamp 1679581782
transform 1 0 3264 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_35
timestamp 1679581782
transform 1 0 3936 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_42
timestamp 1679581782
transform 1 0 4608 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_49
timestamp 1679581782
transform 1 0 5280 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_56
timestamp 1679581782
transform 1 0 5952 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_63
timestamp 1679581782
transform 1 0 6624 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_70
timestamp 1679581782
transform 1 0 7296 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_77
timestamp 1679581782
transform 1 0 7968 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_84
timestamp 1679581782
transform 1 0 8640 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_91
timestamp 1679581782
transform 1 0 9312 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_98
timestamp 1679581782
transform 1 0 9984 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_105
timestamp 1679581782
transform 1 0 10656 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_112
timestamp 1679581782
transform 1 0 11328 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_119
timestamp 1679581782
transform 1 0 12000 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_126
timestamp 1679581782
transform 1 0 12672 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_133
timestamp 1679581782
transform 1 0 13344 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_140
timestamp 1679581782
transform 1 0 14016 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_147
timestamp 1679581782
transform 1 0 14688 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_154
timestamp 1679581782
transform 1 0 15360 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_161
timestamp 1679581782
transform 1 0 16032 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_168
timestamp 1679581782
transform 1 0 16704 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_175
timestamp 1679581782
transform 1 0 17376 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_182
timestamp 1679581782
transform 1 0 18048 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_189
timestamp 1679581782
transform 1 0 18720 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_196
timestamp 1679581782
transform 1 0 19392 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_203
timestamp 1679581782
transform 1 0 20064 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_210
timestamp 1679581782
transform 1 0 20736 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_217
timestamp 1679581782
transform 1 0 21408 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_224
timestamp 1679581782
transform 1 0 22080 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_231
timestamp 1679581782
transform 1 0 22752 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_238
timestamp 1679581782
transform 1 0 23424 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_245
timestamp 1679581782
transform 1 0 24096 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_252
timestamp 1679581782
transform 1 0 24768 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_259
timestamp 1679581782
transform 1 0 25440 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_266
timestamp 1679581782
transform 1 0 26112 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_273
timestamp 1679581782
transform 1 0 26784 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_280
timestamp 1679581782
transform 1 0 27456 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_287
timestamp 1679581782
transform 1 0 28128 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_294
timestamp 1679581782
transform 1 0 28800 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_301
timestamp 1679581782
transform 1 0 29472 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_308
timestamp 1679581782
transform 1 0 30144 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_315
timestamp 1679581782
transform 1 0 30816 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_322
timestamp 1679581782
transform 1 0 31488 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_329
timestamp 1679581782
transform 1 0 32160 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_336
timestamp 1679581782
transform 1 0 32832 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_343
timestamp 1679581782
transform 1 0 33504 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_350
timestamp 1679581782
transform 1 0 34176 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_357
timestamp 1679581782
transform 1 0 34848 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_364
timestamp 1679581782
transform 1 0 35520 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_371
timestamp 1679581782
transform 1 0 36192 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_378
timestamp 1679581782
transform 1 0 36864 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_385
timestamp 1679581782
transform 1 0 37536 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_392
timestamp 1679581782
transform 1 0 38208 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_399
timestamp 1679581782
transform 1 0 38880 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_406
timestamp 1679581782
transform 1 0 39552 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_413
timestamp 1679581782
transform 1 0 40224 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_420
timestamp 1679581782
transform 1 0 40896 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_427
timestamp 1679581782
transform 1 0 41568 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_434
timestamp 1679581782
transform 1 0 42240 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_441
timestamp 1679581782
transform 1 0 42912 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_448
timestamp 1679581782
transform 1 0 43584 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_455
timestamp 1679581782
transform 1 0 44256 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_462
timestamp 1679581782
transform 1 0 44928 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_469
timestamp 1679581782
transform 1 0 45600 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_476
timestamp 1679581782
transform 1 0 46272 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_483
timestamp 1679581782
transform 1 0 46944 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_490
timestamp 1679581782
transform 1 0 47616 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_497
timestamp 1679581782
transform 1 0 48288 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_504
timestamp 1679581782
transform 1 0 48960 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_511
timestamp 1679581782
transform 1 0 49632 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_518
timestamp 1679581782
transform 1 0 50304 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_525
timestamp 1679581782
transform 1 0 50976 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_532
timestamp 1679581782
transform 1 0 51648 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_539
timestamp 1679581782
transform 1 0 52320 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_546
timestamp 1679581782
transform 1 0 52992 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_553
timestamp 1679581782
transform 1 0 53664 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_560
timestamp 1679581782
transform 1 0 54336 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_567
timestamp 1679581782
transform 1 0 55008 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_574
timestamp 1679581782
transform 1 0 55680 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_581
timestamp 1679581782
transform 1 0 56352 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_588
timestamp 1679581782
transform 1 0 57024 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_595
timestamp 1679581782
transform 1 0 57696 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_602
timestamp 1679581782
transform 1 0 58368 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_609
timestamp 1679581782
transform 1 0 59040 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_616
timestamp 1679581782
transform 1 0 59712 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_623
timestamp 1679581782
transform 1 0 60384 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_630
timestamp 1679581782
transform 1 0 61056 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_637
timestamp 1679581782
transform 1 0 61728 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_644
timestamp 1679581782
transform 1 0 62400 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_651
timestamp 1679581782
transform 1 0 63072 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_658
timestamp 1679581782
transform 1 0 63744 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_665
timestamp 1679581782
transform 1 0 64416 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_672
timestamp 1679581782
transform 1 0 65088 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_679
timestamp 1679581782
transform 1 0 65760 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_686
timestamp 1679581782
transform 1 0 66432 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_693
timestamp 1679581782
transform 1 0 67104 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_700
timestamp 1679581782
transform 1 0 67776 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_707
timestamp 1679581782
transform 1 0 68448 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_714
timestamp 1679581782
transform 1 0 69120 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_721
timestamp 1679581782
transform 1 0 69792 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_728
timestamp 1679581782
transform 1 0 70464 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_735
timestamp 1679581782
transform 1 0 71136 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_742
timestamp 1679581782
transform 1 0 71808 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_749
timestamp 1679581782
transform 1 0 72480 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_756
timestamp 1679581782
transform 1 0 73152 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_763
timestamp 1679581782
transform 1 0 73824 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_770
timestamp 1679581782
transform 1 0 74496 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_777
timestamp 1679581782
transform 1 0 75168 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_784
timestamp 1679581782
transform 1 0 75840 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_791
timestamp 1679581782
transform 1 0 76512 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_798
timestamp 1679581782
transform 1 0 77184 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_805
timestamp 1679581782
transform 1 0 77856 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_812
timestamp 1679581782
transform 1 0 78528 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_819
timestamp 1679581782
transform 1 0 79200 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_826
timestamp 1679581782
transform 1 0 79872 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_833
timestamp 1679581782
transform 1 0 80544 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_840
timestamp 1679581782
transform 1 0 81216 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_847
timestamp 1679581782
transform 1 0 81888 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_854
timestamp 1679581782
transform 1 0 82560 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_861
timestamp 1679581782
transform 1 0 83232 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_868
timestamp 1679581782
transform 1 0 83904 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_875
timestamp 1679581782
transform 1 0 84576 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_882
timestamp 1679581782
transform 1 0 85248 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_889
timestamp 1679581782
transform 1 0 85920 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_896
timestamp 1679581782
transform 1 0 86592 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_903
timestamp 1679581782
transform 1 0 87264 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_910
timestamp 1679581782
transform 1 0 87936 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_917
timestamp 1679581782
transform 1 0 88608 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_924
timestamp 1679581782
transform 1 0 89280 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_931
timestamp 1679581782
transform 1 0 89952 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_938
timestamp 1679581782
transform 1 0 90624 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_945
timestamp 1679581782
transform 1 0 91296 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_952
timestamp 1679581782
transform 1 0 91968 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_959
timestamp 1679581782
transform 1 0 92640 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_966
timestamp 1679581782
transform 1 0 93312 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_973
timestamp 1679581782
transform 1 0 93984 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_980
timestamp 1679581782
transform 1 0 94656 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_987
timestamp 1679581782
transform 1 0 95328 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_994
timestamp 1679581782
transform 1 0 96000 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_1001
timestamp 1679581782
transform 1 0 96672 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_1008
timestamp 1679581782
transform 1 0 97344 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_1015
timestamp 1679581782
transform 1 0 98016 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_1022
timestamp 1679581782
transform 1 0 98688 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_0
timestamp 1679581782
transform 1 0 576 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_7
timestamp 1679581782
transform 1 0 1248 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_14
timestamp 1679581782
transform 1 0 1920 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_21
timestamp 1679581782
transform 1 0 2592 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_28
timestamp 1679581782
transform 1 0 3264 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_35
timestamp 1679581782
transform 1 0 3936 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_42
timestamp 1679581782
transform 1 0 4608 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_49
timestamp 1679581782
transform 1 0 5280 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_56
timestamp 1679581782
transform 1 0 5952 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_63
timestamp 1679581782
transform 1 0 6624 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_70
timestamp 1679581782
transform 1 0 7296 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_77
timestamp 1679581782
transform 1 0 7968 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_84
timestamp 1679581782
transform 1 0 8640 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_91
timestamp 1679581782
transform 1 0 9312 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_98
timestamp 1679581782
transform 1 0 9984 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_105
timestamp 1679581782
transform 1 0 10656 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_112
timestamp 1679581782
transform 1 0 11328 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_119
timestamp 1679581782
transform 1 0 12000 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_126
timestamp 1679581782
transform 1 0 12672 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_133
timestamp 1679581782
transform 1 0 13344 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_140
timestamp 1679581782
transform 1 0 14016 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_147
timestamp 1679581782
transform 1 0 14688 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_154
timestamp 1679581782
transform 1 0 15360 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_161
timestamp 1679581782
transform 1 0 16032 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_168
timestamp 1679581782
transform 1 0 16704 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_175
timestamp 1679581782
transform 1 0 17376 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_182
timestamp 1679581782
transform 1 0 18048 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_189
timestamp 1679581782
transform 1 0 18720 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_196
timestamp 1679581782
transform 1 0 19392 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_203
timestamp 1679581782
transform 1 0 20064 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_210
timestamp 1679581782
transform 1 0 20736 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_217
timestamp 1679581782
transform 1 0 21408 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_224
timestamp 1679581782
transform 1 0 22080 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_231
timestamp 1679581782
transform 1 0 22752 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_238
timestamp 1679581782
transform 1 0 23424 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_245
timestamp 1679581782
transform 1 0 24096 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_252
timestamp 1679581782
transform 1 0 24768 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_259
timestamp 1679581782
transform 1 0 25440 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_266
timestamp 1679581782
transform 1 0 26112 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_273
timestamp 1679581782
transform 1 0 26784 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_280
timestamp 1679581782
transform 1 0 27456 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_287
timestamp 1679581782
transform 1 0 28128 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_294
timestamp 1679581782
transform 1 0 28800 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_301
timestamp 1679581782
transform 1 0 29472 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_308
timestamp 1679581782
transform 1 0 30144 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_315
timestamp 1679581782
transform 1 0 30816 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_322
timestamp 1679581782
transform 1 0 31488 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_329
timestamp 1679581782
transform 1 0 32160 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_336
timestamp 1679581782
transform 1 0 32832 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_343
timestamp 1679581782
transform 1 0 33504 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_350
timestamp 1679581782
transform 1 0 34176 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_357
timestamp 1679581782
transform 1 0 34848 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_364
timestamp 1679581782
transform 1 0 35520 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_371
timestamp 1679581782
transform 1 0 36192 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_378
timestamp 1679581782
transform 1 0 36864 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_385
timestamp 1679581782
transform 1 0 37536 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_392
timestamp 1679581782
transform 1 0 38208 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_399
timestamp 1679581782
transform 1 0 38880 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_406
timestamp 1679581782
transform 1 0 39552 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_413
timestamp 1679581782
transform 1 0 40224 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_420
timestamp 1679581782
transform 1 0 40896 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_427
timestamp 1679581782
transform 1 0 41568 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_434
timestamp 1679581782
transform 1 0 42240 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_441
timestamp 1679581782
transform 1 0 42912 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_448
timestamp 1679581782
transform 1 0 43584 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_455
timestamp 1679581782
transform 1 0 44256 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_462
timestamp 1679581782
transform 1 0 44928 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_469
timestamp 1679581782
transform 1 0 45600 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_476
timestamp 1679581782
transform 1 0 46272 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_483
timestamp 1679581782
transform 1 0 46944 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_490
timestamp 1679581782
transform 1 0 47616 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_497
timestamp 1679581782
transform 1 0 48288 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_504
timestamp 1679581782
transform 1 0 48960 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_511
timestamp 1679581782
transform 1 0 49632 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_518
timestamp 1679581782
transform 1 0 50304 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_525
timestamp 1679581782
transform 1 0 50976 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_532
timestamp 1679581782
transform 1 0 51648 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_539
timestamp 1679581782
transform 1 0 52320 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_546
timestamp 1679581782
transform 1 0 52992 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_553
timestamp 1679581782
transform 1 0 53664 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_560
timestamp 1679581782
transform 1 0 54336 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_567
timestamp 1679581782
transform 1 0 55008 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_574
timestamp 1679581782
transform 1 0 55680 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_581
timestamp 1679581782
transform 1 0 56352 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_588
timestamp 1679581782
transform 1 0 57024 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_595
timestamp 1679581782
transform 1 0 57696 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_602
timestamp 1679581782
transform 1 0 58368 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_609
timestamp 1679581782
transform 1 0 59040 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_616
timestamp 1679581782
transform 1 0 59712 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_623
timestamp 1679581782
transform 1 0 60384 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_630
timestamp 1679581782
transform 1 0 61056 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_637
timestamp 1679581782
transform 1 0 61728 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_644
timestamp 1679581782
transform 1 0 62400 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_651
timestamp 1679581782
transform 1 0 63072 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_658
timestamp 1679581782
transform 1 0 63744 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_665
timestamp 1679581782
transform 1 0 64416 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_672
timestamp 1679581782
transform 1 0 65088 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_679
timestamp 1679581782
transform 1 0 65760 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_686
timestamp 1679581782
transform 1 0 66432 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_693
timestamp 1679581782
transform 1 0 67104 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_700
timestamp 1679581782
transform 1 0 67776 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_707
timestamp 1679581782
transform 1 0 68448 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_714
timestamp 1679581782
transform 1 0 69120 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_721
timestamp 1679581782
transform 1 0 69792 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_728
timestamp 1679581782
transform 1 0 70464 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_735
timestamp 1679581782
transform 1 0 71136 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_742
timestamp 1679581782
transform 1 0 71808 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_749
timestamp 1679581782
transform 1 0 72480 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_756
timestamp 1679581782
transform 1 0 73152 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_763
timestamp 1679581782
transform 1 0 73824 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_770
timestamp 1679581782
transform 1 0 74496 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_777
timestamp 1679581782
transform 1 0 75168 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_784
timestamp 1679581782
transform 1 0 75840 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_791
timestamp 1679581782
transform 1 0 76512 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_798
timestamp 1679581782
transform 1 0 77184 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_805
timestamp 1679581782
transform 1 0 77856 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_812
timestamp 1679581782
transform 1 0 78528 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_819
timestamp 1679581782
transform 1 0 79200 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_826
timestamp 1679581782
transform 1 0 79872 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_833
timestamp 1679581782
transform 1 0 80544 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_840
timestamp 1679581782
transform 1 0 81216 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_847
timestamp 1679581782
transform 1 0 81888 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_854
timestamp 1679581782
transform 1 0 82560 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_861
timestamp 1679581782
transform 1 0 83232 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_868
timestamp 1679581782
transform 1 0 83904 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_875
timestamp 1679581782
transform 1 0 84576 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_882
timestamp 1679581782
transform 1 0 85248 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_889
timestamp 1679581782
transform 1 0 85920 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_896
timestamp 1679581782
transform 1 0 86592 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_903
timestamp 1679581782
transform 1 0 87264 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_910
timestamp 1679581782
transform 1 0 87936 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_917
timestamp 1679581782
transform 1 0 88608 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_924
timestamp 1679581782
transform 1 0 89280 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_931
timestamp 1679581782
transform 1 0 89952 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_938
timestamp 1679581782
transform 1 0 90624 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_945
timestamp 1679581782
transform 1 0 91296 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_952
timestamp 1679581782
transform 1 0 91968 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_959
timestamp 1679581782
transform 1 0 92640 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_966
timestamp 1679581782
transform 1 0 93312 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_973
timestamp 1679581782
transform 1 0 93984 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_980
timestamp 1679581782
transform 1 0 94656 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_987
timestamp 1679581782
transform 1 0 95328 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_994
timestamp 1679581782
transform 1 0 96000 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_1001
timestamp 1679581782
transform 1 0 96672 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_1008
timestamp 1679581782
transform 1 0 97344 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_1015
timestamp 1679581782
transform 1 0 98016 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_1022
timestamp 1679581782
transform 1 0 98688 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_4
timestamp 1679581782
transform 1 0 960 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_11
timestamp 1679581782
transform 1 0 1632 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_18
timestamp 1679581782
transform 1 0 2304 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_25
timestamp 1679581782
transform 1 0 2976 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_32
timestamp 1679581782
transform 1 0 3648 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_39
timestamp 1679581782
transform 1 0 4320 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_46
timestamp 1679581782
transform 1 0 4992 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_53
timestamp 1679581782
transform 1 0 5664 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_60
timestamp 1679581782
transform 1 0 6336 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_67
timestamp 1679581782
transform 1 0 7008 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_74
timestamp 1679581782
transform 1 0 7680 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_81
timestamp 1679581782
transform 1 0 8352 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_88
timestamp 1679581782
transform 1 0 9024 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_95
timestamp 1679581782
transform 1 0 9696 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_102
timestamp 1679581782
transform 1 0 10368 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_109
timestamp 1679581782
transform 1 0 11040 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_116
timestamp 1679581782
transform 1 0 11712 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_123
timestamp 1679581782
transform 1 0 12384 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_130
timestamp 1679581782
transform 1 0 13056 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_137
timestamp 1679581782
transform 1 0 13728 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_144
timestamp 1679581782
transform 1 0 14400 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_151
timestamp 1679581782
transform 1 0 15072 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_158
timestamp 1679581782
transform 1 0 15744 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_165
timestamp 1679581782
transform 1 0 16416 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_172
timestamp 1679581782
transform 1 0 17088 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_179
timestamp 1679581782
transform 1 0 17760 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_186
timestamp 1679581782
transform 1 0 18432 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_193
timestamp 1679581782
transform 1 0 19104 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_200
timestamp 1679581782
transform 1 0 19776 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_207
timestamp 1679581782
transform 1 0 20448 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_214
timestamp 1679581782
transform 1 0 21120 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_221
timestamp 1679581782
transform 1 0 21792 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_228
timestamp 1679581782
transform 1 0 22464 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_235
timestamp 1679581782
transform 1 0 23136 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_242
timestamp 1679581782
transform 1 0 23808 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_249
timestamp 1679581782
transform 1 0 24480 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_256
timestamp 1679581782
transform 1 0 25152 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_263
timestamp 1679581782
transform 1 0 25824 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_270
timestamp 1679581782
transform 1 0 26496 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_277
timestamp 1679581782
transform 1 0 27168 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_284
timestamp 1679581782
transform 1 0 27840 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_291
timestamp 1679581782
transform 1 0 28512 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_298
timestamp 1679581782
transform 1 0 29184 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_305
timestamp 1679581782
transform 1 0 29856 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_312
timestamp 1679581782
transform 1 0 30528 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_319
timestamp 1679581782
transform 1 0 31200 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_326
timestamp 1679581782
transform 1 0 31872 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_333
timestamp 1679581782
transform 1 0 32544 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_340
timestamp 1679581782
transform 1 0 33216 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_347
timestamp 1679581782
transform 1 0 33888 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_354
timestamp 1679581782
transform 1 0 34560 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_361
timestamp 1679581782
transform 1 0 35232 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_368
timestamp 1679581782
transform 1 0 35904 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_375
timestamp 1679581782
transform 1 0 36576 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_382
timestamp 1679581782
transform 1 0 37248 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_389
timestamp 1679581782
transform 1 0 37920 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_396
timestamp 1679581782
transform 1 0 38592 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_403
timestamp 1679581782
transform 1 0 39264 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_410
timestamp 1679581782
transform 1 0 39936 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_417
timestamp 1679581782
transform 1 0 40608 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_424
timestamp 1679581782
transform 1 0 41280 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_431
timestamp 1679581782
transform 1 0 41952 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_438
timestamp 1679581782
transform 1 0 42624 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_445
timestamp 1679581782
transform 1 0 43296 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_452
timestamp 1679581782
transform 1 0 43968 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_459
timestamp 1679581782
transform 1 0 44640 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_466
timestamp 1679581782
transform 1 0 45312 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_473
timestamp 1679581782
transform 1 0 45984 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_480
timestamp 1679581782
transform 1 0 46656 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_487
timestamp 1679581782
transform 1 0 47328 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_494
timestamp 1679581782
transform 1 0 48000 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_501
timestamp 1679581782
transform 1 0 48672 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_508
timestamp 1679581782
transform 1 0 49344 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_515
timestamp 1679581782
transform 1 0 50016 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_522
timestamp 1679581782
transform 1 0 50688 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_529
timestamp 1679581782
transform 1 0 51360 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_536
timestamp 1679581782
transform 1 0 52032 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_543
timestamp 1679581782
transform 1 0 52704 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_550
timestamp 1679581782
transform 1 0 53376 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_557
timestamp 1679581782
transform 1 0 54048 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_564
timestamp 1679581782
transform 1 0 54720 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_571
timestamp 1679581782
transform 1 0 55392 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_578
timestamp 1679581782
transform 1 0 56064 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_585
timestamp 1679581782
transform 1 0 56736 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_592
timestamp 1679581782
transform 1 0 57408 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_599
timestamp 1679581782
transform 1 0 58080 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_606
timestamp 1679581782
transform 1 0 58752 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_613
timestamp 1679581782
transform 1 0 59424 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_620
timestamp 1679581782
transform 1 0 60096 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_627
timestamp 1679581782
transform 1 0 60768 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_634
timestamp 1679581782
transform 1 0 61440 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_641
timestamp 1679581782
transform 1 0 62112 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_648
timestamp 1679581782
transform 1 0 62784 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_655
timestamp 1679581782
transform 1 0 63456 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_662
timestamp 1679581782
transform 1 0 64128 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_669
timestamp 1679581782
transform 1 0 64800 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_676
timestamp 1679581782
transform 1 0 65472 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_683
timestamp 1679581782
transform 1 0 66144 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_690
timestamp 1679581782
transform 1 0 66816 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_697
timestamp 1679581782
transform 1 0 67488 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_704
timestamp 1679581782
transform 1 0 68160 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_711
timestamp 1679581782
transform 1 0 68832 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_718
timestamp 1679581782
transform 1 0 69504 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_725
timestamp 1679581782
transform 1 0 70176 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_732
timestamp 1679581782
transform 1 0 70848 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_739
timestamp 1679581782
transform 1 0 71520 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_746
timestamp 1679581782
transform 1 0 72192 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_753
timestamp 1679581782
transform 1 0 72864 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_760
timestamp 1679581782
transform 1 0 73536 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_767
timestamp 1679581782
transform 1 0 74208 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_774
timestamp 1679581782
transform 1 0 74880 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_781
timestamp 1679581782
transform 1 0 75552 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_788
timestamp 1679581782
transform 1 0 76224 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_795
timestamp 1679581782
transform 1 0 76896 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_802
timestamp 1679581782
transform 1 0 77568 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_809
timestamp 1679581782
transform 1 0 78240 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_816
timestamp 1679581782
transform 1 0 78912 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_823
timestamp 1679581782
transform 1 0 79584 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_830
timestamp 1679581782
transform 1 0 80256 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_837
timestamp 1679581782
transform 1 0 80928 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_844
timestamp 1679581782
transform 1 0 81600 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_851
timestamp 1679581782
transform 1 0 82272 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_858
timestamp 1679581782
transform 1 0 82944 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_865
timestamp 1679581782
transform 1 0 83616 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_872
timestamp 1679581782
transform 1 0 84288 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_879
timestamp 1679581782
transform 1 0 84960 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_886
timestamp 1679581782
transform 1 0 85632 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_893
timestamp 1679581782
transform 1 0 86304 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_900
timestamp 1679581782
transform 1 0 86976 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_907
timestamp 1679581782
transform 1 0 87648 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_914
timestamp 1679581782
transform 1 0 88320 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_921
timestamp 1679581782
transform 1 0 88992 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_928
timestamp 1679581782
transform 1 0 89664 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_935
timestamp 1679581782
transform 1 0 90336 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_942
timestamp 1679581782
transform 1 0 91008 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_949
timestamp 1679581782
transform 1 0 91680 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_956
timestamp 1679581782
transform 1 0 92352 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_963
timestamp 1679581782
transform 1 0 93024 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_970
timestamp 1679581782
transform 1 0 93696 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_977
timestamp 1679581782
transform 1 0 94368 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_984
timestamp 1679581782
transform 1 0 95040 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_991
timestamp 1679581782
transform 1 0 95712 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_998
timestamp 1679581782
transform 1 0 96384 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_1005
timestamp 1679581782
transform 1 0 97056 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_1012
timestamp 1679581782
transform 1 0 97728 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_1019
timestamp 1679581782
transform 1 0 98400 0 1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_20_1026
timestamp 1677580104
transform 1 0 99072 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_1028
timestamp 1677579658
transform 1 0 99264 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_0
timestamp 1679581782
transform 1 0 576 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_7
timestamp 1679581782
transform 1 0 1248 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_14
timestamp 1679581782
transform 1 0 1920 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_21
timestamp 1679581782
transform 1 0 2592 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_28
timestamp 1679581782
transform 1 0 3264 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_35
timestamp 1679581782
transform 1 0 3936 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_42
timestamp 1679581782
transform 1 0 4608 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_49
timestamp 1679581782
transform 1 0 5280 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_56
timestamp 1679581782
transform 1 0 5952 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_63
timestamp 1679581782
transform 1 0 6624 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_70
timestamp 1679581782
transform 1 0 7296 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_77
timestamp 1679581782
transform 1 0 7968 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_84
timestamp 1679581782
transform 1 0 8640 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_91
timestamp 1679581782
transform 1 0 9312 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_98
timestamp 1679581782
transform 1 0 9984 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_105
timestamp 1679581782
transform 1 0 10656 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_112
timestamp 1679581782
transform 1 0 11328 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_119
timestamp 1679581782
transform 1 0 12000 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_126
timestamp 1679581782
transform 1 0 12672 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_133
timestamp 1679581782
transform 1 0 13344 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_140
timestamp 1679581782
transform 1 0 14016 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_147
timestamp 1679581782
transform 1 0 14688 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_154
timestamp 1679581782
transform 1 0 15360 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_161
timestamp 1679581782
transform 1 0 16032 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_168
timestamp 1679581782
transform 1 0 16704 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_175
timestamp 1679581782
transform 1 0 17376 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_182
timestamp 1679581782
transform 1 0 18048 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_189
timestamp 1679581782
transform 1 0 18720 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_196
timestamp 1679581782
transform 1 0 19392 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_203
timestamp 1679581782
transform 1 0 20064 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_210
timestamp 1679581782
transform 1 0 20736 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_217
timestamp 1679581782
transform 1 0 21408 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_224
timestamp 1679581782
transform 1 0 22080 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_231
timestamp 1679581782
transform 1 0 22752 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_238
timestamp 1679581782
transform 1 0 23424 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_245
timestamp 1679581782
transform 1 0 24096 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_252
timestamp 1679581782
transform 1 0 24768 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_259
timestamp 1679581782
transform 1 0 25440 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_266
timestamp 1679581782
transform 1 0 26112 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_273
timestamp 1679581782
transform 1 0 26784 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_280
timestamp 1679581782
transform 1 0 27456 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_287
timestamp 1679581782
transform 1 0 28128 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_294
timestamp 1679581782
transform 1 0 28800 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_301
timestamp 1679581782
transform 1 0 29472 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_308
timestamp 1679581782
transform 1 0 30144 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_315
timestamp 1679581782
transform 1 0 30816 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_322
timestamp 1679581782
transform 1 0 31488 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_329
timestamp 1679581782
transform 1 0 32160 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_336
timestamp 1679581782
transform 1 0 32832 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_343
timestamp 1679581782
transform 1 0 33504 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_350
timestamp 1679581782
transform 1 0 34176 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_357
timestamp 1679581782
transform 1 0 34848 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_364
timestamp 1679581782
transform 1 0 35520 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_371
timestamp 1679581782
transform 1 0 36192 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_378
timestamp 1679581782
transform 1 0 36864 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_385
timestamp 1679581782
transform 1 0 37536 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_392
timestamp 1679581782
transform 1 0 38208 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_399
timestamp 1679581782
transform 1 0 38880 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_406
timestamp 1679581782
transform 1 0 39552 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_413
timestamp 1679581782
transform 1 0 40224 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_420
timestamp 1679581782
transform 1 0 40896 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_427
timestamp 1679581782
transform 1 0 41568 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_434
timestamp 1679581782
transform 1 0 42240 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_441
timestamp 1679581782
transform 1 0 42912 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_448
timestamp 1679581782
transform 1 0 43584 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_455
timestamp 1679581782
transform 1 0 44256 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_462
timestamp 1679581782
transform 1 0 44928 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_469
timestamp 1679581782
transform 1 0 45600 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_476
timestamp 1679581782
transform 1 0 46272 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_483
timestamp 1679581782
transform 1 0 46944 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_490
timestamp 1679581782
transform 1 0 47616 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_497
timestamp 1679581782
transform 1 0 48288 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_504
timestamp 1679581782
transform 1 0 48960 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_511
timestamp 1679581782
transform 1 0 49632 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_518
timestamp 1679581782
transform 1 0 50304 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_525
timestamp 1679581782
transform 1 0 50976 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_532
timestamp 1679581782
transform 1 0 51648 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_539
timestamp 1679581782
transform 1 0 52320 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_546
timestamp 1679581782
transform 1 0 52992 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_553
timestamp 1679581782
transform 1 0 53664 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_560
timestamp 1679581782
transform 1 0 54336 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_567
timestamp 1679581782
transform 1 0 55008 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_574
timestamp 1679581782
transform 1 0 55680 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_581
timestamp 1679581782
transform 1 0 56352 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_588
timestamp 1679581782
transform 1 0 57024 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_595
timestamp 1679581782
transform 1 0 57696 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_602
timestamp 1679581782
transform 1 0 58368 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_609
timestamp 1679581782
transform 1 0 59040 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_616
timestamp 1679581782
transform 1 0 59712 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_623
timestamp 1679581782
transform 1 0 60384 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_630
timestamp 1679581782
transform 1 0 61056 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_637
timestamp 1679581782
transform 1 0 61728 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_644
timestamp 1679581782
transform 1 0 62400 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_651
timestamp 1679581782
transform 1 0 63072 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_658
timestamp 1679581782
transform 1 0 63744 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_665
timestamp 1679581782
transform 1 0 64416 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_672
timestamp 1679581782
transform 1 0 65088 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_679
timestamp 1679581782
transform 1 0 65760 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_686
timestamp 1679581782
transform 1 0 66432 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_693
timestamp 1679581782
transform 1 0 67104 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_700
timestamp 1679581782
transform 1 0 67776 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_707
timestamp 1679581782
transform 1 0 68448 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_714
timestamp 1679581782
transform 1 0 69120 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_721
timestamp 1679581782
transform 1 0 69792 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_728
timestamp 1679581782
transform 1 0 70464 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_735
timestamp 1679581782
transform 1 0 71136 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_742
timestamp 1679581782
transform 1 0 71808 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_749
timestamp 1679581782
transform 1 0 72480 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_756
timestamp 1679581782
transform 1 0 73152 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_763
timestamp 1679581782
transform 1 0 73824 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_770
timestamp 1679581782
transform 1 0 74496 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_777
timestamp 1679581782
transform 1 0 75168 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_784
timestamp 1679581782
transform 1 0 75840 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_791
timestamp 1679581782
transform 1 0 76512 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_798
timestamp 1679581782
transform 1 0 77184 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_805
timestamp 1679581782
transform 1 0 77856 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_812
timestamp 1679581782
transform 1 0 78528 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_819
timestamp 1679581782
transform 1 0 79200 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_826
timestamp 1679581782
transform 1 0 79872 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_833
timestamp 1679581782
transform 1 0 80544 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_840
timestamp 1679581782
transform 1 0 81216 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_847
timestamp 1679581782
transform 1 0 81888 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_854
timestamp 1679581782
transform 1 0 82560 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_861
timestamp 1679581782
transform 1 0 83232 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_868
timestamp 1679581782
transform 1 0 83904 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_875
timestamp 1679581782
transform 1 0 84576 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_882
timestamp 1679581782
transform 1 0 85248 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_889
timestamp 1679581782
transform 1 0 85920 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_896
timestamp 1679581782
transform 1 0 86592 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_903
timestamp 1679581782
transform 1 0 87264 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_910
timestamp 1679581782
transform 1 0 87936 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_917
timestamp 1679581782
transform 1 0 88608 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_924
timestamp 1679581782
transform 1 0 89280 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_931
timestamp 1679581782
transform 1 0 89952 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_938
timestamp 1679581782
transform 1 0 90624 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_945
timestamp 1679581782
transform 1 0 91296 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_952
timestamp 1679581782
transform 1 0 91968 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_959
timestamp 1679581782
transform 1 0 92640 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_966
timestamp 1679581782
transform 1 0 93312 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_973
timestamp 1679581782
transform 1 0 93984 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_980
timestamp 1679581782
transform 1 0 94656 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_987
timestamp 1679581782
transform 1 0 95328 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_994
timestamp 1679581782
transform 1 0 96000 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_1001
timestamp 1679581782
transform 1 0 96672 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_1008
timestamp 1679581782
transform 1 0 97344 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_1015
timestamp 1679581782
transform 1 0 98016 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_1022
timestamp 1679581782
transform 1 0 98688 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_4
timestamp 1679581782
transform 1 0 960 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_11
timestamp 1679581782
transform 1 0 1632 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_18
timestamp 1679581782
transform 1 0 2304 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_25
timestamp 1679581782
transform 1 0 2976 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_32
timestamp 1679581782
transform 1 0 3648 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_39
timestamp 1679581782
transform 1 0 4320 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_46
timestamp 1679581782
transform 1 0 4992 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_53
timestamp 1679581782
transform 1 0 5664 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_60
timestamp 1679581782
transform 1 0 6336 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_67
timestamp 1679581782
transform 1 0 7008 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_74
timestamp 1679581782
transform 1 0 7680 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_81
timestamp 1679581782
transform 1 0 8352 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_88
timestamp 1679581782
transform 1 0 9024 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_95
timestamp 1679581782
transform 1 0 9696 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_102
timestamp 1679581782
transform 1 0 10368 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_109
timestamp 1679581782
transform 1 0 11040 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_116
timestamp 1679581782
transform 1 0 11712 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_123
timestamp 1679581782
transform 1 0 12384 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_130
timestamp 1679581782
transform 1 0 13056 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_137
timestamp 1679581782
transform 1 0 13728 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_144
timestamp 1679581782
transform 1 0 14400 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_151
timestamp 1679581782
transform 1 0 15072 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_158
timestamp 1679581782
transform 1 0 15744 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_165
timestamp 1679581782
transform 1 0 16416 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_172
timestamp 1679581782
transform 1 0 17088 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_179
timestamp 1679581782
transform 1 0 17760 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_186
timestamp 1679581782
transform 1 0 18432 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_193
timestamp 1679581782
transform 1 0 19104 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_200
timestamp 1679581782
transform 1 0 19776 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_207
timestamp 1679581782
transform 1 0 20448 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_214
timestamp 1679581782
transform 1 0 21120 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_221
timestamp 1679581782
transform 1 0 21792 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_228
timestamp 1679581782
transform 1 0 22464 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_235
timestamp 1679581782
transform 1 0 23136 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_242
timestamp 1679581782
transform 1 0 23808 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_249
timestamp 1679581782
transform 1 0 24480 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_256
timestamp 1679581782
transform 1 0 25152 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_263
timestamp 1679581782
transform 1 0 25824 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_270
timestamp 1679581782
transform 1 0 26496 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_277
timestamp 1679581782
transform 1 0 27168 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_284
timestamp 1679581782
transform 1 0 27840 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_291
timestamp 1679581782
transform 1 0 28512 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_298
timestamp 1679581782
transform 1 0 29184 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_305
timestamp 1679581782
transform 1 0 29856 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_312
timestamp 1679581782
transform 1 0 30528 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_319
timestamp 1679581782
transform 1 0 31200 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_326
timestamp 1679581782
transform 1 0 31872 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_333
timestamp 1679581782
transform 1 0 32544 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_340
timestamp 1679581782
transform 1 0 33216 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_347
timestamp 1679581782
transform 1 0 33888 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_354
timestamp 1679581782
transform 1 0 34560 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_361
timestamp 1679581782
transform 1 0 35232 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_368
timestamp 1679581782
transform 1 0 35904 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_375
timestamp 1679581782
transform 1 0 36576 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_382
timestamp 1679581782
transform 1 0 37248 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_389
timestamp 1679581782
transform 1 0 37920 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_396
timestamp 1679581782
transform 1 0 38592 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_403
timestamp 1679581782
transform 1 0 39264 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_410
timestamp 1679581782
transform 1 0 39936 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_417
timestamp 1679581782
transform 1 0 40608 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_424
timestamp 1679581782
transform 1 0 41280 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_431
timestamp 1679581782
transform 1 0 41952 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_438
timestamp 1679581782
transform 1 0 42624 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_445
timestamp 1679581782
transform 1 0 43296 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_452
timestamp 1679581782
transform 1 0 43968 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_459
timestamp 1679581782
transform 1 0 44640 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_466
timestamp 1679581782
transform 1 0 45312 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_473
timestamp 1679581782
transform 1 0 45984 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_480
timestamp 1679581782
transform 1 0 46656 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_487
timestamp 1679581782
transform 1 0 47328 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_494
timestamp 1679581782
transform 1 0 48000 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_501
timestamp 1679581782
transform 1 0 48672 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_508
timestamp 1679581782
transform 1 0 49344 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_515
timestamp 1679581782
transform 1 0 50016 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_522
timestamp 1679581782
transform 1 0 50688 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_529
timestamp 1679581782
transform 1 0 51360 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_536
timestamp 1679581782
transform 1 0 52032 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_543
timestamp 1679581782
transform 1 0 52704 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_550
timestamp 1679581782
transform 1 0 53376 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_557
timestamp 1679581782
transform 1 0 54048 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_564
timestamp 1679581782
transform 1 0 54720 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_571
timestamp 1679581782
transform 1 0 55392 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_578
timestamp 1679581782
transform 1 0 56064 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_585
timestamp 1679581782
transform 1 0 56736 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_592
timestamp 1679581782
transform 1 0 57408 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_599
timestamp 1679581782
transform 1 0 58080 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_606
timestamp 1679581782
transform 1 0 58752 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_613
timestamp 1679581782
transform 1 0 59424 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_620
timestamp 1679581782
transform 1 0 60096 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_627
timestamp 1679581782
transform 1 0 60768 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_634
timestamp 1679581782
transform 1 0 61440 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_641
timestamp 1679581782
transform 1 0 62112 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_648
timestamp 1679581782
transform 1 0 62784 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_655
timestamp 1679581782
transform 1 0 63456 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_662
timestamp 1679581782
transform 1 0 64128 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_669
timestamp 1679581782
transform 1 0 64800 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_676
timestamp 1679581782
transform 1 0 65472 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_683
timestamp 1679581782
transform 1 0 66144 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_690
timestamp 1679581782
transform 1 0 66816 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_697
timestamp 1679581782
transform 1 0 67488 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_704
timestamp 1679581782
transform 1 0 68160 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_711
timestamp 1679581782
transform 1 0 68832 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_718
timestamp 1679581782
transform 1 0 69504 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_725
timestamp 1679581782
transform 1 0 70176 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_732
timestamp 1679581782
transform 1 0 70848 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_739
timestamp 1679581782
transform 1 0 71520 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_746
timestamp 1679581782
transform 1 0 72192 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_753
timestamp 1679581782
transform 1 0 72864 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_760
timestamp 1679581782
transform 1 0 73536 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_767
timestamp 1679581782
transform 1 0 74208 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_774
timestamp 1679581782
transform 1 0 74880 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_781
timestamp 1679581782
transform 1 0 75552 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_788
timestamp 1679581782
transform 1 0 76224 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_795
timestamp 1679581782
transform 1 0 76896 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_802
timestamp 1679581782
transform 1 0 77568 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_809
timestamp 1679581782
transform 1 0 78240 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_816
timestamp 1679581782
transform 1 0 78912 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_823
timestamp 1679581782
transform 1 0 79584 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_830
timestamp 1679581782
transform 1 0 80256 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_837
timestamp 1679581782
transform 1 0 80928 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_844
timestamp 1679581782
transform 1 0 81600 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_851
timestamp 1679581782
transform 1 0 82272 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_858
timestamp 1679581782
transform 1 0 82944 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_865
timestamp 1679581782
transform 1 0 83616 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_872
timestamp 1679581782
transform 1 0 84288 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_879
timestamp 1679581782
transform 1 0 84960 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_886
timestamp 1679581782
transform 1 0 85632 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_893
timestamp 1679581782
transform 1 0 86304 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_900
timestamp 1679581782
transform 1 0 86976 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_907
timestamp 1679581782
transform 1 0 87648 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_914
timestamp 1679581782
transform 1 0 88320 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_921
timestamp 1679581782
transform 1 0 88992 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_928
timestamp 1679581782
transform 1 0 89664 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_935
timestamp 1679581782
transform 1 0 90336 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_942
timestamp 1679581782
transform 1 0 91008 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_949
timestamp 1679581782
transform 1 0 91680 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_956
timestamp 1679581782
transform 1 0 92352 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_963
timestamp 1679581782
transform 1 0 93024 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_970
timestamp 1679581782
transform 1 0 93696 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_977
timestamp 1679581782
transform 1 0 94368 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_984
timestamp 1679581782
transform 1 0 95040 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_991
timestamp 1679581782
transform 1 0 95712 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_998
timestamp 1679581782
transform 1 0 96384 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_1005
timestamp 1679581782
transform 1 0 97056 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_1012
timestamp 1679581782
transform 1 0 97728 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_1019
timestamp 1679581782
transform 1 0 98400 0 1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_22_1026
timestamp 1677580104
transform 1 0 99072 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_1028
timestamp 1677579658
transform 1 0 99264 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_0
timestamp 1679581782
transform 1 0 576 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_7
timestamp 1679581782
transform 1 0 1248 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_14
timestamp 1679581782
transform 1 0 1920 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_21
timestamp 1679581782
transform 1 0 2592 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_28
timestamp 1679581782
transform 1 0 3264 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_35
timestamp 1679581782
transform 1 0 3936 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_42
timestamp 1679581782
transform 1 0 4608 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_49
timestamp 1679581782
transform 1 0 5280 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_56
timestamp 1679581782
transform 1 0 5952 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_63
timestamp 1679581782
transform 1 0 6624 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_70
timestamp 1679581782
transform 1 0 7296 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_77
timestamp 1679581782
transform 1 0 7968 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_84
timestamp 1679581782
transform 1 0 8640 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_91
timestamp 1679581782
transform 1 0 9312 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_98
timestamp 1679581782
transform 1 0 9984 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_105
timestamp 1679581782
transform 1 0 10656 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_112
timestamp 1679581782
transform 1 0 11328 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_119
timestamp 1679581782
transform 1 0 12000 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_126
timestamp 1679581782
transform 1 0 12672 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_133
timestamp 1679581782
transform 1 0 13344 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_140
timestamp 1679581782
transform 1 0 14016 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_147
timestamp 1679581782
transform 1 0 14688 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_154
timestamp 1679581782
transform 1 0 15360 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_161
timestamp 1679581782
transform 1 0 16032 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_168
timestamp 1679581782
transform 1 0 16704 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_175
timestamp 1679581782
transform 1 0 17376 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_182
timestamp 1679581782
transform 1 0 18048 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_189
timestamp 1679581782
transform 1 0 18720 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_196
timestamp 1679581782
transform 1 0 19392 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_203
timestamp 1679581782
transform 1 0 20064 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_210
timestamp 1679581782
transform 1 0 20736 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_217
timestamp 1679581782
transform 1 0 21408 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_224
timestamp 1679581782
transform 1 0 22080 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_231
timestamp 1679581782
transform 1 0 22752 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_238
timestamp 1679581782
transform 1 0 23424 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_245
timestamp 1679581782
transform 1 0 24096 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_252
timestamp 1679581782
transform 1 0 24768 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_259
timestamp 1679581782
transform 1 0 25440 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_266
timestamp 1679581782
transform 1 0 26112 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_273
timestamp 1679581782
transform 1 0 26784 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_280
timestamp 1679581782
transform 1 0 27456 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_287
timestamp 1679581782
transform 1 0 28128 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_294
timestamp 1679581782
transform 1 0 28800 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_301
timestamp 1679581782
transform 1 0 29472 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_308
timestamp 1679581782
transform 1 0 30144 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_315
timestamp 1679581782
transform 1 0 30816 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_322
timestamp 1679581782
transform 1 0 31488 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_329
timestamp 1679581782
transform 1 0 32160 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_336
timestamp 1679581782
transform 1 0 32832 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_343
timestamp 1679581782
transform 1 0 33504 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_350
timestamp 1679581782
transform 1 0 34176 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_357
timestamp 1679581782
transform 1 0 34848 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_364
timestamp 1679581782
transform 1 0 35520 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_371
timestamp 1679581782
transform 1 0 36192 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_378
timestamp 1679581782
transform 1 0 36864 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_385
timestamp 1679581782
transform 1 0 37536 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_392
timestamp 1679581782
transform 1 0 38208 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_399
timestamp 1679581782
transform 1 0 38880 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_406
timestamp 1679581782
transform 1 0 39552 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_413
timestamp 1679581782
transform 1 0 40224 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_420
timestamp 1679581782
transform 1 0 40896 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_427
timestamp 1679581782
transform 1 0 41568 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_434
timestamp 1679581782
transform 1 0 42240 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_441
timestamp 1679581782
transform 1 0 42912 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_448
timestamp 1679581782
transform 1 0 43584 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_455
timestamp 1679581782
transform 1 0 44256 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_462
timestamp 1679581782
transform 1 0 44928 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_469
timestamp 1679581782
transform 1 0 45600 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_476
timestamp 1679581782
transform 1 0 46272 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_483
timestamp 1679581782
transform 1 0 46944 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_490
timestamp 1679581782
transform 1 0 47616 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_497
timestamp 1679581782
transform 1 0 48288 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_504
timestamp 1679581782
transform 1 0 48960 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_511
timestamp 1679581782
transform 1 0 49632 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_518
timestamp 1679581782
transform 1 0 50304 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_525
timestamp 1679581782
transform 1 0 50976 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_532
timestamp 1679581782
transform 1 0 51648 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_539
timestamp 1679581782
transform 1 0 52320 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_546
timestamp 1679581782
transform 1 0 52992 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_553
timestamp 1679581782
transform 1 0 53664 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_560
timestamp 1679581782
transform 1 0 54336 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_567
timestamp 1679581782
transform 1 0 55008 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_574
timestamp 1679581782
transform 1 0 55680 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_581
timestamp 1679581782
transform 1 0 56352 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_588
timestamp 1679581782
transform 1 0 57024 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_595
timestamp 1679581782
transform 1 0 57696 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_602
timestamp 1679581782
transform 1 0 58368 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_609
timestamp 1679581782
transform 1 0 59040 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_616
timestamp 1679581782
transform 1 0 59712 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_623
timestamp 1679581782
transform 1 0 60384 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_630
timestamp 1679581782
transform 1 0 61056 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_637
timestamp 1679581782
transform 1 0 61728 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_644
timestamp 1679581782
transform 1 0 62400 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_651
timestamp 1679581782
transform 1 0 63072 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_658
timestamp 1679581782
transform 1 0 63744 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_665
timestamp 1679581782
transform 1 0 64416 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_672
timestamp 1679581782
transform 1 0 65088 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_679
timestamp 1679581782
transform 1 0 65760 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_686
timestamp 1679581782
transform 1 0 66432 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_693
timestamp 1679581782
transform 1 0 67104 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_700
timestamp 1679581782
transform 1 0 67776 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_707
timestamp 1679581782
transform 1 0 68448 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_714
timestamp 1679581782
transform 1 0 69120 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_721
timestamp 1679581782
transform 1 0 69792 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_728
timestamp 1679581782
transform 1 0 70464 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_735
timestamp 1679581782
transform 1 0 71136 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_742
timestamp 1679581782
transform 1 0 71808 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_749
timestamp 1679581782
transform 1 0 72480 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_756
timestamp 1679581782
transform 1 0 73152 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_763
timestamp 1679581782
transform 1 0 73824 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_770
timestamp 1679581782
transform 1 0 74496 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_777
timestamp 1679581782
transform 1 0 75168 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_784
timestamp 1679581782
transform 1 0 75840 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_791
timestamp 1679581782
transform 1 0 76512 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_798
timestamp 1679581782
transform 1 0 77184 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_805
timestamp 1679581782
transform 1 0 77856 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_812
timestamp 1679581782
transform 1 0 78528 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_819
timestamp 1679581782
transform 1 0 79200 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_826
timestamp 1679581782
transform 1 0 79872 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_833
timestamp 1679581782
transform 1 0 80544 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_840
timestamp 1679581782
transform 1 0 81216 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_847
timestamp 1679581782
transform 1 0 81888 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_854
timestamp 1679581782
transform 1 0 82560 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_861
timestamp 1679581782
transform 1 0 83232 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_868
timestamp 1679581782
transform 1 0 83904 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_875
timestamp 1679581782
transform 1 0 84576 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_882
timestamp 1679581782
transform 1 0 85248 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_889
timestamp 1679581782
transform 1 0 85920 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_896
timestamp 1679581782
transform 1 0 86592 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_903
timestamp 1679581782
transform 1 0 87264 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_910
timestamp 1679581782
transform 1 0 87936 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_917
timestamp 1679581782
transform 1 0 88608 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_924
timestamp 1679581782
transform 1 0 89280 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_931
timestamp 1679581782
transform 1 0 89952 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_938
timestamp 1679581782
transform 1 0 90624 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_945
timestamp 1679581782
transform 1 0 91296 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_952
timestamp 1679581782
transform 1 0 91968 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_959
timestamp 1679581782
transform 1 0 92640 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_966
timestamp 1679581782
transform 1 0 93312 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_973
timestamp 1679581782
transform 1 0 93984 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_980
timestamp 1679581782
transform 1 0 94656 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_987
timestamp 1679581782
transform 1 0 95328 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_994
timestamp 1679581782
transform 1 0 96000 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_1001
timestamp 1679581782
transform 1 0 96672 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_1008
timestamp 1679581782
transform 1 0 97344 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_1015
timestamp 1679581782
transform 1 0 98016 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_1022
timestamp 1679581782
transform 1 0 98688 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_4
timestamp 1679581782
transform 1 0 960 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_11
timestamp 1679581782
transform 1 0 1632 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_18
timestamp 1679581782
transform 1 0 2304 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_25
timestamp 1679581782
transform 1 0 2976 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_32
timestamp 1679581782
transform 1 0 3648 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_39
timestamp 1679581782
transform 1 0 4320 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_46
timestamp 1679581782
transform 1 0 4992 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_53
timestamp 1679581782
transform 1 0 5664 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_60
timestamp 1679581782
transform 1 0 6336 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_67
timestamp 1679581782
transform 1 0 7008 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_74
timestamp 1679581782
transform 1 0 7680 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_81
timestamp 1679581782
transform 1 0 8352 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_88
timestamp 1679581782
transform 1 0 9024 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_95
timestamp 1679581782
transform 1 0 9696 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_102
timestamp 1679581782
transform 1 0 10368 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_109
timestamp 1679581782
transform 1 0 11040 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_116
timestamp 1679581782
transform 1 0 11712 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_123
timestamp 1679581782
transform 1 0 12384 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_130
timestamp 1679581782
transform 1 0 13056 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_137
timestamp 1679581782
transform 1 0 13728 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_144
timestamp 1679581782
transform 1 0 14400 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_151
timestamp 1679581782
transform 1 0 15072 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_158
timestamp 1679581782
transform 1 0 15744 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_165
timestamp 1679581782
transform 1 0 16416 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_172
timestamp 1679581782
transform 1 0 17088 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_179
timestamp 1679581782
transform 1 0 17760 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_186
timestamp 1679581782
transform 1 0 18432 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_193
timestamp 1679581782
transform 1 0 19104 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_200
timestamp 1679581782
transform 1 0 19776 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_207
timestamp 1679581782
transform 1 0 20448 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_214
timestamp 1679581782
transform 1 0 21120 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_221
timestamp 1679581782
transform 1 0 21792 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_228
timestamp 1679581782
transform 1 0 22464 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_235
timestamp 1679581782
transform 1 0 23136 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_242
timestamp 1679581782
transform 1 0 23808 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_249
timestamp 1679581782
transform 1 0 24480 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_256
timestamp 1679581782
transform 1 0 25152 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_263
timestamp 1679581782
transform 1 0 25824 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_270
timestamp 1679581782
transform 1 0 26496 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_277
timestamp 1679581782
transform 1 0 27168 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_284
timestamp 1679581782
transform 1 0 27840 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_291
timestamp 1679581782
transform 1 0 28512 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_298
timestamp 1679581782
transform 1 0 29184 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_305
timestamp 1679581782
transform 1 0 29856 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_312
timestamp 1679581782
transform 1 0 30528 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_319
timestamp 1679581782
transform 1 0 31200 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_326
timestamp 1679581782
transform 1 0 31872 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_333
timestamp 1679581782
transform 1 0 32544 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_340
timestamp 1679581782
transform 1 0 33216 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_347
timestamp 1679581782
transform 1 0 33888 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_354
timestamp 1679581782
transform 1 0 34560 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_361
timestamp 1679581782
transform 1 0 35232 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_368
timestamp 1679581782
transform 1 0 35904 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_375
timestamp 1679581782
transform 1 0 36576 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_382
timestamp 1679581782
transform 1 0 37248 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_389
timestamp 1679581782
transform 1 0 37920 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_396
timestamp 1679581782
transform 1 0 38592 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_403
timestamp 1679581782
transform 1 0 39264 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_410
timestamp 1679581782
transform 1 0 39936 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_417
timestamp 1679581782
transform 1 0 40608 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_424
timestamp 1679581782
transform 1 0 41280 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_431
timestamp 1679581782
transform 1 0 41952 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_438
timestamp 1679581782
transform 1 0 42624 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_445
timestamp 1679581782
transform 1 0 43296 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_452
timestamp 1679581782
transform 1 0 43968 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_459
timestamp 1679581782
transform 1 0 44640 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_466
timestamp 1679581782
transform 1 0 45312 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_473
timestamp 1679581782
transform 1 0 45984 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_480
timestamp 1679581782
transform 1 0 46656 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_487
timestamp 1679581782
transform 1 0 47328 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_494
timestamp 1679581782
transform 1 0 48000 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_501
timestamp 1679581782
transform 1 0 48672 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_508
timestamp 1679581782
transform 1 0 49344 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_515
timestamp 1679581782
transform 1 0 50016 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_522
timestamp 1679581782
transform 1 0 50688 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_529
timestamp 1679581782
transform 1 0 51360 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_536
timestamp 1679581782
transform 1 0 52032 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_543
timestamp 1679581782
transform 1 0 52704 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_550
timestamp 1679581782
transform 1 0 53376 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_557
timestamp 1679581782
transform 1 0 54048 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_564
timestamp 1679581782
transform 1 0 54720 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_571
timestamp 1679581782
transform 1 0 55392 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_578
timestamp 1679581782
transform 1 0 56064 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_585
timestamp 1679581782
transform 1 0 56736 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_592
timestamp 1679581782
transform 1 0 57408 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_599
timestamp 1679581782
transform 1 0 58080 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_606
timestamp 1679581782
transform 1 0 58752 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_613
timestamp 1679581782
transform 1 0 59424 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_620
timestamp 1679581782
transform 1 0 60096 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_627
timestamp 1679581782
transform 1 0 60768 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_634
timestamp 1679581782
transform 1 0 61440 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_641
timestamp 1679581782
transform 1 0 62112 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_648
timestamp 1679581782
transform 1 0 62784 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_655
timestamp 1679581782
transform 1 0 63456 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_662
timestamp 1679581782
transform 1 0 64128 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_669
timestamp 1679581782
transform 1 0 64800 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_676
timestamp 1679581782
transform 1 0 65472 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_683
timestamp 1679581782
transform 1 0 66144 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_690
timestamp 1679581782
transform 1 0 66816 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_697
timestamp 1679581782
transform 1 0 67488 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_704
timestamp 1679581782
transform 1 0 68160 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_711
timestamp 1679581782
transform 1 0 68832 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_718
timestamp 1679581782
transform 1 0 69504 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_725
timestamp 1679581782
transform 1 0 70176 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_732
timestamp 1679581782
transform 1 0 70848 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_739
timestamp 1679581782
transform 1 0 71520 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_746
timestamp 1679581782
transform 1 0 72192 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_753
timestamp 1679581782
transform 1 0 72864 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_760
timestamp 1679581782
transform 1 0 73536 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_767
timestamp 1679581782
transform 1 0 74208 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_774
timestamp 1679581782
transform 1 0 74880 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_781
timestamp 1679581782
transform 1 0 75552 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_788
timestamp 1679581782
transform 1 0 76224 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_795
timestamp 1679581782
transform 1 0 76896 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_802
timestamp 1679581782
transform 1 0 77568 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_809
timestamp 1679581782
transform 1 0 78240 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_816
timestamp 1679581782
transform 1 0 78912 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_823
timestamp 1679581782
transform 1 0 79584 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_830
timestamp 1679581782
transform 1 0 80256 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_837
timestamp 1679581782
transform 1 0 80928 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_844
timestamp 1679581782
transform 1 0 81600 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_851
timestamp 1679581782
transform 1 0 82272 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_858
timestamp 1679581782
transform 1 0 82944 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_865
timestamp 1679581782
transform 1 0 83616 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_872
timestamp 1679581782
transform 1 0 84288 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_879
timestamp 1679581782
transform 1 0 84960 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_886
timestamp 1679581782
transform 1 0 85632 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_893
timestamp 1679581782
transform 1 0 86304 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_900
timestamp 1679581782
transform 1 0 86976 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_907
timestamp 1679581782
transform 1 0 87648 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_914
timestamp 1679581782
transform 1 0 88320 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_921
timestamp 1679581782
transform 1 0 88992 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_928
timestamp 1679581782
transform 1 0 89664 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_935
timestamp 1679581782
transform 1 0 90336 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_942
timestamp 1679581782
transform 1 0 91008 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_949
timestamp 1679581782
transform 1 0 91680 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_956
timestamp 1679581782
transform 1 0 92352 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_963
timestamp 1679581782
transform 1 0 93024 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_970
timestamp 1679581782
transform 1 0 93696 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_977
timestamp 1679581782
transform 1 0 94368 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_984
timestamp 1679581782
transform 1 0 95040 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_991
timestamp 1679581782
transform 1 0 95712 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_998
timestamp 1679581782
transform 1 0 96384 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_1005
timestamp 1679581782
transform 1 0 97056 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_1012
timestamp 1679581782
transform 1 0 97728 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_1019
timestamp 1679581782
transform 1 0 98400 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_24_1026
timestamp 1677580104
transform 1 0 99072 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_1028
timestamp 1677579658
transform 1 0 99264 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_0
timestamp 1679581782
transform 1 0 576 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_7
timestamp 1679581782
transform 1 0 1248 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_14
timestamp 1679581782
transform 1 0 1920 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_21
timestamp 1679581782
transform 1 0 2592 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_28
timestamp 1679581782
transform 1 0 3264 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_35
timestamp 1679581782
transform 1 0 3936 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_42
timestamp 1679581782
transform 1 0 4608 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_49
timestamp 1679581782
transform 1 0 5280 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_56
timestamp 1679581782
transform 1 0 5952 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_63
timestamp 1679581782
transform 1 0 6624 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_70
timestamp 1679581782
transform 1 0 7296 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_77
timestamp 1679581782
transform 1 0 7968 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_84
timestamp 1679581782
transform 1 0 8640 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_91
timestamp 1679581782
transform 1 0 9312 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_98
timestamp 1679581782
transform 1 0 9984 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_105
timestamp 1679581782
transform 1 0 10656 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_112
timestamp 1679581782
transform 1 0 11328 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_119
timestamp 1679581782
transform 1 0 12000 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_126
timestamp 1679581782
transform 1 0 12672 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_133
timestamp 1679581782
transform 1 0 13344 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_140
timestamp 1679581782
transform 1 0 14016 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_147
timestamp 1679581782
transform 1 0 14688 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_154
timestamp 1679581782
transform 1 0 15360 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_161
timestamp 1679581782
transform 1 0 16032 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_168
timestamp 1679581782
transform 1 0 16704 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_175
timestamp 1679581782
transform 1 0 17376 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_182
timestamp 1679581782
transform 1 0 18048 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_189
timestamp 1679581782
transform 1 0 18720 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_196
timestamp 1679581782
transform 1 0 19392 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_203
timestamp 1679581782
transform 1 0 20064 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_210
timestamp 1679581782
transform 1 0 20736 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_217
timestamp 1679581782
transform 1 0 21408 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_224
timestamp 1679581782
transform 1 0 22080 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_231
timestamp 1679581782
transform 1 0 22752 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_238
timestamp 1679581782
transform 1 0 23424 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_245
timestamp 1679581782
transform 1 0 24096 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_252
timestamp 1679581782
transform 1 0 24768 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_259
timestamp 1679581782
transform 1 0 25440 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_266
timestamp 1679581782
transform 1 0 26112 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_273
timestamp 1679581782
transform 1 0 26784 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_280
timestamp 1679581782
transform 1 0 27456 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_287
timestamp 1679581782
transform 1 0 28128 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_294
timestamp 1679581782
transform 1 0 28800 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_301
timestamp 1679581782
transform 1 0 29472 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_308
timestamp 1679581782
transform 1 0 30144 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_315
timestamp 1679581782
transform 1 0 30816 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_322
timestamp 1679581782
transform 1 0 31488 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_329
timestamp 1679581782
transform 1 0 32160 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_336
timestamp 1679581782
transform 1 0 32832 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_343
timestamp 1679581782
transform 1 0 33504 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_350
timestamp 1679581782
transform 1 0 34176 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_357
timestamp 1679581782
transform 1 0 34848 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_364
timestamp 1679581782
transform 1 0 35520 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_371
timestamp 1679581782
transform 1 0 36192 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_378
timestamp 1679581782
transform 1 0 36864 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_385
timestamp 1679581782
transform 1 0 37536 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_392
timestamp 1679581782
transform 1 0 38208 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_399
timestamp 1679581782
transform 1 0 38880 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_406
timestamp 1679581782
transform 1 0 39552 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_413
timestamp 1679581782
transform 1 0 40224 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_420
timestamp 1679581782
transform 1 0 40896 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_427
timestamp 1679581782
transform 1 0 41568 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_434
timestamp 1679581782
transform 1 0 42240 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_441
timestamp 1679581782
transform 1 0 42912 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_448
timestamp 1679581782
transform 1 0 43584 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_455
timestamp 1679581782
transform 1 0 44256 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_462
timestamp 1679581782
transform 1 0 44928 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_469
timestamp 1679581782
transform 1 0 45600 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_476
timestamp 1679581782
transform 1 0 46272 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_483
timestamp 1679581782
transform 1 0 46944 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_490
timestamp 1679581782
transform 1 0 47616 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_497
timestamp 1679581782
transform 1 0 48288 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_504
timestamp 1679581782
transform 1 0 48960 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_511
timestamp 1679581782
transform 1 0 49632 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_518
timestamp 1679581782
transform 1 0 50304 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_525
timestamp 1679581782
transform 1 0 50976 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_532
timestamp 1679581782
transform 1 0 51648 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_539
timestamp 1679581782
transform 1 0 52320 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_546
timestamp 1679581782
transform 1 0 52992 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_553
timestamp 1679581782
transform 1 0 53664 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_560
timestamp 1679581782
transform 1 0 54336 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_567
timestamp 1679581782
transform 1 0 55008 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_574
timestamp 1679581782
transform 1 0 55680 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_581
timestamp 1679581782
transform 1 0 56352 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_588
timestamp 1679581782
transform 1 0 57024 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_595
timestamp 1679581782
transform 1 0 57696 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_602
timestamp 1679581782
transform 1 0 58368 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_609
timestamp 1679581782
transform 1 0 59040 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_616
timestamp 1679581782
transform 1 0 59712 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_623
timestamp 1679581782
transform 1 0 60384 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_630
timestamp 1679581782
transform 1 0 61056 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_637
timestamp 1679581782
transform 1 0 61728 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_644
timestamp 1679581782
transform 1 0 62400 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_651
timestamp 1679581782
transform 1 0 63072 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_658
timestamp 1679581782
transform 1 0 63744 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_665
timestamp 1679581782
transform 1 0 64416 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_672
timestamp 1679581782
transform 1 0 65088 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_679
timestamp 1679581782
transform 1 0 65760 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_686
timestamp 1679581782
transform 1 0 66432 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_693
timestamp 1679581782
transform 1 0 67104 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_700
timestamp 1679581782
transform 1 0 67776 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_707
timestamp 1679581782
transform 1 0 68448 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_714
timestamp 1679581782
transform 1 0 69120 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_721
timestamp 1679581782
transform 1 0 69792 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_728
timestamp 1679581782
transform 1 0 70464 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_735
timestamp 1679581782
transform 1 0 71136 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_742
timestamp 1679581782
transform 1 0 71808 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_749
timestamp 1679581782
transform 1 0 72480 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_756
timestamp 1679581782
transform 1 0 73152 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_763
timestamp 1679581782
transform 1 0 73824 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_770
timestamp 1679581782
transform 1 0 74496 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_777
timestamp 1679581782
transform 1 0 75168 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_784
timestamp 1679581782
transform 1 0 75840 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_791
timestamp 1679581782
transform 1 0 76512 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_798
timestamp 1679581782
transform 1 0 77184 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_805
timestamp 1679581782
transform 1 0 77856 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_812
timestamp 1679581782
transform 1 0 78528 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_819
timestamp 1679581782
transform 1 0 79200 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_826
timestamp 1679581782
transform 1 0 79872 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_833
timestamp 1679581782
transform 1 0 80544 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_840
timestamp 1679581782
transform 1 0 81216 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_847
timestamp 1679581782
transform 1 0 81888 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_854
timestamp 1679581782
transform 1 0 82560 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_861
timestamp 1679581782
transform 1 0 83232 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_868
timestamp 1679581782
transform 1 0 83904 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_875
timestamp 1679581782
transform 1 0 84576 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_882
timestamp 1679581782
transform 1 0 85248 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_889
timestamp 1679581782
transform 1 0 85920 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_896
timestamp 1679581782
transform 1 0 86592 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_903
timestamp 1679581782
transform 1 0 87264 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_910
timestamp 1679581782
transform 1 0 87936 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_917
timestamp 1679581782
transform 1 0 88608 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_924
timestamp 1679581782
transform 1 0 89280 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_931
timestamp 1679581782
transform 1 0 89952 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_938
timestamp 1679581782
transform 1 0 90624 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_945
timestamp 1679581782
transform 1 0 91296 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_952
timestamp 1679581782
transform 1 0 91968 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_959
timestamp 1679581782
transform 1 0 92640 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_966
timestamp 1679581782
transform 1 0 93312 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_973
timestamp 1679581782
transform 1 0 93984 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_980
timestamp 1679581782
transform 1 0 94656 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_987
timestamp 1679581782
transform 1 0 95328 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_994
timestamp 1679581782
transform 1 0 96000 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_1001
timestamp 1679581782
transform 1 0 96672 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_1008
timestamp 1679581782
transform 1 0 97344 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_1015
timestamp 1679581782
transform 1 0 98016 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_1022
timestamp 1679581782
transform 1 0 98688 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_0
timestamp 1679581782
transform 1 0 576 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_7
timestamp 1679581782
transform 1 0 1248 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_14
timestamp 1679581782
transform 1 0 1920 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_21
timestamp 1679581782
transform 1 0 2592 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_28
timestamp 1679581782
transform 1 0 3264 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_35
timestamp 1679581782
transform 1 0 3936 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_42
timestamp 1679581782
transform 1 0 4608 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_49
timestamp 1679581782
transform 1 0 5280 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_56
timestamp 1679581782
transform 1 0 5952 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_63
timestamp 1679581782
transform 1 0 6624 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_70
timestamp 1679581782
transform 1 0 7296 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_77
timestamp 1679581782
transform 1 0 7968 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_84
timestamp 1679581782
transform 1 0 8640 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_91
timestamp 1679581782
transform 1 0 9312 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_98
timestamp 1679581782
transform 1 0 9984 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_105
timestamp 1679581782
transform 1 0 10656 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_112
timestamp 1679581782
transform 1 0 11328 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_119
timestamp 1679581782
transform 1 0 12000 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_126
timestamp 1679581782
transform 1 0 12672 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_133
timestamp 1679581782
transform 1 0 13344 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_140
timestamp 1679581782
transform 1 0 14016 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_147
timestamp 1679581782
transform 1 0 14688 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_154
timestamp 1679581782
transform 1 0 15360 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_161
timestamp 1679581782
transform 1 0 16032 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_168
timestamp 1679581782
transform 1 0 16704 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_175
timestamp 1679581782
transform 1 0 17376 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_182
timestamp 1679581782
transform 1 0 18048 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_189
timestamp 1679581782
transform 1 0 18720 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_196
timestamp 1679581782
transform 1 0 19392 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_203
timestamp 1679581782
transform 1 0 20064 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_210
timestamp 1679581782
transform 1 0 20736 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_217
timestamp 1679581782
transform 1 0 21408 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_224
timestamp 1679581782
transform 1 0 22080 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_231
timestamp 1679581782
transform 1 0 22752 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_238
timestamp 1679581782
transform 1 0 23424 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_245
timestamp 1679581782
transform 1 0 24096 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_252
timestamp 1679581782
transform 1 0 24768 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_259
timestamp 1679581782
transform 1 0 25440 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_266
timestamp 1679581782
transform 1 0 26112 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_273
timestamp 1679581782
transform 1 0 26784 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_280
timestamp 1679581782
transform 1 0 27456 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_287
timestamp 1679581782
transform 1 0 28128 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_294
timestamp 1679581782
transform 1 0 28800 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_301
timestamp 1679581782
transform 1 0 29472 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_308
timestamp 1679581782
transform 1 0 30144 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_315
timestamp 1679581782
transform 1 0 30816 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_322
timestamp 1679581782
transform 1 0 31488 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_329
timestamp 1679581782
transform 1 0 32160 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_336
timestamp 1679581782
transform 1 0 32832 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_343
timestamp 1679581782
transform 1 0 33504 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_350
timestamp 1679581782
transform 1 0 34176 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_357
timestamp 1679581782
transform 1 0 34848 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_364
timestamp 1679581782
transform 1 0 35520 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_371
timestamp 1679581782
transform 1 0 36192 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_378
timestamp 1679581782
transform 1 0 36864 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_385
timestamp 1679581782
transform 1 0 37536 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_392
timestamp 1679581782
transform 1 0 38208 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_399
timestamp 1679581782
transform 1 0 38880 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_406
timestamp 1679581782
transform 1 0 39552 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_413
timestamp 1679581782
transform 1 0 40224 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_420
timestamp 1679581782
transform 1 0 40896 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_427
timestamp 1679581782
transform 1 0 41568 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_434
timestamp 1679581782
transform 1 0 42240 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_441
timestamp 1679581782
transform 1 0 42912 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_448
timestamp 1679581782
transform 1 0 43584 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_455
timestamp 1679581782
transform 1 0 44256 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_462
timestamp 1679581782
transform 1 0 44928 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_469
timestamp 1679581782
transform 1 0 45600 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_476
timestamp 1679581782
transform 1 0 46272 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_483
timestamp 1679581782
transform 1 0 46944 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_490
timestamp 1679581782
transform 1 0 47616 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_497
timestamp 1679581782
transform 1 0 48288 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_504
timestamp 1679581782
transform 1 0 48960 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_511
timestamp 1679581782
transform 1 0 49632 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_518
timestamp 1679581782
transform 1 0 50304 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_525
timestamp 1679581782
transform 1 0 50976 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_532
timestamp 1679581782
transform 1 0 51648 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_539
timestamp 1679581782
transform 1 0 52320 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_546
timestamp 1679581782
transform 1 0 52992 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_553
timestamp 1679581782
transform 1 0 53664 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_560
timestamp 1679581782
transform 1 0 54336 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_567
timestamp 1679581782
transform 1 0 55008 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_574
timestamp 1679581782
transform 1 0 55680 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_581
timestamp 1679581782
transform 1 0 56352 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_588
timestamp 1679581782
transform 1 0 57024 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_595
timestamp 1679581782
transform 1 0 57696 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_602
timestamp 1679581782
transform 1 0 58368 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_609
timestamp 1679581782
transform 1 0 59040 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_616
timestamp 1679581782
transform 1 0 59712 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_623
timestamp 1679581782
transform 1 0 60384 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_630
timestamp 1679581782
transform 1 0 61056 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_637
timestamp 1679581782
transform 1 0 61728 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_644
timestamp 1679581782
transform 1 0 62400 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_651
timestamp 1679581782
transform 1 0 63072 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_658
timestamp 1679581782
transform 1 0 63744 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_665
timestamp 1679581782
transform 1 0 64416 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_672
timestamp 1679581782
transform 1 0 65088 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_679
timestamp 1679581782
transform 1 0 65760 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_686
timestamp 1679581782
transform 1 0 66432 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_693
timestamp 1679581782
transform 1 0 67104 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_700
timestamp 1679581782
transform 1 0 67776 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_707
timestamp 1679581782
transform 1 0 68448 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_714
timestamp 1679581782
transform 1 0 69120 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_721
timestamp 1679581782
transform 1 0 69792 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_728
timestamp 1679581782
transform 1 0 70464 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_735
timestamp 1679581782
transform 1 0 71136 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_742
timestamp 1679581782
transform 1 0 71808 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_749
timestamp 1679581782
transform 1 0 72480 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_756
timestamp 1679581782
transform 1 0 73152 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_763
timestamp 1679581782
transform 1 0 73824 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_770
timestamp 1679581782
transform 1 0 74496 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_777
timestamp 1679581782
transform 1 0 75168 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_784
timestamp 1679581782
transform 1 0 75840 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_791
timestamp 1679581782
transform 1 0 76512 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_798
timestamp 1679581782
transform 1 0 77184 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_805
timestamp 1679581782
transform 1 0 77856 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_812
timestamp 1679581782
transform 1 0 78528 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_819
timestamp 1679581782
transform 1 0 79200 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_826
timestamp 1679581782
transform 1 0 79872 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_833
timestamp 1679581782
transform 1 0 80544 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_840
timestamp 1679581782
transform 1 0 81216 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_847
timestamp 1679581782
transform 1 0 81888 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_854
timestamp 1679581782
transform 1 0 82560 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_861
timestamp 1679581782
transform 1 0 83232 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_868
timestamp 1679581782
transform 1 0 83904 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_875
timestamp 1679581782
transform 1 0 84576 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_882
timestamp 1679581782
transform 1 0 85248 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_889
timestamp 1679581782
transform 1 0 85920 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_896
timestamp 1679581782
transform 1 0 86592 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_903
timestamp 1679581782
transform 1 0 87264 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_910
timestamp 1679581782
transform 1 0 87936 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_917
timestamp 1679581782
transform 1 0 88608 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_924
timestamp 1679581782
transform 1 0 89280 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_931
timestamp 1679581782
transform 1 0 89952 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_938
timestamp 1679581782
transform 1 0 90624 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_945
timestamp 1679581782
transform 1 0 91296 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_952
timestamp 1679581782
transform 1 0 91968 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_959
timestamp 1679581782
transform 1 0 92640 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_966
timestamp 1679581782
transform 1 0 93312 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_973
timestamp 1679581782
transform 1 0 93984 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_980
timestamp 1679581782
transform 1 0 94656 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_987
timestamp 1679581782
transform 1 0 95328 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_994
timestamp 1679581782
transform 1 0 96000 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1001
timestamp 1679581782
transform 1 0 96672 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1008
timestamp 1679581782
transform 1 0 97344 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1015
timestamp 1679581782
transform 1 0 98016 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1022
timestamp 1679581782
transform 1 0 98688 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_4
timestamp 1679581782
transform 1 0 960 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_11
timestamp 1679581782
transform 1 0 1632 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_18
timestamp 1679581782
transform 1 0 2304 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_25
timestamp 1679581782
transform 1 0 2976 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_32
timestamp 1679581782
transform 1 0 3648 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_39
timestamp 1679581782
transform 1 0 4320 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_46
timestamp 1679581782
transform 1 0 4992 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_53
timestamp 1679581782
transform 1 0 5664 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_60
timestamp 1679581782
transform 1 0 6336 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_67
timestamp 1679581782
transform 1 0 7008 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_74
timestamp 1679581782
transform 1 0 7680 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_81
timestamp 1679581782
transform 1 0 8352 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_88
timestamp 1679581782
transform 1 0 9024 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_95
timestamp 1679581782
transform 1 0 9696 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_102
timestamp 1679581782
transform 1 0 10368 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_109
timestamp 1679581782
transform 1 0 11040 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_116
timestamp 1679581782
transform 1 0 11712 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_123
timestamp 1679581782
transform 1 0 12384 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_130
timestamp 1679581782
transform 1 0 13056 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_137
timestamp 1679581782
transform 1 0 13728 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_144
timestamp 1679581782
transform 1 0 14400 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_151
timestamp 1679581782
transform 1 0 15072 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_158
timestamp 1679581782
transform 1 0 15744 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_165
timestamp 1679581782
transform 1 0 16416 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_172
timestamp 1679581782
transform 1 0 17088 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_179
timestamp 1679581782
transform 1 0 17760 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_186
timestamp 1679581782
transform 1 0 18432 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_193
timestamp 1679581782
transform 1 0 19104 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_200
timestamp 1679581782
transform 1 0 19776 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_207
timestamp 1679581782
transform 1 0 20448 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_214
timestamp 1679581782
transform 1 0 21120 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_221
timestamp 1679581782
transform 1 0 21792 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_228
timestamp 1679581782
transform 1 0 22464 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_235
timestamp 1679581782
transform 1 0 23136 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_242
timestamp 1679581782
transform 1 0 23808 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_249
timestamp 1679581782
transform 1 0 24480 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_256
timestamp 1679581782
transform 1 0 25152 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_263
timestamp 1679581782
transform 1 0 25824 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_270
timestamp 1679581782
transform 1 0 26496 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_277
timestamp 1679581782
transform 1 0 27168 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_284
timestamp 1679581782
transform 1 0 27840 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_291
timestamp 1679581782
transform 1 0 28512 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_298
timestamp 1679581782
transform 1 0 29184 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_305
timestamp 1679581782
transform 1 0 29856 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_312
timestamp 1679581782
transform 1 0 30528 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_319
timestamp 1679581782
transform 1 0 31200 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_326
timestamp 1679581782
transform 1 0 31872 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_333
timestamp 1679581782
transform 1 0 32544 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_340
timestamp 1679581782
transform 1 0 33216 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_347
timestamp 1679581782
transform 1 0 33888 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_354
timestamp 1679581782
transform 1 0 34560 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_361
timestamp 1679581782
transform 1 0 35232 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_368
timestamp 1679581782
transform 1 0 35904 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_375
timestamp 1679581782
transform 1 0 36576 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_382
timestamp 1679581782
transform 1 0 37248 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_389
timestamp 1679581782
transform 1 0 37920 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_396
timestamp 1679581782
transform 1 0 38592 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_403
timestamp 1679581782
transform 1 0 39264 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_410
timestamp 1679581782
transform 1 0 39936 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_417
timestamp 1679581782
transform 1 0 40608 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_424
timestamp 1679581782
transform 1 0 41280 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_431
timestamp 1679581782
transform 1 0 41952 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_438
timestamp 1679581782
transform 1 0 42624 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_445
timestamp 1679581782
transform 1 0 43296 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_452
timestamp 1679581782
transform 1 0 43968 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_459
timestamp 1679581782
transform 1 0 44640 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_466
timestamp 1679581782
transform 1 0 45312 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_473
timestamp 1679581782
transform 1 0 45984 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_480
timestamp 1679581782
transform 1 0 46656 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_487
timestamp 1679581782
transform 1 0 47328 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_494
timestamp 1679581782
transform 1 0 48000 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_501
timestamp 1679581782
transform 1 0 48672 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_508
timestamp 1679581782
transform 1 0 49344 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_515
timestamp 1679581782
transform 1 0 50016 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_522
timestamp 1679581782
transform 1 0 50688 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_529
timestamp 1679581782
transform 1 0 51360 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_536
timestamp 1679581782
transform 1 0 52032 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_543
timestamp 1679581782
transform 1 0 52704 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_550
timestamp 1679581782
transform 1 0 53376 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_557
timestamp 1679581782
transform 1 0 54048 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_564
timestamp 1679581782
transform 1 0 54720 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_571
timestamp 1679581782
transform 1 0 55392 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_578
timestamp 1679581782
transform 1 0 56064 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_585
timestamp 1679581782
transform 1 0 56736 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_592
timestamp 1679581782
transform 1 0 57408 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_599
timestamp 1679581782
transform 1 0 58080 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_606
timestamp 1679581782
transform 1 0 58752 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_613
timestamp 1679581782
transform 1 0 59424 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_620
timestamp 1679581782
transform 1 0 60096 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_627
timestamp 1679581782
transform 1 0 60768 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_634
timestamp 1679581782
transform 1 0 61440 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_641
timestamp 1679581782
transform 1 0 62112 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_648
timestamp 1679581782
transform 1 0 62784 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_655
timestamp 1679581782
transform 1 0 63456 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_662
timestamp 1679581782
transform 1 0 64128 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_669
timestamp 1679581782
transform 1 0 64800 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_676
timestamp 1679581782
transform 1 0 65472 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_683
timestamp 1679581782
transform 1 0 66144 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_690
timestamp 1679581782
transform 1 0 66816 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_697
timestamp 1679581782
transform 1 0 67488 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_704
timestamp 1679581782
transform 1 0 68160 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_711
timestamp 1679581782
transform 1 0 68832 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_718
timestamp 1679581782
transform 1 0 69504 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_725
timestamp 1679581782
transform 1 0 70176 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_732
timestamp 1679581782
transform 1 0 70848 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_739
timestamp 1679581782
transform 1 0 71520 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_746
timestamp 1679581782
transform 1 0 72192 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_753
timestamp 1679581782
transform 1 0 72864 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_760
timestamp 1679581782
transform 1 0 73536 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_767
timestamp 1679581782
transform 1 0 74208 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_774
timestamp 1679581782
transform 1 0 74880 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_781
timestamp 1679581782
transform 1 0 75552 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_788
timestamp 1679581782
transform 1 0 76224 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_795
timestamp 1679581782
transform 1 0 76896 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_802
timestamp 1679581782
transform 1 0 77568 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_809
timestamp 1679581782
transform 1 0 78240 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_816
timestamp 1679581782
transform 1 0 78912 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_823
timestamp 1679581782
transform 1 0 79584 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_830
timestamp 1679581782
transform 1 0 80256 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_837
timestamp 1679581782
transform 1 0 80928 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_844
timestamp 1679581782
transform 1 0 81600 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_851
timestamp 1679581782
transform 1 0 82272 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_858
timestamp 1679581782
transform 1 0 82944 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_865
timestamp 1679581782
transform 1 0 83616 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_872
timestamp 1679581782
transform 1 0 84288 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_879
timestamp 1679581782
transform 1 0 84960 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_886
timestamp 1679581782
transform 1 0 85632 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_893
timestamp 1679581782
transform 1 0 86304 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_900
timestamp 1679581782
transform 1 0 86976 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_907
timestamp 1679581782
transform 1 0 87648 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_914
timestamp 1679581782
transform 1 0 88320 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_921
timestamp 1679581782
transform 1 0 88992 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_928
timestamp 1679581782
transform 1 0 89664 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_935
timestamp 1679581782
transform 1 0 90336 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_942
timestamp 1679581782
transform 1 0 91008 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_949
timestamp 1679581782
transform 1 0 91680 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_956
timestamp 1679581782
transform 1 0 92352 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_963
timestamp 1679581782
transform 1 0 93024 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_970
timestamp 1679581782
transform 1 0 93696 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_977
timestamp 1679581782
transform 1 0 94368 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_984
timestamp 1679581782
transform 1 0 95040 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_991
timestamp 1679581782
transform 1 0 95712 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_998
timestamp 1679581782
transform 1 0 96384 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1005
timestamp 1679581782
transform 1 0 97056 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1012
timestamp 1679581782
transform 1 0 97728 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1019
timestamp 1679581782
transform 1 0 98400 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_27_1026
timestamp 1677580104
transform 1 0 99072 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_1028
timestamp 1677579658
transform 1 0 99264 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_0
timestamp 1679581782
transform 1 0 576 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_7
timestamp 1679581782
transform 1 0 1248 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_14
timestamp 1679581782
transform 1 0 1920 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_21
timestamp 1679581782
transform 1 0 2592 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_28
timestamp 1679581782
transform 1 0 3264 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_35
timestamp 1679581782
transform 1 0 3936 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_42
timestamp 1679581782
transform 1 0 4608 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_49
timestamp 1679581782
transform 1 0 5280 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_56
timestamp 1679581782
transform 1 0 5952 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_63
timestamp 1679581782
transform 1 0 6624 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_70
timestamp 1679581782
transform 1 0 7296 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_77
timestamp 1679581782
transform 1 0 7968 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_84
timestamp 1679581782
transform 1 0 8640 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_91
timestamp 1679581782
transform 1 0 9312 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_98
timestamp 1679581782
transform 1 0 9984 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_105
timestamp 1679581782
transform 1 0 10656 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_112
timestamp 1679581782
transform 1 0 11328 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_119
timestamp 1679581782
transform 1 0 12000 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_126
timestamp 1679581782
transform 1 0 12672 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_133
timestamp 1679581782
transform 1 0 13344 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_140
timestamp 1679581782
transform 1 0 14016 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_147
timestamp 1679581782
transform 1 0 14688 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_154
timestamp 1679581782
transform 1 0 15360 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_161
timestamp 1679581782
transform 1 0 16032 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_168
timestamp 1679581782
transform 1 0 16704 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_175
timestamp 1679581782
transform 1 0 17376 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_182
timestamp 1679581782
transform 1 0 18048 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_189
timestamp 1679581782
transform 1 0 18720 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_196
timestamp 1679581782
transform 1 0 19392 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_203
timestamp 1679581782
transform 1 0 20064 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_210
timestamp 1679581782
transform 1 0 20736 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_217
timestamp 1679581782
transform 1 0 21408 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_224
timestamp 1679581782
transform 1 0 22080 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_231
timestamp 1679581782
transform 1 0 22752 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_238
timestamp 1679581782
transform 1 0 23424 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_245
timestamp 1679581782
transform 1 0 24096 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_252
timestamp 1679581782
transform 1 0 24768 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_259
timestamp 1679581782
transform 1 0 25440 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_266
timestamp 1679581782
transform 1 0 26112 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_273
timestamp 1679581782
transform 1 0 26784 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_280
timestamp 1679581782
transform 1 0 27456 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_287
timestamp 1679581782
transform 1 0 28128 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_294
timestamp 1679581782
transform 1 0 28800 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_301
timestamp 1679581782
transform 1 0 29472 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_308
timestamp 1679581782
transform 1 0 30144 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_315
timestamp 1679581782
transform 1 0 30816 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_322
timestamp 1679581782
transform 1 0 31488 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_329
timestamp 1679581782
transform 1 0 32160 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_336
timestamp 1679581782
transform 1 0 32832 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_343
timestamp 1679581782
transform 1 0 33504 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_350
timestamp 1679581782
transform 1 0 34176 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_357
timestamp 1679581782
transform 1 0 34848 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_364
timestamp 1679581782
transform 1 0 35520 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_371
timestamp 1679581782
transform 1 0 36192 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_378
timestamp 1679581782
transform 1 0 36864 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_385
timestamp 1679581782
transform 1 0 37536 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_392
timestamp 1679581782
transform 1 0 38208 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_399
timestamp 1679581782
transform 1 0 38880 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_406
timestamp 1679581782
transform 1 0 39552 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_413
timestamp 1679581782
transform 1 0 40224 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_420
timestamp 1679581782
transform 1 0 40896 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_427
timestamp 1679581782
transform 1 0 41568 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_434
timestamp 1679581782
transform 1 0 42240 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_441
timestamp 1679581782
transform 1 0 42912 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_448
timestamp 1679581782
transform 1 0 43584 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_455
timestamp 1679581782
transform 1 0 44256 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_462
timestamp 1679581782
transform 1 0 44928 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_469
timestamp 1679581782
transform 1 0 45600 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_476
timestamp 1679581782
transform 1 0 46272 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_483
timestamp 1679581782
transform 1 0 46944 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_490
timestamp 1679581782
transform 1 0 47616 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_497
timestamp 1679581782
transform 1 0 48288 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_504
timestamp 1679581782
transform 1 0 48960 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_511
timestamp 1679581782
transform 1 0 49632 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_518
timestamp 1679581782
transform 1 0 50304 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_525
timestamp 1679581782
transform 1 0 50976 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_532
timestamp 1679581782
transform 1 0 51648 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_539
timestamp 1679581782
transform 1 0 52320 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_546
timestamp 1679581782
transform 1 0 52992 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_553
timestamp 1679581782
transform 1 0 53664 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_560
timestamp 1679581782
transform 1 0 54336 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_567
timestamp 1679581782
transform 1 0 55008 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_574
timestamp 1679581782
transform 1 0 55680 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_581
timestamp 1679581782
transform 1 0 56352 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_588
timestamp 1679581782
transform 1 0 57024 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_595
timestamp 1679581782
transform 1 0 57696 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_602
timestamp 1679581782
transform 1 0 58368 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_609
timestamp 1679581782
transform 1 0 59040 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_616
timestamp 1679581782
transform 1 0 59712 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_623
timestamp 1679581782
transform 1 0 60384 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_630
timestamp 1679581782
transform 1 0 61056 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_637
timestamp 1679581782
transform 1 0 61728 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_644
timestamp 1679581782
transform 1 0 62400 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_651
timestamp 1679581782
transform 1 0 63072 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_658
timestamp 1679581782
transform 1 0 63744 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_665
timestamp 1679581782
transform 1 0 64416 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_672
timestamp 1679581782
transform 1 0 65088 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_679
timestamp 1679581782
transform 1 0 65760 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_686
timestamp 1679581782
transform 1 0 66432 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_693
timestamp 1679581782
transform 1 0 67104 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_700
timestamp 1679581782
transform 1 0 67776 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_707
timestamp 1679581782
transform 1 0 68448 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_714
timestamp 1679581782
transform 1 0 69120 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_721
timestamp 1679581782
transform 1 0 69792 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_728
timestamp 1679581782
transform 1 0 70464 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_735
timestamp 1679581782
transform 1 0 71136 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_742
timestamp 1679581782
transform 1 0 71808 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_749
timestamp 1679581782
transform 1 0 72480 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_756
timestamp 1679581782
transform 1 0 73152 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_763
timestamp 1679581782
transform 1 0 73824 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_770
timestamp 1679581782
transform 1 0 74496 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_777
timestamp 1679581782
transform 1 0 75168 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_784
timestamp 1679581782
transform 1 0 75840 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_791
timestamp 1679581782
transform 1 0 76512 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_798
timestamp 1679581782
transform 1 0 77184 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_805
timestamp 1679581782
transform 1 0 77856 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_812
timestamp 1679581782
transform 1 0 78528 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_819
timestamp 1679581782
transform 1 0 79200 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_826
timestamp 1679581782
transform 1 0 79872 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_833
timestamp 1679581782
transform 1 0 80544 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_840
timestamp 1679581782
transform 1 0 81216 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_847
timestamp 1679581782
transform 1 0 81888 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_854
timestamp 1679581782
transform 1 0 82560 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_861
timestamp 1679581782
transform 1 0 83232 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_868
timestamp 1679581782
transform 1 0 83904 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_875
timestamp 1679581782
transform 1 0 84576 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_882
timestamp 1679581782
transform 1 0 85248 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_889
timestamp 1679581782
transform 1 0 85920 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_896
timestamp 1679581782
transform 1 0 86592 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_903
timestamp 1679581782
transform 1 0 87264 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_910
timestamp 1679581782
transform 1 0 87936 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_917
timestamp 1679581782
transform 1 0 88608 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_924
timestamp 1679581782
transform 1 0 89280 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_931
timestamp 1679581782
transform 1 0 89952 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_938
timestamp 1679581782
transform 1 0 90624 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_945
timestamp 1679581782
transform 1 0 91296 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_952
timestamp 1679581782
transform 1 0 91968 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_959
timestamp 1679581782
transform 1 0 92640 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_966
timestamp 1679581782
transform 1 0 93312 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_973
timestamp 1679581782
transform 1 0 93984 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_980
timestamp 1679581782
transform 1 0 94656 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_987
timestamp 1679581782
transform 1 0 95328 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_994
timestamp 1679581782
transform 1 0 96000 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_1001
timestamp 1679581782
transform 1 0 96672 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_1008
timestamp 1679581782
transform 1 0 97344 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_1015
timestamp 1679581782
transform 1 0 98016 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_1022
timestamp 1679581782
transform 1 0 98688 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_4
timestamp 1679581782
transform 1 0 960 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_11
timestamp 1679581782
transform 1 0 1632 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_18
timestamp 1679581782
transform 1 0 2304 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_25
timestamp 1679581782
transform 1 0 2976 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_32
timestamp 1679581782
transform 1 0 3648 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_39
timestamp 1679581782
transform 1 0 4320 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_46
timestamp 1679581782
transform 1 0 4992 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_53
timestamp 1679581782
transform 1 0 5664 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_60
timestamp 1679581782
transform 1 0 6336 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_67
timestamp 1679581782
transform 1 0 7008 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_74
timestamp 1679581782
transform 1 0 7680 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_81
timestamp 1679581782
transform 1 0 8352 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_88
timestamp 1679581782
transform 1 0 9024 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_95
timestamp 1679581782
transform 1 0 9696 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_102
timestamp 1679581782
transform 1 0 10368 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_109
timestamp 1679581782
transform 1 0 11040 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_116
timestamp 1679581782
transform 1 0 11712 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_123
timestamp 1679581782
transform 1 0 12384 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_130
timestamp 1679581782
transform 1 0 13056 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_137
timestamp 1679581782
transform 1 0 13728 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_144
timestamp 1679581782
transform 1 0 14400 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_151
timestamp 1679581782
transform 1 0 15072 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_158
timestamp 1679581782
transform 1 0 15744 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_165
timestamp 1679581782
transform 1 0 16416 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_172
timestamp 1679581782
transform 1 0 17088 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_179
timestamp 1679581782
transform 1 0 17760 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_186
timestamp 1679581782
transform 1 0 18432 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_193
timestamp 1679581782
transform 1 0 19104 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_200
timestamp 1679581782
transform 1 0 19776 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_207
timestamp 1679581782
transform 1 0 20448 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_214
timestamp 1679581782
transform 1 0 21120 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_221
timestamp 1679581782
transform 1 0 21792 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_228
timestamp 1679581782
transform 1 0 22464 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_235
timestamp 1679581782
transform 1 0 23136 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_242
timestamp 1679581782
transform 1 0 23808 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_249
timestamp 1679581782
transform 1 0 24480 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_256
timestamp 1679581782
transform 1 0 25152 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_263
timestamp 1679581782
transform 1 0 25824 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_270
timestamp 1679581782
transform 1 0 26496 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_277
timestamp 1679581782
transform 1 0 27168 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_284
timestamp 1679581782
transform 1 0 27840 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_291
timestamp 1679581782
transform 1 0 28512 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_298
timestamp 1679581782
transform 1 0 29184 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_305
timestamp 1679581782
transform 1 0 29856 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_312
timestamp 1679581782
transform 1 0 30528 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_319
timestamp 1679581782
transform 1 0 31200 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_326
timestamp 1679581782
transform 1 0 31872 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_333
timestamp 1679581782
transform 1 0 32544 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_340
timestamp 1679581782
transform 1 0 33216 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_347
timestamp 1679581782
transform 1 0 33888 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_354
timestamp 1679581782
transform 1 0 34560 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_361
timestamp 1679581782
transform 1 0 35232 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_368
timestamp 1679581782
transform 1 0 35904 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_375
timestamp 1679581782
transform 1 0 36576 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_382
timestamp 1679581782
transform 1 0 37248 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_389
timestamp 1679581782
transform 1 0 37920 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_396
timestamp 1679581782
transform 1 0 38592 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_403
timestamp 1679581782
transform 1 0 39264 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_410
timestamp 1679581782
transform 1 0 39936 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_417
timestamp 1679581782
transform 1 0 40608 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_424
timestamp 1679581782
transform 1 0 41280 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_431
timestamp 1679581782
transform 1 0 41952 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_438
timestamp 1679581782
transform 1 0 42624 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_445
timestamp 1679581782
transform 1 0 43296 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_452
timestamp 1679581782
transform 1 0 43968 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_459
timestamp 1679581782
transform 1 0 44640 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_466
timestamp 1679581782
transform 1 0 45312 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_473
timestamp 1679581782
transform 1 0 45984 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_480
timestamp 1679581782
transform 1 0 46656 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_487
timestamp 1679581782
transform 1 0 47328 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_494
timestamp 1679581782
transform 1 0 48000 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_501
timestamp 1679581782
transform 1 0 48672 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_508
timestamp 1679581782
transform 1 0 49344 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_515
timestamp 1679581782
transform 1 0 50016 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_522
timestamp 1679581782
transform 1 0 50688 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_529
timestamp 1679581782
transform 1 0 51360 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_536
timestamp 1679581782
transform 1 0 52032 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_543
timestamp 1679581782
transform 1 0 52704 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_550
timestamp 1679581782
transform 1 0 53376 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_557
timestamp 1679581782
transform 1 0 54048 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_564
timestamp 1679581782
transform 1 0 54720 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_571
timestamp 1679581782
transform 1 0 55392 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_578
timestamp 1679581782
transform 1 0 56064 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_585
timestamp 1679581782
transform 1 0 56736 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_592
timestamp 1679581782
transform 1 0 57408 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_599
timestamp 1679581782
transform 1 0 58080 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_606
timestamp 1679581782
transform 1 0 58752 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_613
timestamp 1679581782
transform 1 0 59424 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_620
timestamp 1679581782
transform 1 0 60096 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_627
timestamp 1679581782
transform 1 0 60768 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_634
timestamp 1679581782
transform 1 0 61440 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_641
timestamp 1679581782
transform 1 0 62112 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_648
timestamp 1679581782
transform 1 0 62784 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_655
timestamp 1679581782
transform 1 0 63456 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_662
timestamp 1679581782
transform 1 0 64128 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_669
timestamp 1679581782
transform 1 0 64800 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_676
timestamp 1679581782
transform 1 0 65472 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_683
timestamp 1679581782
transform 1 0 66144 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_690
timestamp 1679581782
transform 1 0 66816 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_697
timestamp 1679581782
transform 1 0 67488 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_704
timestamp 1679581782
transform 1 0 68160 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_711
timestamp 1679581782
transform 1 0 68832 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_718
timestamp 1679581782
transform 1 0 69504 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_725
timestamp 1679581782
transform 1 0 70176 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_732
timestamp 1679581782
transform 1 0 70848 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_739
timestamp 1679581782
transform 1 0 71520 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_746
timestamp 1679581782
transform 1 0 72192 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_753
timestamp 1679581782
transform 1 0 72864 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_760
timestamp 1679581782
transform 1 0 73536 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_767
timestamp 1679581782
transform 1 0 74208 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_774
timestamp 1679581782
transform 1 0 74880 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_781
timestamp 1679581782
transform 1 0 75552 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_788
timestamp 1679581782
transform 1 0 76224 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_795
timestamp 1679581782
transform 1 0 76896 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_802
timestamp 1679581782
transform 1 0 77568 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_809
timestamp 1679581782
transform 1 0 78240 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_816
timestamp 1679581782
transform 1 0 78912 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_823
timestamp 1679581782
transform 1 0 79584 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_830
timestamp 1679581782
transform 1 0 80256 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_837
timestamp 1679581782
transform 1 0 80928 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_844
timestamp 1679581782
transform 1 0 81600 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_851
timestamp 1679581782
transform 1 0 82272 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_858
timestamp 1679581782
transform 1 0 82944 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_865
timestamp 1679581782
transform 1 0 83616 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_872
timestamp 1679581782
transform 1 0 84288 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_879
timestamp 1679581782
transform 1 0 84960 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_886
timestamp 1679581782
transform 1 0 85632 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_893
timestamp 1679581782
transform 1 0 86304 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_900
timestamp 1679581782
transform 1 0 86976 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_907
timestamp 1679581782
transform 1 0 87648 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_914
timestamp 1679581782
transform 1 0 88320 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_921
timestamp 1679581782
transform 1 0 88992 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_928
timestamp 1679581782
transform 1 0 89664 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_935
timestamp 1679581782
transform 1 0 90336 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_942
timestamp 1679581782
transform 1 0 91008 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_949
timestamp 1679581782
transform 1 0 91680 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_956
timestamp 1679581782
transform 1 0 92352 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_963
timestamp 1679581782
transform 1 0 93024 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_970
timestamp 1679581782
transform 1 0 93696 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_977
timestamp 1679581782
transform 1 0 94368 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_984
timestamp 1679581782
transform 1 0 95040 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_991
timestamp 1679581782
transform 1 0 95712 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_998
timestamp 1679581782
transform 1 0 96384 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_1005
timestamp 1679581782
transform 1 0 97056 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_1012
timestamp 1679581782
transform 1 0 97728 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_1019
timestamp 1679581782
transform 1 0 98400 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_29_1026
timestamp 1677580104
transform 1 0 99072 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_1028
timestamp 1677579658
transform 1 0 99264 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_0
timestamp 1679581782
transform 1 0 576 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_7
timestamp 1679581782
transform 1 0 1248 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_14
timestamp 1679581782
transform 1 0 1920 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_21
timestamp 1679581782
transform 1 0 2592 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_28
timestamp 1679581782
transform 1 0 3264 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_35
timestamp 1679581782
transform 1 0 3936 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_42
timestamp 1679581782
transform 1 0 4608 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_49
timestamp 1679581782
transform 1 0 5280 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_56
timestamp 1679581782
transform 1 0 5952 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_63
timestamp 1679581782
transform 1 0 6624 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_70
timestamp 1679581782
transform 1 0 7296 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_77
timestamp 1679581782
transform 1 0 7968 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_84
timestamp 1679581782
transform 1 0 8640 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_91
timestamp 1679581782
transform 1 0 9312 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_98
timestamp 1679581782
transform 1 0 9984 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_105
timestamp 1679581782
transform 1 0 10656 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_112
timestamp 1679581782
transform 1 0 11328 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_119
timestamp 1679581782
transform 1 0 12000 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_126
timestamp 1679581782
transform 1 0 12672 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_133
timestamp 1679581782
transform 1 0 13344 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_140
timestamp 1679581782
transform 1 0 14016 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_147
timestamp 1679581782
transform 1 0 14688 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_154
timestamp 1679581782
transform 1 0 15360 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_161
timestamp 1679581782
transform 1 0 16032 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_168
timestamp 1679581782
transform 1 0 16704 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_175
timestamp 1679581782
transform 1 0 17376 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_182
timestamp 1679581782
transform 1 0 18048 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_189
timestamp 1679581782
transform 1 0 18720 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_196
timestamp 1679581782
transform 1 0 19392 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_203
timestamp 1679581782
transform 1 0 20064 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_210
timestamp 1679581782
transform 1 0 20736 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_217
timestamp 1679581782
transform 1 0 21408 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_224
timestamp 1679581782
transform 1 0 22080 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_231
timestamp 1679581782
transform 1 0 22752 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_238
timestamp 1679581782
transform 1 0 23424 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_245
timestamp 1679581782
transform 1 0 24096 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_252
timestamp 1679581782
transform 1 0 24768 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_259
timestamp 1679581782
transform 1 0 25440 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_266
timestamp 1679581782
transform 1 0 26112 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_273
timestamp 1679581782
transform 1 0 26784 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_280
timestamp 1679581782
transform 1 0 27456 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_287
timestamp 1679581782
transform 1 0 28128 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_294
timestamp 1679581782
transform 1 0 28800 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_301
timestamp 1679581782
transform 1 0 29472 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_308
timestamp 1679581782
transform 1 0 30144 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_315
timestamp 1679581782
transform 1 0 30816 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_322
timestamp 1679581782
transform 1 0 31488 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_329
timestamp 1679581782
transform 1 0 32160 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_336
timestamp 1679581782
transform 1 0 32832 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_343
timestamp 1679581782
transform 1 0 33504 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_350
timestamp 1679581782
transform 1 0 34176 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_357
timestamp 1679581782
transform 1 0 34848 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_364
timestamp 1679581782
transform 1 0 35520 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_371
timestamp 1679581782
transform 1 0 36192 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_378
timestamp 1679581782
transform 1 0 36864 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_385
timestamp 1679581782
transform 1 0 37536 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_392
timestamp 1679581782
transform 1 0 38208 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_399
timestamp 1679581782
transform 1 0 38880 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_406
timestamp 1679581782
transform 1 0 39552 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_413
timestamp 1679581782
transform 1 0 40224 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_420
timestamp 1679581782
transform 1 0 40896 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_427
timestamp 1679581782
transform 1 0 41568 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_434
timestamp 1679581782
transform 1 0 42240 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_441
timestamp 1679581782
transform 1 0 42912 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_448
timestamp 1679581782
transform 1 0 43584 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_455
timestamp 1679581782
transform 1 0 44256 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_462
timestamp 1679581782
transform 1 0 44928 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_469
timestamp 1679581782
transform 1 0 45600 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_476
timestamp 1679581782
transform 1 0 46272 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_483
timestamp 1679581782
transform 1 0 46944 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_490
timestamp 1679581782
transform 1 0 47616 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_497
timestamp 1679581782
transform 1 0 48288 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_504
timestamp 1679581782
transform 1 0 48960 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_511
timestamp 1679581782
transform 1 0 49632 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_518
timestamp 1679581782
transform 1 0 50304 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_525
timestamp 1679581782
transform 1 0 50976 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_532
timestamp 1679581782
transform 1 0 51648 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_539
timestamp 1679581782
transform 1 0 52320 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_546
timestamp 1679581782
transform 1 0 52992 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_553
timestamp 1679581782
transform 1 0 53664 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_560
timestamp 1679581782
transform 1 0 54336 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_567
timestamp 1679581782
transform 1 0 55008 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_574
timestamp 1679581782
transform 1 0 55680 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_581
timestamp 1679581782
transform 1 0 56352 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_588
timestamp 1679581782
transform 1 0 57024 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_595
timestamp 1679581782
transform 1 0 57696 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_602
timestamp 1679581782
transform 1 0 58368 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_609
timestamp 1679581782
transform 1 0 59040 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_616
timestamp 1679581782
transform 1 0 59712 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_623
timestamp 1679581782
transform 1 0 60384 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_630
timestamp 1679581782
transform 1 0 61056 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_637
timestamp 1679581782
transform 1 0 61728 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_644
timestamp 1679581782
transform 1 0 62400 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_651
timestamp 1679581782
transform 1 0 63072 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_658
timestamp 1679581782
transform 1 0 63744 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_665
timestamp 1679581782
transform 1 0 64416 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_672
timestamp 1679581782
transform 1 0 65088 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_679
timestamp 1679581782
transform 1 0 65760 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_686
timestamp 1679581782
transform 1 0 66432 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_693
timestamp 1679581782
transform 1 0 67104 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_700
timestamp 1679581782
transform 1 0 67776 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_707
timestamp 1679581782
transform 1 0 68448 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_714
timestamp 1679581782
transform 1 0 69120 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_721
timestamp 1679581782
transform 1 0 69792 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_728
timestamp 1679581782
transform 1 0 70464 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_735
timestamp 1679581782
transform 1 0 71136 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_742
timestamp 1679581782
transform 1 0 71808 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_749
timestamp 1679581782
transform 1 0 72480 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_756
timestamp 1679581782
transform 1 0 73152 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_763
timestamp 1679581782
transform 1 0 73824 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_770
timestamp 1679581782
transform 1 0 74496 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_777
timestamp 1679581782
transform 1 0 75168 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_784
timestamp 1679581782
transform 1 0 75840 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_791
timestamp 1679581782
transform 1 0 76512 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_798
timestamp 1679581782
transform 1 0 77184 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_805
timestamp 1679581782
transform 1 0 77856 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_812
timestamp 1679581782
transform 1 0 78528 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_819
timestamp 1679581782
transform 1 0 79200 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_826
timestamp 1679581782
transform 1 0 79872 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_833
timestamp 1679581782
transform 1 0 80544 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_840
timestamp 1679581782
transform 1 0 81216 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_847
timestamp 1679581782
transform 1 0 81888 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_854
timestamp 1679581782
transform 1 0 82560 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_861
timestamp 1679581782
transform 1 0 83232 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_868
timestamp 1679581782
transform 1 0 83904 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_875
timestamp 1679581782
transform 1 0 84576 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_882
timestamp 1679581782
transform 1 0 85248 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_889
timestamp 1679581782
transform 1 0 85920 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_896
timestamp 1679581782
transform 1 0 86592 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_903
timestamp 1679581782
transform 1 0 87264 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_910
timestamp 1679581782
transform 1 0 87936 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_917
timestamp 1679581782
transform 1 0 88608 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_924
timestamp 1679581782
transform 1 0 89280 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_931
timestamp 1679581782
transform 1 0 89952 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_938
timestamp 1679581782
transform 1 0 90624 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_945
timestamp 1679581782
transform 1 0 91296 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_952
timestamp 1679581782
transform 1 0 91968 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_959
timestamp 1679581782
transform 1 0 92640 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_966
timestamp 1679581782
transform 1 0 93312 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_973
timestamp 1679581782
transform 1 0 93984 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_980
timestamp 1679581782
transform 1 0 94656 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_987
timestamp 1679581782
transform 1 0 95328 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_994
timestamp 1679581782
transform 1 0 96000 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_1001
timestamp 1679581782
transform 1 0 96672 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_1008
timestamp 1679581782
transform 1 0 97344 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_1015
timestamp 1679581782
transform 1 0 98016 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_1022
timestamp 1679581782
transform 1 0 98688 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_0
timestamp 1679581782
transform 1 0 576 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_7
timestamp 1679581782
transform 1 0 1248 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_14
timestamp 1679581782
transform 1 0 1920 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_21
timestamp 1679581782
transform 1 0 2592 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_28
timestamp 1679581782
transform 1 0 3264 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_35
timestamp 1679581782
transform 1 0 3936 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_42
timestamp 1679581782
transform 1 0 4608 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_49
timestamp 1679581782
transform 1 0 5280 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_56
timestamp 1679581782
transform 1 0 5952 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_63
timestamp 1679581782
transform 1 0 6624 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_70
timestamp 1679581782
transform 1 0 7296 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_77
timestamp 1679581782
transform 1 0 7968 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_84
timestamp 1679581782
transform 1 0 8640 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_91
timestamp 1679581782
transform 1 0 9312 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_98
timestamp 1679581782
transform 1 0 9984 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_105
timestamp 1679581782
transform 1 0 10656 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_112
timestamp 1679581782
transform 1 0 11328 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_119
timestamp 1679581782
transform 1 0 12000 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_126
timestamp 1679581782
transform 1 0 12672 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_133
timestamp 1679581782
transform 1 0 13344 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_140
timestamp 1679581782
transform 1 0 14016 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_147
timestamp 1679581782
transform 1 0 14688 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_154
timestamp 1679581782
transform 1 0 15360 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_161
timestamp 1679581782
transform 1 0 16032 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_168
timestamp 1679581782
transform 1 0 16704 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_175
timestamp 1679581782
transform 1 0 17376 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_182
timestamp 1679581782
transform 1 0 18048 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_189
timestamp 1679581782
transform 1 0 18720 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_196
timestamp 1679581782
transform 1 0 19392 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_203
timestamp 1679581782
transform 1 0 20064 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_210
timestamp 1679581782
transform 1 0 20736 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_217
timestamp 1679581782
transform 1 0 21408 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_224
timestamp 1679581782
transform 1 0 22080 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_231
timestamp 1679581782
transform 1 0 22752 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_238
timestamp 1679581782
transform 1 0 23424 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_245
timestamp 1679581782
transform 1 0 24096 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_252
timestamp 1679581782
transform 1 0 24768 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_259
timestamp 1679581782
transform 1 0 25440 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_266
timestamp 1679581782
transform 1 0 26112 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_273
timestamp 1679581782
transform 1 0 26784 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_280
timestamp 1679581782
transform 1 0 27456 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_287
timestamp 1679581782
transform 1 0 28128 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_294
timestamp 1679581782
transform 1 0 28800 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_301
timestamp 1679581782
transform 1 0 29472 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_308
timestamp 1679581782
transform 1 0 30144 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_315
timestamp 1679581782
transform 1 0 30816 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_322
timestamp 1679581782
transform 1 0 31488 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_329
timestamp 1679581782
transform 1 0 32160 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_336
timestamp 1679581782
transform 1 0 32832 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_343
timestamp 1679581782
transform 1 0 33504 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_350
timestamp 1679581782
transform 1 0 34176 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_357
timestamp 1679581782
transform 1 0 34848 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_364
timestamp 1679581782
transform 1 0 35520 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_371
timestamp 1679581782
transform 1 0 36192 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_378
timestamp 1679581782
transform 1 0 36864 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_385
timestamp 1679581782
transform 1 0 37536 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_392
timestamp 1679581782
transform 1 0 38208 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_399
timestamp 1679581782
transform 1 0 38880 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_406
timestamp 1679581782
transform 1 0 39552 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_413
timestamp 1679581782
transform 1 0 40224 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_420
timestamp 1679581782
transform 1 0 40896 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_427
timestamp 1679581782
transform 1 0 41568 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_434
timestamp 1679581782
transform 1 0 42240 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_441
timestamp 1679581782
transform 1 0 42912 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_448
timestamp 1679581782
transform 1 0 43584 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_455
timestamp 1679581782
transform 1 0 44256 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_462
timestamp 1679581782
transform 1 0 44928 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_469
timestamp 1679581782
transform 1 0 45600 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_476
timestamp 1679581782
transform 1 0 46272 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_483
timestamp 1679581782
transform 1 0 46944 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_490
timestamp 1679581782
transform 1 0 47616 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_497
timestamp 1679581782
transform 1 0 48288 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_504
timestamp 1679581782
transform 1 0 48960 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_511
timestamp 1679581782
transform 1 0 49632 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_518
timestamp 1679581782
transform 1 0 50304 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_525
timestamp 1679581782
transform 1 0 50976 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_532
timestamp 1679581782
transform 1 0 51648 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_539
timestamp 1679581782
transform 1 0 52320 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_546
timestamp 1679581782
transform 1 0 52992 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_553
timestamp 1679581782
transform 1 0 53664 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_560
timestamp 1679581782
transform 1 0 54336 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_567
timestamp 1679581782
transform 1 0 55008 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_574
timestamp 1679581782
transform 1 0 55680 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_581
timestamp 1679581782
transform 1 0 56352 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_588
timestamp 1679581782
transform 1 0 57024 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_595
timestamp 1679581782
transform 1 0 57696 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_602
timestamp 1679581782
transform 1 0 58368 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_609
timestamp 1679581782
transform 1 0 59040 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_616
timestamp 1679581782
transform 1 0 59712 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_623
timestamp 1679581782
transform 1 0 60384 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_630
timestamp 1679581782
transform 1 0 61056 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_637
timestamp 1679581782
transform 1 0 61728 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_644
timestamp 1679581782
transform 1 0 62400 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_651
timestamp 1679581782
transform 1 0 63072 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_658
timestamp 1679581782
transform 1 0 63744 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_665
timestamp 1679581782
transform 1 0 64416 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_672
timestamp 1679581782
transform 1 0 65088 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_679
timestamp 1679581782
transform 1 0 65760 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_686
timestamp 1679581782
transform 1 0 66432 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_693
timestamp 1679581782
transform 1 0 67104 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_700
timestamp 1679581782
transform 1 0 67776 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_707
timestamp 1679581782
transform 1 0 68448 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_714
timestamp 1679581782
transform 1 0 69120 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_721
timestamp 1679581782
transform 1 0 69792 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_728
timestamp 1679581782
transform 1 0 70464 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_735
timestamp 1679581782
transform 1 0 71136 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_742
timestamp 1679581782
transform 1 0 71808 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_749
timestamp 1679581782
transform 1 0 72480 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_756
timestamp 1679581782
transform 1 0 73152 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_763
timestamp 1679581782
transform 1 0 73824 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_770
timestamp 1679581782
transform 1 0 74496 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_777
timestamp 1679581782
transform 1 0 75168 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_784
timestamp 1679581782
transform 1 0 75840 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_791
timestamp 1679581782
transform 1 0 76512 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_798
timestamp 1679581782
transform 1 0 77184 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_805
timestamp 1679581782
transform 1 0 77856 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_812
timestamp 1679581782
transform 1 0 78528 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_819
timestamp 1679581782
transform 1 0 79200 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_826
timestamp 1679581782
transform 1 0 79872 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_833
timestamp 1679581782
transform 1 0 80544 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_840
timestamp 1679581782
transform 1 0 81216 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_847
timestamp 1679581782
transform 1 0 81888 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_854
timestamp 1679581782
transform 1 0 82560 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_861
timestamp 1679581782
transform 1 0 83232 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_868
timestamp 1679581782
transform 1 0 83904 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_875
timestamp 1679581782
transform 1 0 84576 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_882
timestamp 1679581782
transform 1 0 85248 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_889
timestamp 1679581782
transform 1 0 85920 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_896
timestamp 1679581782
transform 1 0 86592 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_903
timestamp 1679581782
transform 1 0 87264 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_910
timestamp 1679581782
transform 1 0 87936 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_917
timestamp 1679581782
transform 1 0 88608 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_924
timestamp 1679581782
transform 1 0 89280 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_931
timestamp 1679581782
transform 1 0 89952 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_938
timestamp 1679581782
transform 1 0 90624 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_945
timestamp 1679581782
transform 1 0 91296 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_952
timestamp 1679581782
transform 1 0 91968 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_959
timestamp 1679581782
transform 1 0 92640 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_966
timestamp 1679581782
transform 1 0 93312 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_973
timestamp 1679581782
transform 1 0 93984 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_980
timestamp 1679581782
transform 1 0 94656 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_987
timestamp 1679581782
transform 1 0 95328 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_994
timestamp 1679581782
transform 1 0 96000 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_1001
timestamp 1679581782
transform 1 0 96672 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_1008
timestamp 1679581782
transform 1 0 97344 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_1015
timestamp 1679581782
transform 1 0 98016 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_1022
timestamp 1679581782
transform 1 0 98688 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_4
timestamp 1679581782
transform 1 0 960 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_11
timestamp 1679581782
transform 1 0 1632 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_18
timestamp 1679581782
transform 1 0 2304 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_25
timestamp 1679581782
transform 1 0 2976 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_32
timestamp 1679581782
transform 1 0 3648 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_39
timestamp 1679581782
transform 1 0 4320 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_46
timestamp 1679581782
transform 1 0 4992 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_53
timestamp 1679581782
transform 1 0 5664 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_60
timestamp 1679581782
transform 1 0 6336 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_67
timestamp 1679581782
transform 1 0 7008 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_74
timestamp 1679581782
transform 1 0 7680 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_81
timestamp 1679581782
transform 1 0 8352 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_88
timestamp 1679581782
transform 1 0 9024 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_95
timestamp 1679581782
transform 1 0 9696 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_102
timestamp 1679581782
transform 1 0 10368 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_109
timestamp 1679581782
transform 1 0 11040 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_116
timestamp 1679581782
transform 1 0 11712 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_123
timestamp 1679581782
transform 1 0 12384 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_130
timestamp 1679581782
transform 1 0 13056 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_137
timestamp 1679581782
transform 1 0 13728 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_144
timestamp 1679581782
transform 1 0 14400 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_151
timestamp 1679581782
transform 1 0 15072 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_158
timestamp 1679581782
transform 1 0 15744 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_165
timestamp 1679581782
transform 1 0 16416 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_172
timestamp 1679581782
transform 1 0 17088 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_179
timestamp 1679581782
transform 1 0 17760 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_186
timestamp 1679581782
transform 1 0 18432 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_193
timestamp 1679581782
transform 1 0 19104 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_200
timestamp 1679581782
transform 1 0 19776 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_207
timestamp 1679581782
transform 1 0 20448 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_214
timestamp 1679581782
transform 1 0 21120 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_221
timestamp 1679581782
transform 1 0 21792 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_228
timestamp 1679581782
transform 1 0 22464 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_235
timestamp 1679581782
transform 1 0 23136 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_242
timestamp 1679581782
transform 1 0 23808 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_249
timestamp 1679581782
transform 1 0 24480 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_256
timestamp 1679581782
transform 1 0 25152 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_263
timestamp 1679581782
transform 1 0 25824 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_270
timestamp 1679581782
transform 1 0 26496 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_277
timestamp 1679581782
transform 1 0 27168 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_284
timestamp 1679581782
transform 1 0 27840 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_291
timestamp 1679581782
transform 1 0 28512 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_298
timestamp 1679581782
transform 1 0 29184 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_305
timestamp 1679581782
transform 1 0 29856 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_312
timestamp 1679581782
transform 1 0 30528 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_319
timestamp 1679581782
transform 1 0 31200 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_326
timestamp 1679581782
transform 1 0 31872 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_333
timestamp 1679581782
transform 1 0 32544 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_340
timestamp 1679581782
transform 1 0 33216 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_347
timestamp 1679581782
transform 1 0 33888 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_354
timestamp 1679581782
transform 1 0 34560 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_361
timestamp 1679581782
transform 1 0 35232 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_368
timestamp 1679581782
transform 1 0 35904 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_375
timestamp 1679581782
transform 1 0 36576 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_382
timestamp 1679581782
transform 1 0 37248 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_389
timestamp 1679581782
transform 1 0 37920 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_396
timestamp 1679581782
transform 1 0 38592 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_403
timestamp 1679581782
transform 1 0 39264 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_410
timestamp 1679581782
transform 1 0 39936 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_417
timestamp 1679581782
transform 1 0 40608 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_424
timestamp 1679581782
transform 1 0 41280 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_431
timestamp 1679581782
transform 1 0 41952 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_438
timestamp 1679581782
transform 1 0 42624 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_445
timestamp 1679581782
transform 1 0 43296 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_452
timestamp 1679581782
transform 1 0 43968 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_459
timestamp 1679581782
transform 1 0 44640 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_466
timestamp 1679581782
transform 1 0 45312 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_473
timestamp 1679581782
transform 1 0 45984 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_480
timestamp 1679581782
transform 1 0 46656 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_487
timestamp 1679581782
transform 1 0 47328 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_494
timestamp 1679581782
transform 1 0 48000 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_501
timestamp 1679581782
transform 1 0 48672 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_508
timestamp 1679581782
transform 1 0 49344 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_515
timestamp 1679581782
transform 1 0 50016 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_522
timestamp 1679581782
transform 1 0 50688 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_529
timestamp 1679581782
transform 1 0 51360 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_536
timestamp 1679581782
transform 1 0 52032 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_543
timestamp 1679581782
transform 1 0 52704 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_550
timestamp 1679581782
transform 1 0 53376 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_557
timestamp 1679581782
transform 1 0 54048 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_564
timestamp 1679581782
transform 1 0 54720 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_571
timestamp 1679581782
transform 1 0 55392 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_578
timestamp 1679581782
transform 1 0 56064 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_585
timestamp 1679581782
transform 1 0 56736 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_592
timestamp 1679581782
transform 1 0 57408 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_599
timestamp 1679581782
transform 1 0 58080 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_606
timestamp 1679581782
transform 1 0 58752 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_613
timestamp 1679581782
transform 1 0 59424 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_620
timestamp 1679581782
transform 1 0 60096 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_627
timestamp 1679581782
transform 1 0 60768 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_634
timestamp 1679581782
transform 1 0 61440 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_641
timestamp 1679581782
transform 1 0 62112 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_648
timestamp 1679581782
transform 1 0 62784 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_655
timestamp 1679581782
transform 1 0 63456 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_662
timestamp 1679581782
transform 1 0 64128 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_669
timestamp 1679581782
transform 1 0 64800 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_676
timestamp 1679581782
transform 1 0 65472 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_683
timestamp 1679581782
transform 1 0 66144 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_690
timestamp 1679581782
transform 1 0 66816 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_697
timestamp 1679581782
transform 1 0 67488 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_704
timestamp 1679581782
transform 1 0 68160 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_711
timestamp 1679581782
transform 1 0 68832 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_718
timestamp 1679581782
transform 1 0 69504 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_725
timestamp 1679581782
transform 1 0 70176 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_732
timestamp 1679581782
transform 1 0 70848 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_739
timestamp 1679581782
transform 1 0 71520 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_746
timestamp 1679581782
transform 1 0 72192 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_753
timestamp 1679581782
transform 1 0 72864 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_760
timestamp 1679581782
transform 1 0 73536 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_767
timestamp 1679581782
transform 1 0 74208 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_774
timestamp 1679581782
transform 1 0 74880 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_781
timestamp 1679581782
transform 1 0 75552 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_788
timestamp 1679581782
transform 1 0 76224 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_795
timestamp 1679581782
transform 1 0 76896 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_802
timestamp 1679581782
transform 1 0 77568 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_809
timestamp 1679581782
transform 1 0 78240 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_816
timestamp 1679581782
transform 1 0 78912 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_823
timestamp 1679581782
transform 1 0 79584 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_830
timestamp 1679581782
transform 1 0 80256 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_837
timestamp 1679581782
transform 1 0 80928 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_844
timestamp 1679581782
transform 1 0 81600 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_851
timestamp 1679581782
transform 1 0 82272 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_858
timestamp 1679581782
transform 1 0 82944 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_865
timestamp 1679581782
transform 1 0 83616 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_872
timestamp 1679581782
transform 1 0 84288 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_879
timestamp 1679581782
transform 1 0 84960 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_886
timestamp 1679581782
transform 1 0 85632 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_893
timestamp 1679581782
transform 1 0 86304 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_900
timestamp 1679581782
transform 1 0 86976 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_907
timestamp 1679581782
transform 1 0 87648 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_914
timestamp 1679581782
transform 1 0 88320 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_921
timestamp 1679581782
transform 1 0 88992 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_928
timestamp 1679581782
transform 1 0 89664 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_935
timestamp 1679581782
transform 1 0 90336 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_942
timestamp 1679581782
transform 1 0 91008 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_949
timestamp 1679581782
transform 1 0 91680 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_956
timestamp 1679581782
transform 1 0 92352 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_963
timestamp 1679581782
transform 1 0 93024 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_970
timestamp 1679581782
transform 1 0 93696 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_977
timestamp 1679581782
transform 1 0 94368 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_984
timestamp 1679581782
transform 1 0 95040 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_991
timestamp 1679581782
transform 1 0 95712 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_998
timestamp 1679581782
transform 1 0 96384 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_1005
timestamp 1679581782
transform 1 0 97056 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_1012
timestamp 1679581782
transform 1 0 97728 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_1019
timestamp 1679581782
transform 1 0 98400 0 1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_32_1026
timestamp 1677580104
transform 1 0 99072 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_1028
timestamp 1677579658
transform 1 0 99264 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_0
timestamp 1679581782
transform 1 0 576 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_7
timestamp 1679581782
transform 1 0 1248 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_14
timestamp 1679581782
transform 1 0 1920 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_21
timestamp 1679581782
transform 1 0 2592 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_28
timestamp 1679581782
transform 1 0 3264 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_35
timestamp 1679581782
transform 1 0 3936 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_42
timestamp 1679581782
transform 1 0 4608 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_49
timestamp 1679581782
transform 1 0 5280 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_56
timestamp 1679581782
transform 1 0 5952 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_63
timestamp 1679581782
transform 1 0 6624 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_70
timestamp 1679581782
transform 1 0 7296 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_77
timestamp 1679581782
transform 1 0 7968 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_84
timestamp 1679581782
transform 1 0 8640 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_91
timestamp 1679581782
transform 1 0 9312 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_98
timestamp 1679581782
transform 1 0 9984 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_105
timestamp 1679581782
transform 1 0 10656 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_112
timestamp 1679581782
transform 1 0 11328 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_119
timestamp 1679581782
transform 1 0 12000 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_126
timestamp 1679581782
transform 1 0 12672 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_133
timestamp 1679581782
transform 1 0 13344 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_140
timestamp 1679581782
transform 1 0 14016 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_147
timestamp 1679581782
transform 1 0 14688 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_154
timestamp 1679581782
transform 1 0 15360 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_161
timestamp 1679581782
transform 1 0 16032 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_168
timestamp 1679581782
transform 1 0 16704 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_175
timestamp 1679581782
transform 1 0 17376 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_182
timestamp 1679581782
transform 1 0 18048 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_189
timestamp 1679581782
transform 1 0 18720 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_196
timestamp 1679581782
transform 1 0 19392 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_203
timestamp 1679581782
transform 1 0 20064 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_210
timestamp 1679581782
transform 1 0 20736 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_217
timestamp 1679581782
transform 1 0 21408 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_224
timestamp 1679581782
transform 1 0 22080 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_231
timestamp 1679581782
transform 1 0 22752 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_238
timestamp 1679581782
transform 1 0 23424 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_245
timestamp 1679581782
transform 1 0 24096 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_252
timestamp 1679581782
transform 1 0 24768 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_259
timestamp 1679581782
transform 1 0 25440 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_266
timestamp 1679581782
transform 1 0 26112 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_273
timestamp 1679581782
transform 1 0 26784 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_280
timestamp 1679581782
transform 1 0 27456 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_287
timestamp 1679581782
transform 1 0 28128 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_294
timestamp 1679581782
transform 1 0 28800 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_301
timestamp 1679581782
transform 1 0 29472 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_308
timestamp 1679581782
transform 1 0 30144 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_315
timestamp 1679581782
transform 1 0 30816 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_322
timestamp 1679581782
transform 1 0 31488 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_329
timestamp 1679581782
transform 1 0 32160 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_336
timestamp 1679581782
transform 1 0 32832 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_343
timestamp 1679581782
transform 1 0 33504 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_350
timestamp 1679581782
transform 1 0 34176 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_357
timestamp 1679581782
transform 1 0 34848 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_364
timestamp 1679581782
transform 1 0 35520 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_371
timestamp 1679581782
transform 1 0 36192 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_378
timestamp 1679581782
transform 1 0 36864 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_385
timestamp 1679581782
transform 1 0 37536 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_392
timestamp 1679581782
transform 1 0 38208 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_399
timestamp 1679581782
transform 1 0 38880 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_406
timestamp 1679581782
transform 1 0 39552 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_413
timestamp 1679581782
transform 1 0 40224 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_420
timestamp 1679581782
transform 1 0 40896 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_427
timestamp 1679581782
transform 1 0 41568 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_434
timestamp 1679581782
transform 1 0 42240 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_441
timestamp 1679581782
transform 1 0 42912 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_448
timestamp 1679581782
transform 1 0 43584 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_455
timestamp 1679581782
transform 1 0 44256 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_462
timestamp 1679581782
transform 1 0 44928 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_469
timestamp 1679581782
transform 1 0 45600 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_476
timestamp 1679581782
transform 1 0 46272 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_483
timestamp 1679581782
transform 1 0 46944 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_490
timestamp 1679581782
transform 1 0 47616 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_497
timestamp 1679581782
transform 1 0 48288 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_504
timestamp 1679581782
transform 1 0 48960 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_511
timestamp 1679581782
transform 1 0 49632 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_518
timestamp 1679581782
transform 1 0 50304 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_525
timestamp 1679581782
transform 1 0 50976 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_532
timestamp 1679581782
transform 1 0 51648 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_539
timestamp 1679581782
transform 1 0 52320 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_546
timestamp 1679581782
transform 1 0 52992 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_553
timestamp 1679581782
transform 1 0 53664 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_560
timestamp 1679581782
transform 1 0 54336 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_567
timestamp 1679581782
transform 1 0 55008 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_574
timestamp 1679581782
transform 1 0 55680 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_581
timestamp 1679581782
transform 1 0 56352 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_588
timestamp 1679581782
transform 1 0 57024 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_595
timestamp 1679581782
transform 1 0 57696 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_602
timestamp 1679581782
transform 1 0 58368 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_609
timestamp 1679581782
transform 1 0 59040 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_616
timestamp 1679581782
transform 1 0 59712 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_623
timestamp 1679581782
transform 1 0 60384 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_630
timestamp 1679581782
transform 1 0 61056 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_637
timestamp 1679581782
transform 1 0 61728 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_644
timestamp 1679581782
transform 1 0 62400 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_651
timestamp 1679581782
transform 1 0 63072 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_658
timestamp 1679581782
transform 1 0 63744 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_665
timestamp 1679581782
transform 1 0 64416 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_672
timestamp 1679581782
transform 1 0 65088 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_679
timestamp 1679581782
transform 1 0 65760 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_686
timestamp 1679581782
transform 1 0 66432 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_693
timestamp 1679581782
transform 1 0 67104 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_700
timestamp 1679581782
transform 1 0 67776 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_707
timestamp 1679581782
transform 1 0 68448 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_714
timestamp 1679581782
transform 1 0 69120 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_721
timestamp 1679581782
transform 1 0 69792 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_728
timestamp 1679581782
transform 1 0 70464 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_735
timestamp 1679581782
transform 1 0 71136 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_742
timestamp 1679581782
transform 1 0 71808 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_749
timestamp 1679581782
transform 1 0 72480 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_756
timestamp 1679581782
transform 1 0 73152 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_763
timestamp 1679581782
transform 1 0 73824 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_770
timestamp 1679581782
transform 1 0 74496 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_777
timestamp 1679581782
transform 1 0 75168 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_784
timestamp 1679581782
transform 1 0 75840 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_791
timestamp 1679581782
transform 1 0 76512 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_798
timestamp 1679581782
transform 1 0 77184 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_805
timestamp 1679581782
transform 1 0 77856 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_812
timestamp 1679581782
transform 1 0 78528 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_819
timestamp 1679581782
transform 1 0 79200 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_826
timestamp 1679581782
transform 1 0 79872 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_833
timestamp 1679581782
transform 1 0 80544 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_840
timestamp 1679581782
transform 1 0 81216 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_847
timestamp 1679581782
transform 1 0 81888 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_854
timestamp 1679581782
transform 1 0 82560 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_861
timestamp 1679581782
transform 1 0 83232 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_868
timestamp 1679581782
transform 1 0 83904 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_875
timestamp 1679581782
transform 1 0 84576 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_882
timestamp 1679581782
transform 1 0 85248 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_889
timestamp 1679581782
transform 1 0 85920 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_896
timestamp 1679581782
transform 1 0 86592 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_903
timestamp 1679581782
transform 1 0 87264 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_910
timestamp 1679581782
transform 1 0 87936 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_917
timestamp 1679581782
transform 1 0 88608 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_924
timestamp 1679581782
transform 1 0 89280 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_931
timestamp 1679581782
transform 1 0 89952 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_938
timestamp 1679581782
transform 1 0 90624 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_945
timestamp 1679581782
transform 1 0 91296 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_952
timestamp 1679581782
transform 1 0 91968 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_959
timestamp 1679581782
transform 1 0 92640 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_966
timestamp 1679581782
transform 1 0 93312 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_973
timestamp 1679581782
transform 1 0 93984 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_980
timestamp 1679581782
transform 1 0 94656 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_987
timestamp 1679581782
transform 1 0 95328 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_994
timestamp 1679581782
transform 1 0 96000 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_1001
timestamp 1679581782
transform 1 0 96672 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_1008
timestamp 1679581782
transform 1 0 97344 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_1015
timestamp 1679581782
transform 1 0 98016 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_1022
timestamp 1679581782
transform 1 0 98688 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_4
timestamp 1679581782
transform 1 0 960 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_11
timestamp 1679581782
transform 1 0 1632 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_18
timestamp 1679581782
transform 1 0 2304 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_25
timestamp 1679581782
transform 1 0 2976 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_32
timestamp 1679581782
transform 1 0 3648 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_39
timestamp 1679581782
transform 1 0 4320 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_46
timestamp 1679581782
transform 1 0 4992 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_53
timestamp 1679581782
transform 1 0 5664 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_60
timestamp 1679581782
transform 1 0 6336 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_67
timestamp 1679581782
transform 1 0 7008 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_74
timestamp 1679581782
transform 1 0 7680 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_81
timestamp 1679581782
transform 1 0 8352 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_88
timestamp 1679581782
transform 1 0 9024 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_95
timestamp 1679581782
transform 1 0 9696 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_102
timestamp 1679581782
transform 1 0 10368 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_109
timestamp 1679581782
transform 1 0 11040 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_116
timestamp 1679581782
transform 1 0 11712 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_123
timestamp 1679581782
transform 1 0 12384 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_130
timestamp 1679581782
transform 1 0 13056 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_137
timestamp 1679581782
transform 1 0 13728 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_144
timestamp 1679581782
transform 1 0 14400 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_151
timestamp 1679581782
transform 1 0 15072 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_158
timestamp 1679581782
transform 1 0 15744 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_165
timestamp 1679581782
transform 1 0 16416 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_172
timestamp 1679581782
transform 1 0 17088 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_179
timestamp 1679581782
transform 1 0 17760 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_186
timestamp 1679581782
transform 1 0 18432 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_193
timestamp 1679581782
transform 1 0 19104 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_200
timestamp 1679581782
transform 1 0 19776 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_207
timestamp 1679581782
transform 1 0 20448 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_214
timestamp 1679581782
transform 1 0 21120 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_221
timestamp 1679581782
transform 1 0 21792 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_228
timestamp 1679581782
transform 1 0 22464 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_235
timestamp 1679581782
transform 1 0 23136 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_242
timestamp 1679581782
transform 1 0 23808 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_249
timestamp 1679581782
transform 1 0 24480 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_256
timestamp 1679581782
transform 1 0 25152 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_263
timestamp 1679581782
transform 1 0 25824 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_270
timestamp 1679581782
transform 1 0 26496 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_277
timestamp 1679581782
transform 1 0 27168 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_284
timestamp 1679581782
transform 1 0 27840 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_291
timestamp 1679581782
transform 1 0 28512 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_298
timestamp 1679581782
transform 1 0 29184 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_305
timestamp 1679581782
transform 1 0 29856 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_312
timestamp 1679581782
transform 1 0 30528 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_319
timestamp 1679581782
transform 1 0 31200 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_326
timestamp 1679581782
transform 1 0 31872 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_333
timestamp 1679581782
transform 1 0 32544 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_340
timestamp 1679581782
transform 1 0 33216 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_347
timestamp 1679581782
transform 1 0 33888 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_354
timestamp 1679581782
transform 1 0 34560 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_361
timestamp 1679581782
transform 1 0 35232 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_368
timestamp 1679581782
transform 1 0 35904 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_375
timestamp 1679581782
transform 1 0 36576 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_382
timestamp 1679581782
transform 1 0 37248 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_389
timestamp 1679581782
transform 1 0 37920 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_396
timestamp 1679581782
transform 1 0 38592 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_403
timestamp 1679581782
transform 1 0 39264 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_410
timestamp 1679581782
transform 1 0 39936 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_417
timestamp 1679581782
transform 1 0 40608 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_424
timestamp 1679581782
transform 1 0 41280 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_431
timestamp 1679581782
transform 1 0 41952 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_438
timestamp 1679581782
transform 1 0 42624 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_445
timestamp 1679581782
transform 1 0 43296 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_452
timestamp 1679581782
transform 1 0 43968 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_459
timestamp 1679581782
transform 1 0 44640 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_466
timestamp 1679581782
transform 1 0 45312 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_473
timestamp 1679581782
transform 1 0 45984 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_480
timestamp 1679581782
transform 1 0 46656 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_487
timestamp 1679581782
transform 1 0 47328 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_494
timestamp 1679581782
transform 1 0 48000 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_501
timestamp 1679581782
transform 1 0 48672 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_508
timestamp 1679581782
transform 1 0 49344 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_515
timestamp 1679581782
transform 1 0 50016 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_522
timestamp 1679581782
transform 1 0 50688 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_529
timestamp 1679581782
transform 1 0 51360 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_536
timestamp 1679581782
transform 1 0 52032 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_543
timestamp 1679581782
transform 1 0 52704 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_550
timestamp 1679581782
transform 1 0 53376 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_557
timestamp 1679581782
transform 1 0 54048 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_564
timestamp 1679581782
transform 1 0 54720 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_571
timestamp 1679581782
transform 1 0 55392 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_578
timestamp 1679581782
transform 1 0 56064 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_585
timestamp 1679581782
transform 1 0 56736 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_592
timestamp 1679581782
transform 1 0 57408 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_599
timestamp 1679581782
transform 1 0 58080 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_606
timestamp 1679581782
transform 1 0 58752 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_613
timestamp 1679581782
transform 1 0 59424 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_620
timestamp 1679581782
transform 1 0 60096 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_627
timestamp 1679581782
transform 1 0 60768 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_634
timestamp 1679581782
transform 1 0 61440 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_641
timestamp 1679581782
transform 1 0 62112 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_648
timestamp 1679581782
transform 1 0 62784 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_655
timestamp 1679581782
transform 1 0 63456 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_662
timestamp 1679581782
transform 1 0 64128 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_669
timestamp 1679581782
transform 1 0 64800 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_676
timestamp 1679581782
transform 1 0 65472 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_683
timestamp 1679581782
transform 1 0 66144 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_690
timestamp 1679581782
transform 1 0 66816 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_697
timestamp 1679581782
transform 1 0 67488 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_704
timestamp 1679581782
transform 1 0 68160 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_711
timestamp 1679581782
transform 1 0 68832 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_718
timestamp 1679581782
transform 1 0 69504 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_725
timestamp 1679581782
transform 1 0 70176 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_732
timestamp 1679581782
transform 1 0 70848 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_739
timestamp 1679581782
transform 1 0 71520 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_746
timestamp 1679581782
transform 1 0 72192 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_753
timestamp 1679581782
transform 1 0 72864 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_760
timestamp 1679581782
transform 1 0 73536 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_767
timestamp 1679581782
transform 1 0 74208 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_774
timestamp 1679581782
transform 1 0 74880 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_781
timestamp 1679581782
transform 1 0 75552 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_788
timestamp 1679581782
transform 1 0 76224 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_795
timestamp 1679581782
transform 1 0 76896 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_802
timestamp 1679581782
transform 1 0 77568 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_809
timestamp 1679581782
transform 1 0 78240 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_816
timestamp 1679581782
transform 1 0 78912 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_823
timestamp 1679581782
transform 1 0 79584 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_830
timestamp 1679581782
transform 1 0 80256 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_837
timestamp 1679581782
transform 1 0 80928 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_844
timestamp 1679581782
transform 1 0 81600 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_851
timestamp 1679581782
transform 1 0 82272 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_858
timestamp 1679581782
transform 1 0 82944 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_865
timestamp 1679581782
transform 1 0 83616 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_872
timestamp 1679581782
transform 1 0 84288 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_879
timestamp 1679581782
transform 1 0 84960 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_886
timestamp 1679581782
transform 1 0 85632 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_893
timestamp 1679581782
transform 1 0 86304 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_900
timestamp 1679581782
transform 1 0 86976 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_907
timestamp 1679581782
transform 1 0 87648 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_914
timestamp 1679581782
transform 1 0 88320 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_921
timestamp 1679581782
transform 1 0 88992 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_928
timestamp 1679581782
transform 1 0 89664 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_935
timestamp 1679581782
transform 1 0 90336 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_942
timestamp 1679581782
transform 1 0 91008 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_949
timestamp 1679581782
transform 1 0 91680 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_956
timestamp 1679581782
transform 1 0 92352 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_963
timestamp 1679581782
transform 1 0 93024 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_970
timestamp 1679581782
transform 1 0 93696 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_977
timestamp 1679581782
transform 1 0 94368 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_984
timestamp 1679581782
transform 1 0 95040 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_991
timestamp 1679581782
transform 1 0 95712 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_998
timestamp 1679581782
transform 1 0 96384 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_1005
timestamp 1679581782
transform 1 0 97056 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_1012
timestamp 1679581782
transform 1 0 97728 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_1019
timestamp 1679581782
transform 1 0 98400 0 1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_34_1026
timestamp 1677580104
transform 1 0 99072 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_1028
timestamp 1677579658
transform 1 0 99264 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_0
timestamp 1679581782
transform 1 0 576 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_7
timestamp 1679581782
transform 1 0 1248 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_14
timestamp 1679581782
transform 1 0 1920 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_21
timestamp 1679581782
transform 1 0 2592 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_28
timestamp 1679581782
transform 1 0 3264 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_35
timestamp 1679581782
transform 1 0 3936 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_42
timestamp 1679581782
transform 1 0 4608 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_49
timestamp 1679581782
transform 1 0 5280 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_56
timestamp 1679581782
transform 1 0 5952 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_63
timestamp 1679581782
transform 1 0 6624 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_70
timestamp 1679581782
transform 1 0 7296 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_77
timestamp 1679581782
transform 1 0 7968 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_84
timestamp 1679581782
transform 1 0 8640 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_91
timestamp 1679581782
transform 1 0 9312 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_98
timestamp 1679581782
transform 1 0 9984 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_105
timestamp 1679581782
transform 1 0 10656 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_112
timestamp 1679581782
transform 1 0 11328 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_119
timestamp 1679581782
transform 1 0 12000 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_126
timestamp 1679581782
transform 1 0 12672 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_133
timestamp 1679581782
transform 1 0 13344 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_140
timestamp 1679581782
transform 1 0 14016 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_147
timestamp 1679581782
transform 1 0 14688 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_154
timestamp 1679581782
transform 1 0 15360 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_161
timestamp 1679581782
transform 1 0 16032 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_168
timestamp 1679581782
transform 1 0 16704 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_175
timestamp 1679581782
transform 1 0 17376 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_182
timestamp 1679581782
transform 1 0 18048 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_189
timestamp 1679581782
transform 1 0 18720 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_196
timestamp 1679581782
transform 1 0 19392 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_203
timestamp 1679581782
transform 1 0 20064 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_210
timestamp 1679581782
transform 1 0 20736 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_217
timestamp 1679581782
transform 1 0 21408 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_224
timestamp 1679581782
transform 1 0 22080 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_231
timestamp 1679581782
transform 1 0 22752 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_238
timestamp 1679581782
transform 1 0 23424 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_245
timestamp 1679581782
transform 1 0 24096 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_252
timestamp 1679581782
transform 1 0 24768 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_259
timestamp 1679581782
transform 1 0 25440 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_266
timestamp 1679581782
transform 1 0 26112 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_273
timestamp 1679581782
transform 1 0 26784 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_280
timestamp 1679581782
transform 1 0 27456 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_287
timestamp 1679581782
transform 1 0 28128 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_294
timestamp 1679581782
transform 1 0 28800 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_301
timestamp 1679581782
transform 1 0 29472 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_308
timestamp 1679581782
transform 1 0 30144 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_315
timestamp 1679581782
transform 1 0 30816 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_322
timestamp 1679581782
transform 1 0 31488 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_329
timestamp 1679581782
transform 1 0 32160 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_336
timestamp 1679581782
transform 1 0 32832 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_343
timestamp 1679581782
transform 1 0 33504 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_350
timestamp 1679581782
transform 1 0 34176 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_357
timestamp 1679581782
transform 1 0 34848 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_364
timestamp 1679581782
transform 1 0 35520 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_371
timestamp 1679581782
transform 1 0 36192 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_378
timestamp 1679581782
transform 1 0 36864 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_385
timestamp 1679581782
transform 1 0 37536 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_392
timestamp 1679581782
transform 1 0 38208 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_399
timestamp 1679581782
transform 1 0 38880 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_406
timestamp 1679581782
transform 1 0 39552 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_413
timestamp 1679581782
transform 1 0 40224 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_420
timestamp 1679581782
transform 1 0 40896 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_427
timestamp 1679581782
transform 1 0 41568 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_434
timestamp 1679581782
transform 1 0 42240 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_441
timestamp 1679581782
transform 1 0 42912 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_448
timestamp 1679581782
transform 1 0 43584 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_455
timestamp 1679581782
transform 1 0 44256 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_462
timestamp 1679581782
transform 1 0 44928 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_469
timestamp 1679581782
transform 1 0 45600 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_476
timestamp 1679581782
transform 1 0 46272 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_483
timestamp 1679581782
transform 1 0 46944 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_490
timestamp 1679581782
transform 1 0 47616 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_497
timestamp 1679581782
transform 1 0 48288 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_504
timestamp 1679581782
transform 1 0 48960 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_511
timestamp 1679581782
transform 1 0 49632 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_518
timestamp 1679581782
transform 1 0 50304 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_525
timestamp 1679581782
transform 1 0 50976 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_532
timestamp 1679581782
transform 1 0 51648 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_539
timestamp 1679581782
transform 1 0 52320 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_546
timestamp 1679581782
transform 1 0 52992 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_553
timestamp 1679581782
transform 1 0 53664 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_560
timestamp 1679581782
transform 1 0 54336 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_567
timestamp 1679581782
transform 1 0 55008 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_574
timestamp 1679581782
transform 1 0 55680 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_581
timestamp 1679581782
transform 1 0 56352 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_588
timestamp 1679581782
transform 1 0 57024 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_595
timestamp 1679581782
transform 1 0 57696 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_602
timestamp 1679581782
transform 1 0 58368 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_609
timestamp 1679581782
transform 1 0 59040 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_616
timestamp 1679581782
transform 1 0 59712 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_623
timestamp 1679581782
transform 1 0 60384 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_630
timestamp 1679581782
transform 1 0 61056 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_637
timestamp 1679581782
transform 1 0 61728 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_644
timestamp 1679581782
transform 1 0 62400 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_651
timestamp 1679581782
transform 1 0 63072 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_658
timestamp 1679581782
transform 1 0 63744 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_665
timestamp 1679581782
transform 1 0 64416 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_672
timestamp 1679581782
transform 1 0 65088 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_679
timestamp 1679581782
transform 1 0 65760 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_686
timestamp 1679581782
transform 1 0 66432 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_693
timestamp 1679581782
transform 1 0 67104 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_700
timestamp 1679581782
transform 1 0 67776 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_707
timestamp 1679581782
transform 1 0 68448 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_714
timestamp 1679581782
transform 1 0 69120 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_721
timestamp 1679581782
transform 1 0 69792 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_728
timestamp 1679581782
transform 1 0 70464 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_735
timestamp 1679581782
transform 1 0 71136 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_742
timestamp 1679581782
transform 1 0 71808 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_749
timestamp 1679581782
transform 1 0 72480 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_756
timestamp 1679581782
transform 1 0 73152 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_763
timestamp 1679581782
transform 1 0 73824 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_770
timestamp 1679581782
transform 1 0 74496 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_777
timestamp 1679581782
transform 1 0 75168 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_784
timestamp 1679581782
transform 1 0 75840 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_791
timestamp 1679581782
transform 1 0 76512 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_798
timestamp 1679581782
transform 1 0 77184 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_805
timestamp 1679581782
transform 1 0 77856 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_812
timestamp 1679581782
transform 1 0 78528 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_819
timestamp 1679581782
transform 1 0 79200 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_826
timestamp 1679581782
transform 1 0 79872 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_833
timestamp 1679581782
transform 1 0 80544 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_840
timestamp 1679581782
transform 1 0 81216 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_847
timestamp 1679581782
transform 1 0 81888 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_854
timestamp 1679581782
transform 1 0 82560 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_861
timestamp 1679581782
transform 1 0 83232 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_868
timestamp 1679581782
transform 1 0 83904 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_875
timestamp 1679581782
transform 1 0 84576 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_882
timestamp 1679581782
transform 1 0 85248 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_889
timestamp 1679581782
transform 1 0 85920 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_896
timestamp 1679581782
transform 1 0 86592 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_903
timestamp 1679581782
transform 1 0 87264 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_910
timestamp 1679581782
transform 1 0 87936 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_917
timestamp 1679581782
transform 1 0 88608 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_924
timestamp 1679581782
transform 1 0 89280 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_931
timestamp 1679581782
transform 1 0 89952 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_938
timestamp 1679581782
transform 1 0 90624 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_945
timestamp 1679581782
transform 1 0 91296 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_952
timestamp 1679581782
transform 1 0 91968 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_959
timestamp 1679581782
transform 1 0 92640 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_966
timestamp 1679581782
transform 1 0 93312 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_973
timestamp 1679581782
transform 1 0 93984 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_980
timestamp 1679581782
transform 1 0 94656 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_987
timestamp 1679581782
transform 1 0 95328 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_994
timestamp 1679581782
transform 1 0 96000 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_1001
timestamp 1679581782
transform 1 0 96672 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_1008
timestamp 1679581782
transform 1 0 97344 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_1015
timestamp 1679581782
transform 1 0 98016 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_1022
timestamp 1679581782
transform 1 0 98688 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_0
timestamp 1679581782
transform 1 0 576 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_7
timestamp 1679581782
transform 1 0 1248 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_14
timestamp 1679581782
transform 1 0 1920 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_21
timestamp 1679581782
transform 1 0 2592 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_28
timestamp 1679581782
transform 1 0 3264 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_35
timestamp 1679581782
transform 1 0 3936 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_42
timestamp 1679581782
transform 1 0 4608 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_49
timestamp 1679581782
transform 1 0 5280 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_56
timestamp 1679581782
transform 1 0 5952 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_63
timestamp 1679581782
transform 1 0 6624 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_70
timestamp 1679581782
transform 1 0 7296 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_77
timestamp 1679581782
transform 1 0 7968 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_84
timestamp 1679581782
transform 1 0 8640 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_91
timestamp 1679581782
transform 1 0 9312 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_98
timestamp 1679581782
transform 1 0 9984 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_105
timestamp 1679581782
transform 1 0 10656 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_112
timestamp 1679581782
transform 1 0 11328 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_119
timestamp 1679581782
transform 1 0 12000 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_126
timestamp 1679581782
transform 1 0 12672 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_133
timestamp 1679581782
transform 1 0 13344 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_140
timestamp 1679581782
transform 1 0 14016 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_147
timestamp 1679581782
transform 1 0 14688 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_154
timestamp 1679581782
transform 1 0 15360 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_161
timestamp 1679581782
transform 1 0 16032 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_168
timestamp 1679581782
transform 1 0 16704 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_175
timestamp 1679581782
transform 1 0 17376 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_182
timestamp 1679581782
transform 1 0 18048 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_189
timestamp 1679581782
transform 1 0 18720 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_196
timestamp 1679581782
transform 1 0 19392 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_203
timestamp 1679581782
transform 1 0 20064 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_210
timestamp 1679581782
transform 1 0 20736 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_217
timestamp 1679581782
transform 1 0 21408 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_224
timestamp 1679581782
transform 1 0 22080 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_231
timestamp 1679581782
transform 1 0 22752 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_238
timestamp 1679581782
transform 1 0 23424 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_245
timestamp 1679581782
transform 1 0 24096 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_252
timestamp 1679581782
transform 1 0 24768 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_259
timestamp 1679581782
transform 1 0 25440 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_266
timestamp 1679581782
transform 1 0 26112 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_273
timestamp 1679581782
transform 1 0 26784 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_280
timestamp 1679581782
transform 1 0 27456 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_287
timestamp 1679581782
transform 1 0 28128 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_294
timestamp 1679581782
transform 1 0 28800 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_301
timestamp 1679581782
transform 1 0 29472 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_308
timestamp 1679581782
transform 1 0 30144 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_315
timestamp 1679581782
transform 1 0 30816 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_322
timestamp 1679581782
transform 1 0 31488 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_329
timestamp 1679581782
transform 1 0 32160 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_336
timestamp 1679581782
transform 1 0 32832 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_343
timestamp 1679581782
transform 1 0 33504 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_350
timestamp 1679581782
transform 1 0 34176 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_357
timestamp 1679581782
transform 1 0 34848 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_364
timestamp 1679581782
transform 1 0 35520 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_371
timestamp 1679581782
transform 1 0 36192 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_378
timestamp 1679581782
transform 1 0 36864 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_385
timestamp 1679581782
transform 1 0 37536 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_392
timestamp 1679581782
transform 1 0 38208 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_399
timestamp 1679581782
transform 1 0 38880 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_406
timestamp 1679581782
transform 1 0 39552 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_413
timestamp 1679581782
transform 1 0 40224 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_420
timestamp 1679581782
transform 1 0 40896 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_427
timestamp 1679581782
transform 1 0 41568 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_434
timestamp 1679581782
transform 1 0 42240 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_441
timestamp 1679581782
transform 1 0 42912 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_448
timestamp 1679581782
transform 1 0 43584 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_455
timestamp 1679581782
transform 1 0 44256 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_462
timestamp 1679581782
transform 1 0 44928 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_469
timestamp 1679581782
transform 1 0 45600 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_476
timestamp 1679581782
transform 1 0 46272 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_483
timestamp 1679581782
transform 1 0 46944 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_490
timestamp 1679581782
transform 1 0 47616 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_497
timestamp 1679581782
transform 1 0 48288 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_504
timestamp 1679581782
transform 1 0 48960 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_511
timestamp 1679581782
transform 1 0 49632 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_518
timestamp 1679581782
transform 1 0 50304 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_525
timestamp 1679581782
transform 1 0 50976 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_532
timestamp 1679581782
transform 1 0 51648 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_539
timestamp 1679581782
transform 1 0 52320 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_546
timestamp 1679581782
transform 1 0 52992 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_553
timestamp 1679581782
transform 1 0 53664 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_560
timestamp 1679581782
transform 1 0 54336 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_567
timestamp 1679581782
transform 1 0 55008 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_574
timestamp 1679581782
transform 1 0 55680 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_581
timestamp 1679581782
transform 1 0 56352 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_588
timestamp 1679581782
transform 1 0 57024 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_595
timestamp 1679581782
transform 1 0 57696 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_602
timestamp 1679581782
transform 1 0 58368 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_609
timestamp 1679581782
transform 1 0 59040 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_616
timestamp 1679581782
transform 1 0 59712 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_623
timestamp 1679581782
transform 1 0 60384 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_630
timestamp 1679581782
transform 1 0 61056 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_637
timestamp 1679581782
transform 1 0 61728 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_644
timestamp 1679581782
transform 1 0 62400 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_651
timestamp 1679581782
transform 1 0 63072 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_658
timestamp 1679581782
transform 1 0 63744 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_665
timestamp 1679581782
transform 1 0 64416 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_672
timestamp 1679581782
transform 1 0 65088 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_679
timestamp 1679581782
transform 1 0 65760 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_686
timestamp 1679581782
transform 1 0 66432 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_693
timestamp 1679581782
transform 1 0 67104 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_700
timestamp 1679581782
transform 1 0 67776 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_707
timestamp 1679581782
transform 1 0 68448 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_714
timestamp 1679581782
transform 1 0 69120 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_721
timestamp 1679581782
transform 1 0 69792 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_728
timestamp 1679581782
transform 1 0 70464 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_735
timestamp 1679581782
transform 1 0 71136 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_742
timestamp 1679581782
transform 1 0 71808 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_749
timestamp 1679581782
transform 1 0 72480 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_756
timestamp 1679581782
transform 1 0 73152 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_763
timestamp 1679581782
transform 1 0 73824 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_770
timestamp 1679581782
transform 1 0 74496 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_777
timestamp 1679581782
transform 1 0 75168 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_784
timestamp 1679581782
transform 1 0 75840 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_791
timestamp 1679581782
transform 1 0 76512 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_798
timestamp 1679581782
transform 1 0 77184 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_805
timestamp 1679581782
transform 1 0 77856 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_812
timestamp 1679581782
transform 1 0 78528 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_819
timestamp 1679581782
transform 1 0 79200 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_826
timestamp 1679581782
transform 1 0 79872 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_833
timestamp 1679581782
transform 1 0 80544 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_840
timestamp 1679581782
transform 1 0 81216 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_847
timestamp 1679581782
transform 1 0 81888 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_854
timestamp 1679581782
transform 1 0 82560 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_861
timestamp 1679581782
transform 1 0 83232 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_868
timestamp 1679581782
transform 1 0 83904 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_875
timestamp 1679581782
transform 1 0 84576 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_882
timestamp 1679581782
transform 1 0 85248 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_889
timestamp 1679581782
transform 1 0 85920 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_896
timestamp 1679581782
transform 1 0 86592 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_903
timestamp 1679581782
transform 1 0 87264 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_910
timestamp 1679581782
transform 1 0 87936 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_917
timestamp 1679581782
transform 1 0 88608 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_924
timestamp 1679581782
transform 1 0 89280 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_931
timestamp 1679581782
transform 1 0 89952 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_938
timestamp 1679581782
transform 1 0 90624 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_945
timestamp 1679581782
transform 1 0 91296 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_952
timestamp 1679581782
transform 1 0 91968 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_959
timestamp 1679581782
transform 1 0 92640 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_966
timestamp 1679581782
transform 1 0 93312 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_973
timestamp 1679581782
transform 1 0 93984 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_980
timestamp 1679581782
transform 1 0 94656 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_987
timestamp 1679581782
transform 1 0 95328 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_994
timestamp 1679581782
transform 1 0 96000 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_1001
timestamp 1679581782
transform 1 0 96672 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_1008
timestamp 1679581782
transform 1 0 97344 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_1015
timestamp 1679581782
transform 1 0 98016 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_1022
timestamp 1679581782
transform 1 0 98688 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_4
timestamp 1679581782
transform 1 0 960 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_11
timestamp 1679581782
transform 1 0 1632 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_18
timestamp 1679581782
transform 1 0 2304 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_25
timestamp 1679581782
transform 1 0 2976 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_32
timestamp 1679581782
transform 1 0 3648 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_39
timestamp 1679581782
transform 1 0 4320 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_46
timestamp 1679581782
transform 1 0 4992 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_53
timestamp 1679581782
transform 1 0 5664 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_60
timestamp 1679581782
transform 1 0 6336 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_67
timestamp 1679581782
transform 1 0 7008 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_74
timestamp 1679581782
transform 1 0 7680 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_81
timestamp 1679581782
transform 1 0 8352 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_88
timestamp 1679581782
transform 1 0 9024 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_95
timestamp 1679581782
transform 1 0 9696 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_102
timestamp 1679581782
transform 1 0 10368 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_109
timestamp 1679581782
transform 1 0 11040 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_116
timestamp 1679581782
transform 1 0 11712 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_123
timestamp 1679581782
transform 1 0 12384 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_130
timestamp 1679581782
transform 1 0 13056 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_137
timestamp 1679581782
transform 1 0 13728 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_144
timestamp 1679581782
transform 1 0 14400 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_151
timestamp 1679581782
transform 1 0 15072 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_158
timestamp 1679581782
transform 1 0 15744 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_165
timestamp 1679581782
transform 1 0 16416 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_172
timestamp 1679581782
transform 1 0 17088 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_179
timestamp 1679581782
transform 1 0 17760 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_186
timestamp 1679581782
transform 1 0 18432 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_193
timestamp 1679581782
transform 1 0 19104 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_200
timestamp 1679581782
transform 1 0 19776 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_207
timestamp 1679581782
transform 1 0 20448 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_214
timestamp 1679581782
transform 1 0 21120 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_221
timestamp 1679581782
transform 1 0 21792 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_228
timestamp 1679581782
transform 1 0 22464 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_235
timestamp 1679581782
transform 1 0 23136 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_242
timestamp 1679581782
transform 1 0 23808 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_249
timestamp 1679581782
transform 1 0 24480 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_256
timestamp 1679581782
transform 1 0 25152 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_263
timestamp 1679581782
transform 1 0 25824 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_270
timestamp 1679581782
transform 1 0 26496 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_277
timestamp 1679581782
transform 1 0 27168 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_284
timestamp 1679581782
transform 1 0 27840 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_291
timestamp 1679581782
transform 1 0 28512 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_298
timestamp 1679581782
transform 1 0 29184 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_305
timestamp 1679581782
transform 1 0 29856 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_312
timestamp 1679581782
transform 1 0 30528 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_319
timestamp 1679581782
transform 1 0 31200 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_326
timestamp 1679581782
transform 1 0 31872 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_333
timestamp 1679581782
transform 1 0 32544 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_340
timestamp 1679581782
transform 1 0 33216 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_347
timestamp 1679581782
transform 1 0 33888 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_354
timestamp 1679581782
transform 1 0 34560 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_361
timestamp 1679581782
transform 1 0 35232 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_368
timestamp 1679581782
transform 1 0 35904 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_375
timestamp 1679581782
transform 1 0 36576 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_382
timestamp 1679581782
transform 1 0 37248 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_389
timestamp 1679581782
transform 1 0 37920 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_396
timestamp 1679581782
transform 1 0 38592 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_403
timestamp 1679581782
transform 1 0 39264 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_410
timestamp 1679581782
transform 1 0 39936 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_417
timestamp 1679581782
transform 1 0 40608 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_424
timestamp 1679581782
transform 1 0 41280 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_431
timestamp 1679581782
transform 1 0 41952 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_438
timestamp 1679581782
transform 1 0 42624 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_445
timestamp 1679581782
transform 1 0 43296 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_452
timestamp 1679581782
transform 1 0 43968 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_459
timestamp 1679581782
transform 1 0 44640 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_466
timestamp 1679581782
transform 1 0 45312 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_473
timestamp 1679581782
transform 1 0 45984 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_480
timestamp 1679581782
transform 1 0 46656 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_487
timestamp 1679581782
transform 1 0 47328 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_494
timestamp 1679581782
transform 1 0 48000 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_501
timestamp 1679581782
transform 1 0 48672 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_508
timestamp 1679581782
transform 1 0 49344 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_515
timestamp 1679581782
transform 1 0 50016 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_522
timestamp 1679581782
transform 1 0 50688 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_529
timestamp 1679581782
transform 1 0 51360 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_536
timestamp 1679581782
transform 1 0 52032 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_543
timestamp 1679581782
transform 1 0 52704 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_550
timestamp 1679581782
transform 1 0 53376 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_557
timestamp 1679581782
transform 1 0 54048 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_564
timestamp 1679581782
transform 1 0 54720 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_571
timestamp 1679581782
transform 1 0 55392 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_578
timestamp 1679581782
transform 1 0 56064 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_585
timestamp 1679581782
transform 1 0 56736 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_592
timestamp 1679581782
transform 1 0 57408 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_599
timestamp 1679581782
transform 1 0 58080 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_606
timestamp 1679581782
transform 1 0 58752 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_613
timestamp 1679581782
transform 1 0 59424 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_620
timestamp 1679581782
transform 1 0 60096 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_627
timestamp 1679581782
transform 1 0 60768 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_634
timestamp 1679581782
transform 1 0 61440 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_641
timestamp 1679581782
transform 1 0 62112 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_648
timestamp 1679581782
transform 1 0 62784 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_655
timestamp 1679581782
transform 1 0 63456 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_662
timestamp 1679581782
transform 1 0 64128 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_669
timestamp 1679581782
transform 1 0 64800 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_676
timestamp 1679581782
transform 1 0 65472 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_683
timestamp 1679581782
transform 1 0 66144 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_690
timestamp 1679581782
transform 1 0 66816 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_697
timestamp 1679581782
transform 1 0 67488 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_704
timestamp 1679581782
transform 1 0 68160 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_711
timestamp 1679581782
transform 1 0 68832 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_718
timestamp 1679581782
transform 1 0 69504 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_725
timestamp 1679581782
transform 1 0 70176 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_732
timestamp 1679581782
transform 1 0 70848 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_739
timestamp 1679581782
transform 1 0 71520 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_746
timestamp 1679581782
transform 1 0 72192 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_753
timestamp 1679581782
transform 1 0 72864 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_760
timestamp 1679581782
transform 1 0 73536 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_767
timestamp 1679581782
transform 1 0 74208 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_774
timestamp 1679581782
transform 1 0 74880 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_781
timestamp 1679581782
transform 1 0 75552 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_788
timestamp 1679581782
transform 1 0 76224 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_795
timestamp 1679581782
transform 1 0 76896 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_802
timestamp 1679581782
transform 1 0 77568 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_809
timestamp 1679581782
transform 1 0 78240 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_816
timestamp 1679581782
transform 1 0 78912 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_823
timestamp 1679581782
transform 1 0 79584 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_830
timestamp 1679581782
transform 1 0 80256 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_837
timestamp 1679581782
transform 1 0 80928 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_844
timestamp 1679581782
transform 1 0 81600 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_851
timestamp 1679581782
transform 1 0 82272 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_858
timestamp 1679581782
transform 1 0 82944 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_865
timestamp 1679581782
transform 1 0 83616 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_872
timestamp 1679581782
transform 1 0 84288 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_879
timestamp 1679581782
transform 1 0 84960 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_886
timestamp 1679581782
transform 1 0 85632 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_893
timestamp 1679581782
transform 1 0 86304 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_900
timestamp 1679581782
transform 1 0 86976 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_907
timestamp 1679581782
transform 1 0 87648 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_914
timestamp 1679581782
transform 1 0 88320 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_921
timestamp 1679581782
transform 1 0 88992 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_928
timestamp 1679581782
transform 1 0 89664 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_935
timestamp 1679581782
transform 1 0 90336 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_942
timestamp 1679581782
transform 1 0 91008 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_949
timestamp 1679581782
transform 1 0 91680 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_956
timestamp 1679581782
transform 1 0 92352 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_963
timestamp 1679581782
transform 1 0 93024 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_970
timestamp 1679581782
transform 1 0 93696 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_977
timestamp 1679581782
transform 1 0 94368 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_984
timestamp 1679581782
transform 1 0 95040 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_991
timestamp 1679581782
transform 1 0 95712 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_998
timestamp 1679581782
transform 1 0 96384 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_1005
timestamp 1679581782
transform 1 0 97056 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_1012
timestamp 1679581782
transform 1 0 97728 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_1019
timestamp 1679581782
transform 1 0 98400 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_37_1026
timestamp 1677580104
transform 1 0 99072 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_1028
timestamp 1677579658
transform 1 0 99264 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_0
timestamp 1679581782
transform 1 0 576 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_7
timestamp 1679581782
transform 1 0 1248 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_14
timestamp 1679581782
transform 1 0 1920 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_21
timestamp 1679581782
transform 1 0 2592 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_28
timestamp 1679581782
transform 1 0 3264 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_35
timestamp 1679581782
transform 1 0 3936 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_42
timestamp 1679581782
transform 1 0 4608 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_49
timestamp 1679581782
transform 1 0 5280 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_56
timestamp 1679581782
transform 1 0 5952 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_63
timestamp 1679581782
transform 1 0 6624 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_70
timestamp 1679581782
transform 1 0 7296 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_77
timestamp 1679581782
transform 1 0 7968 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_84
timestamp 1679581782
transform 1 0 8640 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_91
timestamp 1679581782
transform 1 0 9312 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_98
timestamp 1679581782
transform 1 0 9984 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_105
timestamp 1679581782
transform 1 0 10656 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_112
timestamp 1679581782
transform 1 0 11328 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_119
timestamp 1679581782
transform 1 0 12000 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_126
timestamp 1679581782
transform 1 0 12672 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_133
timestamp 1679581782
transform 1 0 13344 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_140
timestamp 1679581782
transform 1 0 14016 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_147
timestamp 1679581782
transform 1 0 14688 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_154
timestamp 1679581782
transform 1 0 15360 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_161
timestamp 1679581782
transform 1 0 16032 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_168
timestamp 1679581782
transform 1 0 16704 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_175
timestamp 1679581782
transform 1 0 17376 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_182
timestamp 1679581782
transform 1 0 18048 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_189
timestamp 1679581782
transform 1 0 18720 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_196
timestamp 1679581782
transform 1 0 19392 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_203
timestamp 1679581782
transform 1 0 20064 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_210
timestamp 1679581782
transform 1 0 20736 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_217
timestamp 1679581782
transform 1 0 21408 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_224
timestamp 1679581782
transform 1 0 22080 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_231
timestamp 1679581782
transform 1 0 22752 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_238
timestamp 1679581782
transform 1 0 23424 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_245
timestamp 1679581782
transform 1 0 24096 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_252
timestamp 1679581782
transform 1 0 24768 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_259
timestamp 1679581782
transform 1 0 25440 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_266
timestamp 1679581782
transform 1 0 26112 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_273
timestamp 1679581782
transform 1 0 26784 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_280
timestamp 1679581782
transform 1 0 27456 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_287
timestamp 1679581782
transform 1 0 28128 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_294
timestamp 1679581782
transform 1 0 28800 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_301
timestamp 1679581782
transform 1 0 29472 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_308
timestamp 1679581782
transform 1 0 30144 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_315
timestamp 1679581782
transform 1 0 30816 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_322
timestamp 1679581782
transform 1 0 31488 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_329
timestamp 1679581782
transform 1 0 32160 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_336
timestamp 1679581782
transform 1 0 32832 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_343
timestamp 1679581782
transform 1 0 33504 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_350
timestamp 1679581782
transform 1 0 34176 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_357
timestamp 1679581782
transform 1 0 34848 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_364
timestamp 1679581782
transform 1 0 35520 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_371
timestamp 1679581782
transform 1 0 36192 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_378
timestamp 1679581782
transform 1 0 36864 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_385
timestamp 1679581782
transform 1 0 37536 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_392
timestamp 1679581782
transform 1 0 38208 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_399
timestamp 1679581782
transform 1 0 38880 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_406
timestamp 1679581782
transform 1 0 39552 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_413
timestamp 1679581782
transform 1 0 40224 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_420
timestamp 1679581782
transform 1 0 40896 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_427
timestamp 1679581782
transform 1 0 41568 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_434
timestamp 1679581782
transform 1 0 42240 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_441
timestamp 1679581782
transform 1 0 42912 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_448
timestamp 1679581782
transform 1 0 43584 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_455
timestamp 1679581782
transform 1 0 44256 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_462
timestamp 1679581782
transform 1 0 44928 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_469
timestamp 1679581782
transform 1 0 45600 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_476
timestamp 1679581782
transform 1 0 46272 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_483
timestamp 1679581782
transform 1 0 46944 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_490
timestamp 1679581782
transform 1 0 47616 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_497
timestamp 1679581782
transform 1 0 48288 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_504
timestamp 1679581782
transform 1 0 48960 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_511
timestamp 1679581782
transform 1 0 49632 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_518
timestamp 1679581782
transform 1 0 50304 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_525
timestamp 1679581782
transform 1 0 50976 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_532
timestamp 1679581782
transform 1 0 51648 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_539
timestamp 1679581782
transform 1 0 52320 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_546
timestamp 1679581782
transform 1 0 52992 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_553
timestamp 1679581782
transform 1 0 53664 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_560
timestamp 1679581782
transform 1 0 54336 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_567
timestamp 1679581782
transform 1 0 55008 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_574
timestamp 1679581782
transform 1 0 55680 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_581
timestamp 1679581782
transform 1 0 56352 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_588
timestamp 1679581782
transform 1 0 57024 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_595
timestamp 1679581782
transform 1 0 57696 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_602
timestamp 1679581782
transform 1 0 58368 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_609
timestamp 1679581782
transform 1 0 59040 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_616
timestamp 1679581782
transform 1 0 59712 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_623
timestamp 1679581782
transform 1 0 60384 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_630
timestamp 1679581782
transform 1 0 61056 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_637
timestamp 1679581782
transform 1 0 61728 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_644
timestamp 1679581782
transform 1 0 62400 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_651
timestamp 1679581782
transform 1 0 63072 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_658
timestamp 1679581782
transform 1 0 63744 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_665
timestamp 1679581782
transform 1 0 64416 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_672
timestamp 1679581782
transform 1 0 65088 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_679
timestamp 1679581782
transform 1 0 65760 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_686
timestamp 1679581782
transform 1 0 66432 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_693
timestamp 1679581782
transform 1 0 67104 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_700
timestamp 1679581782
transform 1 0 67776 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_707
timestamp 1679581782
transform 1 0 68448 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_714
timestamp 1679581782
transform 1 0 69120 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_721
timestamp 1679581782
transform 1 0 69792 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_728
timestamp 1679581782
transform 1 0 70464 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_735
timestamp 1679581782
transform 1 0 71136 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_742
timestamp 1679581782
transform 1 0 71808 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_749
timestamp 1679581782
transform 1 0 72480 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_756
timestamp 1679581782
transform 1 0 73152 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_763
timestamp 1679581782
transform 1 0 73824 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_770
timestamp 1679581782
transform 1 0 74496 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_777
timestamp 1679581782
transform 1 0 75168 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_784
timestamp 1679581782
transform 1 0 75840 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_791
timestamp 1679581782
transform 1 0 76512 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_798
timestamp 1679581782
transform 1 0 77184 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_805
timestamp 1679581782
transform 1 0 77856 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_812
timestamp 1679581782
transform 1 0 78528 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_819
timestamp 1679581782
transform 1 0 79200 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_826
timestamp 1679581782
transform 1 0 79872 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_833
timestamp 1679581782
transform 1 0 80544 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_840
timestamp 1679581782
transform 1 0 81216 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_847
timestamp 1679581782
transform 1 0 81888 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_854
timestamp 1679581782
transform 1 0 82560 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_861
timestamp 1679581782
transform 1 0 83232 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_868
timestamp 1679581782
transform 1 0 83904 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_875
timestamp 1679581782
transform 1 0 84576 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_882
timestamp 1679581782
transform 1 0 85248 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_889
timestamp 1679581782
transform 1 0 85920 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_896
timestamp 1679581782
transform 1 0 86592 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_903
timestamp 1679581782
transform 1 0 87264 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_910
timestamp 1679581782
transform 1 0 87936 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_917
timestamp 1679581782
transform 1 0 88608 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_924
timestamp 1679581782
transform 1 0 89280 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_931
timestamp 1679581782
transform 1 0 89952 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_938
timestamp 1679581782
transform 1 0 90624 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_945
timestamp 1679581782
transform 1 0 91296 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_952
timestamp 1679581782
transform 1 0 91968 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_959
timestamp 1679581782
transform 1 0 92640 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_966
timestamp 1679581782
transform 1 0 93312 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_973
timestamp 1679581782
transform 1 0 93984 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_980
timestamp 1679581782
transform 1 0 94656 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_987
timestamp 1679581782
transform 1 0 95328 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_994
timestamp 1679581782
transform 1 0 96000 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_1001
timestamp 1679581782
transform 1 0 96672 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_1008
timestamp 1679581782
transform 1 0 97344 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_1015
timestamp 1679581782
transform 1 0 98016 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_1022
timestamp 1679581782
transform 1 0 98688 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_4
timestamp 1679581782
transform 1 0 960 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_11
timestamp 1679581782
transform 1 0 1632 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_18
timestamp 1679581782
transform 1 0 2304 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_25
timestamp 1679581782
transform 1 0 2976 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_32
timestamp 1679581782
transform 1 0 3648 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_39
timestamp 1679581782
transform 1 0 4320 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_46
timestamp 1679581782
transform 1 0 4992 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_53
timestamp 1679581782
transform 1 0 5664 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_60
timestamp 1679581782
transform 1 0 6336 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_67
timestamp 1679581782
transform 1 0 7008 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_74
timestamp 1679581782
transform 1 0 7680 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_81
timestamp 1679581782
transform 1 0 8352 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_88
timestamp 1679581782
transform 1 0 9024 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_95
timestamp 1679581782
transform 1 0 9696 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_102
timestamp 1679581782
transform 1 0 10368 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_109
timestamp 1679581782
transform 1 0 11040 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_116
timestamp 1679581782
transform 1 0 11712 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_123
timestamp 1679581782
transform 1 0 12384 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_130
timestamp 1679581782
transform 1 0 13056 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_137
timestamp 1679581782
transform 1 0 13728 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_144
timestamp 1679581782
transform 1 0 14400 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_151
timestamp 1679581782
transform 1 0 15072 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_158
timestamp 1679581782
transform 1 0 15744 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_165
timestamp 1679581782
transform 1 0 16416 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_172
timestamp 1679581782
transform 1 0 17088 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_179
timestamp 1679581782
transform 1 0 17760 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_186
timestamp 1679581782
transform 1 0 18432 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_193
timestamp 1679581782
transform 1 0 19104 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_200
timestamp 1679581782
transform 1 0 19776 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_207
timestamp 1679581782
transform 1 0 20448 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_214
timestamp 1679581782
transform 1 0 21120 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_221
timestamp 1679581782
transform 1 0 21792 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_228
timestamp 1679581782
transform 1 0 22464 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_235
timestamp 1679581782
transform 1 0 23136 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_242
timestamp 1679581782
transform 1 0 23808 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_249
timestamp 1679581782
transform 1 0 24480 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_256
timestamp 1679581782
transform 1 0 25152 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_263
timestamp 1679581782
transform 1 0 25824 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_270
timestamp 1679581782
transform 1 0 26496 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_277
timestamp 1679581782
transform 1 0 27168 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_284
timestamp 1679581782
transform 1 0 27840 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_291
timestamp 1679581782
transform 1 0 28512 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_298
timestamp 1679581782
transform 1 0 29184 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_305
timestamp 1679581782
transform 1 0 29856 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_312
timestamp 1679581782
transform 1 0 30528 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_319
timestamp 1679581782
transform 1 0 31200 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_326
timestamp 1679581782
transform 1 0 31872 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_333
timestamp 1679581782
transform 1 0 32544 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_340
timestamp 1679581782
transform 1 0 33216 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_347
timestamp 1679581782
transform 1 0 33888 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_354
timestamp 1679581782
transform 1 0 34560 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_361
timestamp 1679581782
transform 1 0 35232 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_368
timestamp 1679581782
transform 1 0 35904 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_375
timestamp 1679581782
transform 1 0 36576 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_382
timestamp 1679581782
transform 1 0 37248 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_389
timestamp 1679581782
transform 1 0 37920 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_396
timestamp 1679581782
transform 1 0 38592 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_403
timestamp 1679581782
transform 1 0 39264 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_410
timestamp 1679581782
transform 1 0 39936 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_417
timestamp 1679581782
transform 1 0 40608 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_424
timestamp 1679581782
transform 1 0 41280 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_431
timestamp 1679581782
transform 1 0 41952 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_438
timestamp 1679581782
transform 1 0 42624 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_445
timestamp 1679581782
transform 1 0 43296 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_452
timestamp 1679581782
transform 1 0 43968 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_459
timestamp 1679581782
transform 1 0 44640 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_466
timestamp 1679581782
transform 1 0 45312 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_473
timestamp 1679581782
transform 1 0 45984 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_480
timestamp 1679581782
transform 1 0 46656 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_487
timestamp 1679581782
transform 1 0 47328 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_494
timestamp 1679581782
transform 1 0 48000 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_501
timestamp 1679581782
transform 1 0 48672 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_508
timestamp 1679581782
transform 1 0 49344 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_515
timestamp 1679581782
transform 1 0 50016 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_522
timestamp 1679581782
transform 1 0 50688 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_529
timestamp 1679581782
transform 1 0 51360 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_536
timestamp 1679581782
transform 1 0 52032 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_543
timestamp 1679581782
transform 1 0 52704 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_550
timestamp 1679581782
transform 1 0 53376 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_557
timestamp 1679581782
transform 1 0 54048 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_564
timestamp 1679581782
transform 1 0 54720 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_571
timestamp 1679581782
transform 1 0 55392 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_578
timestamp 1679581782
transform 1 0 56064 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_585
timestamp 1679581782
transform 1 0 56736 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_592
timestamp 1679581782
transform 1 0 57408 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_599
timestamp 1679581782
transform 1 0 58080 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_606
timestamp 1679581782
transform 1 0 58752 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_613
timestamp 1679581782
transform 1 0 59424 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_620
timestamp 1679581782
transform 1 0 60096 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_627
timestamp 1679581782
transform 1 0 60768 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_634
timestamp 1679581782
transform 1 0 61440 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_641
timestamp 1679581782
transform 1 0 62112 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_648
timestamp 1679581782
transform 1 0 62784 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_655
timestamp 1679581782
transform 1 0 63456 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_662
timestamp 1679581782
transform 1 0 64128 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_669
timestamp 1679581782
transform 1 0 64800 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_676
timestamp 1679581782
transform 1 0 65472 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_683
timestamp 1679581782
transform 1 0 66144 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_690
timestamp 1679581782
transform 1 0 66816 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_697
timestamp 1679581782
transform 1 0 67488 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_704
timestamp 1679581782
transform 1 0 68160 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_711
timestamp 1679581782
transform 1 0 68832 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_718
timestamp 1679581782
transform 1 0 69504 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_725
timestamp 1679581782
transform 1 0 70176 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_732
timestamp 1679581782
transform 1 0 70848 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_739
timestamp 1679581782
transform 1 0 71520 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_746
timestamp 1679581782
transform 1 0 72192 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_753
timestamp 1679581782
transform 1 0 72864 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_760
timestamp 1679581782
transform 1 0 73536 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_767
timestamp 1679581782
transform 1 0 74208 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_774
timestamp 1679581782
transform 1 0 74880 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_781
timestamp 1679581782
transform 1 0 75552 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_788
timestamp 1679581782
transform 1 0 76224 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_795
timestamp 1679581782
transform 1 0 76896 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_802
timestamp 1679581782
transform 1 0 77568 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_809
timestamp 1679581782
transform 1 0 78240 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_816
timestamp 1679581782
transform 1 0 78912 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_823
timestamp 1679581782
transform 1 0 79584 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_830
timestamp 1679581782
transform 1 0 80256 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_837
timestamp 1679581782
transform 1 0 80928 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_844
timestamp 1679581782
transform 1 0 81600 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_851
timestamp 1679581782
transform 1 0 82272 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_858
timestamp 1679581782
transform 1 0 82944 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_865
timestamp 1679581782
transform 1 0 83616 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_872
timestamp 1679581782
transform 1 0 84288 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_879
timestamp 1679581782
transform 1 0 84960 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_886
timestamp 1679581782
transform 1 0 85632 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_893
timestamp 1679581782
transform 1 0 86304 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_900
timestamp 1679581782
transform 1 0 86976 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_907
timestamp 1679581782
transform 1 0 87648 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_914
timestamp 1679581782
transform 1 0 88320 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_921
timestamp 1679581782
transform 1 0 88992 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_928
timestamp 1679581782
transform 1 0 89664 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_935
timestamp 1679581782
transform 1 0 90336 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_942
timestamp 1679581782
transform 1 0 91008 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_949
timestamp 1679581782
transform 1 0 91680 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_956
timestamp 1679581782
transform 1 0 92352 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_963
timestamp 1679581782
transform 1 0 93024 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_970
timestamp 1679581782
transform 1 0 93696 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_977
timestamp 1679581782
transform 1 0 94368 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_984
timestamp 1679581782
transform 1 0 95040 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_991
timestamp 1679581782
transform 1 0 95712 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_998
timestamp 1679581782
transform 1 0 96384 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_1005
timestamp 1679581782
transform 1 0 97056 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_1012
timestamp 1679581782
transform 1 0 97728 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_1019
timestamp 1679581782
transform 1 0 98400 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_39_1026
timestamp 1677580104
transform 1 0 99072 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_1028
timestamp 1677579658
transform 1 0 99264 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_0
timestamp 1679581782
transform 1 0 576 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_7
timestamp 1679581782
transform 1 0 1248 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_14
timestamp 1679581782
transform 1 0 1920 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_21
timestamp 1679581782
transform 1 0 2592 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_28
timestamp 1679581782
transform 1 0 3264 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_35
timestamp 1679581782
transform 1 0 3936 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_42
timestamp 1679581782
transform 1 0 4608 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_49
timestamp 1679581782
transform 1 0 5280 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_56
timestamp 1679581782
transform 1 0 5952 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_63
timestamp 1679581782
transform 1 0 6624 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_70
timestamp 1679581782
transform 1 0 7296 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_77
timestamp 1679581782
transform 1 0 7968 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_84
timestamp 1679581782
transform 1 0 8640 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_91
timestamp 1679581782
transform 1 0 9312 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_98
timestamp 1679581782
transform 1 0 9984 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_105
timestamp 1679581782
transform 1 0 10656 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_112
timestamp 1679581782
transform 1 0 11328 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_119
timestamp 1679581782
transform 1 0 12000 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_126
timestamp 1679581782
transform 1 0 12672 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_133
timestamp 1679581782
transform 1 0 13344 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_140
timestamp 1679581782
transform 1 0 14016 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_147
timestamp 1679581782
transform 1 0 14688 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_154
timestamp 1679581782
transform 1 0 15360 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_161
timestamp 1679581782
transform 1 0 16032 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_168
timestamp 1679581782
transform 1 0 16704 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_175
timestamp 1679581782
transform 1 0 17376 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_182
timestamp 1679581782
transform 1 0 18048 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_189
timestamp 1679581782
transform 1 0 18720 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_196
timestamp 1679581782
transform 1 0 19392 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_203
timestamp 1679581782
transform 1 0 20064 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_210
timestamp 1679581782
transform 1 0 20736 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_217
timestamp 1679581782
transform 1 0 21408 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_224
timestamp 1679581782
transform 1 0 22080 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_231
timestamp 1679581782
transform 1 0 22752 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_238
timestamp 1679581782
transform 1 0 23424 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_245
timestamp 1679581782
transform 1 0 24096 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_252
timestamp 1679581782
transform 1 0 24768 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_259
timestamp 1679581782
transform 1 0 25440 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_266
timestamp 1679581782
transform 1 0 26112 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_273
timestamp 1679581782
transform 1 0 26784 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_280
timestamp 1679581782
transform 1 0 27456 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_287
timestamp 1679581782
transform 1 0 28128 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_294
timestamp 1679581782
transform 1 0 28800 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_301
timestamp 1679581782
transform 1 0 29472 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_308
timestamp 1679581782
transform 1 0 30144 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_315
timestamp 1679581782
transform 1 0 30816 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_322
timestamp 1679581782
transform 1 0 31488 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_329
timestamp 1679581782
transform 1 0 32160 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_336
timestamp 1679581782
transform 1 0 32832 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_343
timestamp 1679581782
transform 1 0 33504 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_350
timestamp 1679581782
transform 1 0 34176 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_357
timestamp 1679581782
transform 1 0 34848 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_364
timestamp 1679581782
transform 1 0 35520 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_371
timestamp 1679581782
transform 1 0 36192 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_378
timestamp 1679581782
transform 1 0 36864 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_385
timestamp 1679581782
transform 1 0 37536 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_392
timestamp 1679581782
transform 1 0 38208 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_399
timestamp 1679581782
transform 1 0 38880 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_406
timestamp 1679581782
transform 1 0 39552 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_413
timestamp 1679581782
transform 1 0 40224 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_420
timestamp 1679581782
transform 1 0 40896 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_427
timestamp 1679581782
transform 1 0 41568 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_434
timestamp 1679581782
transform 1 0 42240 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_441
timestamp 1679581782
transform 1 0 42912 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_448
timestamp 1679581782
transform 1 0 43584 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_455
timestamp 1679581782
transform 1 0 44256 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_462
timestamp 1679581782
transform 1 0 44928 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_469
timestamp 1679581782
transform 1 0 45600 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_476
timestamp 1679581782
transform 1 0 46272 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_483
timestamp 1679581782
transform 1 0 46944 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_490
timestamp 1679581782
transform 1 0 47616 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_497
timestamp 1679581782
transform 1 0 48288 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_504
timestamp 1679581782
transform 1 0 48960 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_511
timestamp 1679581782
transform 1 0 49632 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_518
timestamp 1679581782
transform 1 0 50304 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_525
timestamp 1679581782
transform 1 0 50976 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_532
timestamp 1679581782
transform 1 0 51648 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_539
timestamp 1679581782
transform 1 0 52320 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_546
timestamp 1679581782
transform 1 0 52992 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_553
timestamp 1679581782
transform 1 0 53664 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_560
timestamp 1679581782
transform 1 0 54336 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_567
timestamp 1679581782
transform 1 0 55008 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_574
timestamp 1679581782
transform 1 0 55680 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_581
timestamp 1679581782
transform 1 0 56352 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_588
timestamp 1679581782
transform 1 0 57024 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_595
timestamp 1679581782
transform 1 0 57696 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_602
timestamp 1679581782
transform 1 0 58368 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_609
timestamp 1679581782
transform 1 0 59040 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_616
timestamp 1679581782
transform 1 0 59712 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_623
timestamp 1679581782
transform 1 0 60384 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_630
timestamp 1679581782
transform 1 0 61056 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_637
timestamp 1679581782
transform 1 0 61728 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_644
timestamp 1679581782
transform 1 0 62400 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_651
timestamp 1679581782
transform 1 0 63072 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_658
timestamp 1679581782
transform 1 0 63744 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_665
timestamp 1679581782
transform 1 0 64416 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_672
timestamp 1679581782
transform 1 0 65088 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_679
timestamp 1679581782
transform 1 0 65760 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_686
timestamp 1679581782
transform 1 0 66432 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_693
timestamp 1679581782
transform 1 0 67104 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_700
timestamp 1679581782
transform 1 0 67776 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_707
timestamp 1679581782
transform 1 0 68448 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_714
timestamp 1679581782
transform 1 0 69120 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_721
timestamp 1679581782
transform 1 0 69792 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_728
timestamp 1679581782
transform 1 0 70464 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_735
timestamp 1679581782
transform 1 0 71136 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_742
timestamp 1679581782
transform 1 0 71808 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_749
timestamp 1679581782
transform 1 0 72480 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_756
timestamp 1679581782
transform 1 0 73152 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_763
timestamp 1679581782
transform 1 0 73824 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_770
timestamp 1679581782
transform 1 0 74496 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_777
timestamp 1679581782
transform 1 0 75168 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_784
timestamp 1679581782
transform 1 0 75840 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_791
timestamp 1679581782
transform 1 0 76512 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_798
timestamp 1679581782
transform 1 0 77184 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_805
timestamp 1679581782
transform 1 0 77856 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_812
timestamp 1679581782
transform 1 0 78528 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_819
timestamp 1679581782
transform 1 0 79200 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_826
timestamp 1679581782
transform 1 0 79872 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_833
timestamp 1679581782
transform 1 0 80544 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_840
timestamp 1679581782
transform 1 0 81216 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_847
timestamp 1679581782
transform 1 0 81888 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_854
timestamp 1679581782
transform 1 0 82560 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_861
timestamp 1679581782
transform 1 0 83232 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_868
timestamp 1679581782
transform 1 0 83904 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_875
timestamp 1679581782
transform 1 0 84576 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_882
timestamp 1679581782
transform 1 0 85248 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_889
timestamp 1679581782
transform 1 0 85920 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_896
timestamp 1679581782
transform 1 0 86592 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_903
timestamp 1679581782
transform 1 0 87264 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_910
timestamp 1679581782
transform 1 0 87936 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_917
timestamp 1679581782
transform 1 0 88608 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_924
timestamp 1679581782
transform 1 0 89280 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_931
timestamp 1679581782
transform 1 0 89952 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_938
timestamp 1679581782
transform 1 0 90624 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_945
timestamp 1679581782
transform 1 0 91296 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_952
timestamp 1679581782
transform 1 0 91968 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_959
timestamp 1679581782
transform 1 0 92640 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_966
timestamp 1679581782
transform 1 0 93312 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_973
timestamp 1679581782
transform 1 0 93984 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_980
timestamp 1679581782
transform 1 0 94656 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_987
timestamp 1679581782
transform 1 0 95328 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_994
timestamp 1679581782
transform 1 0 96000 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_1001
timestamp 1679581782
transform 1 0 96672 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_1008
timestamp 1679581782
transform 1 0 97344 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_1015
timestamp 1679581782
transform 1 0 98016 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_1022
timestamp 1679581782
transform 1 0 98688 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_0
timestamp 1679581782
transform 1 0 576 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_7
timestamp 1679581782
transform 1 0 1248 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_14
timestamp 1679581782
transform 1 0 1920 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_21
timestamp 1679581782
transform 1 0 2592 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_28
timestamp 1679581782
transform 1 0 3264 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_35
timestamp 1679581782
transform 1 0 3936 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_42
timestamp 1679581782
transform 1 0 4608 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_49
timestamp 1679581782
transform 1 0 5280 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_56
timestamp 1679581782
transform 1 0 5952 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_63
timestamp 1679581782
transform 1 0 6624 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_70
timestamp 1679581782
transform 1 0 7296 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_77
timestamp 1679581782
transform 1 0 7968 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_84
timestamp 1679581782
transform 1 0 8640 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_91
timestamp 1679581782
transform 1 0 9312 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_98
timestamp 1679581782
transform 1 0 9984 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_105
timestamp 1679581782
transform 1 0 10656 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_112
timestamp 1679581782
transform 1 0 11328 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_119
timestamp 1679581782
transform 1 0 12000 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_126
timestamp 1679581782
transform 1 0 12672 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_133
timestamp 1679581782
transform 1 0 13344 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_140
timestamp 1679581782
transform 1 0 14016 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_147
timestamp 1679581782
transform 1 0 14688 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_154
timestamp 1679581782
transform 1 0 15360 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_161
timestamp 1679581782
transform 1 0 16032 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_168
timestamp 1679581782
transform 1 0 16704 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_175
timestamp 1679581782
transform 1 0 17376 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_182
timestamp 1679581782
transform 1 0 18048 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_189
timestamp 1679581782
transform 1 0 18720 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_196
timestamp 1679581782
transform 1 0 19392 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_203
timestamp 1679581782
transform 1 0 20064 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_210
timestamp 1679581782
transform 1 0 20736 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_217
timestamp 1679581782
transform 1 0 21408 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_224
timestamp 1679581782
transform 1 0 22080 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_231
timestamp 1679581782
transform 1 0 22752 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_238
timestamp 1679581782
transform 1 0 23424 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_245
timestamp 1679581782
transform 1 0 24096 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_252
timestamp 1679581782
transform 1 0 24768 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_259
timestamp 1679581782
transform 1 0 25440 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_266
timestamp 1679581782
transform 1 0 26112 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_273
timestamp 1679581782
transform 1 0 26784 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_280
timestamp 1679581782
transform 1 0 27456 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_287
timestamp 1679581782
transform 1 0 28128 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_294
timestamp 1679581782
transform 1 0 28800 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_301
timestamp 1679581782
transform 1 0 29472 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_308
timestamp 1679581782
transform 1 0 30144 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_315
timestamp 1679581782
transform 1 0 30816 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_322
timestamp 1679581782
transform 1 0 31488 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_329
timestamp 1679581782
transform 1 0 32160 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_336
timestamp 1679581782
transform 1 0 32832 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_343
timestamp 1679581782
transform 1 0 33504 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_350
timestamp 1679581782
transform 1 0 34176 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_357
timestamp 1679581782
transform 1 0 34848 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_364
timestamp 1679581782
transform 1 0 35520 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_371
timestamp 1679581782
transform 1 0 36192 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_378
timestamp 1679581782
transform 1 0 36864 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_385
timestamp 1679581782
transform 1 0 37536 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_392
timestamp 1679581782
transform 1 0 38208 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_399
timestamp 1679581782
transform 1 0 38880 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_406
timestamp 1679581782
transform 1 0 39552 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_413
timestamp 1679581782
transform 1 0 40224 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_420
timestamp 1679581782
transform 1 0 40896 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_427
timestamp 1679581782
transform 1 0 41568 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_434
timestamp 1679581782
transform 1 0 42240 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_441
timestamp 1679581782
transform 1 0 42912 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_448
timestamp 1679581782
transform 1 0 43584 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_455
timestamp 1679581782
transform 1 0 44256 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_462
timestamp 1679581782
transform 1 0 44928 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_469
timestamp 1679581782
transform 1 0 45600 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_476
timestamp 1679581782
transform 1 0 46272 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_483
timestamp 1679581782
transform 1 0 46944 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_490
timestamp 1679581782
transform 1 0 47616 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_497
timestamp 1679581782
transform 1 0 48288 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_504
timestamp 1679581782
transform 1 0 48960 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_511
timestamp 1679581782
transform 1 0 49632 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_518
timestamp 1679581782
transform 1 0 50304 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_525
timestamp 1679581782
transform 1 0 50976 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_532
timestamp 1679581782
transform 1 0 51648 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_539
timestamp 1679581782
transform 1 0 52320 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_546
timestamp 1679581782
transform 1 0 52992 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_553
timestamp 1679581782
transform 1 0 53664 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_560
timestamp 1679581782
transform 1 0 54336 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_567
timestamp 1679581782
transform 1 0 55008 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_574
timestamp 1679581782
transform 1 0 55680 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_581
timestamp 1679581782
transform 1 0 56352 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_588
timestamp 1679581782
transform 1 0 57024 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_595
timestamp 1679581782
transform 1 0 57696 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_602
timestamp 1679581782
transform 1 0 58368 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_609
timestamp 1679581782
transform 1 0 59040 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_616
timestamp 1679581782
transform 1 0 59712 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_623
timestamp 1679581782
transform 1 0 60384 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_630
timestamp 1679581782
transform 1 0 61056 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_637
timestamp 1679581782
transform 1 0 61728 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_644
timestamp 1679581782
transform 1 0 62400 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_651
timestamp 1679581782
transform 1 0 63072 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_658
timestamp 1679581782
transform 1 0 63744 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_665
timestamp 1679581782
transform 1 0 64416 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_672
timestamp 1679581782
transform 1 0 65088 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_679
timestamp 1679581782
transform 1 0 65760 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_686
timestamp 1679581782
transform 1 0 66432 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_693
timestamp 1679581782
transform 1 0 67104 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_700
timestamp 1679581782
transform 1 0 67776 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_707
timestamp 1679581782
transform 1 0 68448 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_714
timestamp 1679581782
transform 1 0 69120 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_721
timestamp 1679581782
transform 1 0 69792 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_728
timestamp 1679581782
transform 1 0 70464 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_735
timestamp 1679581782
transform 1 0 71136 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_742
timestamp 1679581782
transform 1 0 71808 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_749
timestamp 1679581782
transform 1 0 72480 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_756
timestamp 1679581782
transform 1 0 73152 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_763
timestamp 1679581782
transform 1 0 73824 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_770
timestamp 1679581782
transform 1 0 74496 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_777
timestamp 1679581782
transform 1 0 75168 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_784
timestamp 1679581782
transform 1 0 75840 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_791
timestamp 1679581782
transform 1 0 76512 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_798
timestamp 1679581782
transform 1 0 77184 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_805
timestamp 1679581782
transform 1 0 77856 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_812
timestamp 1679581782
transform 1 0 78528 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_819
timestamp 1679581782
transform 1 0 79200 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_826
timestamp 1679581782
transform 1 0 79872 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_833
timestamp 1679581782
transform 1 0 80544 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_840
timestamp 1679581782
transform 1 0 81216 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_847
timestamp 1679581782
transform 1 0 81888 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_854
timestamp 1679581782
transform 1 0 82560 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_861
timestamp 1679581782
transform 1 0 83232 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_868
timestamp 1679581782
transform 1 0 83904 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_875
timestamp 1679581782
transform 1 0 84576 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_882
timestamp 1679581782
transform 1 0 85248 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_889
timestamp 1679581782
transform 1 0 85920 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_896
timestamp 1679581782
transform 1 0 86592 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_903
timestamp 1679581782
transform 1 0 87264 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_910
timestamp 1679581782
transform 1 0 87936 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_917
timestamp 1679581782
transform 1 0 88608 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_924
timestamp 1679581782
transform 1 0 89280 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_931
timestamp 1679581782
transform 1 0 89952 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_938
timestamp 1679581782
transform 1 0 90624 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_945
timestamp 1679581782
transform 1 0 91296 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_952
timestamp 1679581782
transform 1 0 91968 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_959
timestamp 1679581782
transform 1 0 92640 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_966
timestamp 1679581782
transform 1 0 93312 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_973
timestamp 1679581782
transform 1 0 93984 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_980
timestamp 1679581782
transform 1 0 94656 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_987
timestamp 1679581782
transform 1 0 95328 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_994
timestamp 1679581782
transform 1 0 96000 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_1001
timestamp 1679581782
transform 1 0 96672 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_1008
timestamp 1679581782
transform 1 0 97344 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_1015
timestamp 1679581782
transform 1 0 98016 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_1022
timestamp 1679581782
transform 1 0 98688 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_4
timestamp 1679581782
transform 1 0 960 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_11
timestamp 1679581782
transform 1 0 1632 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_18
timestamp 1679581782
transform 1 0 2304 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_25
timestamp 1679581782
transform 1 0 2976 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_32
timestamp 1679581782
transform 1 0 3648 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_39
timestamp 1679581782
transform 1 0 4320 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_46
timestamp 1679581782
transform 1 0 4992 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_53
timestamp 1679581782
transform 1 0 5664 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_60
timestamp 1679581782
transform 1 0 6336 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_67
timestamp 1679581782
transform 1 0 7008 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_74
timestamp 1679581782
transform 1 0 7680 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_81
timestamp 1679581782
transform 1 0 8352 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_88
timestamp 1679581782
transform 1 0 9024 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_95
timestamp 1679581782
transform 1 0 9696 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_102
timestamp 1679581782
transform 1 0 10368 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_109
timestamp 1679581782
transform 1 0 11040 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_116
timestamp 1679581782
transform 1 0 11712 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_123
timestamp 1679581782
transform 1 0 12384 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_130
timestamp 1679581782
transform 1 0 13056 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_137
timestamp 1679581782
transform 1 0 13728 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_144
timestamp 1679581782
transform 1 0 14400 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_151
timestamp 1679581782
transform 1 0 15072 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_158
timestamp 1679581782
transform 1 0 15744 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_165
timestamp 1679581782
transform 1 0 16416 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_172
timestamp 1679581782
transform 1 0 17088 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_179
timestamp 1679581782
transform 1 0 17760 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_186
timestamp 1679581782
transform 1 0 18432 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_193
timestamp 1679581782
transform 1 0 19104 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_200
timestamp 1679581782
transform 1 0 19776 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_207
timestamp 1679581782
transform 1 0 20448 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_214
timestamp 1679581782
transform 1 0 21120 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_221
timestamp 1679581782
transform 1 0 21792 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_228
timestamp 1679581782
transform 1 0 22464 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_235
timestamp 1679581782
transform 1 0 23136 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_242
timestamp 1679581782
transform 1 0 23808 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_249
timestamp 1679581782
transform 1 0 24480 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_256
timestamp 1679581782
transform 1 0 25152 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_263
timestamp 1679581782
transform 1 0 25824 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_270
timestamp 1679581782
transform 1 0 26496 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_277
timestamp 1679581782
transform 1 0 27168 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_284
timestamp 1679581782
transform 1 0 27840 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_291
timestamp 1679581782
transform 1 0 28512 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_298
timestamp 1679581782
transform 1 0 29184 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_305
timestamp 1679581782
transform 1 0 29856 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_312
timestamp 1679581782
transform 1 0 30528 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_319
timestamp 1679581782
transform 1 0 31200 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_326
timestamp 1679581782
transform 1 0 31872 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_333
timestamp 1679581782
transform 1 0 32544 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_340
timestamp 1679581782
transform 1 0 33216 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_347
timestamp 1679581782
transform 1 0 33888 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_354
timestamp 1679581782
transform 1 0 34560 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_361
timestamp 1679581782
transform 1 0 35232 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_368
timestamp 1679581782
transform 1 0 35904 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_375
timestamp 1679581782
transform 1 0 36576 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_382
timestamp 1679581782
transform 1 0 37248 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_389
timestamp 1679581782
transform 1 0 37920 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_396
timestamp 1679581782
transform 1 0 38592 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_403
timestamp 1679581782
transform 1 0 39264 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_410
timestamp 1679581782
transform 1 0 39936 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_417
timestamp 1679581782
transform 1 0 40608 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_424
timestamp 1679581782
transform 1 0 41280 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_431
timestamp 1679581782
transform 1 0 41952 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_438
timestamp 1679581782
transform 1 0 42624 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_445
timestamp 1679581782
transform 1 0 43296 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_452
timestamp 1679581782
transform 1 0 43968 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_459
timestamp 1679581782
transform 1 0 44640 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_466
timestamp 1679581782
transform 1 0 45312 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_473
timestamp 1679581782
transform 1 0 45984 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_480
timestamp 1679581782
transform 1 0 46656 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_487
timestamp 1679581782
transform 1 0 47328 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_494
timestamp 1679581782
transform 1 0 48000 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_501
timestamp 1679581782
transform 1 0 48672 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_508
timestamp 1679581782
transform 1 0 49344 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_515
timestamp 1679581782
transform 1 0 50016 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_522
timestamp 1679581782
transform 1 0 50688 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_529
timestamp 1679581782
transform 1 0 51360 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_536
timestamp 1679581782
transform 1 0 52032 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_543
timestamp 1679581782
transform 1 0 52704 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_550
timestamp 1679581782
transform 1 0 53376 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_557
timestamp 1679581782
transform 1 0 54048 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_564
timestamp 1679581782
transform 1 0 54720 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_571
timestamp 1679581782
transform 1 0 55392 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_578
timestamp 1679581782
transform 1 0 56064 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_585
timestamp 1679581782
transform 1 0 56736 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_592
timestamp 1679581782
transform 1 0 57408 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_599
timestamp 1679581782
transform 1 0 58080 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_606
timestamp 1679581782
transform 1 0 58752 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_613
timestamp 1679581782
transform 1 0 59424 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_620
timestamp 1679581782
transform 1 0 60096 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_627
timestamp 1679581782
transform 1 0 60768 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_634
timestamp 1679581782
transform 1 0 61440 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_641
timestamp 1679581782
transform 1 0 62112 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_648
timestamp 1679581782
transform 1 0 62784 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_655
timestamp 1679581782
transform 1 0 63456 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_662
timestamp 1679581782
transform 1 0 64128 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_669
timestamp 1679581782
transform 1 0 64800 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_676
timestamp 1679581782
transform 1 0 65472 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_683
timestamp 1679581782
transform 1 0 66144 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_690
timestamp 1679581782
transform 1 0 66816 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_697
timestamp 1679581782
transform 1 0 67488 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_704
timestamp 1679581782
transform 1 0 68160 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_711
timestamp 1679581782
transform 1 0 68832 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_718
timestamp 1679581782
transform 1 0 69504 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_725
timestamp 1679581782
transform 1 0 70176 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_732
timestamp 1679581782
transform 1 0 70848 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_739
timestamp 1679581782
transform 1 0 71520 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_746
timestamp 1679581782
transform 1 0 72192 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_753
timestamp 1679581782
transform 1 0 72864 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_760
timestamp 1679581782
transform 1 0 73536 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_767
timestamp 1679581782
transform 1 0 74208 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_774
timestamp 1679581782
transform 1 0 74880 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_781
timestamp 1679581782
transform 1 0 75552 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_788
timestamp 1679581782
transform 1 0 76224 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_795
timestamp 1679581782
transform 1 0 76896 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_802
timestamp 1679581782
transform 1 0 77568 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_809
timestamp 1679581782
transform 1 0 78240 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_816
timestamp 1679581782
transform 1 0 78912 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_823
timestamp 1679581782
transform 1 0 79584 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_830
timestamp 1679581782
transform 1 0 80256 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_837
timestamp 1679581782
transform 1 0 80928 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_844
timestamp 1679581782
transform 1 0 81600 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_851
timestamp 1679581782
transform 1 0 82272 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_858
timestamp 1679581782
transform 1 0 82944 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_865
timestamp 1679581782
transform 1 0 83616 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_872
timestamp 1679581782
transform 1 0 84288 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_879
timestamp 1679581782
transform 1 0 84960 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_886
timestamp 1679581782
transform 1 0 85632 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_893
timestamp 1679581782
transform 1 0 86304 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_900
timestamp 1679581782
transform 1 0 86976 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_907
timestamp 1679581782
transform 1 0 87648 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_914
timestamp 1679581782
transform 1 0 88320 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_921
timestamp 1679581782
transform 1 0 88992 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_928
timestamp 1679581782
transform 1 0 89664 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_935
timestamp 1679581782
transform 1 0 90336 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_942
timestamp 1679581782
transform 1 0 91008 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_949
timestamp 1679581782
transform 1 0 91680 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_956
timestamp 1679581782
transform 1 0 92352 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_963
timestamp 1679581782
transform 1 0 93024 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_970
timestamp 1679581782
transform 1 0 93696 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_977
timestamp 1679581782
transform 1 0 94368 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_984
timestamp 1679581782
transform 1 0 95040 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_991
timestamp 1679581782
transform 1 0 95712 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_998
timestamp 1679581782
transform 1 0 96384 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_1005
timestamp 1679581782
transform 1 0 97056 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_1012
timestamp 1679581782
transform 1 0 97728 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_1019
timestamp 1679581782
transform 1 0 98400 0 1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_42_1026
timestamp 1677580104
transform 1 0 99072 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_1028
timestamp 1677579658
transform 1 0 99264 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_0
timestamp 1679581782
transform 1 0 576 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_7
timestamp 1679581782
transform 1 0 1248 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_14
timestamp 1679581782
transform 1 0 1920 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_21
timestamp 1679581782
transform 1 0 2592 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_28
timestamp 1679581782
transform 1 0 3264 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_35
timestamp 1679581782
transform 1 0 3936 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_42
timestamp 1679581782
transform 1 0 4608 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_49
timestamp 1679581782
transform 1 0 5280 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_56
timestamp 1679581782
transform 1 0 5952 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_63
timestamp 1679581782
transform 1 0 6624 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_70
timestamp 1679581782
transform 1 0 7296 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_77
timestamp 1679581782
transform 1 0 7968 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_84
timestamp 1679581782
transform 1 0 8640 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_91
timestamp 1679581782
transform 1 0 9312 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_98
timestamp 1679581782
transform 1 0 9984 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_105
timestamp 1679581782
transform 1 0 10656 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_112
timestamp 1679581782
transform 1 0 11328 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_119
timestamp 1679581782
transform 1 0 12000 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_126
timestamp 1679581782
transform 1 0 12672 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_133
timestamp 1679581782
transform 1 0 13344 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_140
timestamp 1679581782
transform 1 0 14016 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_147
timestamp 1679581782
transform 1 0 14688 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_154
timestamp 1679581782
transform 1 0 15360 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_161
timestamp 1679581782
transform 1 0 16032 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_168
timestamp 1679581782
transform 1 0 16704 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_175
timestamp 1679581782
transform 1 0 17376 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_182
timestamp 1679581782
transform 1 0 18048 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_189
timestamp 1679581782
transform 1 0 18720 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_196
timestamp 1679581782
transform 1 0 19392 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_203
timestamp 1679581782
transform 1 0 20064 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_210
timestamp 1679581782
transform 1 0 20736 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_217
timestamp 1679581782
transform 1 0 21408 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_224
timestamp 1679581782
transform 1 0 22080 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_231
timestamp 1679581782
transform 1 0 22752 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_238
timestamp 1679581782
transform 1 0 23424 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_245
timestamp 1679581782
transform 1 0 24096 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_252
timestamp 1679581782
transform 1 0 24768 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_259
timestamp 1679581782
transform 1 0 25440 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_266
timestamp 1679581782
transform 1 0 26112 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_273
timestamp 1679581782
transform 1 0 26784 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_280
timestamp 1679581782
transform 1 0 27456 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_287
timestamp 1679581782
transform 1 0 28128 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_294
timestamp 1679581782
transform 1 0 28800 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_301
timestamp 1679581782
transform 1 0 29472 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_308
timestamp 1679581782
transform 1 0 30144 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_315
timestamp 1679581782
transform 1 0 30816 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_322
timestamp 1679581782
transform 1 0 31488 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_329
timestamp 1679581782
transform 1 0 32160 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_336
timestamp 1679581782
transform 1 0 32832 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_343
timestamp 1679581782
transform 1 0 33504 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_350
timestamp 1679581782
transform 1 0 34176 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_357
timestamp 1679581782
transform 1 0 34848 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_364
timestamp 1679581782
transform 1 0 35520 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_371
timestamp 1679581782
transform 1 0 36192 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_378
timestamp 1679581782
transform 1 0 36864 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_385
timestamp 1679581782
transform 1 0 37536 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_392
timestamp 1679581782
transform 1 0 38208 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_399
timestamp 1679581782
transform 1 0 38880 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_406
timestamp 1679581782
transform 1 0 39552 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_413
timestamp 1679581782
transform 1 0 40224 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_420
timestamp 1679581782
transform 1 0 40896 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_427
timestamp 1679581782
transform 1 0 41568 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_434
timestamp 1679581782
transform 1 0 42240 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_441
timestamp 1679581782
transform 1 0 42912 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_448
timestamp 1679581782
transform 1 0 43584 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_455
timestamp 1679581782
transform 1 0 44256 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_462
timestamp 1679581782
transform 1 0 44928 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_469
timestamp 1679581782
transform 1 0 45600 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_476
timestamp 1679581782
transform 1 0 46272 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_483
timestamp 1679581782
transform 1 0 46944 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_490
timestamp 1679581782
transform 1 0 47616 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_497
timestamp 1679581782
transform 1 0 48288 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_504
timestamp 1679581782
transform 1 0 48960 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_511
timestamp 1679581782
transform 1 0 49632 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_518
timestamp 1679581782
transform 1 0 50304 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_525
timestamp 1679581782
transform 1 0 50976 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_532
timestamp 1679581782
transform 1 0 51648 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_539
timestamp 1679581782
transform 1 0 52320 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_546
timestamp 1679581782
transform 1 0 52992 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_553
timestamp 1679581782
transform 1 0 53664 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_560
timestamp 1679581782
transform 1 0 54336 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_567
timestamp 1679581782
transform 1 0 55008 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_574
timestamp 1679581782
transform 1 0 55680 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_581
timestamp 1679581782
transform 1 0 56352 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_588
timestamp 1679581782
transform 1 0 57024 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_595
timestamp 1679581782
transform 1 0 57696 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_602
timestamp 1679581782
transform 1 0 58368 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_609
timestamp 1679581782
transform 1 0 59040 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_616
timestamp 1679581782
transform 1 0 59712 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_623
timestamp 1679581782
transform 1 0 60384 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_630
timestamp 1679581782
transform 1 0 61056 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_637
timestamp 1679581782
transform 1 0 61728 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_644
timestamp 1679581782
transform 1 0 62400 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_651
timestamp 1679581782
transform 1 0 63072 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_658
timestamp 1679581782
transform 1 0 63744 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_665
timestamp 1679581782
transform 1 0 64416 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_672
timestamp 1679581782
transform 1 0 65088 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_679
timestamp 1679581782
transform 1 0 65760 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_686
timestamp 1679581782
transform 1 0 66432 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_693
timestamp 1679581782
transform 1 0 67104 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_700
timestamp 1679581782
transform 1 0 67776 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_707
timestamp 1679581782
transform 1 0 68448 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_714
timestamp 1679581782
transform 1 0 69120 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_721
timestamp 1679581782
transform 1 0 69792 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_728
timestamp 1679581782
transform 1 0 70464 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_735
timestamp 1679581782
transform 1 0 71136 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_742
timestamp 1679581782
transform 1 0 71808 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_749
timestamp 1679581782
transform 1 0 72480 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_756
timestamp 1679581782
transform 1 0 73152 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_763
timestamp 1679581782
transform 1 0 73824 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_770
timestamp 1679581782
transform 1 0 74496 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_777
timestamp 1679581782
transform 1 0 75168 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_784
timestamp 1679581782
transform 1 0 75840 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_791
timestamp 1679581782
transform 1 0 76512 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_798
timestamp 1679581782
transform 1 0 77184 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_805
timestamp 1679581782
transform 1 0 77856 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_812
timestamp 1679581782
transform 1 0 78528 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_819
timestamp 1679581782
transform 1 0 79200 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_826
timestamp 1679581782
transform 1 0 79872 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_833
timestamp 1679581782
transform 1 0 80544 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_840
timestamp 1679581782
transform 1 0 81216 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_847
timestamp 1679581782
transform 1 0 81888 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_854
timestamp 1679581782
transform 1 0 82560 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_861
timestamp 1679581782
transform 1 0 83232 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_868
timestamp 1679581782
transform 1 0 83904 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_875
timestamp 1679581782
transform 1 0 84576 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_882
timestamp 1679581782
transform 1 0 85248 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_889
timestamp 1679581782
transform 1 0 85920 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_896
timestamp 1679581782
transform 1 0 86592 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_903
timestamp 1679581782
transform 1 0 87264 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_910
timestamp 1679581782
transform 1 0 87936 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_917
timestamp 1679581782
transform 1 0 88608 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_924
timestamp 1679581782
transform 1 0 89280 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_931
timestamp 1679581782
transform 1 0 89952 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_938
timestamp 1679581782
transform 1 0 90624 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_945
timestamp 1679581782
transform 1 0 91296 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_952
timestamp 1679581782
transform 1 0 91968 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_959
timestamp 1679581782
transform 1 0 92640 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_966
timestamp 1679581782
transform 1 0 93312 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_973
timestamp 1679581782
transform 1 0 93984 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_980
timestamp 1679581782
transform 1 0 94656 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_987
timestamp 1679581782
transform 1 0 95328 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_994
timestamp 1679581782
transform 1 0 96000 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_1001
timestamp 1679581782
transform 1 0 96672 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_1008
timestamp 1679581782
transform 1 0 97344 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_1015
timestamp 1679581782
transform 1 0 98016 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_1022
timestamp 1679581782
transform 1 0 98688 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_4
timestamp 1679581782
transform 1 0 960 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_11
timestamp 1679581782
transform 1 0 1632 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_18
timestamp 1679581782
transform 1 0 2304 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_25
timestamp 1679581782
transform 1 0 2976 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_32
timestamp 1679581782
transform 1 0 3648 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_39
timestamp 1679581782
transform 1 0 4320 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_46
timestamp 1679581782
transform 1 0 4992 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_53
timestamp 1679581782
transform 1 0 5664 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_60
timestamp 1679581782
transform 1 0 6336 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_67
timestamp 1679581782
transform 1 0 7008 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_74
timestamp 1679581782
transform 1 0 7680 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_81
timestamp 1679581782
transform 1 0 8352 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_88
timestamp 1679581782
transform 1 0 9024 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_95
timestamp 1679581782
transform 1 0 9696 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_102
timestamp 1679581782
transform 1 0 10368 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_109
timestamp 1679581782
transform 1 0 11040 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_116
timestamp 1679581782
transform 1 0 11712 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_123
timestamp 1679581782
transform 1 0 12384 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_130
timestamp 1679581782
transform 1 0 13056 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_137
timestamp 1679581782
transform 1 0 13728 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_144
timestamp 1679581782
transform 1 0 14400 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_151
timestamp 1679581782
transform 1 0 15072 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_158
timestamp 1679581782
transform 1 0 15744 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_165
timestamp 1679581782
transform 1 0 16416 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_172
timestamp 1679581782
transform 1 0 17088 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_179
timestamp 1679581782
transform 1 0 17760 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_186
timestamp 1679581782
transform 1 0 18432 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_193
timestamp 1679581782
transform 1 0 19104 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_200
timestamp 1679581782
transform 1 0 19776 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_207
timestamp 1679581782
transform 1 0 20448 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_214
timestamp 1679581782
transform 1 0 21120 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_221
timestamp 1679581782
transform 1 0 21792 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_228
timestamp 1679581782
transform 1 0 22464 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_235
timestamp 1679581782
transform 1 0 23136 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_242
timestamp 1679581782
transform 1 0 23808 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_249
timestamp 1679581782
transform 1 0 24480 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_256
timestamp 1679581782
transform 1 0 25152 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_263
timestamp 1679581782
transform 1 0 25824 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_270
timestamp 1679581782
transform 1 0 26496 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_277
timestamp 1679581782
transform 1 0 27168 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_284
timestamp 1679581782
transform 1 0 27840 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_291
timestamp 1679581782
transform 1 0 28512 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_298
timestamp 1679581782
transform 1 0 29184 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_305
timestamp 1679581782
transform 1 0 29856 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_312
timestamp 1679581782
transform 1 0 30528 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_319
timestamp 1679581782
transform 1 0 31200 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_326
timestamp 1679581782
transform 1 0 31872 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_333
timestamp 1679581782
transform 1 0 32544 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_340
timestamp 1679581782
transform 1 0 33216 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_347
timestamp 1679581782
transform 1 0 33888 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_354
timestamp 1679581782
transform 1 0 34560 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_361
timestamp 1679581782
transform 1 0 35232 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_368
timestamp 1679581782
transform 1 0 35904 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_375
timestamp 1679581782
transform 1 0 36576 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_382
timestamp 1679581782
transform 1 0 37248 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_389
timestamp 1679581782
transform 1 0 37920 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_396
timestamp 1679581782
transform 1 0 38592 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_403
timestamp 1679581782
transform 1 0 39264 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_410
timestamp 1679581782
transform 1 0 39936 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_417
timestamp 1679581782
transform 1 0 40608 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_424
timestamp 1679581782
transform 1 0 41280 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_431
timestamp 1679581782
transform 1 0 41952 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_438
timestamp 1679581782
transform 1 0 42624 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_445
timestamp 1679581782
transform 1 0 43296 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_452
timestamp 1679581782
transform 1 0 43968 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_459
timestamp 1679581782
transform 1 0 44640 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_466
timestamp 1679581782
transform 1 0 45312 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_473
timestamp 1679581782
transform 1 0 45984 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_480
timestamp 1679581782
transform 1 0 46656 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_487
timestamp 1679581782
transform 1 0 47328 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_494
timestamp 1679581782
transform 1 0 48000 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_501
timestamp 1679581782
transform 1 0 48672 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_508
timestamp 1679581782
transform 1 0 49344 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_515
timestamp 1679581782
transform 1 0 50016 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_522
timestamp 1679581782
transform 1 0 50688 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_529
timestamp 1679581782
transform 1 0 51360 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_536
timestamp 1679581782
transform 1 0 52032 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_543
timestamp 1679581782
transform 1 0 52704 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_550
timestamp 1679581782
transform 1 0 53376 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_557
timestamp 1679581782
transform 1 0 54048 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_564
timestamp 1679581782
transform 1 0 54720 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_571
timestamp 1679581782
transform 1 0 55392 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_578
timestamp 1679581782
transform 1 0 56064 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_585
timestamp 1679581782
transform 1 0 56736 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_592
timestamp 1679581782
transform 1 0 57408 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_599
timestamp 1679581782
transform 1 0 58080 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_606
timestamp 1679581782
transform 1 0 58752 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_613
timestamp 1679581782
transform 1 0 59424 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_620
timestamp 1679581782
transform 1 0 60096 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_627
timestamp 1679581782
transform 1 0 60768 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_634
timestamp 1679581782
transform 1 0 61440 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_641
timestamp 1679581782
transform 1 0 62112 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_648
timestamp 1679581782
transform 1 0 62784 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_655
timestamp 1679581782
transform 1 0 63456 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_662
timestamp 1679581782
transform 1 0 64128 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_669
timestamp 1679581782
transform 1 0 64800 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_676
timestamp 1679581782
transform 1 0 65472 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_683
timestamp 1679581782
transform 1 0 66144 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_690
timestamp 1679581782
transform 1 0 66816 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_697
timestamp 1679581782
transform 1 0 67488 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_704
timestamp 1679581782
transform 1 0 68160 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_711
timestamp 1679581782
transform 1 0 68832 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_718
timestamp 1679581782
transform 1 0 69504 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_725
timestamp 1679581782
transform 1 0 70176 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_732
timestamp 1679581782
transform 1 0 70848 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_739
timestamp 1679581782
transform 1 0 71520 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_746
timestamp 1679581782
transform 1 0 72192 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_753
timestamp 1679581782
transform 1 0 72864 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_760
timestamp 1679581782
transform 1 0 73536 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_767
timestamp 1679581782
transform 1 0 74208 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_774
timestamp 1679581782
transform 1 0 74880 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_781
timestamp 1679581782
transform 1 0 75552 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_788
timestamp 1679581782
transform 1 0 76224 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_795
timestamp 1679581782
transform 1 0 76896 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_802
timestamp 1679581782
transform 1 0 77568 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_809
timestamp 1679581782
transform 1 0 78240 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_816
timestamp 1679581782
transform 1 0 78912 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_823
timestamp 1679581782
transform 1 0 79584 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_830
timestamp 1679581782
transform 1 0 80256 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_837
timestamp 1679581782
transform 1 0 80928 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_844
timestamp 1679581782
transform 1 0 81600 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_851
timestamp 1679581782
transform 1 0 82272 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_858
timestamp 1679581782
transform 1 0 82944 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_865
timestamp 1679581782
transform 1 0 83616 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_872
timestamp 1679581782
transform 1 0 84288 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_879
timestamp 1679581782
transform 1 0 84960 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_886
timestamp 1679581782
transform 1 0 85632 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_893
timestamp 1679581782
transform 1 0 86304 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_900
timestamp 1679581782
transform 1 0 86976 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_907
timestamp 1679581782
transform 1 0 87648 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_914
timestamp 1679581782
transform 1 0 88320 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_921
timestamp 1679581782
transform 1 0 88992 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_928
timestamp 1679581782
transform 1 0 89664 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_935
timestamp 1679581782
transform 1 0 90336 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_942
timestamp 1679581782
transform 1 0 91008 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_949
timestamp 1679581782
transform 1 0 91680 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_956
timestamp 1679581782
transform 1 0 92352 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_963
timestamp 1679581782
transform 1 0 93024 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_970
timestamp 1679581782
transform 1 0 93696 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_977
timestamp 1679581782
transform 1 0 94368 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_984
timestamp 1679581782
transform 1 0 95040 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_991
timestamp 1679581782
transform 1 0 95712 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_998
timestamp 1679581782
transform 1 0 96384 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_1005
timestamp 1679581782
transform 1 0 97056 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_1012
timestamp 1679581782
transform 1 0 97728 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_1019
timestamp 1679581782
transform 1 0 98400 0 1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_44_1026
timestamp 1677580104
transform 1 0 99072 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_1028
timestamp 1677579658
transform 1 0 99264 0 1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_45_0
timestamp 1679581782
transform 1 0 576 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_7
timestamp 1679581782
transform 1 0 1248 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_14
timestamp 1679581782
transform 1 0 1920 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_21
timestamp 1679581782
transform 1 0 2592 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_28
timestamp 1679581782
transform 1 0 3264 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_35
timestamp 1679581782
transform 1 0 3936 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_42
timestamp 1679581782
transform 1 0 4608 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_49
timestamp 1679581782
transform 1 0 5280 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_56
timestamp 1679581782
transform 1 0 5952 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_63
timestamp 1679581782
transform 1 0 6624 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_70
timestamp 1679581782
transform 1 0 7296 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_77
timestamp 1679581782
transform 1 0 7968 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_84
timestamp 1679581782
transform 1 0 8640 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_91
timestamp 1679581782
transform 1 0 9312 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_98
timestamp 1679581782
transform 1 0 9984 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_105
timestamp 1679581782
transform 1 0 10656 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_112
timestamp 1679581782
transform 1 0 11328 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_119
timestamp 1679581782
transform 1 0 12000 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_126
timestamp 1679581782
transform 1 0 12672 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_133
timestamp 1679581782
transform 1 0 13344 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_140
timestamp 1679581782
transform 1 0 14016 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_147
timestamp 1679581782
transform 1 0 14688 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_154
timestamp 1679581782
transform 1 0 15360 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_161
timestamp 1679581782
transform 1 0 16032 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_168
timestamp 1679581782
transform 1 0 16704 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_175
timestamp 1679581782
transform 1 0 17376 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_182
timestamp 1679581782
transform 1 0 18048 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_189
timestamp 1679581782
transform 1 0 18720 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_196
timestamp 1679581782
transform 1 0 19392 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_203
timestamp 1679581782
transform 1 0 20064 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_210
timestamp 1679581782
transform 1 0 20736 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_217
timestamp 1679581782
transform 1 0 21408 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_224
timestamp 1679581782
transform 1 0 22080 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_231
timestamp 1679581782
transform 1 0 22752 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_238
timestamp 1679581782
transform 1 0 23424 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_245
timestamp 1679581782
transform 1 0 24096 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_252
timestamp 1679581782
transform 1 0 24768 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_259
timestamp 1679581782
transform 1 0 25440 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_266
timestamp 1679581782
transform 1 0 26112 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_273
timestamp 1679581782
transform 1 0 26784 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_280
timestamp 1679581782
transform 1 0 27456 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_287
timestamp 1679581782
transform 1 0 28128 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_294
timestamp 1679581782
transform 1 0 28800 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_301
timestamp 1679581782
transform 1 0 29472 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_308
timestamp 1679581782
transform 1 0 30144 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_315
timestamp 1679581782
transform 1 0 30816 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_322
timestamp 1679581782
transform 1 0 31488 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_329
timestamp 1679581782
transform 1 0 32160 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_336
timestamp 1679581782
transform 1 0 32832 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_343
timestamp 1679581782
transform 1 0 33504 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_350
timestamp 1679581782
transform 1 0 34176 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_357
timestamp 1679581782
transform 1 0 34848 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_364
timestamp 1679581782
transform 1 0 35520 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_371
timestamp 1679581782
transform 1 0 36192 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_378
timestamp 1679581782
transform 1 0 36864 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_385
timestamp 1679581782
transform 1 0 37536 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_392
timestamp 1679581782
transform 1 0 38208 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_399
timestamp 1679581782
transform 1 0 38880 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_406
timestamp 1679581782
transform 1 0 39552 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_413
timestamp 1679581782
transform 1 0 40224 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_420
timestamp 1679581782
transform 1 0 40896 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_427
timestamp 1679581782
transform 1 0 41568 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_434
timestamp 1679581782
transform 1 0 42240 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_441
timestamp 1679581782
transform 1 0 42912 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_448
timestamp 1679581782
transform 1 0 43584 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_455
timestamp 1679581782
transform 1 0 44256 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_462
timestamp 1679581782
transform 1 0 44928 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_469
timestamp 1679581782
transform 1 0 45600 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_476
timestamp 1679581782
transform 1 0 46272 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_483
timestamp 1679581782
transform 1 0 46944 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_490
timestamp 1679581782
transform 1 0 47616 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_497
timestamp 1679581782
transform 1 0 48288 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_504
timestamp 1679581782
transform 1 0 48960 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_511
timestamp 1679581782
transform 1 0 49632 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_518
timestamp 1679581782
transform 1 0 50304 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_525
timestamp 1679581782
transform 1 0 50976 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_532
timestamp 1679581782
transform 1 0 51648 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_539
timestamp 1679581782
transform 1 0 52320 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_546
timestamp 1679581782
transform 1 0 52992 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_553
timestamp 1679581782
transform 1 0 53664 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_560
timestamp 1679581782
transform 1 0 54336 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_567
timestamp 1679581782
transform 1 0 55008 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_574
timestamp 1679581782
transform 1 0 55680 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_581
timestamp 1679581782
transform 1 0 56352 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_588
timestamp 1679581782
transform 1 0 57024 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_595
timestamp 1679581782
transform 1 0 57696 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_602
timestamp 1679581782
transform 1 0 58368 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_609
timestamp 1679581782
transform 1 0 59040 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_616
timestamp 1679581782
transform 1 0 59712 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_623
timestamp 1679581782
transform 1 0 60384 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_630
timestamp 1679581782
transform 1 0 61056 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_637
timestamp 1679581782
transform 1 0 61728 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_644
timestamp 1679581782
transform 1 0 62400 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_651
timestamp 1679581782
transform 1 0 63072 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_658
timestamp 1679581782
transform 1 0 63744 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_665
timestamp 1679581782
transform 1 0 64416 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_672
timestamp 1679581782
transform 1 0 65088 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_679
timestamp 1679581782
transform 1 0 65760 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_686
timestamp 1679581782
transform 1 0 66432 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_693
timestamp 1679581782
transform 1 0 67104 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_700
timestamp 1679581782
transform 1 0 67776 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_707
timestamp 1679581782
transform 1 0 68448 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_714
timestamp 1679581782
transform 1 0 69120 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_721
timestamp 1679581782
transform 1 0 69792 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_728
timestamp 1679581782
transform 1 0 70464 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_735
timestamp 1679581782
transform 1 0 71136 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_742
timestamp 1679581782
transform 1 0 71808 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_749
timestamp 1679581782
transform 1 0 72480 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_756
timestamp 1679581782
transform 1 0 73152 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_763
timestamp 1679581782
transform 1 0 73824 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_770
timestamp 1679581782
transform 1 0 74496 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_777
timestamp 1679581782
transform 1 0 75168 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_784
timestamp 1679581782
transform 1 0 75840 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_791
timestamp 1679581782
transform 1 0 76512 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_798
timestamp 1679581782
transform 1 0 77184 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_805
timestamp 1679581782
transform 1 0 77856 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_812
timestamp 1679581782
transform 1 0 78528 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_819
timestamp 1679581782
transform 1 0 79200 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_826
timestamp 1679581782
transform 1 0 79872 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_833
timestamp 1679581782
transform 1 0 80544 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_840
timestamp 1679581782
transform 1 0 81216 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_847
timestamp 1679581782
transform 1 0 81888 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_854
timestamp 1679581782
transform 1 0 82560 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_861
timestamp 1679581782
transform 1 0 83232 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_868
timestamp 1679581782
transform 1 0 83904 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_875
timestamp 1679581782
transform 1 0 84576 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_882
timestamp 1679581782
transform 1 0 85248 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_889
timestamp 1679581782
transform 1 0 85920 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_896
timestamp 1679581782
transform 1 0 86592 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_903
timestamp 1679581782
transform 1 0 87264 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_910
timestamp 1679581782
transform 1 0 87936 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_917
timestamp 1679581782
transform 1 0 88608 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_924
timestamp 1679581782
transform 1 0 89280 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_931
timestamp 1679581782
transform 1 0 89952 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_938
timestamp 1679581782
transform 1 0 90624 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_945
timestamp 1679581782
transform 1 0 91296 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_952
timestamp 1679581782
transform 1 0 91968 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_959
timestamp 1679581782
transform 1 0 92640 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_966
timestamp 1679581782
transform 1 0 93312 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_973
timestamp 1679581782
transform 1 0 93984 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_980
timestamp 1679581782
transform 1 0 94656 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_987
timestamp 1679581782
transform 1 0 95328 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_994
timestamp 1679581782
transform 1 0 96000 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_1001
timestamp 1679581782
transform 1 0 96672 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_1008
timestamp 1679581782
transform 1 0 97344 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_1015
timestamp 1679581782
transform 1 0 98016 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_1022
timestamp 1679581782
transform 1 0 98688 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_4
timestamp 1679581782
transform 1 0 960 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_11
timestamp 1679581782
transform 1 0 1632 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_18
timestamp 1679581782
transform 1 0 2304 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_25
timestamp 1679581782
transform 1 0 2976 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_32
timestamp 1679581782
transform 1 0 3648 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_39
timestamp 1679581782
transform 1 0 4320 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_46
timestamp 1679581782
transform 1 0 4992 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_53
timestamp 1679581782
transform 1 0 5664 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_60
timestamp 1679581782
transform 1 0 6336 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_67
timestamp 1679581782
transform 1 0 7008 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_74
timestamp 1679581782
transform 1 0 7680 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_81
timestamp 1679581782
transform 1 0 8352 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_88
timestamp 1679581782
transform 1 0 9024 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_95
timestamp 1679581782
transform 1 0 9696 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_102
timestamp 1679581782
transform 1 0 10368 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_109
timestamp 1679581782
transform 1 0 11040 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_116
timestamp 1679581782
transform 1 0 11712 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_123
timestamp 1679581782
transform 1 0 12384 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_130
timestamp 1679581782
transform 1 0 13056 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_137
timestamp 1679581782
transform 1 0 13728 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_144
timestamp 1679581782
transform 1 0 14400 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_151
timestamp 1679581782
transform 1 0 15072 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_158
timestamp 1679581782
transform 1 0 15744 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_165
timestamp 1679581782
transform 1 0 16416 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_172
timestamp 1679581782
transform 1 0 17088 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_179
timestamp 1679581782
transform 1 0 17760 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_186
timestamp 1679581782
transform 1 0 18432 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_193
timestamp 1679581782
transform 1 0 19104 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_200
timestamp 1679581782
transform 1 0 19776 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_207
timestamp 1679581782
transform 1 0 20448 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_214
timestamp 1679581782
transform 1 0 21120 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_221
timestamp 1679581782
transform 1 0 21792 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_228
timestamp 1679581782
transform 1 0 22464 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_235
timestamp 1679581782
transform 1 0 23136 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_242
timestamp 1679581782
transform 1 0 23808 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_249
timestamp 1679581782
transform 1 0 24480 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_256
timestamp 1679581782
transform 1 0 25152 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_263
timestamp 1679581782
transform 1 0 25824 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_270
timestamp 1679581782
transform 1 0 26496 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_277
timestamp 1679581782
transform 1 0 27168 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_284
timestamp 1679581782
transform 1 0 27840 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_291
timestamp 1679581782
transform 1 0 28512 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_298
timestamp 1679581782
transform 1 0 29184 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_305
timestamp 1679581782
transform 1 0 29856 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_312
timestamp 1679581782
transform 1 0 30528 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_319
timestamp 1679581782
transform 1 0 31200 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_326
timestamp 1679581782
transform 1 0 31872 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_333
timestamp 1679581782
transform 1 0 32544 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_340
timestamp 1679581782
transform 1 0 33216 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_347
timestamp 1679581782
transform 1 0 33888 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_354
timestamp 1679581782
transform 1 0 34560 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_361
timestamp 1679581782
transform 1 0 35232 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_368
timestamp 1679581782
transform 1 0 35904 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_375
timestamp 1679581782
transform 1 0 36576 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_382
timestamp 1679581782
transform 1 0 37248 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_389
timestamp 1679581782
transform 1 0 37920 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_396
timestamp 1679581782
transform 1 0 38592 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_403
timestamp 1679581782
transform 1 0 39264 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_410
timestamp 1679581782
transform 1 0 39936 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_417
timestamp 1679581782
transform 1 0 40608 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_424
timestamp 1679581782
transform 1 0 41280 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_431
timestamp 1679581782
transform 1 0 41952 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_438
timestamp 1679581782
transform 1 0 42624 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_445
timestamp 1679581782
transform 1 0 43296 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_452
timestamp 1679581782
transform 1 0 43968 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_459
timestamp 1679581782
transform 1 0 44640 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_466
timestamp 1679581782
transform 1 0 45312 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_473
timestamp 1679581782
transform 1 0 45984 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_480
timestamp 1679581782
transform 1 0 46656 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_487
timestamp 1679581782
transform 1 0 47328 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_494
timestamp 1679581782
transform 1 0 48000 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_501
timestamp 1679581782
transform 1 0 48672 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_508
timestamp 1679581782
transform 1 0 49344 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_515
timestamp 1679581782
transform 1 0 50016 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_522
timestamp 1679581782
transform 1 0 50688 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_529
timestamp 1679581782
transform 1 0 51360 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_536
timestamp 1679581782
transform 1 0 52032 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_543
timestamp 1679581782
transform 1 0 52704 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_550
timestamp 1679581782
transform 1 0 53376 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_557
timestamp 1679581782
transform 1 0 54048 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_564
timestamp 1679581782
transform 1 0 54720 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_571
timestamp 1679581782
transform 1 0 55392 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_578
timestamp 1679581782
transform 1 0 56064 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_585
timestamp 1679581782
transform 1 0 56736 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_592
timestamp 1679581782
transform 1 0 57408 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_599
timestamp 1679581782
transform 1 0 58080 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_606
timestamp 1679581782
transform 1 0 58752 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_613
timestamp 1679581782
transform 1 0 59424 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_620
timestamp 1679581782
transform 1 0 60096 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_627
timestamp 1679581782
transform 1 0 60768 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_634
timestamp 1679581782
transform 1 0 61440 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_641
timestamp 1679581782
transform 1 0 62112 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_648
timestamp 1679581782
transform 1 0 62784 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_655
timestamp 1679581782
transform 1 0 63456 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_662
timestamp 1679581782
transform 1 0 64128 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_669
timestamp 1679581782
transform 1 0 64800 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_676
timestamp 1679581782
transform 1 0 65472 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_683
timestamp 1679581782
transform 1 0 66144 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_690
timestamp 1679581782
transform 1 0 66816 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_697
timestamp 1679581782
transform 1 0 67488 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_704
timestamp 1679581782
transform 1 0 68160 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_711
timestamp 1679581782
transform 1 0 68832 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_718
timestamp 1679581782
transform 1 0 69504 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_725
timestamp 1679581782
transform 1 0 70176 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_732
timestamp 1679581782
transform 1 0 70848 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_739
timestamp 1679581782
transform 1 0 71520 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_746
timestamp 1679581782
transform 1 0 72192 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_753
timestamp 1679581782
transform 1 0 72864 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_760
timestamp 1679581782
transform 1 0 73536 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_767
timestamp 1679581782
transform 1 0 74208 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_774
timestamp 1679581782
transform 1 0 74880 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_781
timestamp 1679581782
transform 1 0 75552 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_788
timestamp 1679581782
transform 1 0 76224 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_795
timestamp 1679581782
transform 1 0 76896 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_802
timestamp 1679581782
transform 1 0 77568 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_809
timestamp 1679581782
transform 1 0 78240 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_816
timestamp 1679581782
transform 1 0 78912 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_823
timestamp 1679581782
transform 1 0 79584 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_830
timestamp 1679581782
transform 1 0 80256 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_837
timestamp 1679581782
transform 1 0 80928 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_844
timestamp 1679581782
transform 1 0 81600 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_851
timestamp 1679581782
transform 1 0 82272 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_858
timestamp 1679581782
transform 1 0 82944 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_865
timestamp 1679581782
transform 1 0 83616 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_872
timestamp 1679581782
transform 1 0 84288 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_879
timestamp 1679581782
transform 1 0 84960 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_886
timestamp 1679581782
transform 1 0 85632 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_893
timestamp 1679581782
transform 1 0 86304 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_900
timestamp 1679581782
transform 1 0 86976 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_907
timestamp 1679581782
transform 1 0 87648 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_914
timestamp 1679581782
transform 1 0 88320 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_921
timestamp 1679581782
transform 1 0 88992 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_928
timestamp 1679581782
transform 1 0 89664 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_935
timestamp 1679581782
transform 1 0 90336 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_942
timestamp 1679581782
transform 1 0 91008 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_949
timestamp 1679581782
transform 1 0 91680 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_956
timestamp 1679581782
transform 1 0 92352 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_963
timestamp 1679581782
transform 1 0 93024 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_970
timestamp 1679581782
transform 1 0 93696 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_977
timestamp 1679581782
transform 1 0 94368 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_984
timestamp 1679581782
transform 1 0 95040 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_991
timestamp 1679581782
transform 1 0 95712 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_998
timestamp 1679581782
transform 1 0 96384 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_1005
timestamp 1679581782
transform 1 0 97056 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_1012
timestamp 1679581782
transform 1 0 97728 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_1019
timestamp 1679581782
transform 1 0 98400 0 1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_46_1026
timestamp 1677580104
transform 1 0 99072 0 1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_46_1028
timestamp 1677579658
transform 1 0 99264 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_47_0
timestamp 1679581782
transform 1 0 576 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_7
timestamp 1679581782
transform 1 0 1248 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_14
timestamp 1679581782
transform 1 0 1920 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_21
timestamp 1679581782
transform 1 0 2592 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_28
timestamp 1679581782
transform 1 0 3264 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_35
timestamp 1679581782
transform 1 0 3936 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_42
timestamp 1679581782
transform 1 0 4608 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_49
timestamp 1679581782
transform 1 0 5280 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_56
timestamp 1679581782
transform 1 0 5952 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_63
timestamp 1679581782
transform 1 0 6624 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_70
timestamp 1679581782
transform 1 0 7296 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_77
timestamp 1679581782
transform 1 0 7968 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_84
timestamp 1679581782
transform 1 0 8640 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_91
timestamp 1679581782
transform 1 0 9312 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_98
timestamp 1679581782
transform 1 0 9984 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_105
timestamp 1679581782
transform 1 0 10656 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_112
timestamp 1679581782
transform 1 0 11328 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_119
timestamp 1679581782
transform 1 0 12000 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_126
timestamp 1679581782
transform 1 0 12672 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_133
timestamp 1679581782
transform 1 0 13344 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_140
timestamp 1679581782
transform 1 0 14016 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_147
timestamp 1679581782
transform 1 0 14688 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_154
timestamp 1679581782
transform 1 0 15360 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_161
timestamp 1679581782
transform 1 0 16032 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_168
timestamp 1679581782
transform 1 0 16704 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_175
timestamp 1679581782
transform 1 0 17376 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_182
timestamp 1679581782
transform 1 0 18048 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_189
timestamp 1679581782
transform 1 0 18720 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_196
timestamp 1679581782
transform 1 0 19392 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_203
timestamp 1679581782
transform 1 0 20064 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_210
timestamp 1679581782
transform 1 0 20736 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_217
timestamp 1679581782
transform 1 0 21408 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_224
timestamp 1679581782
transform 1 0 22080 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_231
timestamp 1679581782
transform 1 0 22752 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_238
timestamp 1679581782
transform 1 0 23424 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_245
timestamp 1679581782
transform 1 0 24096 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_252
timestamp 1679581782
transform 1 0 24768 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_259
timestamp 1679581782
transform 1 0 25440 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_266
timestamp 1679581782
transform 1 0 26112 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_273
timestamp 1679581782
transform 1 0 26784 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_280
timestamp 1679581782
transform 1 0 27456 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_287
timestamp 1679581782
transform 1 0 28128 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_294
timestamp 1679581782
transform 1 0 28800 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_301
timestamp 1679581782
transform 1 0 29472 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_308
timestamp 1679581782
transform 1 0 30144 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_315
timestamp 1679581782
transform 1 0 30816 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_322
timestamp 1679581782
transform 1 0 31488 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_329
timestamp 1679581782
transform 1 0 32160 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_336
timestamp 1679581782
transform 1 0 32832 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_343
timestamp 1679581782
transform 1 0 33504 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_350
timestamp 1679581782
transform 1 0 34176 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_357
timestamp 1679581782
transform 1 0 34848 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_364
timestamp 1679581782
transform 1 0 35520 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_371
timestamp 1679581782
transform 1 0 36192 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_378
timestamp 1679581782
transform 1 0 36864 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_385
timestamp 1679581782
transform 1 0 37536 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_392
timestamp 1679581782
transform 1 0 38208 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_399
timestamp 1679581782
transform 1 0 38880 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_406
timestamp 1679581782
transform 1 0 39552 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_413
timestamp 1679581782
transform 1 0 40224 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_420
timestamp 1679581782
transform 1 0 40896 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_427
timestamp 1679581782
transform 1 0 41568 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_434
timestamp 1679581782
transform 1 0 42240 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_441
timestamp 1679581782
transform 1 0 42912 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_448
timestamp 1679581782
transform 1 0 43584 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_455
timestamp 1679581782
transform 1 0 44256 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_462
timestamp 1679581782
transform 1 0 44928 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_469
timestamp 1679581782
transform 1 0 45600 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_476
timestamp 1679581782
transform 1 0 46272 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_483
timestamp 1679581782
transform 1 0 46944 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_490
timestamp 1679581782
transform 1 0 47616 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_497
timestamp 1679581782
transform 1 0 48288 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_504
timestamp 1679581782
transform 1 0 48960 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_511
timestamp 1679581782
transform 1 0 49632 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_518
timestamp 1679581782
transform 1 0 50304 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_525
timestamp 1679581782
transform 1 0 50976 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_532
timestamp 1679581782
transform 1 0 51648 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_539
timestamp 1679581782
transform 1 0 52320 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_546
timestamp 1679581782
transform 1 0 52992 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_553
timestamp 1679581782
transform 1 0 53664 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_560
timestamp 1679581782
transform 1 0 54336 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_567
timestamp 1679581782
transform 1 0 55008 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_574
timestamp 1679581782
transform 1 0 55680 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_581
timestamp 1679581782
transform 1 0 56352 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_588
timestamp 1679581782
transform 1 0 57024 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_595
timestamp 1679581782
transform 1 0 57696 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_602
timestamp 1679581782
transform 1 0 58368 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_609
timestamp 1679581782
transform 1 0 59040 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_616
timestamp 1679581782
transform 1 0 59712 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_623
timestamp 1679581782
transform 1 0 60384 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_630
timestamp 1679581782
transform 1 0 61056 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_637
timestamp 1679581782
transform 1 0 61728 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_644
timestamp 1679581782
transform 1 0 62400 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_651
timestamp 1679581782
transform 1 0 63072 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_658
timestamp 1679581782
transform 1 0 63744 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_665
timestamp 1679581782
transform 1 0 64416 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_672
timestamp 1679581782
transform 1 0 65088 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_679
timestamp 1679581782
transform 1 0 65760 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_686
timestamp 1679581782
transform 1 0 66432 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_693
timestamp 1679581782
transform 1 0 67104 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_700
timestamp 1679581782
transform 1 0 67776 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_707
timestamp 1679581782
transform 1 0 68448 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_714
timestamp 1679581782
transform 1 0 69120 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_721
timestamp 1679581782
transform 1 0 69792 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_728
timestamp 1679581782
transform 1 0 70464 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_735
timestamp 1679581782
transform 1 0 71136 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_742
timestamp 1679581782
transform 1 0 71808 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_749
timestamp 1679581782
transform 1 0 72480 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_756
timestamp 1679581782
transform 1 0 73152 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_763
timestamp 1679581782
transform 1 0 73824 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_770
timestamp 1679581782
transform 1 0 74496 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_777
timestamp 1679581782
transform 1 0 75168 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_784
timestamp 1679581782
transform 1 0 75840 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_791
timestamp 1679581782
transform 1 0 76512 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_798
timestamp 1679581782
transform 1 0 77184 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_805
timestamp 1679581782
transform 1 0 77856 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_812
timestamp 1679581782
transform 1 0 78528 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_819
timestamp 1679581782
transform 1 0 79200 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_826
timestamp 1679581782
transform 1 0 79872 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_833
timestamp 1679581782
transform 1 0 80544 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_840
timestamp 1679581782
transform 1 0 81216 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_847
timestamp 1679581782
transform 1 0 81888 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_854
timestamp 1679581782
transform 1 0 82560 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_861
timestamp 1679581782
transform 1 0 83232 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_868
timestamp 1679581782
transform 1 0 83904 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_875
timestamp 1679581782
transform 1 0 84576 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_882
timestamp 1679581782
transform 1 0 85248 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_889
timestamp 1679581782
transform 1 0 85920 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_896
timestamp 1679581782
transform 1 0 86592 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_903
timestamp 1679581782
transform 1 0 87264 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_910
timestamp 1679581782
transform 1 0 87936 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_917
timestamp 1679581782
transform 1 0 88608 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_924
timestamp 1679581782
transform 1 0 89280 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_931
timestamp 1679581782
transform 1 0 89952 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_938
timestamp 1679581782
transform 1 0 90624 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_945
timestamp 1679581782
transform 1 0 91296 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_952
timestamp 1679581782
transform 1 0 91968 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_959
timestamp 1679581782
transform 1 0 92640 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_966
timestamp 1679581782
transform 1 0 93312 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_973
timestamp 1679581782
transform 1 0 93984 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_980
timestamp 1679581782
transform 1 0 94656 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_987
timestamp 1679581782
transform 1 0 95328 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_994
timestamp 1679581782
transform 1 0 96000 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_1001
timestamp 1679581782
transform 1 0 96672 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_1008
timestamp 1679581782
transform 1 0 97344 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_1015
timestamp 1679581782
transform 1 0 98016 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_1022
timestamp 1679581782
transform 1 0 98688 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_0
timestamp 1679581782
transform 1 0 576 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_7
timestamp 1679581782
transform 1 0 1248 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_14
timestamp 1679581782
transform 1 0 1920 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_21
timestamp 1679581782
transform 1 0 2592 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_28
timestamp 1679581782
transform 1 0 3264 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_35
timestamp 1679581782
transform 1 0 3936 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_42
timestamp 1679581782
transform 1 0 4608 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_49
timestamp 1679581782
transform 1 0 5280 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_56
timestamp 1679581782
transform 1 0 5952 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_63
timestamp 1679581782
transform 1 0 6624 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_70
timestamp 1679581782
transform 1 0 7296 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_77
timestamp 1679581782
transform 1 0 7968 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_84
timestamp 1679581782
transform 1 0 8640 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_91
timestamp 1679581782
transform 1 0 9312 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_98
timestamp 1679581782
transform 1 0 9984 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_105
timestamp 1679581782
transform 1 0 10656 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_112
timestamp 1679581782
transform 1 0 11328 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_119
timestamp 1679581782
transform 1 0 12000 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_126
timestamp 1679581782
transform 1 0 12672 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_133
timestamp 1679581782
transform 1 0 13344 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_140
timestamp 1679581782
transform 1 0 14016 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_147
timestamp 1679581782
transform 1 0 14688 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_154
timestamp 1679581782
transform 1 0 15360 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_161
timestamp 1679581782
transform 1 0 16032 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_168
timestamp 1679581782
transform 1 0 16704 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_175
timestamp 1679581782
transform 1 0 17376 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_182
timestamp 1679581782
transform 1 0 18048 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_189
timestamp 1679581782
transform 1 0 18720 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_196
timestamp 1679581782
transform 1 0 19392 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_203
timestamp 1679581782
transform 1 0 20064 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_210
timestamp 1679581782
transform 1 0 20736 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_217
timestamp 1679581782
transform 1 0 21408 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_224
timestamp 1679581782
transform 1 0 22080 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_231
timestamp 1679581782
transform 1 0 22752 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_238
timestamp 1679581782
transform 1 0 23424 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_245
timestamp 1679581782
transform 1 0 24096 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_252
timestamp 1679581782
transform 1 0 24768 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_259
timestamp 1679581782
transform 1 0 25440 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_266
timestamp 1679581782
transform 1 0 26112 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_273
timestamp 1679581782
transform 1 0 26784 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_280
timestamp 1679581782
transform 1 0 27456 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_287
timestamp 1679581782
transform 1 0 28128 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_294
timestamp 1679581782
transform 1 0 28800 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_301
timestamp 1679581782
transform 1 0 29472 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_308
timestamp 1679581782
transform 1 0 30144 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_315
timestamp 1679581782
transform 1 0 30816 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_322
timestamp 1679581782
transform 1 0 31488 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_329
timestamp 1679581782
transform 1 0 32160 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_336
timestamp 1679581782
transform 1 0 32832 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_343
timestamp 1679581782
transform 1 0 33504 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_350
timestamp 1679581782
transform 1 0 34176 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_357
timestamp 1679581782
transform 1 0 34848 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_364
timestamp 1679581782
transform 1 0 35520 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_371
timestamp 1679581782
transform 1 0 36192 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_378
timestamp 1679581782
transform 1 0 36864 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_385
timestamp 1679581782
transform 1 0 37536 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_392
timestamp 1679581782
transform 1 0 38208 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_399
timestamp 1679581782
transform 1 0 38880 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_406
timestamp 1679581782
transform 1 0 39552 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_413
timestamp 1679581782
transform 1 0 40224 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_420
timestamp 1679581782
transform 1 0 40896 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_427
timestamp 1679581782
transform 1 0 41568 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_434
timestamp 1679581782
transform 1 0 42240 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_441
timestamp 1679581782
transform 1 0 42912 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_448
timestamp 1679581782
transform 1 0 43584 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_455
timestamp 1679581782
transform 1 0 44256 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_462
timestamp 1679581782
transform 1 0 44928 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_469
timestamp 1679581782
transform 1 0 45600 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_476
timestamp 1679581782
transform 1 0 46272 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_483
timestamp 1679581782
transform 1 0 46944 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_490
timestamp 1679581782
transform 1 0 47616 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_497
timestamp 1679581782
transform 1 0 48288 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_504
timestamp 1679581782
transform 1 0 48960 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_511
timestamp 1679581782
transform 1 0 49632 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_518
timestamp 1679581782
transform 1 0 50304 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_525
timestamp 1679581782
transform 1 0 50976 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_532
timestamp 1679581782
transform 1 0 51648 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_539
timestamp 1679581782
transform 1 0 52320 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_546
timestamp 1679581782
transform 1 0 52992 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_553
timestamp 1679581782
transform 1 0 53664 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_560
timestamp 1679581782
transform 1 0 54336 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_567
timestamp 1679581782
transform 1 0 55008 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_574
timestamp 1679581782
transform 1 0 55680 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_581
timestamp 1679581782
transform 1 0 56352 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_588
timestamp 1679581782
transform 1 0 57024 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_595
timestamp 1679581782
transform 1 0 57696 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_602
timestamp 1679581782
transform 1 0 58368 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_609
timestamp 1679581782
transform 1 0 59040 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_616
timestamp 1679581782
transform 1 0 59712 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_623
timestamp 1679581782
transform 1 0 60384 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_630
timestamp 1679581782
transform 1 0 61056 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_637
timestamp 1679581782
transform 1 0 61728 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_644
timestamp 1679581782
transform 1 0 62400 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_651
timestamp 1679581782
transform 1 0 63072 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_658
timestamp 1679581782
transform 1 0 63744 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_665
timestamp 1679581782
transform 1 0 64416 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_672
timestamp 1679581782
transform 1 0 65088 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_679
timestamp 1679581782
transform 1 0 65760 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_686
timestamp 1679581782
transform 1 0 66432 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_693
timestamp 1679581782
transform 1 0 67104 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_700
timestamp 1679581782
transform 1 0 67776 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_707
timestamp 1679581782
transform 1 0 68448 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_714
timestamp 1679581782
transform 1 0 69120 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_721
timestamp 1679581782
transform 1 0 69792 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_728
timestamp 1679581782
transform 1 0 70464 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_735
timestamp 1679581782
transform 1 0 71136 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_742
timestamp 1679581782
transform 1 0 71808 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_749
timestamp 1679581782
transform 1 0 72480 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_756
timestamp 1679581782
transform 1 0 73152 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_763
timestamp 1679581782
transform 1 0 73824 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_770
timestamp 1679581782
transform 1 0 74496 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_777
timestamp 1679581782
transform 1 0 75168 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_784
timestamp 1679581782
transform 1 0 75840 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_791
timestamp 1679581782
transform 1 0 76512 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_798
timestamp 1679581782
transform 1 0 77184 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_805
timestamp 1679581782
transform 1 0 77856 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_812
timestamp 1679581782
transform 1 0 78528 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_819
timestamp 1679581782
transform 1 0 79200 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_826
timestamp 1679581782
transform 1 0 79872 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_833
timestamp 1679581782
transform 1 0 80544 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_840
timestamp 1679581782
transform 1 0 81216 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_847
timestamp 1679581782
transform 1 0 81888 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_854
timestamp 1679581782
transform 1 0 82560 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_861
timestamp 1679581782
transform 1 0 83232 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_868
timestamp 1679581782
transform 1 0 83904 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_875
timestamp 1679581782
transform 1 0 84576 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_882
timestamp 1679581782
transform 1 0 85248 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_889
timestamp 1679581782
transform 1 0 85920 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_896
timestamp 1679581782
transform 1 0 86592 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_903
timestamp 1679581782
transform 1 0 87264 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_910
timestamp 1679581782
transform 1 0 87936 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_917
timestamp 1679581782
transform 1 0 88608 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_924
timestamp 1679581782
transform 1 0 89280 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_931
timestamp 1679581782
transform 1 0 89952 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_938
timestamp 1679581782
transform 1 0 90624 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_945
timestamp 1679581782
transform 1 0 91296 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_952
timestamp 1679581782
transform 1 0 91968 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_959
timestamp 1679581782
transform 1 0 92640 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_966
timestamp 1679581782
transform 1 0 93312 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_973
timestamp 1679581782
transform 1 0 93984 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_980
timestamp 1679581782
transform 1 0 94656 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_987
timestamp 1679581782
transform 1 0 95328 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_994
timestamp 1679581782
transform 1 0 96000 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_1001
timestamp 1679581782
transform 1 0 96672 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_1008
timestamp 1679581782
transform 1 0 97344 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_1015
timestamp 1679581782
transform 1 0 98016 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_1022
timestamp 1679581782
transform 1 0 98688 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_4
timestamp 1679581782
transform 1 0 960 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_11
timestamp 1679581782
transform 1 0 1632 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_18
timestamp 1679581782
transform 1 0 2304 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_25
timestamp 1679581782
transform 1 0 2976 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_32
timestamp 1679581782
transform 1 0 3648 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_39
timestamp 1679581782
transform 1 0 4320 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_46
timestamp 1679581782
transform 1 0 4992 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_53
timestamp 1679581782
transform 1 0 5664 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_60
timestamp 1679581782
transform 1 0 6336 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_67
timestamp 1679581782
transform 1 0 7008 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_74
timestamp 1679581782
transform 1 0 7680 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_81
timestamp 1679581782
transform 1 0 8352 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_88
timestamp 1679581782
transform 1 0 9024 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_95
timestamp 1679581782
transform 1 0 9696 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_102
timestamp 1679581782
transform 1 0 10368 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_109
timestamp 1679581782
transform 1 0 11040 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_116
timestamp 1679581782
transform 1 0 11712 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_123
timestamp 1679581782
transform 1 0 12384 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_130
timestamp 1679581782
transform 1 0 13056 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_137
timestamp 1679581782
transform 1 0 13728 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_144
timestamp 1679581782
transform 1 0 14400 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_151
timestamp 1679581782
transform 1 0 15072 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_158
timestamp 1679581782
transform 1 0 15744 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_165
timestamp 1679581782
transform 1 0 16416 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_172
timestamp 1679581782
transform 1 0 17088 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_179
timestamp 1679581782
transform 1 0 17760 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_186
timestamp 1679581782
transform 1 0 18432 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_193
timestamp 1679581782
transform 1 0 19104 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_200
timestamp 1679581782
transform 1 0 19776 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_207
timestamp 1679581782
transform 1 0 20448 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_214
timestamp 1679581782
transform 1 0 21120 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_221
timestamp 1679581782
transform 1 0 21792 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_228
timestamp 1679581782
transform 1 0 22464 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_235
timestamp 1679581782
transform 1 0 23136 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_242
timestamp 1679581782
transform 1 0 23808 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_249
timestamp 1679581782
transform 1 0 24480 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_256
timestamp 1679581782
transform 1 0 25152 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_263
timestamp 1679581782
transform 1 0 25824 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_270
timestamp 1679581782
transform 1 0 26496 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_277
timestamp 1679581782
transform 1 0 27168 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_284
timestamp 1679581782
transform 1 0 27840 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_291
timestamp 1679581782
transform 1 0 28512 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_298
timestamp 1679581782
transform 1 0 29184 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_305
timestamp 1679581782
transform 1 0 29856 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_312
timestamp 1679581782
transform 1 0 30528 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_319
timestamp 1679581782
transform 1 0 31200 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_326
timestamp 1679581782
transform 1 0 31872 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_333
timestamp 1679581782
transform 1 0 32544 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_340
timestamp 1679581782
transform 1 0 33216 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_347
timestamp 1679581782
transform 1 0 33888 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_354
timestamp 1679581782
transform 1 0 34560 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_361
timestamp 1679581782
transform 1 0 35232 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_368
timestamp 1679581782
transform 1 0 35904 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_375
timestamp 1679581782
transform 1 0 36576 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_382
timestamp 1679581782
transform 1 0 37248 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_389
timestamp 1679581782
transform 1 0 37920 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_396
timestamp 1679581782
transform 1 0 38592 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_403
timestamp 1679581782
transform 1 0 39264 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_410
timestamp 1679581782
transform 1 0 39936 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_417
timestamp 1679581782
transform 1 0 40608 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_424
timestamp 1679581782
transform 1 0 41280 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_431
timestamp 1679581782
transform 1 0 41952 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_438
timestamp 1679581782
transform 1 0 42624 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_445
timestamp 1679581782
transform 1 0 43296 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_452
timestamp 1679581782
transform 1 0 43968 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_459
timestamp 1679581782
transform 1 0 44640 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_466
timestamp 1679581782
transform 1 0 45312 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_473
timestamp 1679581782
transform 1 0 45984 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_480
timestamp 1679581782
transform 1 0 46656 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_487
timestamp 1679581782
transform 1 0 47328 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_494
timestamp 1679581782
transform 1 0 48000 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_501
timestamp 1679581782
transform 1 0 48672 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_508
timestamp 1679581782
transform 1 0 49344 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_515
timestamp 1679581782
transform 1 0 50016 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_522
timestamp 1679581782
transform 1 0 50688 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_529
timestamp 1679581782
transform 1 0 51360 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_536
timestamp 1679581782
transform 1 0 52032 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_543
timestamp 1679581782
transform 1 0 52704 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_550
timestamp 1679581782
transform 1 0 53376 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_557
timestamp 1679581782
transform 1 0 54048 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_564
timestamp 1679581782
transform 1 0 54720 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_571
timestamp 1679581782
transform 1 0 55392 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_578
timestamp 1679581782
transform 1 0 56064 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_585
timestamp 1679581782
transform 1 0 56736 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_592
timestamp 1679581782
transform 1 0 57408 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_599
timestamp 1679581782
transform 1 0 58080 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_606
timestamp 1679581782
transform 1 0 58752 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_613
timestamp 1679581782
transform 1 0 59424 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_620
timestamp 1679581782
transform 1 0 60096 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_627
timestamp 1679581782
transform 1 0 60768 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_634
timestamp 1679581782
transform 1 0 61440 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_641
timestamp 1679581782
transform 1 0 62112 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_648
timestamp 1679581782
transform 1 0 62784 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_655
timestamp 1679581782
transform 1 0 63456 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_662
timestamp 1679581782
transform 1 0 64128 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_669
timestamp 1679581782
transform 1 0 64800 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_676
timestamp 1679581782
transform 1 0 65472 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_683
timestamp 1679581782
transform 1 0 66144 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_690
timestamp 1679581782
transform 1 0 66816 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_697
timestamp 1679581782
transform 1 0 67488 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_704
timestamp 1679581782
transform 1 0 68160 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_711
timestamp 1679581782
transform 1 0 68832 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_718
timestamp 1679581782
transform 1 0 69504 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_725
timestamp 1679581782
transform 1 0 70176 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_732
timestamp 1679581782
transform 1 0 70848 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_739
timestamp 1679581782
transform 1 0 71520 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_746
timestamp 1679581782
transform 1 0 72192 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_753
timestamp 1679581782
transform 1 0 72864 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_760
timestamp 1679581782
transform 1 0 73536 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_767
timestamp 1679581782
transform 1 0 74208 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_774
timestamp 1679581782
transform 1 0 74880 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_781
timestamp 1679581782
transform 1 0 75552 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_788
timestamp 1679581782
transform 1 0 76224 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_795
timestamp 1679581782
transform 1 0 76896 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_802
timestamp 1679581782
transform 1 0 77568 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_809
timestamp 1679581782
transform 1 0 78240 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_816
timestamp 1679581782
transform 1 0 78912 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_823
timestamp 1679581782
transform 1 0 79584 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_830
timestamp 1679581782
transform 1 0 80256 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_837
timestamp 1679581782
transform 1 0 80928 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_844
timestamp 1679581782
transform 1 0 81600 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_851
timestamp 1679581782
transform 1 0 82272 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_858
timestamp 1679581782
transform 1 0 82944 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_865
timestamp 1679581782
transform 1 0 83616 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_872
timestamp 1679581782
transform 1 0 84288 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_879
timestamp 1679581782
transform 1 0 84960 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_886
timestamp 1679581782
transform 1 0 85632 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_893
timestamp 1679581782
transform 1 0 86304 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_900
timestamp 1679581782
transform 1 0 86976 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_907
timestamp 1679581782
transform 1 0 87648 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_914
timestamp 1679581782
transform 1 0 88320 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_921
timestamp 1679581782
transform 1 0 88992 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_928
timestamp 1679581782
transform 1 0 89664 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_935
timestamp 1679581782
transform 1 0 90336 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_942
timestamp 1679581782
transform 1 0 91008 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_949
timestamp 1679581782
transform 1 0 91680 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_956
timestamp 1679581782
transform 1 0 92352 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_963
timestamp 1679581782
transform 1 0 93024 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_970
timestamp 1679581782
transform 1 0 93696 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_977
timestamp 1679581782
transform 1 0 94368 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_984
timestamp 1679581782
transform 1 0 95040 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_991
timestamp 1679581782
transform 1 0 95712 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_998
timestamp 1679581782
transform 1 0 96384 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_1005
timestamp 1679581782
transform 1 0 97056 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_1012
timestamp 1679581782
transform 1 0 97728 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_1019
timestamp 1679581782
transform 1 0 98400 0 -1 38556
box -48 -56 720 834
use sg13g2_fill_2  FILLER_49_1026
timestamp 1677580104
transform 1 0 99072 0 -1 38556
box -48 -56 240 834
use sg13g2_fill_1  FILLER_49_1028
timestamp 1677579658
transform 1 0 99264 0 -1 38556
box -48 -56 144 834
use sg13g2_decap_8  FILLER_50_0
timestamp 1679581782
transform 1 0 576 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_7
timestamp 1679581782
transform 1 0 1248 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_14
timestamp 1679581782
transform 1 0 1920 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_21
timestamp 1679581782
transform 1 0 2592 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_28
timestamp 1679581782
transform 1 0 3264 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_35
timestamp 1679581782
transform 1 0 3936 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_42
timestamp 1679581782
transform 1 0 4608 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_49
timestamp 1679581782
transform 1 0 5280 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_56
timestamp 1679581782
transform 1 0 5952 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_63
timestamp 1679581782
transform 1 0 6624 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_70
timestamp 1679581782
transform 1 0 7296 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_77
timestamp 1679581782
transform 1 0 7968 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_84
timestamp 1679581782
transform 1 0 8640 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_91
timestamp 1679581782
transform 1 0 9312 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_98
timestamp 1679581782
transform 1 0 9984 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_105
timestamp 1679581782
transform 1 0 10656 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_112
timestamp 1679581782
transform 1 0 11328 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_119
timestamp 1679581782
transform 1 0 12000 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_126
timestamp 1679581782
transform 1 0 12672 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_133
timestamp 1679581782
transform 1 0 13344 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_140
timestamp 1679581782
transform 1 0 14016 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_147
timestamp 1679581782
transform 1 0 14688 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_154
timestamp 1679581782
transform 1 0 15360 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_161
timestamp 1679581782
transform 1 0 16032 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_168
timestamp 1679581782
transform 1 0 16704 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_175
timestamp 1679581782
transform 1 0 17376 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_182
timestamp 1679581782
transform 1 0 18048 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_189
timestamp 1679581782
transform 1 0 18720 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_196
timestamp 1679581782
transform 1 0 19392 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_203
timestamp 1679581782
transform 1 0 20064 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_210
timestamp 1679581782
transform 1 0 20736 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_217
timestamp 1679581782
transform 1 0 21408 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_224
timestamp 1679581782
transform 1 0 22080 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_231
timestamp 1679581782
transform 1 0 22752 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_238
timestamp 1679581782
transform 1 0 23424 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_245
timestamp 1679581782
transform 1 0 24096 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_252
timestamp 1679581782
transform 1 0 24768 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_259
timestamp 1679581782
transform 1 0 25440 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_266
timestamp 1679581782
transform 1 0 26112 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_273
timestamp 1679581782
transform 1 0 26784 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_280
timestamp 1679581782
transform 1 0 27456 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_287
timestamp 1679581782
transform 1 0 28128 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_294
timestamp 1679581782
transform 1 0 28800 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_301
timestamp 1679581782
transform 1 0 29472 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_308
timestamp 1679581782
transform 1 0 30144 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_315
timestamp 1679581782
transform 1 0 30816 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_322
timestamp 1679581782
transform 1 0 31488 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_329
timestamp 1679581782
transform 1 0 32160 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_336
timestamp 1679581782
transform 1 0 32832 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_343
timestamp 1679581782
transform 1 0 33504 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_350
timestamp 1679581782
transform 1 0 34176 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_357
timestamp 1679581782
transform 1 0 34848 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_364
timestamp 1679581782
transform 1 0 35520 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_371
timestamp 1679581782
transform 1 0 36192 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_378
timestamp 1679581782
transform 1 0 36864 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_385
timestamp 1679581782
transform 1 0 37536 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_392
timestamp 1679581782
transform 1 0 38208 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_399
timestamp 1679581782
transform 1 0 38880 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_406
timestamp 1679581782
transform 1 0 39552 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_413
timestamp 1679581782
transform 1 0 40224 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_420
timestamp 1679581782
transform 1 0 40896 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_427
timestamp 1679581782
transform 1 0 41568 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_434
timestamp 1679581782
transform 1 0 42240 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_441
timestamp 1679581782
transform 1 0 42912 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_448
timestamp 1679581782
transform 1 0 43584 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_455
timestamp 1679581782
transform 1 0 44256 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_462
timestamp 1679581782
transform 1 0 44928 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_469
timestamp 1679581782
transform 1 0 45600 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_476
timestamp 1679581782
transform 1 0 46272 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_483
timestamp 1679581782
transform 1 0 46944 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_490
timestamp 1679581782
transform 1 0 47616 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_497
timestamp 1679581782
transform 1 0 48288 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_504
timestamp 1679581782
transform 1 0 48960 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_511
timestamp 1679581782
transform 1 0 49632 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_518
timestamp 1679581782
transform 1 0 50304 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_525
timestamp 1679581782
transform 1 0 50976 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_532
timestamp 1679581782
transform 1 0 51648 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_539
timestamp 1679581782
transform 1 0 52320 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_546
timestamp 1679581782
transform 1 0 52992 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_553
timestamp 1679581782
transform 1 0 53664 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_560
timestamp 1679581782
transform 1 0 54336 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_567
timestamp 1679581782
transform 1 0 55008 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_574
timestamp 1679581782
transform 1 0 55680 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_581
timestamp 1679581782
transform 1 0 56352 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_588
timestamp 1679581782
transform 1 0 57024 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_595
timestamp 1679581782
transform 1 0 57696 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_602
timestamp 1679581782
transform 1 0 58368 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_609
timestamp 1679581782
transform 1 0 59040 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_616
timestamp 1679581782
transform 1 0 59712 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_623
timestamp 1679581782
transform 1 0 60384 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_630
timestamp 1679581782
transform 1 0 61056 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_637
timestamp 1679581782
transform 1 0 61728 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_644
timestamp 1679581782
transform 1 0 62400 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_651
timestamp 1679581782
transform 1 0 63072 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_658
timestamp 1679581782
transform 1 0 63744 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_665
timestamp 1679581782
transform 1 0 64416 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_672
timestamp 1679581782
transform 1 0 65088 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_679
timestamp 1679581782
transform 1 0 65760 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_686
timestamp 1679581782
transform 1 0 66432 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_693
timestamp 1679581782
transform 1 0 67104 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_700
timestamp 1679581782
transform 1 0 67776 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_707
timestamp 1679581782
transform 1 0 68448 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_714
timestamp 1679581782
transform 1 0 69120 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_721
timestamp 1679581782
transform 1 0 69792 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_728
timestamp 1679581782
transform 1 0 70464 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_735
timestamp 1679581782
transform 1 0 71136 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_742
timestamp 1679581782
transform 1 0 71808 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_749
timestamp 1679581782
transform 1 0 72480 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_756
timestamp 1679581782
transform 1 0 73152 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_763
timestamp 1679581782
transform 1 0 73824 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_770
timestamp 1679581782
transform 1 0 74496 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_777
timestamp 1679581782
transform 1 0 75168 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_784
timestamp 1679581782
transform 1 0 75840 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_791
timestamp 1679581782
transform 1 0 76512 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_798
timestamp 1679581782
transform 1 0 77184 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_805
timestamp 1679581782
transform 1 0 77856 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_812
timestamp 1679581782
transform 1 0 78528 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_819
timestamp 1679581782
transform 1 0 79200 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_826
timestamp 1679581782
transform 1 0 79872 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_833
timestamp 1679581782
transform 1 0 80544 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_840
timestamp 1679581782
transform 1 0 81216 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_847
timestamp 1679581782
transform 1 0 81888 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_854
timestamp 1679581782
transform 1 0 82560 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_861
timestamp 1679581782
transform 1 0 83232 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_868
timestamp 1679581782
transform 1 0 83904 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_875
timestamp 1679581782
transform 1 0 84576 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_882
timestamp 1679581782
transform 1 0 85248 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_889
timestamp 1679581782
transform 1 0 85920 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_896
timestamp 1679581782
transform 1 0 86592 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_903
timestamp 1679581782
transform 1 0 87264 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_910
timestamp 1679581782
transform 1 0 87936 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_917
timestamp 1679581782
transform 1 0 88608 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_924
timestamp 1679581782
transform 1 0 89280 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_931
timestamp 1679581782
transform 1 0 89952 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_938
timestamp 1679581782
transform 1 0 90624 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_945
timestamp 1679581782
transform 1 0 91296 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_952
timestamp 1679581782
transform 1 0 91968 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_959
timestamp 1679581782
transform 1 0 92640 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_966
timestamp 1679581782
transform 1 0 93312 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_973
timestamp 1679581782
transform 1 0 93984 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_980
timestamp 1679581782
transform 1 0 94656 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_987
timestamp 1679581782
transform 1 0 95328 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_994
timestamp 1679581782
transform 1 0 96000 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_1001
timestamp 1679581782
transform 1 0 96672 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_1008
timestamp 1679581782
transform 1 0 97344 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_1015
timestamp 1679581782
transform 1 0 98016 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_1022
timestamp 1679581782
transform 1 0 98688 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_4
timestamp 1679581782
transform 1 0 960 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_11
timestamp 1679581782
transform 1 0 1632 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_18
timestamp 1679581782
transform 1 0 2304 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_25
timestamp 1679581782
transform 1 0 2976 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_32
timestamp 1679581782
transform 1 0 3648 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_39
timestamp 1679581782
transform 1 0 4320 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_46
timestamp 1679581782
transform 1 0 4992 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_53
timestamp 1679581782
transform 1 0 5664 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_60
timestamp 1679581782
transform 1 0 6336 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_67
timestamp 1679581782
transform 1 0 7008 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_74
timestamp 1679581782
transform 1 0 7680 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_81
timestamp 1679581782
transform 1 0 8352 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_88
timestamp 1679581782
transform 1 0 9024 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_95
timestamp 1679581782
transform 1 0 9696 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_102
timestamp 1679581782
transform 1 0 10368 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_109
timestamp 1679581782
transform 1 0 11040 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_116
timestamp 1679581782
transform 1 0 11712 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_123
timestamp 1679581782
transform 1 0 12384 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_130
timestamp 1679581782
transform 1 0 13056 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_137
timestamp 1679581782
transform 1 0 13728 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_144
timestamp 1679581782
transform 1 0 14400 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_151
timestamp 1679581782
transform 1 0 15072 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_158
timestamp 1679581782
transform 1 0 15744 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_165
timestamp 1679581782
transform 1 0 16416 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_172
timestamp 1679581782
transform 1 0 17088 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_179
timestamp 1679581782
transform 1 0 17760 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_186
timestamp 1679581782
transform 1 0 18432 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_193
timestamp 1679581782
transform 1 0 19104 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_200
timestamp 1679581782
transform 1 0 19776 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_207
timestamp 1679581782
transform 1 0 20448 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_214
timestamp 1679581782
transform 1 0 21120 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_221
timestamp 1679581782
transform 1 0 21792 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_228
timestamp 1679581782
transform 1 0 22464 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_235
timestamp 1679581782
transform 1 0 23136 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_242
timestamp 1679581782
transform 1 0 23808 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_249
timestamp 1679581782
transform 1 0 24480 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_256
timestamp 1679581782
transform 1 0 25152 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_263
timestamp 1679581782
transform 1 0 25824 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_270
timestamp 1679581782
transform 1 0 26496 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_277
timestamp 1679581782
transform 1 0 27168 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_284
timestamp 1679581782
transform 1 0 27840 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_291
timestamp 1679581782
transform 1 0 28512 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_298
timestamp 1679581782
transform 1 0 29184 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_305
timestamp 1679581782
transform 1 0 29856 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_312
timestamp 1679581782
transform 1 0 30528 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_319
timestamp 1679581782
transform 1 0 31200 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_326
timestamp 1679581782
transform 1 0 31872 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_333
timestamp 1679581782
transform 1 0 32544 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_340
timestamp 1679581782
transform 1 0 33216 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_347
timestamp 1679581782
transform 1 0 33888 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_354
timestamp 1679581782
transform 1 0 34560 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_361
timestamp 1679581782
transform 1 0 35232 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_368
timestamp 1679581782
transform 1 0 35904 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_375
timestamp 1679581782
transform 1 0 36576 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_382
timestamp 1679581782
transform 1 0 37248 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_389
timestamp 1679581782
transform 1 0 37920 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_396
timestamp 1679581782
transform 1 0 38592 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_403
timestamp 1679581782
transform 1 0 39264 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_410
timestamp 1679581782
transform 1 0 39936 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_417
timestamp 1679581782
transform 1 0 40608 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_424
timestamp 1679581782
transform 1 0 41280 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_431
timestamp 1679581782
transform 1 0 41952 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_438
timestamp 1679581782
transform 1 0 42624 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_445
timestamp 1679581782
transform 1 0 43296 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_452
timestamp 1679581782
transform 1 0 43968 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_459
timestamp 1679581782
transform 1 0 44640 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_466
timestamp 1679581782
transform 1 0 45312 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_473
timestamp 1679581782
transform 1 0 45984 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_480
timestamp 1679581782
transform 1 0 46656 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_487
timestamp 1679581782
transform 1 0 47328 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_494
timestamp 1679581782
transform 1 0 48000 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_501
timestamp 1679581782
transform 1 0 48672 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_508
timestamp 1679581782
transform 1 0 49344 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_515
timestamp 1679581782
transform 1 0 50016 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_522
timestamp 1679581782
transform 1 0 50688 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_529
timestamp 1679581782
transform 1 0 51360 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_536
timestamp 1679581782
transform 1 0 52032 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_543
timestamp 1679581782
transform 1 0 52704 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_550
timestamp 1679581782
transform 1 0 53376 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_557
timestamp 1679581782
transform 1 0 54048 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_564
timestamp 1679581782
transform 1 0 54720 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_571
timestamp 1679581782
transform 1 0 55392 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_578
timestamp 1679581782
transform 1 0 56064 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_585
timestamp 1679581782
transform 1 0 56736 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_592
timestamp 1679581782
transform 1 0 57408 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_599
timestamp 1679581782
transform 1 0 58080 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_606
timestamp 1679581782
transform 1 0 58752 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_613
timestamp 1679581782
transform 1 0 59424 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_620
timestamp 1679581782
transform 1 0 60096 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_627
timestamp 1679581782
transform 1 0 60768 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_634
timestamp 1679581782
transform 1 0 61440 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_641
timestamp 1679581782
transform 1 0 62112 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_648
timestamp 1679581782
transform 1 0 62784 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_655
timestamp 1679581782
transform 1 0 63456 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_662
timestamp 1679581782
transform 1 0 64128 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_669
timestamp 1679581782
transform 1 0 64800 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_676
timestamp 1679581782
transform 1 0 65472 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_683
timestamp 1679581782
transform 1 0 66144 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_690
timestamp 1679581782
transform 1 0 66816 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_697
timestamp 1679581782
transform 1 0 67488 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_704
timestamp 1679581782
transform 1 0 68160 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_711
timestamp 1679581782
transform 1 0 68832 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_718
timestamp 1679581782
transform 1 0 69504 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_725
timestamp 1679581782
transform 1 0 70176 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_732
timestamp 1679581782
transform 1 0 70848 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_739
timestamp 1679581782
transform 1 0 71520 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_746
timestamp 1679581782
transform 1 0 72192 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_753
timestamp 1679581782
transform 1 0 72864 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_760
timestamp 1679581782
transform 1 0 73536 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_767
timestamp 1679581782
transform 1 0 74208 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_774
timestamp 1679581782
transform 1 0 74880 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_781
timestamp 1679581782
transform 1 0 75552 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_788
timestamp 1679581782
transform 1 0 76224 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_795
timestamp 1679581782
transform 1 0 76896 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_802
timestamp 1679581782
transform 1 0 77568 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_809
timestamp 1679581782
transform 1 0 78240 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_816
timestamp 1679581782
transform 1 0 78912 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_823
timestamp 1679581782
transform 1 0 79584 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_830
timestamp 1679581782
transform 1 0 80256 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_837
timestamp 1679581782
transform 1 0 80928 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_844
timestamp 1679581782
transform 1 0 81600 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_851
timestamp 1679581782
transform 1 0 82272 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_858
timestamp 1679581782
transform 1 0 82944 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_865
timestamp 1679581782
transform 1 0 83616 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_872
timestamp 1679581782
transform 1 0 84288 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_879
timestamp 1679581782
transform 1 0 84960 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_886
timestamp 1679581782
transform 1 0 85632 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_893
timestamp 1679581782
transform 1 0 86304 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_900
timestamp 1679581782
transform 1 0 86976 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_907
timestamp 1679581782
transform 1 0 87648 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_914
timestamp 1679581782
transform 1 0 88320 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_921
timestamp 1679581782
transform 1 0 88992 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_928
timestamp 1679581782
transform 1 0 89664 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_935
timestamp 1679581782
transform 1 0 90336 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_942
timestamp 1679581782
transform 1 0 91008 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_949
timestamp 1679581782
transform 1 0 91680 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_956
timestamp 1679581782
transform 1 0 92352 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_963
timestamp 1679581782
transform 1 0 93024 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_970
timestamp 1679581782
transform 1 0 93696 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_977
timestamp 1679581782
transform 1 0 94368 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_984
timestamp 1679581782
transform 1 0 95040 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_991
timestamp 1679581782
transform 1 0 95712 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_998
timestamp 1679581782
transform 1 0 96384 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_1005
timestamp 1679581782
transform 1 0 97056 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_1012
timestamp 1679581782
transform 1 0 97728 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_1019
timestamp 1679581782
transform 1 0 98400 0 -1 40068
box -48 -56 720 834
use sg13g2_fill_2  FILLER_51_1026
timestamp 1677580104
transform 1 0 99072 0 -1 40068
box -48 -56 240 834
use sg13g2_fill_1  FILLER_51_1028
timestamp 1677579658
transform 1 0 99264 0 -1 40068
box -48 -56 144 834
use sg13g2_decap_8  FILLER_52_0
timestamp 1679581782
transform 1 0 576 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_7
timestamp 1679581782
transform 1 0 1248 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_14
timestamp 1679581782
transform 1 0 1920 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_21
timestamp 1679581782
transform 1 0 2592 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_28
timestamp 1679581782
transform 1 0 3264 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_35
timestamp 1679581782
transform 1 0 3936 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_42
timestamp 1679581782
transform 1 0 4608 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_49
timestamp 1679581782
transform 1 0 5280 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_56
timestamp 1679581782
transform 1 0 5952 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_63
timestamp 1679581782
transform 1 0 6624 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_70
timestamp 1679581782
transform 1 0 7296 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_77
timestamp 1679581782
transform 1 0 7968 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_84
timestamp 1679581782
transform 1 0 8640 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_91
timestamp 1679581782
transform 1 0 9312 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_98
timestamp 1679581782
transform 1 0 9984 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_105
timestamp 1679581782
transform 1 0 10656 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_112
timestamp 1679581782
transform 1 0 11328 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_119
timestamp 1679581782
transform 1 0 12000 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_126
timestamp 1679581782
transform 1 0 12672 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_133
timestamp 1679581782
transform 1 0 13344 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_140
timestamp 1679581782
transform 1 0 14016 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_147
timestamp 1679581782
transform 1 0 14688 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_154
timestamp 1679581782
transform 1 0 15360 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_161
timestamp 1679581782
transform 1 0 16032 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_168
timestamp 1679581782
transform 1 0 16704 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_175
timestamp 1679581782
transform 1 0 17376 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_182
timestamp 1679581782
transform 1 0 18048 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_189
timestamp 1679581782
transform 1 0 18720 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_196
timestamp 1679581782
transform 1 0 19392 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_203
timestamp 1679581782
transform 1 0 20064 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_210
timestamp 1679581782
transform 1 0 20736 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_217
timestamp 1679581782
transform 1 0 21408 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_224
timestamp 1679581782
transform 1 0 22080 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_231
timestamp 1679581782
transform 1 0 22752 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_238
timestamp 1679581782
transform 1 0 23424 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_245
timestamp 1679581782
transform 1 0 24096 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_252
timestamp 1679581782
transform 1 0 24768 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_259
timestamp 1679581782
transform 1 0 25440 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_266
timestamp 1679581782
transform 1 0 26112 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_273
timestamp 1679581782
transform 1 0 26784 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_280
timestamp 1679581782
transform 1 0 27456 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_287
timestamp 1679581782
transform 1 0 28128 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_294
timestamp 1679581782
transform 1 0 28800 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_301
timestamp 1679581782
transform 1 0 29472 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_308
timestamp 1679581782
transform 1 0 30144 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_315
timestamp 1679581782
transform 1 0 30816 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_322
timestamp 1679581782
transform 1 0 31488 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_329
timestamp 1679581782
transform 1 0 32160 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_336
timestamp 1679581782
transform 1 0 32832 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_343
timestamp 1679581782
transform 1 0 33504 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_350
timestamp 1679581782
transform 1 0 34176 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_357
timestamp 1679581782
transform 1 0 34848 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_364
timestamp 1679581782
transform 1 0 35520 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_371
timestamp 1679581782
transform 1 0 36192 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_378
timestamp 1679581782
transform 1 0 36864 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_385
timestamp 1679581782
transform 1 0 37536 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_392
timestamp 1679581782
transform 1 0 38208 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_399
timestamp 1679581782
transform 1 0 38880 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_406
timestamp 1679581782
transform 1 0 39552 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_413
timestamp 1679581782
transform 1 0 40224 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_420
timestamp 1679581782
transform 1 0 40896 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_427
timestamp 1679581782
transform 1 0 41568 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_434
timestamp 1679581782
transform 1 0 42240 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_441
timestamp 1679581782
transform 1 0 42912 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_448
timestamp 1679581782
transform 1 0 43584 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_455
timestamp 1679581782
transform 1 0 44256 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_462
timestamp 1679581782
transform 1 0 44928 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_469
timestamp 1679581782
transform 1 0 45600 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_476
timestamp 1679581782
transform 1 0 46272 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_483
timestamp 1679581782
transform 1 0 46944 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_490
timestamp 1679581782
transform 1 0 47616 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_497
timestamp 1679581782
transform 1 0 48288 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_504
timestamp 1679581782
transform 1 0 48960 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_511
timestamp 1679581782
transform 1 0 49632 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_518
timestamp 1679581782
transform 1 0 50304 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_525
timestamp 1679581782
transform 1 0 50976 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_532
timestamp 1679581782
transform 1 0 51648 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_539
timestamp 1679581782
transform 1 0 52320 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_546
timestamp 1679581782
transform 1 0 52992 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_553
timestamp 1679581782
transform 1 0 53664 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_560
timestamp 1679581782
transform 1 0 54336 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_567
timestamp 1679581782
transform 1 0 55008 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_574
timestamp 1679581782
transform 1 0 55680 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_581
timestamp 1679581782
transform 1 0 56352 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_588
timestamp 1679581782
transform 1 0 57024 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_595
timestamp 1679581782
transform 1 0 57696 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_602
timestamp 1679581782
transform 1 0 58368 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_609
timestamp 1679581782
transform 1 0 59040 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_616
timestamp 1679581782
transform 1 0 59712 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_623
timestamp 1679581782
transform 1 0 60384 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_630
timestamp 1679581782
transform 1 0 61056 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_637
timestamp 1679581782
transform 1 0 61728 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_644
timestamp 1679581782
transform 1 0 62400 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_651
timestamp 1679581782
transform 1 0 63072 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_658
timestamp 1679581782
transform 1 0 63744 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_665
timestamp 1679581782
transform 1 0 64416 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_672
timestamp 1679581782
transform 1 0 65088 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_679
timestamp 1679581782
transform 1 0 65760 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_686
timestamp 1679581782
transform 1 0 66432 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_693
timestamp 1679581782
transform 1 0 67104 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_700
timestamp 1679581782
transform 1 0 67776 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_707
timestamp 1679581782
transform 1 0 68448 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_714
timestamp 1679581782
transform 1 0 69120 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_721
timestamp 1679581782
transform 1 0 69792 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_728
timestamp 1679581782
transform 1 0 70464 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_735
timestamp 1679581782
transform 1 0 71136 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_742
timestamp 1679581782
transform 1 0 71808 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_749
timestamp 1679581782
transform 1 0 72480 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_756
timestamp 1679581782
transform 1 0 73152 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_763
timestamp 1679581782
transform 1 0 73824 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_770
timestamp 1679581782
transform 1 0 74496 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_777
timestamp 1679581782
transform 1 0 75168 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_784
timestamp 1679581782
transform 1 0 75840 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_791
timestamp 1679581782
transform 1 0 76512 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_798
timestamp 1679581782
transform 1 0 77184 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_805
timestamp 1679581782
transform 1 0 77856 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_812
timestamp 1679581782
transform 1 0 78528 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_819
timestamp 1679581782
transform 1 0 79200 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_826
timestamp 1679581782
transform 1 0 79872 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_833
timestamp 1679581782
transform 1 0 80544 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_840
timestamp 1679581782
transform 1 0 81216 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_847
timestamp 1679581782
transform 1 0 81888 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_854
timestamp 1679581782
transform 1 0 82560 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_861
timestamp 1679581782
transform 1 0 83232 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_868
timestamp 1679581782
transform 1 0 83904 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_875
timestamp 1679581782
transform 1 0 84576 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_882
timestamp 1679581782
transform 1 0 85248 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_889
timestamp 1679581782
transform 1 0 85920 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_896
timestamp 1679581782
transform 1 0 86592 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_903
timestamp 1679581782
transform 1 0 87264 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_910
timestamp 1679581782
transform 1 0 87936 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_917
timestamp 1679581782
transform 1 0 88608 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_924
timestamp 1679581782
transform 1 0 89280 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_931
timestamp 1679581782
transform 1 0 89952 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_938
timestamp 1679581782
transform 1 0 90624 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_945
timestamp 1679581782
transform 1 0 91296 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_952
timestamp 1679581782
transform 1 0 91968 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_959
timestamp 1679581782
transform 1 0 92640 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_966
timestamp 1679581782
transform 1 0 93312 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_973
timestamp 1679581782
transform 1 0 93984 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_980
timestamp 1679581782
transform 1 0 94656 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_987
timestamp 1679581782
transform 1 0 95328 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_994
timestamp 1679581782
transform 1 0 96000 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_1001
timestamp 1679581782
transform 1 0 96672 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_1008
timestamp 1679581782
transform 1 0 97344 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_1015
timestamp 1679581782
transform 1 0 98016 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_1022
timestamp 1679581782
transform 1 0 98688 0 1 40068
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_0
timestamp 1679581782
transform 1 0 576 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_7
timestamp 1679581782
transform 1 0 1248 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_14
timestamp 1679581782
transform 1 0 1920 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_21
timestamp 1679581782
transform 1 0 2592 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_28
timestamp 1679581782
transform 1 0 3264 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_35
timestamp 1679581782
transform 1 0 3936 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_42
timestamp 1679581782
transform 1 0 4608 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_49
timestamp 1679581782
transform 1 0 5280 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_56
timestamp 1679581782
transform 1 0 5952 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_63
timestamp 1679581782
transform 1 0 6624 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_70
timestamp 1679581782
transform 1 0 7296 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_77
timestamp 1679581782
transform 1 0 7968 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_84
timestamp 1679581782
transform 1 0 8640 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_91
timestamp 1679581782
transform 1 0 9312 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_98
timestamp 1679581782
transform 1 0 9984 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_105
timestamp 1679581782
transform 1 0 10656 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_112
timestamp 1679581782
transform 1 0 11328 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_119
timestamp 1679581782
transform 1 0 12000 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_126
timestamp 1679581782
transform 1 0 12672 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_133
timestamp 1679581782
transform 1 0 13344 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_140
timestamp 1679581782
transform 1 0 14016 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_147
timestamp 1679581782
transform 1 0 14688 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_154
timestamp 1679581782
transform 1 0 15360 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_161
timestamp 1679581782
transform 1 0 16032 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_168
timestamp 1679581782
transform 1 0 16704 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_175
timestamp 1679581782
transform 1 0 17376 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_182
timestamp 1679581782
transform 1 0 18048 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_189
timestamp 1679581782
transform 1 0 18720 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_196
timestamp 1679581782
transform 1 0 19392 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_203
timestamp 1679581782
transform 1 0 20064 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_210
timestamp 1679581782
transform 1 0 20736 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_217
timestamp 1679581782
transform 1 0 21408 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_224
timestamp 1679581782
transform 1 0 22080 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_231
timestamp 1679581782
transform 1 0 22752 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_238
timestamp 1679581782
transform 1 0 23424 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_245
timestamp 1679581782
transform 1 0 24096 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_252
timestamp 1679581782
transform 1 0 24768 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_259
timestamp 1679581782
transform 1 0 25440 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_266
timestamp 1679581782
transform 1 0 26112 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_273
timestamp 1679581782
transform 1 0 26784 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_280
timestamp 1679581782
transform 1 0 27456 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_287
timestamp 1679581782
transform 1 0 28128 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_294
timestamp 1679581782
transform 1 0 28800 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_301
timestamp 1679581782
transform 1 0 29472 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_308
timestamp 1679581782
transform 1 0 30144 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_315
timestamp 1679581782
transform 1 0 30816 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_322
timestamp 1679581782
transform 1 0 31488 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_329
timestamp 1679581782
transform 1 0 32160 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_336
timestamp 1679581782
transform 1 0 32832 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_343
timestamp 1679581782
transform 1 0 33504 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_350
timestamp 1679581782
transform 1 0 34176 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_357
timestamp 1679581782
transform 1 0 34848 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_364
timestamp 1679581782
transform 1 0 35520 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_371
timestamp 1679581782
transform 1 0 36192 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_378
timestamp 1679581782
transform 1 0 36864 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_385
timestamp 1679581782
transform 1 0 37536 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_392
timestamp 1679581782
transform 1 0 38208 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_399
timestamp 1679581782
transform 1 0 38880 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_406
timestamp 1679581782
transform 1 0 39552 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_413
timestamp 1679581782
transform 1 0 40224 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_420
timestamp 1679581782
transform 1 0 40896 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_427
timestamp 1679581782
transform 1 0 41568 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_434
timestamp 1679581782
transform 1 0 42240 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_441
timestamp 1679581782
transform 1 0 42912 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_448
timestamp 1679581782
transform 1 0 43584 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_455
timestamp 1679581782
transform 1 0 44256 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_462
timestamp 1679581782
transform 1 0 44928 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_469
timestamp 1679581782
transform 1 0 45600 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_476
timestamp 1679581782
transform 1 0 46272 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_483
timestamp 1679581782
transform 1 0 46944 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_490
timestamp 1679581782
transform 1 0 47616 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_497
timestamp 1679581782
transform 1 0 48288 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_504
timestamp 1679581782
transform 1 0 48960 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_511
timestamp 1679581782
transform 1 0 49632 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_518
timestamp 1679581782
transform 1 0 50304 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_525
timestamp 1679581782
transform 1 0 50976 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_532
timestamp 1679581782
transform 1 0 51648 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_539
timestamp 1679581782
transform 1 0 52320 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_546
timestamp 1679581782
transform 1 0 52992 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_553
timestamp 1679581782
transform 1 0 53664 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_560
timestamp 1679581782
transform 1 0 54336 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_567
timestamp 1679581782
transform 1 0 55008 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_574
timestamp 1679581782
transform 1 0 55680 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_581
timestamp 1679581782
transform 1 0 56352 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_588
timestamp 1679581782
transform 1 0 57024 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_595
timestamp 1679581782
transform 1 0 57696 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_602
timestamp 1679581782
transform 1 0 58368 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_609
timestamp 1679581782
transform 1 0 59040 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_616
timestamp 1679581782
transform 1 0 59712 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_623
timestamp 1679581782
transform 1 0 60384 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_630
timestamp 1679581782
transform 1 0 61056 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_637
timestamp 1679581782
transform 1 0 61728 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_644
timestamp 1679581782
transform 1 0 62400 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_651
timestamp 1679581782
transform 1 0 63072 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_658
timestamp 1679581782
transform 1 0 63744 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_665
timestamp 1679581782
transform 1 0 64416 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_672
timestamp 1679581782
transform 1 0 65088 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_679
timestamp 1679581782
transform 1 0 65760 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_686
timestamp 1679581782
transform 1 0 66432 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_693
timestamp 1679581782
transform 1 0 67104 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_700
timestamp 1679581782
transform 1 0 67776 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_707
timestamp 1679581782
transform 1 0 68448 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_714
timestamp 1679581782
transform 1 0 69120 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_721
timestamp 1679581782
transform 1 0 69792 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_728
timestamp 1679581782
transform 1 0 70464 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_735
timestamp 1679581782
transform 1 0 71136 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_742
timestamp 1679581782
transform 1 0 71808 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_749
timestamp 1679581782
transform 1 0 72480 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_756
timestamp 1679581782
transform 1 0 73152 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_763
timestamp 1679581782
transform 1 0 73824 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_770
timestamp 1679581782
transform 1 0 74496 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_777
timestamp 1679581782
transform 1 0 75168 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_784
timestamp 1679581782
transform 1 0 75840 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_791
timestamp 1679581782
transform 1 0 76512 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_798
timestamp 1679581782
transform 1 0 77184 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_805
timestamp 1679581782
transform 1 0 77856 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_812
timestamp 1679581782
transform 1 0 78528 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_819
timestamp 1679581782
transform 1 0 79200 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_826
timestamp 1679581782
transform 1 0 79872 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_833
timestamp 1679581782
transform 1 0 80544 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_840
timestamp 1679581782
transform 1 0 81216 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_847
timestamp 1679581782
transform 1 0 81888 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_854
timestamp 1679581782
transform 1 0 82560 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_861
timestamp 1679581782
transform 1 0 83232 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_868
timestamp 1679581782
transform 1 0 83904 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_875
timestamp 1679581782
transform 1 0 84576 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_882
timestamp 1679581782
transform 1 0 85248 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_889
timestamp 1679581782
transform 1 0 85920 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_896
timestamp 1679581782
transform 1 0 86592 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_903
timestamp 1679581782
transform 1 0 87264 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_910
timestamp 1679581782
transform 1 0 87936 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_917
timestamp 1679581782
transform 1 0 88608 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_924
timestamp 1679581782
transform 1 0 89280 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_931
timestamp 1679581782
transform 1 0 89952 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_938
timestamp 1679581782
transform 1 0 90624 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_945
timestamp 1679581782
transform 1 0 91296 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_952
timestamp 1679581782
transform 1 0 91968 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_959
timestamp 1679581782
transform 1 0 92640 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_966
timestamp 1679581782
transform 1 0 93312 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_973
timestamp 1679581782
transform 1 0 93984 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_980
timestamp 1679581782
transform 1 0 94656 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_987
timestamp 1679581782
transform 1 0 95328 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_994
timestamp 1679581782
transform 1 0 96000 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_1001
timestamp 1679581782
transform 1 0 96672 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_1008
timestamp 1679581782
transform 1 0 97344 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_1015
timestamp 1679581782
transform 1 0 98016 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_1022
timestamp 1679581782
transform 1 0 98688 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_4
timestamp 1679581782
transform 1 0 960 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_11
timestamp 1679581782
transform 1 0 1632 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_18
timestamp 1679581782
transform 1 0 2304 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_25
timestamp 1679581782
transform 1 0 2976 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_32
timestamp 1679581782
transform 1 0 3648 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_39
timestamp 1679581782
transform 1 0 4320 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_46
timestamp 1679581782
transform 1 0 4992 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_53
timestamp 1679581782
transform 1 0 5664 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_60
timestamp 1679581782
transform 1 0 6336 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_67
timestamp 1679581782
transform 1 0 7008 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_74
timestamp 1679581782
transform 1 0 7680 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_81
timestamp 1679581782
transform 1 0 8352 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_88
timestamp 1679581782
transform 1 0 9024 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_95
timestamp 1679581782
transform 1 0 9696 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_102
timestamp 1679581782
transform 1 0 10368 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_109
timestamp 1679581782
transform 1 0 11040 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_116
timestamp 1679581782
transform 1 0 11712 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_123
timestamp 1679581782
transform 1 0 12384 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_130
timestamp 1679581782
transform 1 0 13056 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_137
timestamp 1679581782
transform 1 0 13728 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_144
timestamp 1679581782
transform 1 0 14400 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_151
timestamp 1679581782
transform 1 0 15072 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_158
timestamp 1679581782
transform 1 0 15744 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_165
timestamp 1679581782
transform 1 0 16416 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_172
timestamp 1679581782
transform 1 0 17088 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_179
timestamp 1679581782
transform 1 0 17760 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_186
timestamp 1679581782
transform 1 0 18432 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_193
timestamp 1679581782
transform 1 0 19104 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_200
timestamp 1679581782
transform 1 0 19776 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_207
timestamp 1679581782
transform 1 0 20448 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_214
timestamp 1679581782
transform 1 0 21120 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_221
timestamp 1679581782
transform 1 0 21792 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_228
timestamp 1679581782
transform 1 0 22464 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_235
timestamp 1679581782
transform 1 0 23136 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_242
timestamp 1679581782
transform 1 0 23808 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_249
timestamp 1679581782
transform 1 0 24480 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_256
timestamp 1679581782
transform 1 0 25152 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_263
timestamp 1679581782
transform 1 0 25824 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_270
timestamp 1679581782
transform 1 0 26496 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_277
timestamp 1679581782
transform 1 0 27168 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_284
timestamp 1679581782
transform 1 0 27840 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_291
timestamp 1679581782
transform 1 0 28512 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_298
timestamp 1679581782
transform 1 0 29184 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_305
timestamp 1679581782
transform 1 0 29856 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_312
timestamp 1679581782
transform 1 0 30528 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_319
timestamp 1679581782
transform 1 0 31200 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_326
timestamp 1679581782
transform 1 0 31872 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_333
timestamp 1679581782
transform 1 0 32544 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_340
timestamp 1679581782
transform 1 0 33216 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_347
timestamp 1679581782
transform 1 0 33888 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_354
timestamp 1679581782
transform 1 0 34560 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_361
timestamp 1679581782
transform 1 0 35232 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_368
timestamp 1679581782
transform 1 0 35904 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_375
timestamp 1679581782
transform 1 0 36576 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_382
timestamp 1679581782
transform 1 0 37248 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_389
timestamp 1679581782
transform 1 0 37920 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_396
timestamp 1679581782
transform 1 0 38592 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_403
timestamp 1679581782
transform 1 0 39264 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_410
timestamp 1679581782
transform 1 0 39936 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_417
timestamp 1679581782
transform 1 0 40608 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_424
timestamp 1679581782
transform 1 0 41280 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_431
timestamp 1679581782
transform 1 0 41952 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_438
timestamp 1679581782
transform 1 0 42624 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_445
timestamp 1679581782
transform 1 0 43296 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_452
timestamp 1679581782
transform 1 0 43968 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_459
timestamp 1679581782
transform 1 0 44640 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_466
timestamp 1679581782
transform 1 0 45312 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_473
timestamp 1679581782
transform 1 0 45984 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_480
timestamp 1679581782
transform 1 0 46656 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_487
timestamp 1679581782
transform 1 0 47328 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_494
timestamp 1679581782
transform 1 0 48000 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_501
timestamp 1679581782
transform 1 0 48672 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_508
timestamp 1679581782
transform 1 0 49344 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_515
timestamp 1679581782
transform 1 0 50016 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_522
timestamp 1679581782
transform 1 0 50688 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_529
timestamp 1679581782
transform 1 0 51360 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_536
timestamp 1679581782
transform 1 0 52032 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_543
timestamp 1679581782
transform 1 0 52704 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_550
timestamp 1679581782
transform 1 0 53376 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_557
timestamp 1679581782
transform 1 0 54048 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_564
timestamp 1679581782
transform 1 0 54720 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_571
timestamp 1679581782
transform 1 0 55392 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_578
timestamp 1679581782
transform 1 0 56064 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_585
timestamp 1679581782
transform 1 0 56736 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_592
timestamp 1679581782
transform 1 0 57408 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_599
timestamp 1679581782
transform 1 0 58080 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_606
timestamp 1679581782
transform 1 0 58752 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_613
timestamp 1679581782
transform 1 0 59424 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_620
timestamp 1679581782
transform 1 0 60096 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_627
timestamp 1679581782
transform 1 0 60768 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_634
timestamp 1679581782
transform 1 0 61440 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_641
timestamp 1679581782
transform 1 0 62112 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_648
timestamp 1679581782
transform 1 0 62784 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_655
timestamp 1679581782
transform 1 0 63456 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_662
timestamp 1679581782
transform 1 0 64128 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_669
timestamp 1679581782
transform 1 0 64800 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_676
timestamp 1679581782
transform 1 0 65472 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_683
timestamp 1679581782
transform 1 0 66144 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_690
timestamp 1679581782
transform 1 0 66816 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_697
timestamp 1679581782
transform 1 0 67488 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_704
timestamp 1679581782
transform 1 0 68160 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_711
timestamp 1679581782
transform 1 0 68832 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_718
timestamp 1679581782
transform 1 0 69504 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_725
timestamp 1679581782
transform 1 0 70176 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_732
timestamp 1679581782
transform 1 0 70848 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_739
timestamp 1679581782
transform 1 0 71520 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_746
timestamp 1679581782
transform 1 0 72192 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_753
timestamp 1679581782
transform 1 0 72864 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_760
timestamp 1679581782
transform 1 0 73536 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_767
timestamp 1679581782
transform 1 0 74208 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_774
timestamp 1679581782
transform 1 0 74880 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_781
timestamp 1679581782
transform 1 0 75552 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_788
timestamp 1679581782
transform 1 0 76224 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_795
timestamp 1679581782
transform 1 0 76896 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_802
timestamp 1679581782
transform 1 0 77568 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_809
timestamp 1679581782
transform 1 0 78240 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_816
timestamp 1679581782
transform 1 0 78912 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_823
timestamp 1679581782
transform 1 0 79584 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_830
timestamp 1679581782
transform 1 0 80256 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_837
timestamp 1679581782
transform 1 0 80928 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_844
timestamp 1679581782
transform 1 0 81600 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_851
timestamp 1679581782
transform 1 0 82272 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_858
timestamp 1679581782
transform 1 0 82944 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_865
timestamp 1679581782
transform 1 0 83616 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_872
timestamp 1679581782
transform 1 0 84288 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_879
timestamp 1679581782
transform 1 0 84960 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_886
timestamp 1679581782
transform 1 0 85632 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_893
timestamp 1679581782
transform 1 0 86304 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_900
timestamp 1679581782
transform 1 0 86976 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_907
timestamp 1679581782
transform 1 0 87648 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_914
timestamp 1679581782
transform 1 0 88320 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_921
timestamp 1679581782
transform 1 0 88992 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_928
timestamp 1679581782
transform 1 0 89664 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_935
timestamp 1679581782
transform 1 0 90336 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_942
timestamp 1679581782
transform 1 0 91008 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_949
timestamp 1679581782
transform 1 0 91680 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_956
timestamp 1679581782
transform 1 0 92352 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_963
timestamp 1679581782
transform 1 0 93024 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_970
timestamp 1679581782
transform 1 0 93696 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_977
timestamp 1679581782
transform 1 0 94368 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_984
timestamp 1679581782
transform 1 0 95040 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_991
timestamp 1679581782
transform 1 0 95712 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_998
timestamp 1679581782
transform 1 0 96384 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_1005
timestamp 1679581782
transform 1 0 97056 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_1012
timestamp 1679581782
transform 1 0 97728 0 1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_1019
timestamp 1679581782
transform 1 0 98400 0 1 41580
box -48 -56 720 834
use sg13g2_fill_2  FILLER_54_1026
timestamp 1677580104
transform 1 0 99072 0 1 41580
box -48 -56 240 834
use sg13g2_fill_1  FILLER_54_1028
timestamp 1677579658
transform 1 0 99264 0 1 41580
box -48 -56 144 834
use sg13g2_decap_8  FILLER_55_0
timestamp 1679581782
transform 1 0 576 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_7
timestamp 1679581782
transform 1 0 1248 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_14
timestamp 1679581782
transform 1 0 1920 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_21
timestamp 1679581782
transform 1 0 2592 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_28
timestamp 1679581782
transform 1 0 3264 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_35
timestamp 1679581782
transform 1 0 3936 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_42
timestamp 1679581782
transform 1 0 4608 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_49
timestamp 1679581782
transform 1 0 5280 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_56
timestamp 1679581782
transform 1 0 5952 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_63
timestamp 1679581782
transform 1 0 6624 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_70
timestamp 1679581782
transform 1 0 7296 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_77
timestamp 1679581782
transform 1 0 7968 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_84
timestamp 1679581782
transform 1 0 8640 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_91
timestamp 1679581782
transform 1 0 9312 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_98
timestamp 1679581782
transform 1 0 9984 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_105
timestamp 1679581782
transform 1 0 10656 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_112
timestamp 1679581782
transform 1 0 11328 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_119
timestamp 1679581782
transform 1 0 12000 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_126
timestamp 1679581782
transform 1 0 12672 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_133
timestamp 1679581782
transform 1 0 13344 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_140
timestamp 1679581782
transform 1 0 14016 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_147
timestamp 1679581782
transform 1 0 14688 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_154
timestamp 1679581782
transform 1 0 15360 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_161
timestamp 1679581782
transform 1 0 16032 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_168
timestamp 1679581782
transform 1 0 16704 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_175
timestamp 1679581782
transform 1 0 17376 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_182
timestamp 1679581782
transform 1 0 18048 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_189
timestamp 1679581782
transform 1 0 18720 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_196
timestamp 1679581782
transform 1 0 19392 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_203
timestamp 1679581782
transform 1 0 20064 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_210
timestamp 1679581782
transform 1 0 20736 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_217
timestamp 1679581782
transform 1 0 21408 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_224
timestamp 1679581782
transform 1 0 22080 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_231
timestamp 1679581782
transform 1 0 22752 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_238
timestamp 1679581782
transform 1 0 23424 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_245
timestamp 1679581782
transform 1 0 24096 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_252
timestamp 1679581782
transform 1 0 24768 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_259
timestamp 1679581782
transform 1 0 25440 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_266
timestamp 1679581782
transform 1 0 26112 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_273
timestamp 1679581782
transform 1 0 26784 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_280
timestamp 1679581782
transform 1 0 27456 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_287
timestamp 1679581782
transform 1 0 28128 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_294
timestamp 1679581782
transform 1 0 28800 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_301
timestamp 1679581782
transform 1 0 29472 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_308
timestamp 1679581782
transform 1 0 30144 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_315
timestamp 1679581782
transform 1 0 30816 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_322
timestamp 1679581782
transform 1 0 31488 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_329
timestamp 1679581782
transform 1 0 32160 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_336
timestamp 1679581782
transform 1 0 32832 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_343
timestamp 1679581782
transform 1 0 33504 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_350
timestamp 1679581782
transform 1 0 34176 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_357
timestamp 1679581782
transform 1 0 34848 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_364
timestamp 1679581782
transform 1 0 35520 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_371
timestamp 1679581782
transform 1 0 36192 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_378
timestamp 1679581782
transform 1 0 36864 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_385
timestamp 1679581782
transform 1 0 37536 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_392
timestamp 1679581782
transform 1 0 38208 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_399
timestamp 1679581782
transform 1 0 38880 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_406
timestamp 1679581782
transform 1 0 39552 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_413
timestamp 1679581782
transform 1 0 40224 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_420
timestamp 1679581782
transform 1 0 40896 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_427
timestamp 1679581782
transform 1 0 41568 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_434
timestamp 1679581782
transform 1 0 42240 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_441
timestamp 1679581782
transform 1 0 42912 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_448
timestamp 1679581782
transform 1 0 43584 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_455
timestamp 1679581782
transform 1 0 44256 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_462
timestamp 1679581782
transform 1 0 44928 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_469
timestamp 1679581782
transform 1 0 45600 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_476
timestamp 1679581782
transform 1 0 46272 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_483
timestamp 1679581782
transform 1 0 46944 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_490
timestamp 1679581782
transform 1 0 47616 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_497
timestamp 1679581782
transform 1 0 48288 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_504
timestamp 1679581782
transform 1 0 48960 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_511
timestamp 1679581782
transform 1 0 49632 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_518
timestamp 1679581782
transform 1 0 50304 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_525
timestamp 1679581782
transform 1 0 50976 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_532
timestamp 1679581782
transform 1 0 51648 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_539
timestamp 1679581782
transform 1 0 52320 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_546
timestamp 1679581782
transform 1 0 52992 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_553
timestamp 1679581782
transform 1 0 53664 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_560
timestamp 1679581782
transform 1 0 54336 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_567
timestamp 1679581782
transform 1 0 55008 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_574
timestamp 1679581782
transform 1 0 55680 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_581
timestamp 1679581782
transform 1 0 56352 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_588
timestamp 1679581782
transform 1 0 57024 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_595
timestamp 1679581782
transform 1 0 57696 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_602
timestamp 1679581782
transform 1 0 58368 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_609
timestamp 1679581782
transform 1 0 59040 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_616
timestamp 1679581782
transform 1 0 59712 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_623
timestamp 1679581782
transform 1 0 60384 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_630
timestamp 1679581782
transform 1 0 61056 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_637
timestamp 1679581782
transform 1 0 61728 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_644
timestamp 1679581782
transform 1 0 62400 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_651
timestamp 1679581782
transform 1 0 63072 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_658
timestamp 1679581782
transform 1 0 63744 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_665
timestamp 1679581782
transform 1 0 64416 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_672
timestamp 1679581782
transform 1 0 65088 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_679
timestamp 1679581782
transform 1 0 65760 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_686
timestamp 1679581782
transform 1 0 66432 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_693
timestamp 1679581782
transform 1 0 67104 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_700
timestamp 1679581782
transform 1 0 67776 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_707
timestamp 1679581782
transform 1 0 68448 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_714
timestamp 1679581782
transform 1 0 69120 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_721
timestamp 1679581782
transform 1 0 69792 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_728
timestamp 1679581782
transform 1 0 70464 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_735
timestamp 1679581782
transform 1 0 71136 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_742
timestamp 1679581782
transform 1 0 71808 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_749
timestamp 1679581782
transform 1 0 72480 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_756
timestamp 1679581782
transform 1 0 73152 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_763
timestamp 1679581782
transform 1 0 73824 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_770
timestamp 1679581782
transform 1 0 74496 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_777
timestamp 1679581782
transform 1 0 75168 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_784
timestamp 1679581782
transform 1 0 75840 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_791
timestamp 1679581782
transform 1 0 76512 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_798
timestamp 1679581782
transform 1 0 77184 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_805
timestamp 1679581782
transform 1 0 77856 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_812
timestamp 1679581782
transform 1 0 78528 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_819
timestamp 1679581782
transform 1 0 79200 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_826
timestamp 1679581782
transform 1 0 79872 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_833
timestamp 1679581782
transform 1 0 80544 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_840
timestamp 1679581782
transform 1 0 81216 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_847
timestamp 1679581782
transform 1 0 81888 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_854
timestamp 1679581782
transform 1 0 82560 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_861
timestamp 1679581782
transform 1 0 83232 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_868
timestamp 1679581782
transform 1 0 83904 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_875
timestamp 1679581782
transform 1 0 84576 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_882
timestamp 1679581782
transform 1 0 85248 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_889
timestamp 1679581782
transform 1 0 85920 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_896
timestamp 1679581782
transform 1 0 86592 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_903
timestamp 1679581782
transform 1 0 87264 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_910
timestamp 1679581782
transform 1 0 87936 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_917
timestamp 1679581782
transform 1 0 88608 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_924
timestamp 1679581782
transform 1 0 89280 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_931
timestamp 1679581782
transform 1 0 89952 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_938
timestamp 1679581782
transform 1 0 90624 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_945
timestamp 1679581782
transform 1 0 91296 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_952
timestamp 1679581782
transform 1 0 91968 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_959
timestamp 1679581782
transform 1 0 92640 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_966
timestamp 1679581782
transform 1 0 93312 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_973
timestamp 1679581782
transform 1 0 93984 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_980
timestamp 1679581782
transform 1 0 94656 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_987
timestamp 1679581782
transform 1 0 95328 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_994
timestamp 1679581782
transform 1 0 96000 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_1001
timestamp 1679581782
transform 1 0 96672 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_1008
timestamp 1679581782
transform 1 0 97344 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_1015
timestamp 1679581782
transform 1 0 98016 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_1022
timestamp 1679581782
transform 1 0 98688 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_4
timestamp 1679581782
transform 1 0 960 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_11
timestamp 1679581782
transform 1 0 1632 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_18
timestamp 1679581782
transform 1 0 2304 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_25
timestamp 1679581782
transform 1 0 2976 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_32
timestamp 1679581782
transform 1 0 3648 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_39
timestamp 1679581782
transform 1 0 4320 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_46
timestamp 1679581782
transform 1 0 4992 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_53
timestamp 1679581782
transform 1 0 5664 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_60
timestamp 1679581782
transform 1 0 6336 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_67
timestamp 1679581782
transform 1 0 7008 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_74
timestamp 1679581782
transform 1 0 7680 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_81
timestamp 1679581782
transform 1 0 8352 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_88
timestamp 1679581782
transform 1 0 9024 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_95
timestamp 1679581782
transform 1 0 9696 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_102
timestamp 1679581782
transform 1 0 10368 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_109
timestamp 1679581782
transform 1 0 11040 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_116
timestamp 1679581782
transform 1 0 11712 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_123
timestamp 1679581782
transform 1 0 12384 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_130
timestamp 1679581782
transform 1 0 13056 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_137
timestamp 1679581782
transform 1 0 13728 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_144
timestamp 1679581782
transform 1 0 14400 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_151
timestamp 1679581782
transform 1 0 15072 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_158
timestamp 1679581782
transform 1 0 15744 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_165
timestamp 1679581782
transform 1 0 16416 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_172
timestamp 1679581782
transform 1 0 17088 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_179
timestamp 1679581782
transform 1 0 17760 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_186
timestamp 1679581782
transform 1 0 18432 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_193
timestamp 1679581782
transform 1 0 19104 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_200
timestamp 1679581782
transform 1 0 19776 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_207
timestamp 1679581782
transform 1 0 20448 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_214
timestamp 1679581782
transform 1 0 21120 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_221
timestamp 1679581782
transform 1 0 21792 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_228
timestamp 1679581782
transform 1 0 22464 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_235
timestamp 1679581782
transform 1 0 23136 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_242
timestamp 1679581782
transform 1 0 23808 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_249
timestamp 1679581782
transform 1 0 24480 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_256
timestamp 1679581782
transform 1 0 25152 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_263
timestamp 1679581782
transform 1 0 25824 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_270
timestamp 1679581782
transform 1 0 26496 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_277
timestamp 1679581782
transform 1 0 27168 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_284
timestamp 1679581782
transform 1 0 27840 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_291
timestamp 1679581782
transform 1 0 28512 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_298
timestamp 1679581782
transform 1 0 29184 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_305
timestamp 1679581782
transform 1 0 29856 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_312
timestamp 1679581782
transform 1 0 30528 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_319
timestamp 1679581782
transform 1 0 31200 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_326
timestamp 1679581782
transform 1 0 31872 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_333
timestamp 1679581782
transform 1 0 32544 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_340
timestamp 1679581782
transform 1 0 33216 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_347
timestamp 1679581782
transform 1 0 33888 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_354
timestamp 1679581782
transform 1 0 34560 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_361
timestamp 1679581782
transform 1 0 35232 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_368
timestamp 1679581782
transform 1 0 35904 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_375
timestamp 1679581782
transform 1 0 36576 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_382
timestamp 1679581782
transform 1 0 37248 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_389
timestamp 1679581782
transform 1 0 37920 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_396
timestamp 1679581782
transform 1 0 38592 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_403
timestamp 1679581782
transform 1 0 39264 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_410
timestamp 1679581782
transform 1 0 39936 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_417
timestamp 1679581782
transform 1 0 40608 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_424
timestamp 1679581782
transform 1 0 41280 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_431
timestamp 1679581782
transform 1 0 41952 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_438
timestamp 1679581782
transform 1 0 42624 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_445
timestamp 1679581782
transform 1 0 43296 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_452
timestamp 1679581782
transform 1 0 43968 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_459
timestamp 1679581782
transform 1 0 44640 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_466
timestamp 1679581782
transform 1 0 45312 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_473
timestamp 1679581782
transform 1 0 45984 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_480
timestamp 1679581782
transform 1 0 46656 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_487
timestamp 1679581782
transform 1 0 47328 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_494
timestamp 1679581782
transform 1 0 48000 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_501
timestamp 1679581782
transform 1 0 48672 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_508
timestamp 1679581782
transform 1 0 49344 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_515
timestamp 1679581782
transform 1 0 50016 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_522
timestamp 1679581782
transform 1 0 50688 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_529
timestamp 1679581782
transform 1 0 51360 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_536
timestamp 1679581782
transform 1 0 52032 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_543
timestamp 1679581782
transform 1 0 52704 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_550
timestamp 1679581782
transform 1 0 53376 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_557
timestamp 1679581782
transform 1 0 54048 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_564
timestamp 1679581782
transform 1 0 54720 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_571
timestamp 1679581782
transform 1 0 55392 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_578
timestamp 1679581782
transform 1 0 56064 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_585
timestamp 1679581782
transform 1 0 56736 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_592
timestamp 1679581782
transform 1 0 57408 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_599
timestamp 1679581782
transform 1 0 58080 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_606
timestamp 1679581782
transform 1 0 58752 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_613
timestamp 1679581782
transform 1 0 59424 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_620
timestamp 1679581782
transform 1 0 60096 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_627
timestamp 1679581782
transform 1 0 60768 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_634
timestamp 1679581782
transform 1 0 61440 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_641
timestamp 1679581782
transform 1 0 62112 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_648
timestamp 1679581782
transform 1 0 62784 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_655
timestamp 1679581782
transform 1 0 63456 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_662
timestamp 1679581782
transform 1 0 64128 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_669
timestamp 1679581782
transform 1 0 64800 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_676
timestamp 1679581782
transform 1 0 65472 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_683
timestamp 1679581782
transform 1 0 66144 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_690
timestamp 1679581782
transform 1 0 66816 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_697
timestamp 1679581782
transform 1 0 67488 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_704
timestamp 1679581782
transform 1 0 68160 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_711
timestamp 1679581782
transform 1 0 68832 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_718
timestamp 1679581782
transform 1 0 69504 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_725
timestamp 1679581782
transform 1 0 70176 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_732
timestamp 1679581782
transform 1 0 70848 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_739
timestamp 1679581782
transform 1 0 71520 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_746
timestamp 1679581782
transform 1 0 72192 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_753
timestamp 1679581782
transform 1 0 72864 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_760
timestamp 1679581782
transform 1 0 73536 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_767
timestamp 1679581782
transform 1 0 74208 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_774
timestamp 1679581782
transform 1 0 74880 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_781
timestamp 1679581782
transform 1 0 75552 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_788
timestamp 1679581782
transform 1 0 76224 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_795
timestamp 1679581782
transform 1 0 76896 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_802
timestamp 1679581782
transform 1 0 77568 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_809
timestamp 1679581782
transform 1 0 78240 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_816
timestamp 1679581782
transform 1 0 78912 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_823
timestamp 1679581782
transform 1 0 79584 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_830
timestamp 1679581782
transform 1 0 80256 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_837
timestamp 1679581782
transform 1 0 80928 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_844
timestamp 1679581782
transform 1 0 81600 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_851
timestamp 1679581782
transform 1 0 82272 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_858
timestamp 1679581782
transform 1 0 82944 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_865
timestamp 1679581782
transform 1 0 83616 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_872
timestamp 1679581782
transform 1 0 84288 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_879
timestamp 1679581782
transform 1 0 84960 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_886
timestamp 1679581782
transform 1 0 85632 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_893
timestamp 1679581782
transform 1 0 86304 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_900
timestamp 1679581782
transform 1 0 86976 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_907
timestamp 1679581782
transform 1 0 87648 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_914
timestamp 1679581782
transform 1 0 88320 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_921
timestamp 1679581782
transform 1 0 88992 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_928
timestamp 1679581782
transform 1 0 89664 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_935
timestamp 1679581782
transform 1 0 90336 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_942
timestamp 1679581782
transform 1 0 91008 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_949
timestamp 1679581782
transform 1 0 91680 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_956
timestamp 1679581782
transform 1 0 92352 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_963
timestamp 1679581782
transform 1 0 93024 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_970
timestamp 1679581782
transform 1 0 93696 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_977
timestamp 1679581782
transform 1 0 94368 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_984
timestamp 1679581782
transform 1 0 95040 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_991
timestamp 1679581782
transform 1 0 95712 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_998
timestamp 1679581782
transform 1 0 96384 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_1005
timestamp 1679581782
transform 1 0 97056 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_1012
timestamp 1679581782
transform 1 0 97728 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_1019
timestamp 1679581782
transform 1 0 98400 0 1 43092
box -48 -56 720 834
use sg13g2_fill_2  FILLER_56_1026
timestamp 1677580104
transform 1 0 99072 0 1 43092
box -48 -56 240 834
use sg13g2_fill_1  FILLER_56_1028
timestamp 1677579658
transform 1 0 99264 0 1 43092
box -48 -56 144 834
use sg13g2_decap_8  FILLER_57_0
timestamp 1679581782
transform 1 0 576 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_7
timestamp 1679581782
transform 1 0 1248 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_14
timestamp 1679581782
transform 1 0 1920 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_21
timestamp 1679581782
transform 1 0 2592 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_28
timestamp 1679581782
transform 1 0 3264 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_35
timestamp 1679581782
transform 1 0 3936 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_42
timestamp 1679581782
transform 1 0 4608 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_49
timestamp 1679581782
transform 1 0 5280 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_56
timestamp 1679581782
transform 1 0 5952 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_63
timestamp 1679581782
transform 1 0 6624 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_70
timestamp 1679581782
transform 1 0 7296 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_77
timestamp 1679581782
transform 1 0 7968 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_84
timestamp 1679581782
transform 1 0 8640 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_91
timestamp 1679581782
transform 1 0 9312 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_98
timestamp 1679581782
transform 1 0 9984 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_105
timestamp 1679581782
transform 1 0 10656 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_112
timestamp 1679581782
transform 1 0 11328 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_119
timestamp 1679581782
transform 1 0 12000 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_126
timestamp 1679581782
transform 1 0 12672 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_133
timestamp 1679581782
transform 1 0 13344 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_140
timestamp 1679581782
transform 1 0 14016 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_147
timestamp 1679581782
transform 1 0 14688 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_154
timestamp 1679581782
transform 1 0 15360 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_161
timestamp 1679581782
transform 1 0 16032 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_168
timestamp 1679581782
transform 1 0 16704 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_175
timestamp 1679581782
transform 1 0 17376 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_182
timestamp 1679581782
transform 1 0 18048 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_189
timestamp 1679581782
transform 1 0 18720 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_196
timestamp 1679581782
transform 1 0 19392 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_203
timestamp 1679581782
transform 1 0 20064 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_210
timestamp 1679581782
transform 1 0 20736 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_217
timestamp 1679581782
transform 1 0 21408 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_224
timestamp 1679581782
transform 1 0 22080 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_231
timestamp 1679581782
transform 1 0 22752 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_238
timestamp 1679581782
transform 1 0 23424 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_245
timestamp 1679581782
transform 1 0 24096 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_252
timestamp 1679581782
transform 1 0 24768 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_259
timestamp 1679581782
transform 1 0 25440 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_266
timestamp 1679581782
transform 1 0 26112 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_273
timestamp 1679581782
transform 1 0 26784 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_280
timestamp 1679581782
transform 1 0 27456 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_287
timestamp 1679581782
transform 1 0 28128 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_294
timestamp 1679581782
transform 1 0 28800 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_301
timestamp 1679581782
transform 1 0 29472 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_308
timestamp 1679581782
transform 1 0 30144 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_315
timestamp 1679581782
transform 1 0 30816 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_322
timestamp 1679581782
transform 1 0 31488 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_329
timestamp 1679581782
transform 1 0 32160 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_336
timestamp 1679581782
transform 1 0 32832 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_343
timestamp 1679581782
transform 1 0 33504 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_350
timestamp 1679581782
transform 1 0 34176 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_357
timestamp 1679581782
transform 1 0 34848 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_364
timestamp 1679581782
transform 1 0 35520 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_371
timestamp 1679581782
transform 1 0 36192 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_378
timestamp 1679581782
transform 1 0 36864 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_385
timestamp 1679581782
transform 1 0 37536 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_392
timestamp 1679581782
transform 1 0 38208 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_399
timestamp 1679581782
transform 1 0 38880 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_406
timestamp 1679581782
transform 1 0 39552 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_413
timestamp 1679581782
transform 1 0 40224 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_420
timestamp 1679581782
transform 1 0 40896 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_427
timestamp 1679581782
transform 1 0 41568 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_434
timestamp 1679581782
transform 1 0 42240 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_441
timestamp 1679581782
transform 1 0 42912 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_448
timestamp 1679581782
transform 1 0 43584 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_455
timestamp 1679581782
transform 1 0 44256 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_462
timestamp 1679581782
transform 1 0 44928 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_469
timestamp 1679581782
transform 1 0 45600 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_476
timestamp 1679581782
transform 1 0 46272 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_483
timestamp 1679581782
transform 1 0 46944 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_490
timestamp 1679581782
transform 1 0 47616 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_497
timestamp 1679581782
transform 1 0 48288 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_504
timestamp 1679581782
transform 1 0 48960 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_511
timestamp 1679581782
transform 1 0 49632 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_518
timestamp 1679581782
transform 1 0 50304 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_525
timestamp 1679581782
transform 1 0 50976 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_532
timestamp 1679581782
transform 1 0 51648 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_539
timestamp 1679581782
transform 1 0 52320 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_546
timestamp 1679581782
transform 1 0 52992 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_553
timestamp 1679581782
transform 1 0 53664 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_560
timestamp 1679581782
transform 1 0 54336 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_567
timestamp 1679581782
transform 1 0 55008 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_574
timestamp 1679581782
transform 1 0 55680 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_581
timestamp 1679581782
transform 1 0 56352 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_588
timestamp 1679581782
transform 1 0 57024 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_595
timestamp 1679581782
transform 1 0 57696 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_602
timestamp 1679581782
transform 1 0 58368 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_609
timestamp 1679581782
transform 1 0 59040 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_616
timestamp 1679581782
transform 1 0 59712 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_623
timestamp 1679581782
transform 1 0 60384 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_630
timestamp 1679581782
transform 1 0 61056 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_637
timestamp 1679581782
transform 1 0 61728 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_644
timestamp 1679581782
transform 1 0 62400 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_651
timestamp 1679581782
transform 1 0 63072 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_658
timestamp 1679581782
transform 1 0 63744 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_665
timestamp 1679581782
transform 1 0 64416 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_672
timestamp 1679581782
transform 1 0 65088 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_679
timestamp 1679581782
transform 1 0 65760 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_686
timestamp 1679581782
transform 1 0 66432 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_693
timestamp 1679581782
transform 1 0 67104 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_700
timestamp 1679581782
transform 1 0 67776 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_707
timestamp 1679581782
transform 1 0 68448 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_714
timestamp 1679581782
transform 1 0 69120 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_721
timestamp 1679581782
transform 1 0 69792 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_728
timestamp 1679581782
transform 1 0 70464 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_735
timestamp 1679581782
transform 1 0 71136 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_742
timestamp 1679581782
transform 1 0 71808 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_749
timestamp 1679581782
transform 1 0 72480 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_756
timestamp 1679581782
transform 1 0 73152 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_763
timestamp 1679581782
transform 1 0 73824 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_770
timestamp 1679581782
transform 1 0 74496 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_777
timestamp 1679581782
transform 1 0 75168 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_784
timestamp 1679581782
transform 1 0 75840 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_791
timestamp 1679581782
transform 1 0 76512 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_798
timestamp 1679581782
transform 1 0 77184 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_805
timestamp 1679581782
transform 1 0 77856 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_812
timestamp 1679581782
transform 1 0 78528 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_819
timestamp 1679581782
transform 1 0 79200 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_826
timestamp 1679581782
transform 1 0 79872 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_833
timestamp 1679581782
transform 1 0 80544 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_840
timestamp 1679581782
transform 1 0 81216 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_847
timestamp 1679581782
transform 1 0 81888 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_854
timestamp 1679581782
transform 1 0 82560 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_861
timestamp 1679581782
transform 1 0 83232 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_868
timestamp 1679581782
transform 1 0 83904 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_875
timestamp 1679581782
transform 1 0 84576 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_882
timestamp 1679581782
transform 1 0 85248 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_889
timestamp 1679581782
transform 1 0 85920 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_896
timestamp 1679581782
transform 1 0 86592 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_903
timestamp 1679581782
transform 1 0 87264 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_910
timestamp 1679581782
transform 1 0 87936 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_917
timestamp 1679581782
transform 1 0 88608 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_924
timestamp 1679581782
transform 1 0 89280 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_931
timestamp 1679581782
transform 1 0 89952 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_938
timestamp 1679581782
transform 1 0 90624 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_945
timestamp 1679581782
transform 1 0 91296 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_952
timestamp 1679581782
transform 1 0 91968 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_959
timestamp 1679581782
transform 1 0 92640 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_966
timestamp 1679581782
transform 1 0 93312 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_973
timestamp 1679581782
transform 1 0 93984 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_980
timestamp 1679581782
transform 1 0 94656 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_987
timestamp 1679581782
transform 1 0 95328 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_994
timestamp 1679581782
transform 1 0 96000 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_1001
timestamp 1679581782
transform 1 0 96672 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_1008
timestamp 1679581782
transform 1 0 97344 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_1015
timestamp 1679581782
transform 1 0 98016 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_1022
timestamp 1679581782
transform 1 0 98688 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_0
timestamp 1679581782
transform 1 0 576 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_7
timestamp 1679581782
transform 1 0 1248 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_14
timestamp 1679581782
transform 1 0 1920 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_21
timestamp 1679581782
transform 1 0 2592 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_28
timestamp 1679581782
transform 1 0 3264 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_35
timestamp 1679581782
transform 1 0 3936 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_42
timestamp 1679581782
transform 1 0 4608 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_49
timestamp 1679581782
transform 1 0 5280 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_56
timestamp 1679581782
transform 1 0 5952 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_63
timestamp 1679581782
transform 1 0 6624 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_70
timestamp 1679581782
transform 1 0 7296 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_77
timestamp 1679581782
transform 1 0 7968 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_84
timestamp 1679581782
transform 1 0 8640 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_91
timestamp 1679581782
transform 1 0 9312 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_98
timestamp 1679581782
transform 1 0 9984 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_105
timestamp 1679581782
transform 1 0 10656 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_112
timestamp 1679581782
transform 1 0 11328 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_119
timestamp 1679581782
transform 1 0 12000 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_126
timestamp 1679581782
transform 1 0 12672 0 1 44604
box -48 -56 720 834
use sg13g2_decap_4  FILLER_58_133
timestamp 1679577901
transform 1 0 13344 0 1 44604
box -48 -56 432 834
use sg13g2_fill_2  FILLER_58_137
timestamp 1677580104
transform 1 0 13728 0 1 44604
box -48 -56 240 834
use sg13g2_decap_8  FILLER_58_147
timestamp 1679581782
transform 1 0 14688 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_154
timestamp 1679581782
transform 1 0 15360 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_161
timestamp 1679581782
transform 1 0 16032 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_168
timestamp 1679581782
transform 1 0 16704 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_175
timestamp 1679581782
transform 1 0 17376 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_182
timestamp 1679581782
transform 1 0 18048 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_189
timestamp 1679581782
transform 1 0 18720 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_196
timestamp 1679581782
transform 1 0 19392 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_203
timestamp 1679581782
transform 1 0 20064 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_210
timestamp 1679581782
transform 1 0 20736 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_217
timestamp 1679581782
transform 1 0 21408 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_224
timestamp 1679581782
transform 1 0 22080 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_231
timestamp 1679581782
transform 1 0 22752 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_238
timestamp 1679581782
transform 1 0 23424 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_245
timestamp 1679581782
transform 1 0 24096 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_252
timestamp 1679581782
transform 1 0 24768 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_259
timestamp 1679581782
transform 1 0 25440 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_266
timestamp 1679581782
transform 1 0 26112 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_273
timestamp 1679581782
transform 1 0 26784 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_280
timestamp 1679581782
transform 1 0 27456 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_287
timestamp 1679581782
transform 1 0 28128 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_294
timestamp 1679581782
transform 1 0 28800 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_301
timestamp 1679581782
transform 1 0 29472 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_308
timestamp 1679581782
transform 1 0 30144 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_315
timestamp 1679581782
transform 1 0 30816 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_322
timestamp 1679581782
transform 1 0 31488 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_329
timestamp 1679581782
transform 1 0 32160 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_336
timestamp 1679581782
transform 1 0 32832 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_343
timestamp 1679581782
transform 1 0 33504 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_350
timestamp 1679581782
transform 1 0 34176 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_357
timestamp 1679581782
transform 1 0 34848 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_364
timestamp 1679581782
transform 1 0 35520 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_371
timestamp 1679581782
transform 1 0 36192 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_378
timestamp 1679581782
transform 1 0 36864 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_385
timestamp 1679581782
transform 1 0 37536 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_392
timestamp 1679581782
transform 1 0 38208 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_399
timestamp 1679581782
transform 1 0 38880 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_406
timestamp 1679581782
transform 1 0 39552 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_413
timestamp 1679581782
transform 1 0 40224 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_420
timestamp 1679581782
transform 1 0 40896 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_427
timestamp 1679581782
transform 1 0 41568 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_434
timestamp 1679581782
transform 1 0 42240 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_441
timestamp 1679581782
transform 1 0 42912 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_448
timestamp 1679581782
transform 1 0 43584 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_455
timestamp 1679581782
transform 1 0 44256 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_462
timestamp 1679581782
transform 1 0 44928 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_469
timestamp 1679581782
transform 1 0 45600 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_476
timestamp 1679581782
transform 1 0 46272 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_483
timestamp 1679581782
transform 1 0 46944 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_490
timestamp 1679581782
transform 1 0 47616 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_497
timestamp 1679581782
transform 1 0 48288 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_504
timestamp 1679581782
transform 1 0 48960 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_511
timestamp 1679581782
transform 1 0 49632 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_518
timestamp 1679581782
transform 1 0 50304 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_525
timestamp 1679581782
transform 1 0 50976 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_532
timestamp 1679581782
transform 1 0 51648 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_539
timestamp 1679581782
transform 1 0 52320 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_546
timestamp 1679581782
transform 1 0 52992 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_553
timestamp 1679581782
transform 1 0 53664 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_560
timestamp 1679581782
transform 1 0 54336 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_567
timestamp 1679581782
transform 1 0 55008 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_574
timestamp 1679581782
transform 1 0 55680 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_581
timestamp 1679581782
transform 1 0 56352 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_588
timestamp 1679581782
transform 1 0 57024 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_595
timestamp 1679581782
transform 1 0 57696 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_602
timestamp 1679581782
transform 1 0 58368 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_609
timestamp 1679581782
transform 1 0 59040 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_616
timestamp 1679581782
transform 1 0 59712 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_623
timestamp 1679581782
transform 1 0 60384 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_630
timestamp 1679581782
transform 1 0 61056 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_637
timestamp 1679581782
transform 1 0 61728 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_644
timestamp 1679581782
transform 1 0 62400 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_651
timestamp 1679581782
transform 1 0 63072 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_658
timestamp 1679581782
transform 1 0 63744 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_665
timestamp 1679581782
transform 1 0 64416 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_672
timestamp 1679581782
transform 1 0 65088 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_679
timestamp 1679581782
transform 1 0 65760 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_686
timestamp 1679581782
transform 1 0 66432 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_693
timestamp 1679581782
transform 1 0 67104 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_700
timestamp 1679581782
transform 1 0 67776 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_707
timestamp 1679581782
transform 1 0 68448 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_714
timestamp 1679581782
transform 1 0 69120 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_721
timestamp 1679581782
transform 1 0 69792 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_728
timestamp 1679581782
transform 1 0 70464 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_735
timestamp 1679581782
transform 1 0 71136 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_742
timestamp 1679581782
transform 1 0 71808 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_749
timestamp 1679581782
transform 1 0 72480 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_756
timestamp 1679581782
transform 1 0 73152 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_763
timestamp 1679581782
transform 1 0 73824 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_770
timestamp 1679581782
transform 1 0 74496 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_777
timestamp 1679581782
transform 1 0 75168 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_784
timestamp 1679581782
transform 1 0 75840 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_791
timestamp 1679581782
transform 1 0 76512 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_798
timestamp 1679581782
transform 1 0 77184 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_805
timestamp 1679581782
transform 1 0 77856 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_812
timestamp 1679581782
transform 1 0 78528 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_819
timestamp 1679581782
transform 1 0 79200 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_826
timestamp 1679581782
transform 1 0 79872 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_833
timestamp 1679581782
transform 1 0 80544 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_840
timestamp 1679581782
transform 1 0 81216 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_847
timestamp 1679581782
transform 1 0 81888 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_854
timestamp 1679581782
transform 1 0 82560 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_861
timestamp 1679581782
transform 1 0 83232 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_868
timestamp 1679581782
transform 1 0 83904 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_875
timestamp 1679581782
transform 1 0 84576 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_882
timestamp 1679581782
transform 1 0 85248 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_889
timestamp 1679581782
transform 1 0 85920 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_896
timestamp 1679581782
transform 1 0 86592 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_903
timestamp 1679581782
transform 1 0 87264 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_910
timestamp 1679581782
transform 1 0 87936 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_917
timestamp 1679581782
transform 1 0 88608 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_924
timestamp 1679581782
transform 1 0 89280 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_931
timestamp 1679581782
transform 1 0 89952 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_938
timestamp 1679581782
transform 1 0 90624 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_945
timestamp 1679581782
transform 1 0 91296 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_952
timestamp 1679581782
transform 1 0 91968 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_959
timestamp 1679581782
transform 1 0 92640 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_966
timestamp 1679581782
transform 1 0 93312 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_973
timestamp 1679581782
transform 1 0 93984 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_980
timestamp 1679581782
transform 1 0 94656 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_987
timestamp 1679581782
transform 1 0 95328 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_994
timestamp 1679581782
transform 1 0 96000 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_1001
timestamp 1679581782
transform 1 0 96672 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_1008
timestamp 1679581782
transform 1 0 97344 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_1015
timestamp 1679581782
transform 1 0 98016 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_1022
timestamp 1679581782
transform 1 0 98688 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_4
timestamp 1679581782
transform 1 0 960 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_11
timestamp 1679581782
transform 1 0 1632 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_18
timestamp 1679581782
transform 1 0 2304 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_25
timestamp 1679581782
transform 1 0 2976 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_32
timestamp 1679581782
transform 1 0 3648 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_39
timestamp 1679581782
transform 1 0 4320 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_46
timestamp 1679581782
transform 1 0 4992 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_53
timestamp 1679581782
transform 1 0 5664 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_60
timestamp 1679581782
transform 1 0 6336 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_4  FILLER_59_67
timestamp 1679577901
transform 1 0 7008 0 -1 46116
box -48 -56 432 834
use sg13g2_fill_1  FILLER_59_71
timestamp 1677579658
transform 1 0 7392 0 -1 46116
box -48 -56 144 834
use sg13g2_decap_8  FILLER_59_85
timestamp 1679581782
transform 1 0 8736 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_92
timestamp 1679581782
transform 1 0 9408 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_99
timestamp 1679581782
transform 1 0 10080 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_106
timestamp 1679581782
transform 1 0 10752 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_113
timestamp 1679581782
transform 1 0 11424 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_120
timestamp 1679581782
transform 1 0 12096 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_127
timestamp 1679581782
transform 1 0 12768 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_4  FILLER_59_134
timestamp 1679577901
transform 1 0 13440 0 -1 46116
box -48 -56 432 834
use sg13g2_fill_2  FILLER_59_138
timestamp 1677580104
transform 1 0 13824 0 -1 46116
box -48 -56 240 834
use sg13g2_decap_8  FILLER_59_145
timestamp 1679581782
transform 1 0 14496 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_152
timestamp 1679581782
transform 1 0 15168 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_159
timestamp 1679581782
transform 1 0 15840 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_166
timestamp 1679581782
transform 1 0 16512 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_173
timestamp 1679581782
transform 1 0 17184 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_180
timestamp 1679581782
transform 1 0 17856 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_187
timestamp 1679581782
transform 1 0 18528 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_194
timestamp 1679581782
transform 1 0 19200 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_201
timestamp 1679581782
transform 1 0 19872 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_208
timestamp 1679581782
transform 1 0 20544 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_215
timestamp 1679581782
transform 1 0 21216 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_222
timestamp 1679581782
transform 1 0 21888 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_229
timestamp 1679581782
transform 1 0 22560 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_236
timestamp 1679581782
transform 1 0 23232 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_243
timestamp 1679581782
transform 1 0 23904 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_250
timestamp 1679581782
transform 1 0 24576 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_257
timestamp 1679581782
transform 1 0 25248 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_264
timestamp 1679581782
transform 1 0 25920 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_271
timestamp 1679581782
transform 1 0 26592 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_278
timestamp 1679581782
transform 1 0 27264 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_285
timestamp 1679581782
transform 1 0 27936 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_292
timestamp 1679581782
transform 1 0 28608 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_299
timestamp 1679581782
transform 1 0 29280 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_306
timestamp 1679581782
transform 1 0 29952 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_313
timestamp 1679581782
transform 1 0 30624 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_320
timestamp 1679581782
transform 1 0 31296 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_327
timestamp 1679581782
transform 1 0 31968 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_334
timestamp 1679581782
transform 1 0 32640 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_341
timestamp 1679581782
transform 1 0 33312 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_348
timestamp 1679581782
transform 1 0 33984 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_355
timestamp 1679581782
transform 1 0 34656 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_362
timestamp 1679581782
transform 1 0 35328 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_369
timestamp 1679581782
transform 1 0 36000 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_376
timestamp 1679581782
transform 1 0 36672 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_383
timestamp 1679581782
transform 1 0 37344 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_390
timestamp 1679581782
transform 1 0 38016 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_397
timestamp 1679581782
transform 1 0 38688 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_404
timestamp 1679581782
transform 1 0 39360 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_411
timestamp 1679581782
transform 1 0 40032 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_418
timestamp 1679581782
transform 1 0 40704 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_425
timestamp 1679581782
transform 1 0 41376 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_432
timestamp 1679581782
transform 1 0 42048 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_439
timestamp 1679581782
transform 1 0 42720 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_446
timestamp 1679581782
transform 1 0 43392 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_453
timestamp 1679581782
transform 1 0 44064 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_460
timestamp 1679581782
transform 1 0 44736 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_467
timestamp 1679581782
transform 1 0 45408 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_474
timestamp 1679581782
transform 1 0 46080 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_481
timestamp 1679581782
transform 1 0 46752 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_488
timestamp 1679581782
transform 1 0 47424 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_495
timestamp 1679581782
transform 1 0 48096 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_502
timestamp 1679581782
transform 1 0 48768 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_509
timestamp 1679581782
transform 1 0 49440 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_516
timestamp 1679581782
transform 1 0 50112 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_523
timestamp 1679581782
transform 1 0 50784 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_530
timestamp 1679581782
transform 1 0 51456 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_537
timestamp 1679581782
transform 1 0 52128 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_544
timestamp 1679581782
transform 1 0 52800 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_551
timestamp 1679581782
transform 1 0 53472 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_558
timestamp 1679581782
transform 1 0 54144 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_565
timestamp 1679581782
transform 1 0 54816 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_572
timestamp 1679581782
transform 1 0 55488 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_579
timestamp 1679581782
transform 1 0 56160 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_586
timestamp 1679581782
transform 1 0 56832 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_593
timestamp 1679581782
transform 1 0 57504 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_600
timestamp 1679581782
transform 1 0 58176 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_607
timestamp 1679581782
transform 1 0 58848 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_614
timestamp 1679581782
transform 1 0 59520 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_621
timestamp 1679581782
transform 1 0 60192 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_628
timestamp 1679581782
transform 1 0 60864 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_635
timestamp 1679581782
transform 1 0 61536 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_642
timestamp 1679581782
transform 1 0 62208 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_649
timestamp 1679581782
transform 1 0 62880 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_656
timestamp 1679581782
transform 1 0 63552 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_663
timestamp 1679581782
transform 1 0 64224 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_670
timestamp 1679581782
transform 1 0 64896 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_677
timestamp 1679581782
transform 1 0 65568 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_684
timestamp 1679581782
transform 1 0 66240 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_691
timestamp 1679581782
transform 1 0 66912 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_698
timestamp 1679581782
transform 1 0 67584 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_705
timestamp 1679581782
transform 1 0 68256 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_712
timestamp 1679581782
transform 1 0 68928 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_719
timestamp 1679581782
transform 1 0 69600 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_726
timestamp 1679581782
transform 1 0 70272 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_733
timestamp 1679581782
transform 1 0 70944 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_740
timestamp 1679581782
transform 1 0 71616 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_747
timestamp 1679581782
transform 1 0 72288 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_754
timestamp 1679581782
transform 1 0 72960 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_761
timestamp 1679581782
transform 1 0 73632 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_768
timestamp 1679581782
transform 1 0 74304 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_775
timestamp 1679581782
transform 1 0 74976 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_782
timestamp 1679581782
transform 1 0 75648 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_789
timestamp 1679581782
transform 1 0 76320 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_796
timestamp 1679581782
transform 1 0 76992 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_803
timestamp 1679581782
transform 1 0 77664 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_810
timestamp 1679581782
transform 1 0 78336 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_817
timestamp 1679581782
transform 1 0 79008 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_824
timestamp 1679581782
transform 1 0 79680 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_831
timestamp 1679581782
transform 1 0 80352 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_838
timestamp 1679581782
transform 1 0 81024 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_845
timestamp 1679581782
transform 1 0 81696 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_852
timestamp 1679581782
transform 1 0 82368 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_859
timestamp 1679581782
transform 1 0 83040 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_866
timestamp 1679581782
transform 1 0 83712 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_873
timestamp 1679581782
transform 1 0 84384 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_880
timestamp 1679581782
transform 1 0 85056 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_887
timestamp 1679581782
transform 1 0 85728 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_894
timestamp 1679581782
transform 1 0 86400 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_901
timestamp 1679581782
transform 1 0 87072 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_908
timestamp 1679581782
transform 1 0 87744 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_915
timestamp 1679581782
transform 1 0 88416 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_922
timestamp 1679581782
transform 1 0 89088 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_929
timestamp 1679581782
transform 1 0 89760 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_936
timestamp 1679581782
transform 1 0 90432 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_943
timestamp 1679581782
transform 1 0 91104 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_950
timestamp 1679581782
transform 1 0 91776 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_957
timestamp 1679581782
transform 1 0 92448 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_964
timestamp 1679581782
transform 1 0 93120 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_971
timestamp 1679581782
transform 1 0 93792 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_978
timestamp 1679581782
transform 1 0 94464 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_985
timestamp 1679581782
transform 1 0 95136 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_992
timestamp 1679581782
transform 1 0 95808 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_999
timestamp 1679581782
transform 1 0 96480 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_1006
timestamp 1679581782
transform 1 0 97152 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_1013
timestamp 1679581782
transform 1 0 97824 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_1020
timestamp 1679581782
transform 1 0 98496 0 -1 46116
box -48 -56 720 834
use sg13g2_fill_2  FILLER_59_1027
timestamp 1677580104
transform 1 0 99168 0 -1 46116
box -48 -56 240 834
use sg13g2_decap_8  FILLER_60_0
timestamp 1679581782
transform 1 0 576 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_7
timestamp 1679581782
transform 1 0 1248 0 1 46116
box -48 -56 720 834
use sg13g2_decap_4  FILLER_60_14
timestamp 1679577901
transform 1 0 1920 0 1 46116
box -48 -56 432 834
use sg13g2_fill_2  FILLER_60_18
timestamp 1677580104
transform 1 0 2304 0 1 46116
box -48 -56 240 834
use sg13g2_decap_8  FILLER_60_25
timestamp 1679581782
transform 1 0 2976 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_32
timestamp 1679581782
transform 1 0 3648 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_39
timestamp 1679581782
transform 1 0 4320 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_46
timestamp 1679581782
transform 1 0 4992 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_53
timestamp 1679581782
transform 1 0 5664 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_60
timestamp 1679581782
transform 1 0 6336 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_67
timestamp 1679581782
transform 1 0 7008 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_74
timestamp 1679581782
transform 1 0 7680 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_81
timestamp 1679581782
transform 1 0 8352 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_88
timestamp 1679581782
transform 1 0 9024 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_95
timestamp 1679581782
transform 1 0 9696 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_102
timestamp 1679581782
transform 1 0 10368 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_109
timestamp 1679581782
transform 1 0 11040 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_116
timestamp 1679581782
transform 1 0 11712 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_123
timestamp 1679581782
transform 1 0 12384 0 1 46116
box -48 -56 720 834
use sg13g2_decap_4  FILLER_60_130
timestamp 1679577901
transform 1 0 13056 0 1 46116
box -48 -56 432 834
use sg13g2_fill_2  FILLER_60_134
timestamp 1677580104
transform 1 0 13440 0 1 46116
box -48 -56 240 834
use sg13g2_decap_8  FILLER_60_144
timestamp 1679581782
transform 1 0 14400 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_151
timestamp 1679581782
transform 1 0 15072 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_158
timestamp 1679581782
transform 1 0 15744 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_165
timestamp 1679581782
transform 1 0 16416 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_172
timestamp 1679581782
transform 1 0 17088 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_179
timestamp 1679581782
transform 1 0 17760 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_186
timestamp 1679581782
transform 1 0 18432 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_193
timestamp 1679581782
transform 1 0 19104 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_200
timestamp 1679581782
transform 1 0 19776 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_207
timestamp 1679581782
transform 1 0 20448 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_214
timestamp 1679581782
transform 1 0 21120 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_221
timestamp 1679581782
transform 1 0 21792 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_228
timestamp 1679581782
transform 1 0 22464 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_235
timestamp 1679581782
transform 1 0 23136 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_242
timestamp 1679581782
transform 1 0 23808 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_249
timestamp 1679581782
transform 1 0 24480 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_256
timestamp 1679581782
transform 1 0 25152 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_263
timestamp 1679581782
transform 1 0 25824 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_270
timestamp 1679581782
transform 1 0 26496 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_277
timestamp 1679581782
transform 1 0 27168 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_284
timestamp 1679581782
transform 1 0 27840 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_291
timestamp 1679581782
transform 1 0 28512 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_298
timestamp 1679581782
transform 1 0 29184 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_305
timestamp 1679581782
transform 1 0 29856 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_312
timestamp 1679581782
transform 1 0 30528 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_319
timestamp 1679581782
transform 1 0 31200 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_326
timestamp 1679581782
transform 1 0 31872 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_333
timestamp 1679581782
transform 1 0 32544 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_340
timestamp 1679581782
transform 1 0 33216 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_347
timestamp 1679581782
transform 1 0 33888 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_354
timestamp 1679581782
transform 1 0 34560 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_361
timestamp 1679581782
transform 1 0 35232 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_368
timestamp 1679581782
transform 1 0 35904 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_375
timestamp 1679581782
transform 1 0 36576 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_382
timestamp 1679581782
transform 1 0 37248 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_389
timestamp 1679581782
transform 1 0 37920 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_396
timestamp 1679581782
transform 1 0 38592 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_403
timestamp 1679581782
transform 1 0 39264 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_410
timestamp 1679581782
transform 1 0 39936 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_417
timestamp 1679581782
transform 1 0 40608 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_424
timestamp 1679581782
transform 1 0 41280 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_431
timestamp 1679581782
transform 1 0 41952 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_438
timestamp 1679581782
transform 1 0 42624 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_445
timestamp 1679581782
transform 1 0 43296 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_452
timestamp 1679581782
transform 1 0 43968 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_459
timestamp 1679581782
transform 1 0 44640 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_466
timestamp 1679581782
transform 1 0 45312 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_473
timestamp 1679581782
transform 1 0 45984 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_480
timestamp 1679581782
transform 1 0 46656 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_487
timestamp 1679581782
transform 1 0 47328 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_494
timestamp 1679581782
transform 1 0 48000 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_501
timestamp 1679581782
transform 1 0 48672 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_508
timestamp 1679581782
transform 1 0 49344 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_515
timestamp 1679581782
transform 1 0 50016 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_522
timestamp 1679581782
transform 1 0 50688 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_529
timestamp 1679581782
transform 1 0 51360 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_536
timestamp 1679581782
transform 1 0 52032 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_543
timestamp 1679581782
transform 1 0 52704 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_550
timestamp 1679581782
transform 1 0 53376 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_557
timestamp 1679581782
transform 1 0 54048 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_564
timestamp 1679581782
transform 1 0 54720 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_571
timestamp 1679581782
transform 1 0 55392 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_578
timestamp 1679581782
transform 1 0 56064 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_585
timestamp 1679581782
transform 1 0 56736 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_592
timestamp 1679581782
transform 1 0 57408 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_599
timestamp 1679581782
transform 1 0 58080 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_606
timestamp 1679581782
transform 1 0 58752 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_613
timestamp 1679581782
transform 1 0 59424 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_620
timestamp 1679581782
transform 1 0 60096 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_627
timestamp 1679581782
transform 1 0 60768 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_634
timestamp 1679581782
transform 1 0 61440 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_641
timestamp 1679581782
transform 1 0 62112 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_648
timestamp 1679581782
transform 1 0 62784 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_655
timestamp 1679581782
transform 1 0 63456 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_662
timestamp 1679581782
transform 1 0 64128 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_669
timestamp 1679581782
transform 1 0 64800 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_676
timestamp 1679581782
transform 1 0 65472 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_683
timestamp 1679581782
transform 1 0 66144 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_690
timestamp 1679581782
transform 1 0 66816 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_697
timestamp 1679581782
transform 1 0 67488 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_704
timestamp 1679581782
transform 1 0 68160 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_711
timestamp 1679581782
transform 1 0 68832 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_718
timestamp 1679581782
transform 1 0 69504 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_725
timestamp 1679581782
transform 1 0 70176 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_732
timestamp 1679581782
transform 1 0 70848 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_739
timestamp 1679581782
transform 1 0 71520 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_746
timestamp 1679581782
transform 1 0 72192 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_753
timestamp 1679581782
transform 1 0 72864 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_760
timestamp 1679581782
transform 1 0 73536 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_767
timestamp 1679581782
transform 1 0 74208 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_774
timestamp 1679581782
transform 1 0 74880 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_781
timestamp 1679581782
transform 1 0 75552 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_788
timestamp 1679581782
transform 1 0 76224 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_795
timestamp 1679581782
transform 1 0 76896 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_802
timestamp 1679581782
transform 1 0 77568 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_809
timestamp 1679581782
transform 1 0 78240 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_816
timestamp 1679581782
transform 1 0 78912 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_823
timestamp 1679581782
transform 1 0 79584 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_830
timestamp 1679581782
transform 1 0 80256 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_837
timestamp 1679581782
transform 1 0 80928 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_844
timestamp 1679581782
transform 1 0 81600 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_851
timestamp 1679581782
transform 1 0 82272 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_858
timestamp 1679581782
transform 1 0 82944 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_865
timestamp 1679581782
transform 1 0 83616 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_872
timestamp 1679581782
transform 1 0 84288 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_879
timestamp 1679581782
transform 1 0 84960 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_886
timestamp 1679581782
transform 1 0 85632 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_893
timestamp 1679581782
transform 1 0 86304 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_900
timestamp 1679581782
transform 1 0 86976 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_907
timestamp 1679581782
transform 1 0 87648 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_914
timestamp 1679581782
transform 1 0 88320 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_921
timestamp 1679581782
transform 1 0 88992 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_928
timestamp 1679581782
transform 1 0 89664 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_935
timestamp 1679581782
transform 1 0 90336 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_942
timestamp 1679581782
transform 1 0 91008 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_949
timestamp 1679581782
transform 1 0 91680 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_956
timestamp 1679581782
transform 1 0 92352 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_963
timestamp 1679581782
transform 1 0 93024 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_970
timestamp 1679581782
transform 1 0 93696 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_977
timestamp 1679581782
transform 1 0 94368 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_984
timestamp 1679581782
transform 1 0 95040 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_991
timestamp 1679581782
transform 1 0 95712 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_998
timestamp 1679581782
transform 1 0 96384 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_1005
timestamp 1679581782
transform 1 0 97056 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_1012
timestamp 1679581782
transform 1 0 97728 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_1019
timestamp 1679581782
transform 1 0 98400 0 1 46116
box -48 -56 720 834
use sg13g2_fill_2  FILLER_60_1026
timestamp 1677580104
transform 1 0 99072 0 1 46116
box -48 -56 240 834
use sg13g2_fill_1  FILLER_60_1028
timestamp 1677579658
transform 1 0 99264 0 1 46116
box -48 -56 144 834
use sg13g2_decap_8  FILLER_61_4
timestamp 1679581782
transform 1 0 960 0 -1 47628
box -48 -56 720 834
use sg13g2_fill_2  FILLER_61_11
timestamp 1677580104
transform 1 0 1632 0 -1 47628
box -48 -56 240 834
use sg13g2_fill_1  FILLER_61_13
timestamp 1677579658
transform 1 0 1824 0 -1 47628
box -48 -56 144 834
use sg13g2_decap_4  FILLER_61_27
timestamp 1679577901
transform 1 0 3168 0 -1 47628
box -48 -56 432 834
use sg13g2_fill_1  FILLER_61_31
timestamp 1677579658
transform 1 0 3552 0 -1 47628
box -48 -56 144 834
use sg13g2_decap_8  FILLER_61_37
timestamp 1679581782
transform 1 0 4128 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_44
timestamp 1679581782
transform 1 0 4800 0 -1 47628
box -48 -56 720 834
use sg13g2_fill_2  FILLER_61_68
timestamp 1677580104
transform 1 0 7104 0 -1 47628
box -48 -56 240 834
use sg13g2_decap_8  FILLER_61_74
timestamp 1679581782
transform 1 0 7680 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_81
timestamp 1679581782
transform 1 0 8352 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_88
timestamp 1679581782
transform 1 0 9024 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_95
timestamp 1679581782
transform 1 0 9696 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_102
timestamp 1679581782
transform 1 0 10368 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_109
timestamp 1679581782
transform 1 0 11040 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_116
timestamp 1679581782
transform 1 0 11712 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_123
timestamp 1679581782
transform 1 0 12384 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_151
timestamp 1679581782
transform 1 0 15072 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_158
timestamp 1679581782
transform 1 0 15744 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_165
timestamp 1679581782
transform 1 0 16416 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_172
timestamp 1679581782
transform 1 0 17088 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_179
timestamp 1679581782
transform 1 0 17760 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_186
timestamp 1679581782
transform 1 0 18432 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_193
timestamp 1679581782
transform 1 0 19104 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_200
timestamp 1679581782
transform 1 0 19776 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_207
timestamp 1679581782
transform 1 0 20448 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_214
timestamp 1679581782
transform 1 0 21120 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_221
timestamp 1679581782
transform 1 0 21792 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_228
timestamp 1679581782
transform 1 0 22464 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_235
timestamp 1679581782
transform 1 0 23136 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_242
timestamp 1679581782
transform 1 0 23808 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_249
timestamp 1679581782
transform 1 0 24480 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_256
timestamp 1679581782
transform 1 0 25152 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_263
timestamp 1679581782
transform 1 0 25824 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_270
timestamp 1679581782
transform 1 0 26496 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_277
timestamp 1679581782
transform 1 0 27168 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_284
timestamp 1679581782
transform 1 0 27840 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_291
timestamp 1679581782
transform 1 0 28512 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_298
timestamp 1679581782
transform 1 0 29184 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_305
timestamp 1679581782
transform 1 0 29856 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_312
timestamp 1679581782
transform 1 0 30528 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_319
timestamp 1679581782
transform 1 0 31200 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_326
timestamp 1679581782
transform 1 0 31872 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_333
timestamp 1679581782
transform 1 0 32544 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_340
timestamp 1679581782
transform 1 0 33216 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_347
timestamp 1679581782
transform 1 0 33888 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_354
timestamp 1679581782
transform 1 0 34560 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_361
timestamp 1679581782
transform 1 0 35232 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_368
timestamp 1679581782
transform 1 0 35904 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_375
timestamp 1679581782
transform 1 0 36576 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_382
timestamp 1679581782
transform 1 0 37248 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_389
timestamp 1679581782
transform 1 0 37920 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_396
timestamp 1679581782
transform 1 0 38592 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_403
timestamp 1679581782
transform 1 0 39264 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_410
timestamp 1679581782
transform 1 0 39936 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_417
timestamp 1679581782
transform 1 0 40608 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_424
timestamp 1679581782
transform 1 0 41280 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_431
timestamp 1679581782
transform 1 0 41952 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_438
timestamp 1679581782
transform 1 0 42624 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_445
timestamp 1679581782
transform 1 0 43296 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_452
timestamp 1679581782
transform 1 0 43968 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_459
timestamp 1679581782
transform 1 0 44640 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_466
timestamp 1679581782
transform 1 0 45312 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_473
timestamp 1679581782
transform 1 0 45984 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_480
timestamp 1679581782
transform 1 0 46656 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_487
timestamp 1679581782
transform 1 0 47328 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_494
timestamp 1679581782
transform 1 0 48000 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_501
timestamp 1679581782
transform 1 0 48672 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_508
timestamp 1679581782
transform 1 0 49344 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_515
timestamp 1679581782
transform 1 0 50016 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_522
timestamp 1679581782
transform 1 0 50688 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_529
timestamp 1679581782
transform 1 0 51360 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_536
timestamp 1679581782
transform 1 0 52032 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_543
timestamp 1679581782
transform 1 0 52704 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_550
timestamp 1679581782
transform 1 0 53376 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_557
timestamp 1679581782
transform 1 0 54048 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_564
timestamp 1679581782
transform 1 0 54720 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_571
timestamp 1679581782
transform 1 0 55392 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_578
timestamp 1679581782
transform 1 0 56064 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_585
timestamp 1679581782
transform 1 0 56736 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_592
timestamp 1679581782
transform 1 0 57408 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_599
timestamp 1679581782
transform 1 0 58080 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_606
timestamp 1679581782
transform 1 0 58752 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_613
timestamp 1679581782
transform 1 0 59424 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_620
timestamp 1679581782
transform 1 0 60096 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_627
timestamp 1679581782
transform 1 0 60768 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_634
timestamp 1679581782
transform 1 0 61440 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_641
timestamp 1679581782
transform 1 0 62112 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_648
timestamp 1679581782
transform 1 0 62784 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_655
timestamp 1679581782
transform 1 0 63456 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_662
timestamp 1679581782
transform 1 0 64128 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_669
timestamp 1679581782
transform 1 0 64800 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_676
timestamp 1679581782
transform 1 0 65472 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_683
timestamp 1679581782
transform 1 0 66144 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_690
timestamp 1679581782
transform 1 0 66816 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_697
timestamp 1679581782
transform 1 0 67488 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_704
timestamp 1679581782
transform 1 0 68160 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_711
timestamp 1679581782
transform 1 0 68832 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_718
timestamp 1679581782
transform 1 0 69504 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_725
timestamp 1679581782
transform 1 0 70176 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_732
timestamp 1679581782
transform 1 0 70848 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_739
timestamp 1679581782
transform 1 0 71520 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_746
timestamp 1679581782
transform 1 0 72192 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_753
timestamp 1679581782
transform 1 0 72864 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_760
timestamp 1679581782
transform 1 0 73536 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_767
timestamp 1679581782
transform 1 0 74208 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_774
timestamp 1679581782
transform 1 0 74880 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_781
timestamp 1679581782
transform 1 0 75552 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_788
timestamp 1679581782
transform 1 0 76224 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_795
timestamp 1679581782
transform 1 0 76896 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_802
timestamp 1679581782
transform 1 0 77568 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_809
timestamp 1679581782
transform 1 0 78240 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_816
timestamp 1679581782
transform 1 0 78912 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_823
timestamp 1679581782
transform 1 0 79584 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_830
timestamp 1679581782
transform 1 0 80256 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_837
timestamp 1679581782
transform 1 0 80928 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_844
timestamp 1679581782
transform 1 0 81600 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_851
timestamp 1679581782
transform 1 0 82272 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_858
timestamp 1679581782
transform 1 0 82944 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_865
timestamp 1679581782
transform 1 0 83616 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_872
timestamp 1679581782
transform 1 0 84288 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_879
timestamp 1679581782
transform 1 0 84960 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_886
timestamp 1679581782
transform 1 0 85632 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_893
timestamp 1679581782
transform 1 0 86304 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_900
timestamp 1679581782
transform 1 0 86976 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_907
timestamp 1679581782
transform 1 0 87648 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_914
timestamp 1679581782
transform 1 0 88320 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_921
timestamp 1679581782
transform 1 0 88992 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_928
timestamp 1679581782
transform 1 0 89664 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_935
timestamp 1679581782
transform 1 0 90336 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_942
timestamp 1679581782
transform 1 0 91008 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_949
timestamp 1679581782
transform 1 0 91680 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_956
timestamp 1679581782
transform 1 0 92352 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_963
timestamp 1679581782
transform 1 0 93024 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_970
timestamp 1679581782
transform 1 0 93696 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_977
timestamp 1679581782
transform 1 0 94368 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_984
timestamp 1679581782
transform 1 0 95040 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_991
timestamp 1679581782
transform 1 0 95712 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_998
timestamp 1679581782
transform 1 0 96384 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_1005
timestamp 1679581782
transform 1 0 97056 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_1012
timestamp 1679581782
transform 1 0 97728 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_1019
timestamp 1679581782
transform 1 0 98400 0 -1 47628
box -48 -56 720 834
use sg13g2_fill_2  FILLER_61_1026
timestamp 1677580104
transform 1 0 99072 0 -1 47628
box -48 -56 240 834
use sg13g2_fill_1  FILLER_61_1028
timestamp 1677579658
transform 1 0 99264 0 -1 47628
box -48 -56 144 834
use sg13g2_decap_8  FILLER_62_0
timestamp 1679581782
transform 1 0 576 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_7
timestamp 1679581782
transform 1 0 1248 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_14
timestamp 1679581782
transform 1 0 1920 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_21
timestamp 1679581782
transform 1 0 2592 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_28
timestamp 1679581782
transform 1 0 3264 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_35
timestamp 1679581782
transform 1 0 3936 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_42
timestamp 1679581782
transform 1 0 4608 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_49
timestamp 1679581782
transform 1 0 5280 0 1 47628
box -48 -56 720 834
use sg13g2_fill_1  FILLER_62_56
timestamp 1677579658
transform 1 0 5952 0 1 47628
box -48 -56 144 834
use sg13g2_decap_8  FILLER_62_62
timestamp 1679581782
transform 1 0 6528 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_69
timestamp 1679581782
transform 1 0 7200 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_76
timestamp 1679581782
transform 1 0 7872 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_83
timestamp 1679581782
transform 1 0 8544 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_98
timestamp 1679581782
transform 1 0 9984 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_105
timestamp 1679581782
transform 1 0 10656 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_112
timestamp 1679581782
transform 1 0 11328 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_119
timestamp 1679581782
transform 1 0 12000 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_126
timestamp 1679581782
transform 1 0 12672 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_133
timestamp 1679581782
transform 1 0 13344 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_140
timestamp 1679581782
transform 1 0 14016 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_147
timestamp 1679581782
transform 1 0 14688 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_154
timestamp 1679581782
transform 1 0 15360 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_161
timestamp 1679581782
transform 1 0 16032 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_168
timestamp 1679581782
transform 1 0 16704 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_175
timestamp 1679581782
transform 1 0 17376 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_182
timestamp 1679581782
transform 1 0 18048 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_189
timestamp 1679581782
transform 1 0 18720 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_196
timestamp 1679581782
transform 1 0 19392 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_203
timestamp 1679581782
transform 1 0 20064 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_210
timestamp 1679581782
transform 1 0 20736 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_217
timestamp 1679581782
transform 1 0 21408 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_224
timestamp 1679581782
transform 1 0 22080 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_231
timestamp 1679581782
transform 1 0 22752 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_238
timestamp 1679581782
transform 1 0 23424 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_245
timestamp 1679581782
transform 1 0 24096 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_252
timestamp 1679581782
transform 1 0 24768 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_259
timestamp 1679581782
transform 1 0 25440 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_266
timestamp 1679581782
transform 1 0 26112 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_273
timestamp 1679581782
transform 1 0 26784 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_280
timestamp 1679581782
transform 1 0 27456 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_287
timestamp 1679581782
transform 1 0 28128 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_294
timestamp 1679581782
transform 1 0 28800 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_301
timestamp 1679581782
transform 1 0 29472 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_308
timestamp 1679581782
transform 1 0 30144 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_315
timestamp 1679581782
transform 1 0 30816 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_322
timestamp 1679581782
transform 1 0 31488 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_329
timestamp 1679581782
transform 1 0 32160 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_336
timestamp 1679581782
transform 1 0 32832 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_343
timestamp 1679581782
transform 1 0 33504 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_350
timestamp 1679581782
transform 1 0 34176 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_357
timestamp 1679581782
transform 1 0 34848 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_364
timestamp 1679581782
transform 1 0 35520 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_371
timestamp 1679581782
transform 1 0 36192 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_378
timestamp 1679581782
transform 1 0 36864 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_385
timestamp 1679581782
transform 1 0 37536 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_392
timestamp 1679581782
transform 1 0 38208 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_399
timestamp 1679581782
transform 1 0 38880 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_406
timestamp 1679581782
transform 1 0 39552 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_413
timestamp 1679581782
transform 1 0 40224 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_420
timestamp 1679581782
transform 1 0 40896 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_427
timestamp 1679581782
transform 1 0 41568 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_434
timestamp 1679581782
transform 1 0 42240 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_441
timestamp 1679581782
transform 1 0 42912 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_448
timestamp 1679581782
transform 1 0 43584 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_455
timestamp 1679581782
transform 1 0 44256 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_462
timestamp 1679581782
transform 1 0 44928 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_469
timestamp 1679581782
transform 1 0 45600 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_476
timestamp 1679581782
transform 1 0 46272 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_483
timestamp 1679581782
transform 1 0 46944 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_490
timestamp 1679581782
transform 1 0 47616 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_497
timestamp 1679581782
transform 1 0 48288 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_504
timestamp 1679581782
transform 1 0 48960 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_511
timestamp 1679581782
transform 1 0 49632 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_518
timestamp 1679581782
transform 1 0 50304 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_525
timestamp 1679581782
transform 1 0 50976 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_532
timestamp 1679581782
transform 1 0 51648 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_539
timestamp 1679581782
transform 1 0 52320 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_546
timestamp 1679581782
transform 1 0 52992 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_553
timestamp 1679581782
transform 1 0 53664 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_560
timestamp 1679581782
transform 1 0 54336 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_567
timestamp 1679581782
transform 1 0 55008 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_574
timestamp 1679581782
transform 1 0 55680 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_581
timestamp 1679581782
transform 1 0 56352 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_588
timestamp 1679581782
transform 1 0 57024 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_595
timestamp 1679581782
transform 1 0 57696 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_602
timestamp 1679581782
transform 1 0 58368 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_609
timestamp 1679581782
transform 1 0 59040 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_616
timestamp 1679581782
transform 1 0 59712 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_623
timestamp 1679581782
transform 1 0 60384 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_630
timestamp 1679581782
transform 1 0 61056 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_637
timestamp 1679581782
transform 1 0 61728 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_644
timestamp 1679581782
transform 1 0 62400 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_651
timestamp 1679581782
transform 1 0 63072 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_658
timestamp 1679581782
transform 1 0 63744 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_665
timestamp 1679581782
transform 1 0 64416 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_672
timestamp 1679581782
transform 1 0 65088 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_679
timestamp 1679581782
transform 1 0 65760 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_686
timestamp 1679581782
transform 1 0 66432 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_693
timestamp 1679581782
transform 1 0 67104 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_700
timestamp 1679581782
transform 1 0 67776 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_707
timestamp 1679581782
transform 1 0 68448 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_714
timestamp 1679581782
transform 1 0 69120 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_721
timestamp 1679581782
transform 1 0 69792 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_728
timestamp 1679581782
transform 1 0 70464 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_735
timestamp 1679581782
transform 1 0 71136 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_742
timestamp 1679581782
transform 1 0 71808 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_749
timestamp 1679581782
transform 1 0 72480 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_756
timestamp 1679581782
transform 1 0 73152 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_763
timestamp 1679581782
transform 1 0 73824 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_770
timestamp 1679581782
transform 1 0 74496 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_777
timestamp 1679581782
transform 1 0 75168 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_784
timestamp 1679581782
transform 1 0 75840 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_791
timestamp 1679581782
transform 1 0 76512 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_798
timestamp 1679581782
transform 1 0 77184 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_805
timestamp 1679581782
transform 1 0 77856 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_812
timestamp 1679581782
transform 1 0 78528 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_819
timestamp 1679581782
transform 1 0 79200 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_826
timestamp 1679581782
transform 1 0 79872 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_833
timestamp 1679581782
transform 1 0 80544 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_840
timestamp 1679581782
transform 1 0 81216 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_847
timestamp 1679581782
transform 1 0 81888 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_854
timestamp 1679581782
transform 1 0 82560 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_861
timestamp 1679581782
transform 1 0 83232 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_868
timestamp 1679581782
transform 1 0 83904 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_875
timestamp 1679581782
transform 1 0 84576 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_882
timestamp 1679581782
transform 1 0 85248 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_889
timestamp 1679581782
transform 1 0 85920 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_896
timestamp 1679581782
transform 1 0 86592 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_903
timestamp 1679581782
transform 1 0 87264 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_910
timestamp 1679581782
transform 1 0 87936 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_917
timestamp 1679581782
transform 1 0 88608 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_924
timestamp 1679581782
transform 1 0 89280 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_931
timestamp 1679581782
transform 1 0 89952 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_938
timestamp 1679581782
transform 1 0 90624 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_945
timestamp 1679581782
transform 1 0 91296 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_952
timestamp 1679581782
transform 1 0 91968 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_959
timestamp 1679581782
transform 1 0 92640 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_966
timestamp 1679581782
transform 1 0 93312 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_973
timestamp 1679581782
transform 1 0 93984 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_980
timestamp 1679581782
transform 1 0 94656 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_987
timestamp 1679581782
transform 1 0 95328 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_994
timestamp 1679581782
transform 1 0 96000 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_1001
timestamp 1679581782
transform 1 0 96672 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_1008
timestamp 1679581782
transform 1 0 97344 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_1015
timestamp 1679581782
transform 1 0 98016 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_1022
timestamp 1679581782
transform 1 0 98688 0 1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_0
timestamp 1679581782
transform 1 0 576 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_7
timestamp 1679581782
transform 1 0 1248 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_14
timestamp 1679581782
transform 1 0 1920 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_21
timestamp 1679581782
transform 1 0 2592 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_28
timestamp 1679581782
transform 1 0 3264 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_35
timestamp 1679581782
transform 1 0 3936 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_42
timestamp 1679581782
transform 1 0 4608 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_49
timestamp 1679581782
transform 1 0 5280 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_56
timestamp 1679581782
transform 1 0 5952 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_63
timestamp 1679581782
transform 1 0 6624 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_70
timestamp 1679581782
transform 1 0 7296 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_77
timestamp 1679581782
transform 1 0 7968 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_84
timestamp 1679581782
transform 1 0 8640 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_91
timestamp 1679581782
transform 1 0 9312 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_98
timestamp 1679581782
transform 1 0 9984 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_105
timestamp 1679581782
transform 1 0 10656 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_112
timestamp 1679581782
transform 1 0 11328 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_119
timestamp 1679581782
transform 1 0 12000 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_126
timestamp 1679581782
transform 1 0 12672 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_133
timestamp 1679581782
transform 1 0 13344 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_140
timestamp 1679581782
transform 1 0 14016 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_147
timestamp 1679581782
transform 1 0 14688 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_154
timestamp 1679581782
transform 1 0 15360 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_161
timestamp 1679581782
transform 1 0 16032 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_168
timestamp 1679581782
transform 1 0 16704 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_175
timestamp 1679581782
transform 1 0 17376 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_182
timestamp 1679581782
transform 1 0 18048 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_189
timestamp 1679581782
transform 1 0 18720 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_196
timestamp 1679581782
transform 1 0 19392 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_203
timestamp 1679581782
transform 1 0 20064 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_210
timestamp 1679581782
transform 1 0 20736 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_217
timestamp 1679581782
transform 1 0 21408 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_224
timestamp 1679581782
transform 1 0 22080 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_231
timestamp 1679581782
transform 1 0 22752 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_238
timestamp 1679581782
transform 1 0 23424 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_245
timestamp 1679581782
transform 1 0 24096 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_252
timestamp 1679581782
transform 1 0 24768 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_259
timestamp 1679581782
transform 1 0 25440 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_266
timestamp 1679581782
transform 1 0 26112 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_273
timestamp 1679581782
transform 1 0 26784 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_280
timestamp 1679581782
transform 1 0 27456 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_287
timestamp 1679581782
transform 1 0 28128 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_294
timestamp 1679581782
transform 1 0 28800 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_301
timestamp 1679581782
transform 1 0 29472 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_308
timestamp 1679581782
transform 1 0 30144 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_315
timestamp 1679581782
transform 1 0 30816 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_322
timestamp 1679581782
transform 1 0 31488 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_329
timestamp 1679581782
transform 1 0 32160 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_336
timestamp 1679581782
transform 1 0 32832 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_343
timestamp 1679581782
transform 1 0 33504 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_350
timestamp 1679581782
transform 1 0 34176 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_357
timestamp 1679581782
transform 1 0 34848 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_364
timestamp 1679581782
transform 1 0 35520 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_371
timestamp 1679581782
transform 1 0 36192 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_378
timestamp 1679581782
transform 1 0 36864 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_385
timestamp 1679581782
transform 1 0 37536 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_392
timestamp 1679581782
transform 1 0 38208 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_399
timestamp 1679581782
transform 1 0 38880 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_406
timestamp 1679581782
transform 1 0 39552 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_413
timestamp 1679581782
transform 1 0 40224 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_420
timestamp 1679581782
transform 1 0 40896 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_427
timestamp 1679581782
transform 1 0 41568 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_434
timestamp 1679581782
transform 1 0 42240 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_441
timestamp 1679581782
transform 1 0 42912 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_448
timestamp 1679581782
transform 1 0 43584 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_455
timestamp 1679581782
transform 1 0 44256 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_462
timestamp 1679581782
transform 1 0 44928 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_469
timestamp 1679581782
transform 1 0 45600 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_476
timestamp 1679581782
transform 1 0 46272 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_483
timestamp 1679581782
transform 1 0 46944 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_490
timestamp 1679581782
transform 1 0 47616 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_497
timestamp 1679581782
transform 1 0 48288 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_504
timestamp 1679581782
transform 1 0 48960 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_511
timestamp 1679581782
transform 1 0 49632 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_518
timestamp 1679581782
transform 1 0 50304 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_525
timestamp 1679581782
transform 1 0 50976 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_532
timestamp 1679581782
transform 1 0 51648 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_539
timestamp 1679581782
transform 1 0 52320 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_546
timestamp 1679581782
transform 1 0 52992 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_553
timestamp 1679581782
transform 1 0 53664 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_560
timestamp 1679581782
transform 1 0 54336 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_567
timestamp 1679581782
transform 1 0 55008 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_574
timestamp 1679581782
transform 1 0 55680 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_581
timestamp 1679581782
transform 1 0 56352 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_588
timestamp 1679581782
transform 1 0 57024 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_595
timestamp 1679581782
transform 1 0 57696 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_602
timestamp 1679581782
transform 1 0 58368 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_609
timestamp 1679581782
transform 1 0 59040 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_616
timestamp 1679581782
transform 1 0 59712 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_623
timestamp 1679581782
transform 1 0 60384 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_630
timestamp 1679581782
transform 1 0 61056 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_637
timestamp 1679581782
transform 1 0 61728 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_644
timestamp 1679581782
transform 1 0 62400 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_651
timestamp 1679581782
transform 1 0 63072 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_658
timestamp 1679581782
transform 1 0 63744 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_665
timestamp 1679581782
transform 1 0 64416 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_672
timestamp 1679581782
transform 1 0 65088 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_679
timestamp 1679581782
transform 1 0 65760 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_686
timestamp 1679581782
transform 1 0 66432 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_693
timestamp 1679581782
transform 1 0 67104 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_700
timestamp 1679581782
transform 1 0 67776 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_707
timestamp 1679581782
transform 1 0 68448 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_714
timestamp 1679581782
transform 1 0 69120 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_721
timestamp 1679581782
transform 1 0 69792 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_728
timestamp 1679581782
transform 1 0 70464 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_735
timestamp 1679581782
transform 1 0 71136 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_742
timestamp 1679581782
transform 1 0 71808 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_749
timestamp 1679581782
transform 1 0 72480 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_756
timestamp 1679581782
transform 1 0 73152 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_763
timestamp 1679581782
transform 1 0 73824 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_770
timestamp 1679581782
transform 1 0 74496 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_777
timestamp 1679581782
transform 1 0 75168 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_784
timestamp 1679581782
transform 1 0 75840 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_791
timestamp 1679581782
transform 1 0 76512 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_798
timestamp 1679581782
transform 1 0 77184 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_805
timestamp 1679581782
transform 1 0 77856 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_812
timestamp 1679581782
transform 1 0 78528 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_819
timestamp 1679581782
transform 1 0 79200 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_826
timestamp 1679581782
transform 1 0 79872 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_833
timestamp 1679581782
transform 1 0 80544 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_840
timestamp 1679581782
transform 1 0 81216 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_847
timestamp 1679581782
transform 1 0 81888 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_854
timestamp 1679581782
transform 1 0 82560 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_861
timestamp 1679581782
transform 1 0 83232 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_868
timestamp 1679581782
transform 1 0 83904 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_875
timestamp 1679581782
transform 1 0 84576 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_882
timestamp 1679581782
transform 1 0 85248 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_889
timestamp 1679581782
transform 1 0 85920 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_896
timestamp 1679581782
transform 1 0 86592 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_903
timestamp 1679581782
transform 1 0 87264 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_910
timestamp 1679581782
transform 1 0 87936 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_917
timestamp 1679581782
transform 1 0 88608 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_924
timestamp 1679581782
transform 1 0 89280 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_931
timestamp 1679581782
transform 1 0 89952 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_938
timestamp 1679581782
transform 1 0 90624 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_945
timestamp 1679581782
transform 1 0 91296 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_952
timestamp 1679581782
transform 1 0 91968 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_959
timestamp 1679581782
transform 1 0 92640 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_966
timestamp 1679581782
transform 1 0 93312 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_973
timestamp 1679581782
transform 1 0 93984 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_980
timestamp 1679581782
transform 1 0 94656 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_987
timestamp 1679581782
transform 1 0 95328 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_994
timestamp 1679581782
transform 1 0 96000 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_1001
timestamp 1679581782
transform 1 0 96672 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_1008
timestamp 1679581782
transform 1 0 97344 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_1015
timestamp 1679581782
transform 1 0 98016 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_1022
timestamp 1679581782
transform 1 0 98688 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_4
timestamp 1679581782
transform 1 0 960 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_11
timestamp 1679581782
transform 1 0 1632 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_18
timestamp 1679581782
transform 1 0 2304 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_25
timestamp 1679581782
transform 1 0 2976 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_32
timestamp 1679581782
transform 1 0 3648 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_39
timestamp 1679581782
transform 1 0 4320 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_46
timestamp 1679581782
transform 1 0 4992 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_53
timestamp 1679581782
transform 1 0 5664 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_60
timestamp 1679581782
transform 1 0 6336 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_67
timestamp 1679581782
transform 1 0 7008 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_74
timestamp 1679581782
transform 1 0 7680 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_81
timestamp 1679581782
transform 1 0 8352 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_88
timestamp 1679581782
transform 1 0 9024 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_95
timestamp 1679581782
transform 1 0 9696 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_102
timestamp 1679581782
transform 1 0 10368 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_109
timestamp 1679581782
transform 1 0 11040 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_116
timestamp 1679581782
transform 1 0 11712 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_123
timestamp 1679581782
transform 1 0 12384 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_130
timestamp 1679581782
transform 1 0 13056 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_137
timestamp 1679581782
transform 1 0 13728 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_144
timestamp 1679581782
transform 1 0 14400 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_151
timestamp 1679581782
transform 1 0 15072 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_158
timestamp 1679581782
transform 1 0 15744 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_165
timestamp 1679581782
transform 1 0 16416 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_172
timestamp 1679581782
transform 1 0 17088 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_179
timestamp 1679581782
transform 1 0 17760 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_186
timestamp 1679581782
transform 1 0 18432 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_193
timestamp 1679581782
transform 1 0 19104 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_200
timestamp 1679581782
transform 1 0 19776 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_207
timestamp 1679581782
transform 1 0 20448 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_214
timestamp 1679581782
transform 1 0 21120 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_221
timestamp 1679581782
transform 1 0 21792 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_228
timestamp 1679581782
transform 1 0 22464 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_235
timestamp 1679581782
transform 1 0 23136 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_242
timestamp 1679581782
transform 1 0 23808 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_249
timestamp 1679581782
transform 1 0 24480 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_256
timestamp 1679581782
transform 1 0 25152 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_263
timestamp 1679581782
transform 1 0 25824 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_270
timestamp 1679581782
transform 1 0 26496 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_277
timestamp 1679581782
transform 1 0 27168 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_284
timestamp 1679581782
transform 1 0 27840 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_291
timestamp 1679581782
transform 1 0 28512 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_298
timestamp 1679581782
transform 1 0 29184 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_305
timestamp 1679581782
transform 1 0 29856 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_312
timestamp 1679581782
transform 1 0 30528 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_319
timestamp 1679581782
transform 1 0 31200 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_326
timestamp 1679581782
transform 1 0 31872 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_333
timestamp 1679581782
transform 1 0 32544 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_340
timestamp 1679581782
transform 1 0 33216 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_347
timestamp 1679581782
transform 1 0 33888 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_354
timestamp 1679581782
transform 1 0 34560 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_361
timestamp 1679581782
transform 1 0 35232 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_368
timestamp 1679581782
transform 1 0 35904 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_375
timestamp 1679581782
transform 1 0 36576 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_382
timestamp 1679581782
transform 1 0 37248 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_389
timestamp 1679581782
transform 1 0 37920 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_396
timestamp 1679581782
transform 1 0 38592 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_403
timestamp 1679581782
transform 1 0 39264 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_410
timestamp 1679581782
transform 1 0 39936 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_417
timestamp 1679581782
transform 1 0 40608 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_424
timestamp 1679581782
transform 1 0 41280 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_431
timestamp 1679581782
transform 1 0 41952 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_438
timestamp 1679581782
transform 1 0 42624 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_445
timestamp 1679581782
transform 1 0 43296 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_452
timestamp 1679581782
transform 1 0 43968 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_459
timestamp 1679581782
transform 1 0 44640 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_466
timestamp 1679581782
transform 1 0 45312 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_473
timestamp 1679581782
transform 1 0 45984 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_480
timestamp 1679581782
transform 1 0 46656 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_487
timestamp 1679581782
transform 1 0 47328 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_494
timestamp 1679581782
transform 1 0 48000 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_501
timestamp 1679581782
transform 1 0 48672 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_508
timestamp 1679581782
transform 1 0 49344 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_515
timestamp 1679581782
transform 1 0 50016 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_522
timestamp 1679581782
transform 1 0 50688 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_529
timestamp 1679581782
transform 1 0 51360 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_536
timestamp 1679581782
transform 1 0 52032 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_543
timestamp 1679581782
transform 1 0 52704 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_550
timestamp 1679581782
transform 1 0 53376 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_557
timestamp 1679581782
transform 1 0 54048 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_564
timestamp 1679581782
transform 1 0 54720 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_571
timestamp 1679581782
transform 1 0 55392 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_578
timestamp 1679581782
transform 1 0 56064 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_585
timestamp 1679581782
transform 1 0 56736 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_592
timestamp 1679581782
transform 1 0 57408 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_599
timestamp 1679581782
transform 1 0 58080 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_606
timestamp 1679581782
transform 1 0 58752 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_613
timestamp 1679581782
transform 1 0 59424 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_620
timestamp 1679581782
transform 1 0 60096 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_627
timestamp 1679581782
transform 1 0 60768 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_634
timestamp 1679581782
transform 1 0 61440 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_641
timestamp 1679581782
transform 1 0 62112 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_648
timestamp 1679581782
transform 1 0 62784 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_655
timestamp 1679581782
transform 1 0 63456 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_662
timestamp 1679581782
transform 1 0 64128 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_669
timestamp 1679581782
transform 1 0 64800 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_676
timestamp 1679581782
transform 1 0 65472 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_683
timestamp 1679581782
transform 1 0 66144 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_690
timestamp 1679581782
transform 1 0 66816 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_697
timestamp 1679581782
transform 1 0 67488 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_704
timestamp 1679581782
transform 1 0 68160 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_711
timestamp 1679581782
transform 1 0 68832 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_718
timestamp 1679581782
transform 1 0 69504 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_725
timestamp 1679581782
transform 1 0 70176 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_732
timestamp 1679581782
transform 1 0 70848 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_739
timestamp 1679581782
transform 1 0 71520 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_746
timestamp 1679581782
transform 1 0 72192 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_753
timestamp 1679581782
transform 1 0 72864 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_760
timestamp 1679581782
transform 1 0 73536 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_767
timestamp 1679581782
transform 1 0 74208 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_774
timestamp 1679581782
transform 1 0 74880 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_781
timestamp 1679581782
transform 1 0 75552 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_788
timestamp 1679581782
transform 1 0 76224 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_795
timestamp 1679581782
transform 1 0 76896 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_802
timestamp 1679581782
transform 1 0 77568 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_809
timestamp 1679581782
transform 1 0 78240 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_816
timestamp 1679581782
transform 1 0 78912 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_823
timestamp 1679581782
transform 1 0 79584 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_830
timestamp 1679581782
transform 1 0 80256 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_837
timestamp 1679581782
transform 1 0 80928 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_844
timestamp 1679581782
transform 1 0 81600 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_851
timestamp 1679581782
transform 1 0 82272 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_858
timestamp 1679581782
transform 1 0 82944 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_865
timestamp 1679581782
transform 1 0 83616 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_872
timestamp 1679581782
transform 1 0 84288 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_879
timestamp 1679581782
transform 1 0 84960 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_886
timestamp 1679581782
transform 1 0 85632 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_893
timestamp 1679581782
transform 1 0 86304 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_900
timestamp 1679581782
transform 1 0 86976 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_907
timestamp 1679581782
transform 1 0 87648 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_914
timestamp 1679581782
transform 1 0 88320 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_921
timestamp 1679581782
transform 1 0 88992 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_928
timestamp 1679581782
transform 1 0 89664 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_935
timestamp 1679581782
transform 1 0 90336 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_942
timestamp 1679581782
transform 1 0 91008 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_949
timestamp 1679581782
transform 1 0 91680 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_956
timestamp 1679581782
transform 1 0 92352 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_963
timestamp 1679581782
transform 1 0 93024 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_970
timestamp 1679581782
transform 1 0 93696 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_977
timestamp 1679581782
transform 1 0 94368 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_984
timestamp 1679581782
transform 1 0 95040 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_991
timestamp 1679581782
transform 1 0 95712 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_998
timestamp 1679581782
transform 1 0 96384 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_1005
timestamp 1679581782
transform 1 0 97056 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_1012
timestamp 1679581782
transform 1 0 97728 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_1019
timestamp 1679581782
transform 1 0 98400 0 1 49140
box -48 -56 720 834
use sg13g2_fill_2  FILLER_64_1026
timestamp 1677580104
transform 1 0 99072 0 1 49140
box -48 -56 240 834
use sg13g2_fill_1  FILLER_64_1028
timestamp 1677579658
transform 1 0 99264 0 1 49140
box -48 -56 144 834
use sg13g2_decap_8  FILLER_65_0
timestamp 1679581782
transform 1 0 576 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_7
timestamp 1679581782
transform 1 0 1248 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_14
timestamp 1679581782
transform 1 0 1920 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_21
timestamp 1679581782
transform 1 0 2592 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_28
timestamp 1679581782
transform 1 0 3264 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_35
timestamp 1679581782
transform 1 0 3936 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_42
timestamp 1679581782
transform 1 0 4608 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_49
timestamp 1679581782
transform 1 0 5280 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_56
timestamp 1679581782
transform 1 0 5952 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_63
timestamp 1679581782
transform 1 0 6624 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_70
timestamp 1679581782
transform 1 0 7296 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_77
timestamp 1679581782
transform 1 0 7968 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_84
timestamp 1679581782
transform 1 0 8640 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_91
timestamp 1679581782
transform 1 0 9312 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_98
timestamp 1679581782
transform 1 0 9984 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_105
timestamp 1679581782
transform 1 0 10656 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_112
timestamp 1679581782
transform 1 0 11328 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_119
timestamp 1679581782
transform 1 0 12000 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_126
timestamp 1679581782
transform 1 0 12672 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_133
timestamp 1679581782
transform 1 0 13344 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_140
timestamp 1679581782
transform 1 0 14016 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_147
timestamp 1679581782
transform 1 0 14688 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_154
timestamp 1679581782
transform 1 0 15360 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_161
timestamp 1679581782
transform 1 0 16032 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_168
timestamp 1679581782
transform 1 0 16704 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_175
timestamp 1679581782
transform 1 0 17376 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_182
timestamp 1679581782
transform 1 0 18048 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_189
timestamp 1679581782
transform 1 0 18720 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_196
timestamp 1679581782
transform 1 0 19392 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_203
timestamp 1679581782
transform 1 0 20064 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_210
timestamp 1679581782
transform 1 0 20736 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_217
timestamp 1679581782
transform 1 0 21408 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_224
timestamp 1679581782
transform 1 0 22080 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_231
timestamp 1679581782
transform 1 0 22752 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_238
timestamp 1679581782
transform 1 0 23424 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_245
timestamp 1679581782
transform 1 0 24096 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_252
timestamp 1679581782
transform 1 0 24768 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_259
timestamp 1679581782
transform 1 0 25440 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_266
timestamp 1679581782
transform 1 0 26112 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_273
timestamp 1679581782
transform 1 0 26784 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_280
timestamp 1679581782
transform 1 0 27456 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_287
timestamp 1679581782
transform 1 0 28128 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_294
timestamp 1679581782
transform 1 0 28800 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_301
timestamp 1679581782
transform 1 0 29472 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_308
timestamp 1679581782
transform 1 0 30144 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_315
timestamp 1679581782
transform 1 0 30816 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_322
timestamp 1679581782
transform 1 0 31488 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_329
timestamp 1679581782
transform 1 0 32160 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_336
timestamp 1679581782
transform 1 0 32832 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_343
timestamp 1679581782
transform 1 0 33504 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_350
timestamp 1679581782
transform 1 0 34176 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_357
timestamp 1679581782
transform 1 0 34848 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_364
timestamp 1679581782
transform 1 0 35520 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_371
timestamp 1679581782
transform 1 0 36192 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_378
timestamp 1679581782
transform 1 0 36864 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_385
timestamp 1679581782
transform 1 0 37536 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_392
timestamp 1679581782
transform 1 0 38208 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_399
timestamp 1679581782
transform 1 0 38880 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_406
timestamp 1679581782
transform 1 0 39552 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_413
timestamp 1679581782
transform 1 0 40224 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_420
timestamp 1679581782
transform 1 0 40896 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_427
timestamp 1679581782
transform 1 0 41568 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_434
timestamp 1679581782
transform 1 0 42240 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_441
timestamp 1679581782
transform 1 0 42912 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_448
timestamp 1679581782
transform 1 0 43584 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_455
timestamp 1679581782
transform 1 0 44256 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_462
timestamp 1679581782
transform 1 0 44928 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_469
timestamp 1679581782
transform 1 0 45600 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_476
timestamp 1679581782
transform 1 0 46272 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_483
timestamp 1679581782
transform 1 0 46944 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_490
timestamp 1679581782
transform 1 0 47616 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_497
timestamp 1679581782
transform 1 0 48288 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_504
timestamp 1679581782
transform 1 0 48960 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_511
timestamp 1679581782
transform 1 0 49632 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_518
timestamp 1679581782
transform 1 0 50304 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_525
timestamp 1679581782
transform 1 0 50976 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_532
timestamp 1679581782
transform 1 0 51648 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_539
timestamp 1679581782
transform 1 0 52320 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_546
timestamp 1679581782
transform 1 0 52992 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_553
timestamp 1679581782
transform 1 0 53664 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_560
timestamp 1679581782
transform 1 0 54336 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_567
timestamp 1679581782
transform 1 0 55008 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_574
timestamp 1679581782
transform 1 0 55680 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_581
timestamp 1679581782
transform 1 0 56352 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_588
timestamp 1679581782
transform 1 0 57024 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_595
timestamp 1679581782
transform 1 0 57696 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_602
timestamp 1679581782
transform 1 0 58368 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_609
timestamp 1679581782
transform 1 0 59040 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_616
timestamp 1679581782
transform 1 0 59712 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_623
timestamp 1679581782
transform 1 0 60384 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_630
timestamp 1679581782
transform 1 0 61056 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_637
timestamp 1679581782
transform 1 0 61728 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_644
timestamp 1679581782
transform 1 0 62400 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_651
timestamp 1679581782
transform 1 0 63072 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_658
timestamp 1679581782
transform 1 0 63744 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_665
timestamp 1679581782
transform 1 0 64416 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_672
timestamp 1679581782
transform 1 0 65088 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_679
timestamp 1679581782
transform 1 0 65760 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_686
timestamp 1679581782
transform 1 0 66432 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_693
timestamp 1679581782
transform 1 0 67104 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_700
timestamp 1679581782
transform 1 0 67776 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_707
timestamp 1679581782
transform 1 0 68448 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_714
timestamp 1679581782
transform 1 0 69120 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_721
timestamp 1679581782
transform 1 0 69792 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_728
timestamp 1679581782
transform 1 0 70464 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_735
timestamp 1679581782
transform 1 0 71136 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_742
timestamp 1679581782
transform 1 0 71808 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_749
timestamp 1679581782
transform 1 0 72480 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_756
timestamp 1679581782
transform 1 0 73152 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_763
timestamp 1679581782
transform 1 0 73824 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_770
timestamp 1679581782
transform 1 0 74496 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_777
timestamp 1679581782
transform 1 0 75168 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_784
timestamp 1679581782
transform 1 0 75840 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_791
timestamp 1679581782
transform 1 0 76512 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_798
timestamp 1679581782
transform 1 0 77184 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_805
timestamp 1679581782
transform 1 0 77856 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_812
timestamp 1679581782
transform 1 0 78528 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_819
timestamp 1679581782
transform 1 0 79200 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_826
timestamp 1679581782
transform 1 0 79872 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_833
timestamp 1679581782
transform 1 0 80544 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_840
timestamp 1679581782
transform 1 0 81216 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_847
timestamp 1679581782
transform 1 0 81888 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_854
timestamp 1679581782
transform 1 0 82560 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_861
timestamp 1679581782
transform 1 0 83232 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_868
timestamp 1679581782
transform 1 0 83904 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_875
timestamp 1679581782
transform 1 0 84576 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_882
timestamp 1679581782
transform 1 0 85248 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_889
timestamp 1679581782
transform 1 0 85920 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_896
timestamp 1679581782
transform 1 0 86592 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_903
timestamp 1679581782
transform 1 0 87264 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_910
timestamp 1679581782
transform 1 0 87936 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_917
timestamp 1679581782
transform 1 0 88608 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_924
timestamp 1679581782
transform 1 0 89280 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_931
timestamp 1679581782
transform 1 0 89952 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_938
timestamp 1679581782
transform 1 0 90624 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_945
timestamp 1679581782
transform 1 0 91296 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_952
timestamp 1679581782
transform 1 0 91968 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_959
timestamp 1679581782
transform 1 0 92640 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_966
timestamp 1679581782
transform 1 0 93312 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_973
timestamp 1679581782
transform 1 0 93984 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_980
timestamp 1679581782
transform 1 0 94656 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_987
timestamp 1679581782
transform 1 0 95328 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_994
timestamp 1679581782
transform 1 0 96000 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_1001
timestamp 1679581782
transform 1 0 96672 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_1008
timestamp 1679581782
transform 1 0 97344 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_1015
timestamp 1679581782
transform 1 0 98016 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_1022
timestamp 1679581782
transform 1 0 98688 0 -1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_4
timestamp 1679581782
transform 1 0 960 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_11
timestamp 1679581782
transform 1 0 1632 0 1 50652
box -48 -56 720 834
use sg13g2_fill_1  FILLER_66_18
timestamp 1677579658
transform 1 0 2304 0 1 50652
box -48 -56 144 834
use sg13g2_decap_8  FILLER_66_27
timestamp 1679581782
transform 1 0 3168 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_34
timestamp 1679581782
transform 1 0 3840 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_41
timestamp 1679581782
transform 1 0 4512 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_48
timestamp 1679581782
transform 1 0 5184 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_55
timestamp 1679581782
transform 1 0 5856 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_62
timestamp 1679581782
transform 1 0 6528 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_69
timestamp 1679581782
transform 1 0 7200 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_76
timestamp 1679581782
transform 1 0 7872 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_83
timestamp 1679581782
transform 1 0 8544 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_90
timestamp 1679581782
transform 1 0 9216 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_97
timestamp 1679581782
transform 1 0 9888 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_104
timestamp 1679581782
transform 1 0 10560 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_111
timestamp 1679581782
transform 1 0 11232 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_118
timestamp 1679581782
transform 1 0 11904 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_125
timestamp 1679581782
transform 1 0 12576 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_132
timestamp 1679581782
transform 1 0 13248 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_139
timestamp 1679581782
transform 1 0 13920 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_146
timestamp 1679581782
transform 1 0 14592 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_153
timestamp 1679581782
transform 1 0 15264 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_160
timestamp 1679581782
transform 1 0 15936 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_167
timestamp 1679581782
transform 1 0 16608 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_174
timestamp 1679581782
transform 1 0 17280 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_181
timestamp 1679581782
transform 1 0 17952 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_188
timestamp 1679581782
transform 1 0 18624 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_195
timestamp 1679581782
transform 1 0 19296 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_202
timestamp 1679581782
transform 1 0 19968 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_209
timestamp 1679581782
transform 1 0 20640 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_216
timestamp 1679581782
transform 1 0 21312 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_223
timestamp 1679581782
transform 1 0 21984 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_230
timestamp 1679581782
transform 1 0 22656 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_237
timestamp 1679581782
transform 1 0 23328 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_244
timestamp 1679581782
transform 1 0 24000 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_251
timestamp 1679581782
transform 1 0 24672 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_258
timestamp 1679581782
transform 1 0 25344 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_265
timestamp 1679581782
transform 1 0 26016 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_272
timestamp 1679581782
transform 1 0 26688 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_279
timestamp 1679581782
transform 1 0 27360 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_286
timestamp 1679581782
transform 1 0 28032 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_293
timestamp 1679581782
transform 1 0 28704 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_300
timestamp 1679581782
transform 1 0 29376 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_307
timestamp 1679581782
transform 1 0 30048 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_314
timestamp 1679581782
transform 1 0 30720 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_321
timestamp 1679581782
transform 1 0 31392 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_328
timestamp 1679581782
transform 1 0 32064 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_335
timestamp 1679581782
transform 1 0 32736 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_342
timestamp 1679581782
transform 1 0 33408 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_349
timestamp 1679581782
transform 1 0 34080 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_356
timestamp 1679581782
transform 1 0 34752 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_363
timestamp 1679581782
transform 1 0 35424 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_370
timestamp 1679581782
transform 1 0 36096 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_377
timestamp 1679581782
transform 1 0 36768 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_384
timestamp 1679581782
transform 1 0 37440 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_391
timestamp 1679581782
transform 1 0 38112 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_398
timestamp 1679581782
transform 1 0 38784 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_405
timestamp 1679581782
transform 1 0 39456 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_412
timestamp 1679581782
transform 1 0 40128 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_419
timestamp 1679581782
transform 1 0 40800 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_426
timestamp 1679581782
transform 1 0 41472 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_433
timestamp 1679581782
transform 1 0 42144 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_440
timestamp 1679581782
transform 1 0 42816 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_447
timestamp 1679581782
transform 1 0 43488 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_454
timestamp 1679581782
transform 1 0 44160 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_461
timestamp 1679581782
transform 1 0 44832 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_468
timestamp 1679581782
transform 1 0 45504 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_475
timestamp 1679581782
transform 1 0 46176 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_482
timestamp 1679581782
transform 1 0 46848 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_489
timestamp 1679581782
transform 1 0 47520 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_496
timestamp 1679581782
transform 1 0 48192 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_503
timestamp 1679581782
transform 1 0 48864 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_510
timestamp 1679581782
transform 1 0 49536 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_517
timestamp 1679581782
transform 1 0 50208 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_524
timestamp 1679581782
transform 1 0 50880 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_531
timestamp 1679581782
transform 1 0 51552 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_538
timestamp 1679581782
transform 1 0 52224 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_545
timestamp 1679581782
transform 1 0 52896 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_552
timestamp 1679581782
transform 1 0 53568 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_559
timestamp 1679581782
transform 1 0 54240 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_566
timestamp 1679581782
transform 1 0 54912 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_573
timestamp 1679581782
transform 1 0 55584 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_580
timestamp 1679581782
transform 1 0 56256 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_587
timestamp 1679581782
transform 1 0 56928 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_594
timestamp 1679581782
transform 1 0 57600 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_601
timestamp 1679581782
transform 1 0 58272 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_608
timestamp 1679581782
transform 1 0 58944 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_615
timestamp 1679581782
transform 1 0 59616 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_622
timestamp 1679581782
transform 1 0 60288 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_629
timestamp 1679581782
transform 1 0 60960 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_636
timestamp 1679581782
transform 1 0 61632 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_643
timestamp 1679581782
transform 1 0 62304 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_650
timestamp 1679581782
transform 1 0 62976 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_657
timestamp 1679581782
transform 1 0 63648 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_664
timestamp 1679581782
transform 1 0 64320 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_671
timestamp 1679581782
transform 1 0 64992 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_678
timestamp 1679581782
transform 1 0 65664 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_685
timestamp 1679581782
transform 1 0 66336 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_692
timestamp 1679581782
transform 1 0 67008 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_699
timestamp 1679581782
transform 1 0 67680 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_706
timestamp 1679581782
transform 1 0 68352 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_713
timestamp 1679581782
transform 1 0 69024 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_720
timestamp 1679581782
transform 1 0 69696 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_727
timestamp 1679581782
transform 1 0 70368 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_734
timestamp 1679581782
transform 1 0 71040 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_741
timestamp 1679581782
transform 1 0 71712 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_748
timestamp 1679581782
transform 1 0 72384 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_755
timestamp 1679581782
transform 1 0 73056 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_762
timestamp 1679581782
transform 1 0 73728 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_769
timestamp 1679581782
transform 1 0 74400 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_776
timestamp 1679581782
transform 1 0 75072 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_783
timestamp 1679581782
transform 1 0 75744 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_790
timestamp 1679581782
transform 1 0 76416 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_797
timestamp 1679581782
transform 1 0 77088 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_804
timestamp 1679581782
transform 1 0 77760 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_811
timestamp 1679581782
transform 1 0 78432 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_818
timestamp 1679581782
transform 1 0 79104 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_825
timestamp 1679581782
transform 1 0 79776 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_832
timestamp 1679581782
transform 1 0 80448 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_839
timestamp 1679581782
transform 1 0 81120 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_846
timestamp 1679581782
transform 1 0 81792 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_853
timestamp 1679581782
transform 1 0 82464 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_860
timestamp 1679581782
transform 1 0 83136 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_867
timestamp 1679581782
transform 1 0 83808 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_874
timestamp 1679581782
transform 1 0 84480 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_881
timestamp 1679581782
transform 1 0 85152 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_888
timestamp 1679581782
transform 1 0 85824 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_895
timestamp 1679581782
transform 1 0 86496 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_902
timestamp 1679581782
transform 1 0 87168 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_909
timestamp 1679581782
transform 1 0 87840 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_916
timestamp 1679581782
transform 1 0 88512 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_923
timestamp 1679581782
transform 1 0 89184 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_930
timestamp 1679581782
transform 1 0 89856 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_937
timestamp 1679581782
transform 1 0 90528 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_944
timestamp 1679581782
transform 1 0 91200 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_951
timestamp 1679581782
transform 1 0 91872 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_958
timestamp 1679581782
transform 1 0 92544 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_965
timestamp 1679581782
transform 1 0 93216 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_972
timestamp 1679581782
transform 1 0 93888 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_979
timestamp 1679581782
transform 1 0 94560 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_986
timestamp 1679581782
transform 1 0 95232 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_993
timestamp 1679581782
transform 1 0 95904 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_1000
timestamp 1679581782
transform 1 0 96576 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_1007
timestamp 1679581782
transform 1 0 97248 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_1014
timestamp 1679581782
transform 1 0 97920 0 1 50652
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_1021
timestamp 1679581782
transform 1 0 98592 0 1 50652
box -48 -56 720 834
use sg13g2_fill_1  FILLER_66_1028
timestamp 1677579658
transform 1 0 99264 0 1 50652
box -48 -56 144 834
use sg13g2_decap_8  FILLER_67_0
timestamp 1679581782
transform 1 0 576 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_7
timestamp 1679581782
transform 1 0 1248 0 -1 52164
box -48 -56 720 834
use sg13g2_fill_1  FILLER_67_14
timestamp 1677579658
transform 1 0 1920 0 -1 52164
box -48 -56 144 834
use sg13g2_fill_2  FILLER_67_31
timestamp 1677580104
transform 1 0 3552 0 -1 52164
box -48 -56 240 834
use sg13g2_fill_1  FILLER_67_33
timestamp 1677579658
transform 1 0 3744 0 -1 52164
box -48 -56 144 834
use sg13g2_decap_8  FILLER_67_38
timestamp 1679581782
transform 1 0 4224 0 -1 52164
box -48 -56 720 834
use sg13g2_fill_2  FILLER_67_45
timestamp 1677580104
transform 1 0 4896 0 -1 52164
box -48 -56 240 834
use sg13g2_fill_1  FILLER_67_47
timestamp 1677579658
transform 1 0 5088 0 -1 52164
box -48 -56 144 834
use sg13g2_fill_2  FILLER_67_55
timestamp 1677580104
transform 1 0 5856 0 -1 52164
box -48 -56 240 834
use sg13g2_fill_1  FILLER_67_57
timestamp 1677579658
transform 1 0 6048 0 -1 52164
box -48 -56 144 834
use sg13g2_decap_8  FILLER_67_70
timestamp 1679581782
transform 1 0 7296 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_77
timestamp 1679581782
transform 1 0 7968 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_84
timestamp 1679581782
transform 1 0 8640 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_91
timestamp 1679581782
transform 1 0 9312 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_98
timestamp 1679581782
transform 1 0 9984 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_105
timestamp 1679581782
transform 1 0 10656 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_112
timestamp 1679581782
transform 1 0 11328 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_119
timestamp 1679581782
transform 1 0 12000 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_126
timestamp 1679581782
transform 1 0 12672 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_133
timestamp 1679581782
transform 1 0 13344 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_140
timestamp 1679581782
transform 1 0 14016 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_147
timestamp 1679581782
transform 1 0 14688 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_154
timestamp 1679581782
transform 1 0 15360 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_161
timestamp 1679581782
transform 1 0 16032 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_168
timestamp 1679581782
transform 1 0 16704 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_175
timestamp 1679581782
transform 1 0 17376 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_182
timestamp 1679581782
transform 1 0 18048 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_189
timestamp 1679581782
transform 1 0 18720 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_196
timestamp 1679581782
transform 1 0 19392 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_203
timestamp 1679581782
transform 1 0 20064 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_210
timestamp 1679581782
transform 1 0 20736 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_217
timestamp 1679581782
transform 1 0 21408 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_224
timestamp 1679581782
transform 1 0 22080 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_231
timestamp 1679581782
transform 1 0 22752 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_238
timestamp 1679581782
transform 1 0 23424 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_245
timestamp 1679581782
transform 1 0 24096 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_252
timestamp 1679581782
transform 1 0 24768 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_259
timestamp 1679581782
transform 1 0 25440 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_266
timestamp 1679581782
transform 1 0 26112 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_273
timestamp 1679581782
transform 1 0 26784 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_280
timestamp 1679581782
transform 1 0 27456 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_287
timestamp 1679581782
transform 1 0 28128 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_294
timestamp 1679581782
transform 1 0 28800 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_301
timestamp 1679581782
transform 1 0 29472 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_308
timestamp 1679581782
transform 1 0 30144 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_315
timestamp 1679581782
transform 1 0 30816 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_322
timestamp 1679581782
transform 1 0 31488 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_329
timestamp 1679581782
transform 1 0 32160 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_336
timestamp 1679581782
transform 1 0 32832 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_343
timestamp 1679581782
transform 1 0 33504 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_350
timestamp 1679581782
transform 1 0 34176 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_357
timestamp 1679581782
transform 1 0 34848 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_364
timestamp 1679581782
transform 1 0 35520 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_371
timestamp 1679581782
transform 1 0 36192 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_378
timestamp 1679581782
transform 1 0 36864 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_385
timestamp 1679581782
transform 1 0 37536 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_392
timestamp 1679581782
transform 1 0 38208 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_399
timestamp 1679581782
transform 1 0 38880 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_406
timestamp 1679581782
transform 1 0 39552 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_413
timestamp 1679581782
transform 1 0 40224 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_420
timestamp 1679581782
transform 1 0 40896 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_427
timestamp 1679581782
transform 1 0 41568 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_434
timestamp 1679581782
transform 1 0 42240 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_441
timestamp 1679581782
transform 1 0 42912 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_448
timestamp 1679581782
transform 1 0 43584 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_455
timestamp 1679581782
transform 1 0 44256 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_462
timestamp 1679581782
transform 1 0 44928 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_469
timestamp 1679581782
transform 1 0 45600 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_476
timestamp 1679581782
transform 1 0 46272 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_483
timestamp 1679581782
transform 1 0 46944 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_490
timestamp 1679581782
transform 1 0 47616 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_497
timestamp 1679581782
transform 1 0 48288 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_504
timestamp 1679581782
transform 1 0 48960 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_511
timestamp 1679581782
transform 1 0 49632 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_518
timestamp 1679581782
transform 1 0 50304 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_525
timestamp 1679581782
transform 1 0 50976 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_532
timestamp 1679581782
transform 1 0 51648 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_539
timestamp 1679581782
transform 1 0 52320 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_546
timestamp 1679581782
transform 1 0 52992 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_553
timestamp 1679581782
transform 1 0 53664 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_560
timestamp 1679581782
transform 1 0 54336 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_567
timestamp 1679581782
transform 1 0 55008 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_574
timestamp 1679581782
transform 1 0 55680 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_581
timestamp 1679581782
transform 1 0 56352 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_588
timestamp 1679581782
transform 1 0 57024 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_595
timestamp 1679581782
transform 1 0 57696 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_602
timestamp 1679581782
transform 1 0 58368 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_609
timestamp 1679581782
transform 1 0 59040 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_616
timestamp 1679581782
transform 1 0 59712 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_623
timestamp 1679581782
transform 1 0 60384 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_630
timestamp 1679581782
transform 1 0 61056 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_637
timestamp 1679581782
transform 1 0 61728 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_644
timestamp 1679581782
transform 1 0 62400 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_651
timestamp 1679581782
transform 1 0 63072 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_658
timestamp 1679581782
transform 1 0 63744 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_665
timestamp 1679581782
transform 1 0 64416 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_672
timestamp 1679581782
transform 1 0 65088 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_679
timestamp 1679581782
transform 1 0 65760 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_686
timestamp 1679581782
transform 1 0 66432 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_693
timestamp 1679581782
transform 1 0 67104 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_700
timestamp 1679581782
transform 1 0 67776 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_707
timestamp 1679581782
transform 1 0 68448 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_714
timestamp 1679581782
transform 1 0 69120 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_721
timestamp 1679581782
transform 1 0 69792 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_728
timestamp 1679581782
transform 1 0 70464 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_735
timestamp 1679581782
transform 1 0 71136 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_742
timestamp 1679581782
transform 1 0 71808 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_749
timestamp 1679581782
transform 1 0 72480 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_756
timestamp 1679581782
transform 1 0 73152 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_763
timestamp 1679581782
transform 1 0 73824 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_770
timestamp 1679581782
transform 1 0 74496 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_777
timestamp 1679581782
transform 1 0 75168 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_784
timestamp 1679581782
transform 1 0 75840 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_791
timestamp 1679581782
transform 1 0 76512 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_798
timestamp 1679581782
transform 1 0 77184 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_805
timestamp 1679581782
transform 1 0 77856 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_812
timestamp 1679581782
transform 1 0 78528 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_819
timestamp 1679581782
transform 1 0 79200 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_826
timestamp 1679581782
transform 1 0 79872 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_833
timestamp 1679581782
transform 1 0 80544 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_840
timestamp 1679581782
transform 1 0 81216 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_847
timestamp 1679581782
transform 1 0 81888 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_854
timestamp 1679581782
transform 1 0 82560 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_861
timestamp 1679581782
transform 1 0 83232 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_868
timestamp 1679581782
transform 1 0 83904 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_875
timestamp 1679581782
transform 1 0 84576 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_882
timestamp 1679581782
transform 1 0 85248 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_889
timestamp 1679581782
transform 1 0 85920 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_896
timestamp 1679581782
transform 1 0 86592 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_903
timestamp 1679581782
transform 1 0 87264 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_910
timestamp 1679581782
transform 1 0 87936 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_917
timestamp 1679581782
transform 1 0 88608 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_924
timestamp 1679581782
transform 1 0 89280 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_931
timestamp 1679581782
transform 1 0 89952 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_938
timestamp 1679581782
transform 1 0 90624 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_945
timestamp 1679581782
transform 1 0 91296 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_952
timestamp 1679581782
transform 1 0 91968 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_959
timestamp 1679581782
transform 1 0 92640 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_966
timestamp 1679581782
transform 1 0 93312 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_973
timestamp 1679581782
transform 1 0 93984 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_980
timestamp 1679581782
transform 1 0 94656 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_987
timestamp 1679581782
transform 1 0 95328 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_994
timestamp 1679581782
transform 1 0 96000 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_1001
timestamp 1679581782
transform 1 0 96672 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_1008
timestamp 1679581782
transform 1 0 97344 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_1015
timestamp 1679581782
transform 1 0 98016 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_1022
timestamp 1679581782
transform 1 0 98688 0 -1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_4
timestamp 1679581782
transform 1 0 960 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_11
timestamp 1679581782
transform 1 0 1632 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_18
timestamp 1679581782
transform 1 0 2304 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_25
timestamp 1679581782
transform 1 0 2976 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_32
timestamp 1679581782
transform 1 0 3648 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_39
timestamp 1679581782
transform 1 0 4320 0 1 52164
box -48 -56 720 834
use sg13g2_decap_4  FILLER_68_46
timestamp 1679577901
transform 1 0 4992 0 1 52164
box -48 -56 432 834
use sg13g2_fill_2  FILLER_68_50
timestamp 1677580104
transform 1 0 5376 0 1 52164
box -48 -56 240 834
use sg13g2_decap_8  FILLER_68_68
timestamp 1679581782
transform 1 0 7104 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_75
timestamp 1679581782
transform 1 0 7776 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_82
timestamp 1679581782
transform 1 0 8448 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_89
timestamp 1679581782
transform 1 0 9120 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_96
timestamp 1679581782
transform 1 0 9792 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_103
timestamp 1679581782
transform 1 0 10464 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_110
timestamp 1679581782
transform 1 0 11136 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_117
timestamp 1679581782
transform 1 0 11808 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_124
timestamp 1679581782
transform 1 0 12480 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_131
timestamp 1679581782
transform 1 0 13152 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_138
timestamp 1679581782
transform 1 0 13824 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_145
timestamp 1679581782
transform 1 0 14496 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_152
timestamp 1679581782
transform 1 0 15168 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_159
timestamp 1679581782
transform 1 0 15840 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_166
timestamp 1679581782
transform 1 0 16512 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_173
timestamp 1679581782
transform 1 0 17184 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_180
timestamp 1679581782
transform 1 0 17856 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_187
timestamp 1679581782
transform 1 0 18528 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_194
timestamp 1679581782
transform 1 0 19200 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_201
timestamp 1679581782
transform 1 0 19872 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_208
timestamp 1679581782
transform 1 0 20544 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_215
timestamp 1679581782
transform 1 0 21216 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_222
timestamp 1679581782
transform 1 0 21888 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_229
timestamp 1679581782
transform 1 0 22560 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_236
timestamp 1679581782
transform 1 0 23232 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_243
timestamp 1679581782
transform 1 0 23904 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_250
timestamp 1679581782
transform 1 0 24576 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_257
timestamp 1679581782
transform 1 0 25248 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_264
timestamp 1679581782
transform 1 0 25920 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_271
timestamp 1679581782
transform 1 0 26592 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_278
timestamp 1679581782
transform 1 0 27264 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_285
timestamp 1679581782
transform 1 0 27936 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_292
timestamp 1679581782
transform 1 0 28608 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_299
timestamp 1679581782
transform 1 0 29280 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_306
timestamp 1679581782
transform 1 0 29952 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_313
timestamp 1679581782
transform 1 0 30624 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_320
timestamp 1679581782
transform 1 0 31296 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_327
timestamp 1679581782
transform 1 0 31968 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_334
timestamp 1679581782
transform 1 0 32640 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_341
timestamp 1679581782
transform 1 0 33312 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_348
timestamp 1679581782
transform 1 0 33984 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_355
timestamp 1679581782
transform 1 0 34656 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_362
timestamp 1679581782
transform 1 0 35328 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_369
timestamp 1679581782
transform 1 0 36000 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_376
timestamp 1679581782
transform 1 0 36672 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_383
timestamp 1679581782
transform 1 0 37344 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_390
timestamp 1679581782
transform 1 0 38016 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_397
timestamp 1679581782
transform 1 0 38688 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_404
timestamp 1679581782
transform 1 0 39360 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_411
timestamp 1679581782
transform 1 0 40032 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_418
timestamp 1679581782
transform 1 0 40704 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_425
timestamp 1679581782
transform 1 0 41376 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_432
timestamp 1679581782
transform 1 0 42048 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_439
timestamp 1679581782
transform 1 0 42720 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_446
timestamp 1679581782
transform 1 0 43392 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_453
timestamp 1679581782
transform 1 0 44064 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_460
timestamp 1679581782
transform 1 0 44736 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_467
timestamp 1679581782
transform 1 0 45408 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_474
timestamp 1679581782
transform 1 0 46080 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_481
timestamp 1679581782
transform 1 0 46752 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_488
timestamp 1679581782
transform 1 0 47424 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_495
timestamp 1679581782
transform 1 0 48096 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_502
timestamp 1679581782
transform 1 0 48768 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_509
timestamp 1679581782
transform 1 0 49440 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_516
timestamp 1679581782
transform 1 0 50112 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_523
timestamp 1679581782
transform 1 0 50784 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_530
timestamp 1679581782
transform 1 0 51456 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_537
timestamp 1679581782
transform 1 0 52128 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_544
timestamp 1679581782
transform 1 0 52800 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_551
timestamp 1679581782
transform 1 0 53472 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_558
timestamp 1679581782
transform 1 0 54144 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_565
timestamp 1679581782
transform 1 0 54816 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_572
timestamp 1679581782
transform 1 0 55488 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_579
timestamp 1679581782
transform 1 0 56160 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_586
timestamp 1679581782
transform 1 0 56832 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_593
timestamp 1679581782
transform 1 0 57504 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_600
timestamp 1679581782
transform 1 0 58176 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_607
timestamp 1679581782
transform 1 0 58848 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_614
timestamp 1679581782
transform 1 0 59520 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_621
timestamp 1679581782
transform 1 0 60192 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_628
timestamp 1679581782
transform 1 0 60864 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_635
timestamp 1679581782
transform 1 0 61536 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_642
timestamp 1679581782
transform 1 0 62208 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_649
timestamp 1679581782
transform 1 0 62880 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_656
timestamp 1679581782
transform 1 0 63552 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_663
timestamp 1679581782
transform 1 0 64224 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_670
timestamp 1679581782
transform 1 0 64896 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_677
timestamp 1679581782
transform 1 0 65568 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_684
timestamp 1679581782
transform 1 0 66240 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_691
timestamp 1679581782
transform 1 0 66912 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_698
timestamp 1679581782
transform 1 0 67584 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_705
timestamp 1679581782
transform 1 0 68256 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_712
timestamp 1679581782
transform 1 0 68928 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_719
timestamp 1679581782
transform 1 0 69600 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_726
timestamp 1679581782
transform 1 0 70272 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_733
timestamp 1679581782
transform 1 0 70944 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_740
timestamp 1679581782
transform 1 0 71616 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_747
timestamp 1679581782
transform 1 0 72288 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_754
timestamp 1679581782
transform 1 0 72960 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_761
timestamp 1679581782
transform 1 0 73632 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_768
timestamp 1679581782
transform 1 0 74304 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_775
timestamp 1679581782
transform 1 0 74976 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_782
timestamp 1679581782
transform 1 0 75648 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_789
timestamp 1679581782
transform 1 0 76320 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_796
timestamp 1679581782
transform 1 0 76992 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_803
timestamp 1679581782
transform 1 0 77664 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_810
timestamp 1679581782
transform 1 0 78336 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_817
timestamp 1679581782
transform 1 0 79008 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_824
timestamp 1679581782
transform 1 0 79680 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_831
timestamp 1679581782
transform 1 0 80352 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_838
timestamp 1679581782
transform 1 0 81024 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_845
timestamp 1679581782
transform 1 0 81696 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_852
timestamp 1679581782
transform 1 0 82368 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_859
timestamp 1679581782
transform 1 0 83040 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_866
timestamp 1679581782
transform 1 0 83712 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_873
timestamp 1679581782
transform 1 0 84384 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_880
timestamp 1679581782
transform 1 0 85056 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_887
timestamp 1679581782
transform 1 0 85728 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_894
timestamp 1679581782
transform 1 0 86400 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_901
timestamp 1679581782
transform 1 0 87072 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_908
timestamp 1679581782
transform 1 0 87744 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_915
timestamp 1679581782
transform 1 0 88416 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_922
timestamp 1679581782
transform 1 0 89088 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_929
timestamp 1679581782
transform 1 0 89760 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_936
timestamp 1679581782
transform 1 0 90432 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_943
timestamp 1679581782
transform 1 0 91104 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_950
timestamp 1679581782
transform 1 0 91776 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_957
timestamp 1679581782
transform 1 0 92448 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_964
timestamp 1679581782
transform 1 0 93120 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_971
timestamp 1679581782
transform 1 0 93792 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_978
timestamp 1679581782
transform 1 0 94464 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_985
timestamp 1679581782
transform 1 0 95136 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_992
timestamp 1679581782
transform 1 0 95808 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_999
timestamp 1679581782
transform 1 0 96480 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_1006
timestamp 1679581782
transform 1 0 97152 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_1013
timestamp 1679581782
transform 1 0 97824 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_1020
timestamp 1679581782
transform 1 0 98496 0 1 52164
box -48 -56 720 834
use sg13g2_fill_2  FILLER_68_1027
timestamp 1677580104
transform 1 0 99168 0 1 52164
box -48 -56 240 834
use sg13g2_decap_8  FILLER_69_0
timestamp 1679581782
transform 1 0 576 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_7
timestamp 1679581782
transform 1 0 1248 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_14
timestamp 1679581782
transform 1 0 1920 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_21
timestamp 1679581782
transform 1 0 2592 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_28
timestamp 1679581782
transform 1 0 3264 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_35
timestamp 1679581782
transform 1 0 3936 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_42
timestamp 1679581782
transform 1 0 4608 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_49
timestamp 1679581782
transform 1 0 5280 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_4  FILLER_69_56
timestamp 1679577901
transform 1 0 5952 0 -1 53676
box -48 -56 432 834
use sg13g2_decap_8  FILLER_69_64
timestamp 1679581782
transform 1 0 6720 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_71
timestamp 1679581782
transform 1 0 7392 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_78
timestamp 1679581782
transform 1 0 8064 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_85
timestamp 1679581782
transform 1 0 8736 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_92
timestamp 1679581782
transform 1 0 9408 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_99
timestamp 1679581782
transform 1 0 10080 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_106
timestamp 1679581782
transform 1 0 10752 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_113
timestamp 1679581782
transform 1 0 11424 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_120
timestamp 1679581782
transform 1 0 12096 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_127
timestamp 1679581782
transform 1 0 12768 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_134
timestamp 1679581782
transform 1 0 13440 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_141
timestamp 1679581782
transform 1 0 14112 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_148
timestamp 1679581782
transform 1 0 14784 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_155
timestamp 1679581782
transform 1 0 15456 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_162
timestamp 1679581782
transform 1 0 16128 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_169
timestamp 1679581782
transform 1 0 16800 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_176
timestamp 1679581782
transform 1 0 17472 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_183
timestamp 1679581782
transform 1 0 18144 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_190
timestamp 1679581782
transform 1 0 18816 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_197
timestamp 1679581782
transform 1 0 19488 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_204
timestamp 1679581782
transform 1 0 20160 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_211
timestamp 1679581782
transform 1 0 20832 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_218
timestamp 1679581782
transform 1 0 21504 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_225
timestamp 1679581782
transform 1 0 22176 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_232
timestamp 1679581782
transform 1 0 22848 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_239
timestamp 1679581782
transform 1 0 23520 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_246
timestamp 1679581782
transform 1 0 24192 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_253
timestamp 1679581782
transform 1 0 24864 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_260
timestamp 1679581782
transform 1 0 25536 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_267
timestamp 1679581782
transform 1 0 26208 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_274
timestamp 1679581782
transform 1 0 26880 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_281
timestamp 1679581782
transform 1 0 27552 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_288
timestamp 1679581782
transform 1 0 28224 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_295
timestamp 1679581782
transform 1 0 28896 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_302
timestamp 1679581782
transform 1 0 29568 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_309
timestamp 1679581782
transform 1 0 30240 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_316
timestamp 1679581782
transform 1 0 30912 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_323
timestamp 1679581782
transform 1 0 31584 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_330
timestamp 1679581782
transform 1 0 32256 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_337
timestamp 1679581782
transform 1 0 32928 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_344
timestamp 1679581782
transform 1 0 33600 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_351
timestamp 1679581782
transform 1 0 34272 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_358
timestamp 1679581782
transform 1 0 34944 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_365
timestamp 1679581782
transform 1 0 35616 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_372
timestamp 1679581782
transform 1 0 36288 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_379
timestamp 1679581782
transform 1 0 36960 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_386
timestamp 1679581782
transform 1 0 37632 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_393
timestamp 1679581782
transform 1 0 38304 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_400
timestamp 1679581782
transform 1 0 38976 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_407
timestamp 1679581782
transform 1 0 39648 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_414
timestamp 1679581782
transform 1 0 40320 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_421
timestamp 1679581782
transform 1 0 40992 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_428
timestamp 1679581782
transform 1 0 41664 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_435
timestamp 1679581782
transform 1 0 42336 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_442
timestamp 1679581782
transform 1 0 43008 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_449
timestamp 1679581782
transform 1 0 43680 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_456
timestamp 1679581782
transform 1 0 44352 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_463
timestamp 1679581782
transform 1 0 45024 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_470
timestamp 1679581782
transform 1 0 45696 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_477
timestamp 1679581782
transform 1 0 46368 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_484
timestamp 1679581782
transform 1 0 47040 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_491
timestamp 1679581782
transform 1 0 47712 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_498
timestamp 1679581782
transform 1 0 48384 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_505
timestamp 1679581782
transform 1 0 49056 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_512
timestamp 1679581782
transform 1 0 49728 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_519
timestamp 1679581782
transform 1 0 50400 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_526
timestamp 1679581782
transform 1 0 51072 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_533
timestamp 1679581782
transform 1 0 51744 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_540
timestamp 1679581782
transform 1 0 52416 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_547
timestamp 1679581782
transform 1 0 53088 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_554
timestamp 1679581782
transform 1 0 53760 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_561
timestamp 1679581782
transform 1 0 54432 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_568
timestamp 1679581782
transform 1 0 55104 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_575
timestamp 1679581782
transform 1 0 55776 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_582
timestamp 1679581782
transform 1 0 56448 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_589
timestamp 1679581782
transform 1 0 57120 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_596
timestamp 1679581782
transform 1 0 57792 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_603
timestamp 1679581782
transform 1 0 58464 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_610
timestamp 1679581782
transform 1 0 59136 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_617
timestamp 1679581782
transform 1 0 59808 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_624
timestamp 1679581782
transform 1 0 60480 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_631
timestamp 1679581782
transform 1 0 61152 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_638
timestamp 1679581782
transform 1 0 61824 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_645
timestamp 1679581782
transform 1 0 62496 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_652
timestamp 1679581782
transform 1 0 63168 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_659
timestamp 1679581782
transform 1 0 63840 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_666
timestamp 1679581782
transform 1 0 64512 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_673
timestamp 1679581782
transform 1 0 65184 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_680
timestamp 1679581782
transform 1 0 65856 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_687
timestamp 1679581782
transform 1 0 66528 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_694
timestamp 1679581782
transform 1 0 67200 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_701
timestamp 1679581782
transform 1 0 67872 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_708
timestamp 1679581782
transform 1 0 68544 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_715
timestamp 1679581782
transform 1 0 69216 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_722
timestamp 1679581782
transform 1 0 69888 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_729
timestamp 1679581782
transform 1 0 70560 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_736
timestamp 1679581782
transform 1 0 71232 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_743
timestamp 1679581782
transform 1 0 71904 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_750
timestamp 1679581782
transform 1 0 72576 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_757
timestamp 1679581782
transform 1 0 73248 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_764
timestamp 1679581782
transform 1 0 73920 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_771
timestamp 1679581782
transform 1 0 74592 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_778
timestamp 1679581782
transform 1 0 75264 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_785
timestamp 1679581782
transform 1 0 75936 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_792
timestamp 1679581782
transform 1 0 76608 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_799
timestamp 1679581782
transform 1 0 77280 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_806
timestamp 1679581782
transform 1 0 77952 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_813
timestamp 1679581782
transform 1 0 78624 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_820
timestamp 1679581782
transform 1 0 79296 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_827
timestamp 1679581782
transform 1 0 79968 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_834
timestamp 1679581782
transform 1 0 80640 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_841
timestamp 1679581782
transform 1 0 81312 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_848
timestamp 1679581782
transform 1 0 81984 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_855
timestamp 1679581782
transform 1 0 82656 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_862
timestamp 1679581782
transform 1 0 83328 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_869
timestamp 1679581782
transform 1 0 84000 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_876
timestamp 1679581782
transform 1 0 84672 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_883
timestamp 1679581782
transform 1 0 85344 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_890
timestamp 1679581782
transform 1 0 86016 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_897
timestamp 1679581782
transform 1 0 86688 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_904
timestamp 1679581782
transform 1 0 87360 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_911
timestamp 1679581782
transform 1 0 88032 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_918
timestamp 1679581782
transform 1 0 88704 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_925
timestamp 1679581782
transform 1 0 89376 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_932
timestamp 1679581782
transform 1 0 90048 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_939
timestamp 1679581782
transform 1 0 90720 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_946
timestamp 1679581782
transform 1 0 91392 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_953
timestamp 1679581782
transform 1 0 92064 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_960
timestamp 1679581782
transform 1 0 92736 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_967
timestamp 1679581782
transform 1 0 93408 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_974
timestamp 1679581782
transform 1 0 94080 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_981
timestamp 1679581782
transform 1 0 94752 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_988
timestamp 1679581782
transform 1 0 95424 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_995
timestamp 1679581782
transform 1 0 96096 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_1002
timestamp 1679581782
transform 1 0 96768 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_1009
timestamp 1679581782
transform 1 0 97440 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_1016
timestamp 1679581782
transform 1 0 98112 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_4  FILLER_69_1023
timestamp 1679577901
transform 1 0 98784 0 -1 53676
box -48 -56 432 834
use sg13g2_fill_2  FILLER_69_1027
timestamp 1677580104
transform 1 0 99168 0 -1 53676
box -48 -56 240 834
use sg13g2_decap_8  FILLER_70_0
timestamp 1679581782
transform 1 0 576 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_7
timestamp 1679581782
transform 1 0 1248 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_14
timestamp 1679581782
transform 1 0 1920 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_21
timestamp 1679581782
transform 1 0 2592 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_28
timestamp 1679581782
transform 1 0 3264 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_35
timestamp 1679581782
transform 1 0 3936 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_42
timestamp 1679581782
transform 1 0 4608 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_49
timestamp 1679581782
transform 1 0 5280 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_56
timestamp 1679581782
transform 1 0 5952 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_63
timestamp 1679581782
transform 1 0 6624 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_70
timestamp 1679581782
transform 1 0 7296 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_77
timestamp 1679581782
transform 1 0 7968 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_84
timestamp 1679581782
transform 1 0 8640 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_91
timestamp 1679581782
transform 1 0 9312 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_98
timestamp 1679581782
transform 1 0 9984 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_105
timestamp 1679581782
transform 1 0 10656 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_112
timestamp 1679581782
transform 1 0 11328 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_119
timestamp 1679581782
transform 1 0 12000 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_126
timestamp 1679581782
transform 1 0 12672 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_133
timestamp 1679581782
transform 1 0 13344 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_140
timestamp 1679581782
transform 1 0 14016 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_147
timestamp 1679581782
transform 1 0 14688 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_154
timestamp 1679581782
transform 1 0 15360 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_161
timestamp 1679581782
transform 1 0 16032 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_168
timestamp 1679581782
transform 1 0 16704 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_175
timestamp 1679581782
transform 1 0 17376 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_182
timestamp 1679581782
transform 1 0 18048 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_189
timestamp 1679581782
transform 1 0 18720 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_196
timestamp 1679581782
transform 1 0 19392 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_203
timestamp 1679581782
transform 1 0 20064 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_210
timestamp 1679581782
transform 1 0 20736 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_217
timestamp 1679581782
transform 1 0 21408 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_224
timestamp 1679581782
transform 1 0 22080 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_231
timestamp 1679581782
transform 1 0 22752 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_238
timestamp 1679581782
transform 1 0 23424 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_245
timestamp 1679581782
transform 1 0 24096 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_252
timestamp 1679581782
transform 1 0 24768 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_259
timestamp 1679581782
transform 1 0 25440 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_266
timestamp 1679581782
transform 1 0 26112 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_273
timestamp 1679581782
transform 1 0 26784 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_280
timestamp 1679581782
transform 1 0 27456 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_287
timestamp 1679581782
transform 1 0 28128 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_294
timestamp 1679581782
transform 1 0 28800 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_301
timestamp 1679581782
transform 1 0 29472 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_308
timestamp 1679581782
transform 1 0 30144 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_315
timestamp 1679581782
transform 1 0 30816 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_322
timestamp 1679581782
transform 1 0 31488 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_329
timestamp 1679581782
transform 1 0 32160 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_336
timestamp 1679581782
transform 1 0 32832 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_343
timestamp 1679581782
transform 1 0 33504 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_350
timestamp 1679581782
transform 1 0 34176 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_357
timestamp 1679581782
transform 1 0 34848 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_364
timestamp 1679581782
transform 1 0 35520 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_371
timestamp 1679581782
transform 1 0 36192 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_378
timestamp 1679581782
transform 1 0 36864 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_385
timestamp 1679581782
transform 1 0 37536 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_392
timestamp 1679581782
transform 1 0 38208 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_399
timestamp 1679581782
transform 1 0 38880 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_406
timestamp 1679581782
transform 1 0 39552 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_413
timestamp 1679581782
transform 1 0 40224 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_420
timestamp 1679581782
transform 1 0 40896 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_427
timestamp 1679581782
transform 1 0 41568 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_434
timestamp 1679581782
transform 1 0 42240 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_441
timestamp 1679581782
transform 1 0 42912 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_448
timestamp 1679581782
transform 1 0 43584 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_455
timestamp 1679581782
transform 1 0 44256 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_462
timestamp 1679581782
transform 1 0 44928 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_469
timestamp 1679581782
transform 1 0 45600 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_476
timestamp 1679581782
transform 1 0 46272 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_483
timestamp 1679581782
transform 1 0 46944 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_490
timestamp 1679581782
transform 1 0 47616 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_497
timestamp 1679581782
transform 1 0 48288 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_504
timestamp 1679581782
transform 1 0 48960 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_511
timestamp 1679581782
transform 1 0 49632 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_518
timestamp 1679581782
transform 1 0 50304 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_525
timestamp 1679581782
transform 1 0 50976 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_532
timestamp 1679581782
transform 1 0 51648 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_539
timestamp 1679581782
transform 1 0 52320 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_546
timestamp 1679581782
transform 1 0 52992 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_553
timestamp 1679581782
transform 1 0 53664 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_560
timestamp 1679581782
transform 1 0 54336 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_567
timestamp 1679581782
transform 1 0 55008 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_574
timestamp 1679581782
transform 1 0 55680 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_581
timestamp 1679581782
transform 1 0 56352 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_588
timestamp 1679581782
transform 1 0 57024 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_595
timestamp 1679581782
transform 1 0 57696 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_602
timestamp 1679581782
transform 1 0 58368 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_609
timestamp 1679581782
transform 1 0 59040 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_616
timestamp 1679581782
transform 1 0 59712 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_623
timestamp 1679581782
transform 1 0 60384 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_630
timestamp 1679581782
transform 1 0 61056 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_637
timestamp 1679581782
transform 1 0 61728 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_644
timestamp 1679581782
transform 1 0 62400 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_651
timestamp 1679581782
transform 1 0 63072 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_658
timestamp 1679581782
transform 1 0 63744 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_665
timestamp 1679581782
transform 1 0 64416 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_672
timestamp 1679581782
transform 1 0 65088 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_679
timestamp 1679581782
transform 1 0 65760 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_686
timestamp 1679581782
transform 1 0 66432 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_693
timestamp 1679581782
transform 1 0 67104 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_700
timestamp 1679581782
transform 1 0 67776 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_707
timestamp 1679581782
transform 1 0 68448 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_714
timestamp 1679581782
transform 1 0 69120 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_721
timestamp 1679581782
transform 1 0 69792 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_728
timestamp 1679581782
transform 1 0 70464 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_735
timestamp 1679581782
transform 1 0 71136 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_742
timestamp 1679581782
transform 1 0 71808 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_749
timestamp 1679581782
transform 1 0 72480 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_756
timestamp 1679581782
transform 1 0 73152 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_763
timestamp 1679581782
transform 1 0 73824 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_770
timestamp 1679581782
transform 1 0 74496 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_777
timestamp 1679581782
transform 1 0 75168 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_784
timestamp 1679581782
transform 1 0 75840 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_791
timestamp 1679581782
transform 1 0 76512 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_798
timestamp 1679581782
transform 1 0 77184 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_805
timestamp 1679581782
transform 1 0 77856 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_812
timestamp 1679581782
transform 1 0 78528 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_819
timestamp 1679581782
transform 1 0 79200 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_826
timestamp 1679581782
transform 1 0 79872 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_833
timestamp 1679581782
transform 1 0 80544 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_840
timestamp 1679581782
transform 1 0 81216 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_847
timestamp 1679581782
transform 1 0 81888 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_854
timestamp 1679581782
transform 1 0 82560 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_861
timestamp 1679581782
transform 1 0 83232 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_868
timestamp 1679581782
transform 1 0 83904 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_875
timestamp 1679581782
transform 1 0 84576 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_882
timestamp 1679581782
transform 1 0 85248 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_889
timestamp 1679581782
transform 1 0 85920 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_896
timestamp 1679581782
transform 1 0 86592 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_903
timestamp 1679581782
transform 1 0 87264 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_910
timestamp 1679581782
transform 1 0 87936 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_917
timestamp 1679581782
transform 1 0 88608 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_924
timestamp 1679581782
transform 1 0 89280 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_931
timestamp 1679581782
transform 1 0 89952 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_938
timestamp 1679581782
transform 1 0 90624 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_945
timestamp 1679581782
transform 1 0 91296 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_952
timestamp 1679581782
transform 1 0 91968 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_959
timestamp 1679581782
transform 1 0 92640 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_966
timestamp 1679581782
transform 1 0 93312 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_973
timestamp 1679581782
transform 1 0 93984 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_980
timestamp 1679581782
transform 1 0 94656 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_987
timestamp 1679581782
transform 1 0 95328 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_994
timestamp 1679581782
transform 1 0 96000 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_1001
timestamp 1679581782
transform 1 0 96672 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_1008
timestamp 1679581782
transform 1 0 97344 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_1015
timestamp 1679581782
transform 1 0 98016 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_1022
timestamp 1679581782
transform 1 0 98688 0 1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_4
timestamp 1679581782
transform 1 0 960 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_11
timestamp 1679581782
transform 1 0 1632 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_18
timestamp 1679581782
transform 1 0 2304 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_25
timestamp 1679581782
transform 1 0 2976 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_32
timestamp 1679581782
transform 1 0 3648 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_39
timestamp 1679581782
transform 1 0 4320 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_46
timestamp 1679581782
transform 1 0 4992 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_53
timestamp 1679581782
transform 1 0 5664 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_60
timestamp 1679581782
transform 1 0 6336 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_67
timestamp 1679581782
transform 1 0 7008 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_74
timestamp 1679581782
transform 1 0 7680 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_81
timestamp 1679581782
transform 1 0 8352 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_88
timestamp 1679581782
transform 1 0 9024 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_95
timestamp 1679581782
transform 1 0 9696 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_102
timestamp 1679581782
transform 1 0 10368 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_109
timestamp 1679581782
transform 1 0 11040 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_116
timestamp 1679581782
transform 1 0 11712 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_123
timestamp 1679581782
transform 1 0 12384 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_130
timestamp 1679581782
transform 1 0 13056 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_137
timestamp 1679581782
transform 1 0 13728 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_144
timestamp 1679581782
transform 1 0 14400 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_151
timestamp 1679581782
transform 1 0 15072 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_158
timestamp 1679581782
transform 1 0 15744 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_165
timestamp 1679581782
transform 1 0 16416 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_172
timestamp 1679581782
transform 1 0 17088 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_179
timestamp 1679581782
transform 1 0 17760 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_186
timestamp 1679581782
transform 1 0 18432 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_193
timestamp 1679581782
transform 1 0 19104 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_200
timestamp 1679581782
transform 1 0 19776 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_207
timestamp 1679581782
transform 1 0 20448 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_214
timestamp 1679581782
transform 1 0 21120 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_221
timestamp 1679581782
transform 1 0 21792 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_228
timestamp 1679581782
transform 1 0 22464 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_235
timestamp 1679581782
transform 1 0 23136 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_242
timestamp 1679581782
transform 1 0 23808 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_249
timestamp 1679581782
transform 1 0 24480 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_256
timestamp 1679581782
transform 1 0 25152 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_263
timestamp 1679581782
transform 1 0 25824 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_270
timestamp 1679581782
transform 1 0 26496 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_277
timestamp 1679581782
transform 1 0 27168 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_284
timestamp 1679581782
transform 1 0 27840 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_291
timestamp 1679581782
transform 1 0 28512 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_298
timestamp 1679581782
transform 1 0 29184 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_305
timestamp 1679581782
transform 1 0 29856 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_312
timestamp 1679581782
transform 1 0 30528 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_319
timestamp 1679581782
transform 1 0 31200 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_326
timestamp 1679581782
transform 1 0 31872 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_333
timestamp 1679581782
transform 1 0 32544 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_340
timestamp 1679581782
transform 1 0 33216 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_347
timestamp 1679581782
transform 1 0 33888 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_354
timestamp 1679581782
transform 1 0 34560 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_361
timestamp 1679581782
transform 1 0 35232 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_368
timestamp 1679581782
transform 1 0 35904 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_375
timestamp 1679581782
transform 1 0 36576 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_382
timestamp 1679581782
transform 1 0 37248 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_389
timestamp 1679581782
transform 1 0 37920 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_396
timestamp 1679581782
transform 1 0 38592 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_403
timestamp 1679581782
transform 1 0 39264 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_410
timestamp 1679581782
transform 1 0 39936 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_417
timestamp 1679581782
transform 1 0 40608 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_424
timestamp 1679581782
transform 1 0 41280 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_431
timestamp 1679581782
transform 1 0 41952 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_438
timestamp 1679581782
transform 1 0 42624 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_445
timestamp 1679581782
transform 1 0 43296 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_452
timestamp 1679581782
transform 1 0 43968 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_459
timestamp 1679581782
transform 1 0 44640 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_466
timestamp 1679581782
transform 1 0 45312 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_473
timestamp 1679581782
transform 1 0 45984 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_480
timestamp 1679581782
transform 1 0 46656 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_487
timestamp 1679581782
transform 1 0 47328 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_494
timestamp 1679581782
transform 1 0 48000 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_501
timestamp 1679581782
transform 1 0 48672 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_508
timestamp 1679581782
transform 1 0 49344 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_515
timestamp 1679581782
transform 1 0 50016 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_522
timestamp 1679581782
transform 1 0 50688 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_529
timestamp 1679581782
transform 1 0 51360 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_536
timestamp 1679581782
transform 1 0 52032 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_543
timestamp 1679581782
transform 1 0 52704 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_550
timestamp 1679581782
transform 1 0 53376 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_557
timestamp 1679581782
transform 1 0 54048 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_564
timestamp 1679581782
transform 1 0 54720 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_571
timestamp 1679581782
transform 1 0 55392 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_578
timestamp 1679581782
transform 1 0 56064 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_585
timestamp 1679581782
transform 1 0 56736 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_592
timestamp 1679581782
transform 1 0 57408 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_599
timestamp 1679581782
transform 1 0 58080 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_606
timestamp 1679581782
transform 1 0 58752 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_613
timestamp 1679581782
transform 1 0 59424 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_620
timestamp 1679581782
transform 1 0 60096 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_627
timestamp 1679581782
transform 1 0 60768 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_634
timestamp 1679581782
transform 1 0 61440 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_641
timestamp 1679581782
transform 1 0 62112 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_648
timestamp 1679581782
transform 1 0 62784 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_655
timestamp 1679581782
transform 1 0 63456 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_662
timestamp 1679581782
transform 1 0 64128 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_669
timestamp 1679581782
transform 1 0 64800 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_676
timestamp 1679581782
transform 1 0 65472 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_683
timestamp 1679581782
transform 1 0 66144 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_690
timestamp 1679581782
transform 1 0 66816 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_697
timestamp 1679581782
transform 1 0 67488 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_704
timestamp 1679581782
transform 1 0 68160 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_711
timestamp 1679581782
transform 1 0 68832 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_718
timestamp 1679581782
transform 1 0 69504 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_725
timestamp 1679581782
transform 1 0 70176 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_732
timestamp 1679581782
transform 1 0 70848 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_739
timestamp 1679581782
transform 1 0 71520 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_746
timestamp 1679581782
transform 1 0 72192 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_753
timestamp 1679581782
transform 1 0 72864 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_760
timestamp 1679581782
transform 1 0 73536 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_767
timestamp 1679581782
transform 1 0 74208 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_774
timestamp 1679581782
transform 1 0 74880 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_781
timestamp 1679581782
transform 1 0 75552 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_788
timestamp 1679581782
transform 1 0 76224 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_795
timestamp 1679581782
transform 1 0 76896 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_802
timestamp 1679581782
transform 1 0 77568 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_809
timestamp 1679581782
transform 1 0 78240 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_816
timestamp 1679581782
transform 1 0 78912 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_823
timestamp 1679581782
transform 1 0 79584 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_830
timestamp 1679581782
transform 1 0 80256 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_837
timestamp 1679581782
transform 1 0 80928 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_844
timestamp 1679581782
transform 1 0 81600 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_851
timestamp 1679581782
transform 1 0 82272 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_858
timestamp 1679581782
transform 1 0 82944 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_865
timestamp 1679581782
transform 1 0 83616 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_872
timestamp 1679581782
transform 1 0 84288 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_879
timestamp 1679581782
transform 1 0 84960 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_886
timestamp 1679581782
transform 1 0 85632 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_893
timestamp 1679581782
transform 1 0 86304 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_900
timestamp 1679581782
transform 1 0 86976 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_907
timestamp 1679581782
transform 1 0 87648 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_914
timestamp 1679581782
transform 1 0 88320 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_921
timestamp 1679581782
transform 1 0 88992 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_928
timestamp 1679581782
transform 1 0 89664 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_935
timestamp 1679581782
transform 1 0 90336 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_942
timestamp 1679581782
transform 1 0 91008 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_949
timestamp 1679581782
transform 1 0 91680 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_956
timestamp 1679581782
transform 1 0 92352 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_963
timestamp 1679581782
transform 1 0 93024 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_970
timestamp 1679581782
transform 1 0 93696 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_977
timestamp 1679581782
transform 1 0 94368 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_984
timestamp 1679581782
transform 1 0 95040 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_991
timestamp 1679581782
transform 1 0 95712 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_998
timestamp 1679581782
transform 1 0 96384 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_1005
timestamp 1679581782
transform 1 0 97056 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_1012
timestamp 1679581782
transform 1 0 97728 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_1019
timestamp 1679581782
transform 1 0 98400 0 -1 55188
box -48 -56 720 834
use sg13g2_fill_2  FILLER_71_1026
timestamp 1677580104
transform 1 0 99072 0 -1 55188
box -48 -56 240 834
use sg13g2_fill_1  FILLER_71_1028
timestamp 1677579658
transform 1 0 99264 0 -1 55188
box -48 -56 144 834
use sg13g2_decap_8  FILLER_72_0
timestamp 1679581782
transform 1 0 576 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_7
timestamp 1679581782
transform 1 0 1248 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_14
timestamp 1679581782
transform 1 0 1920 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_21
timestamp 1679581782
transform 1 0 2592 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_28
timestamp 1679581782
transform 1 0 3264 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_35
timestamp 1679581782
transform 1 0 3936 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_42
timestamp 1679581782
transform 1 0 4608 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_49
timestamp 1679581782
transform 1 0 5280 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_56
timestamp 1679581782
transform 1 0 5952 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_63
timestamp 1679581782
transform 1 0 6624 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_70
timestamp 1679581782
transform 1 0 7296 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_77
timestamp 1679581782
transform 1 0 7968 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_84
timestamp 1679581782
transform 1 0 8640 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_91
timestamp 1679581782
transform 1 0 9312 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_98
timestamp 1679581782
transform 1 0 9984 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_105
timestamp 1679581782
transform 1 0 10656 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_112
timestamp 1679581782
transform 1 0 11328 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_119
timestamp 1679581782
transform 1 0 12000 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_126
timestamp 1679581782
transform 1 0 12672 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_133
timestamp 1679581782
transform 1 0 13344 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_140
timestamp 1679581782
transform 1 0 14016 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_147
timestamp 1679581782
transform 1 0 14688 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_154
timestamp 1679581782
transform 1 0 15360 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_161
timestamp 1679581782
transform 1 0 16032 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_168
timestamp 1679581782
transform 1 0 16704 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_175
timestamp 1679581782
transform 1 0 17376 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_182
timestamp 1679581782
transform 1 0 18048 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_189
timestamp 1679581782
transform 1 0 18720 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_196
timestamp 1679581782
transform 1 0 19392 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_203
timestamp 1679581782
transform 1 0 20064 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_210
timestamp 1679581782
transform 1 0 20736 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_217
timestamp 1679581782
transform 1 0 21408 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_224
timestamp 1679581782
transform 1 0 22080 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_231
timestamp 1679581782
transform 1 0 22752 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_238
timestamp 1679581782
transform 1 0 23424 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_245
timestamp 1679581782
transform 1 0 24096 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_252
timestamp 1679581782
transform 1 0 24768 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_259
timestamp 1679581782
transform 1 0 25440 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_266
timestamp 1679581782
transform 1 0 26112 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_273
timestamp 1679581782
transform 1 0 26784 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_280
timestamp 1679581782
transform 1 0 27456 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_287
timestamp 1679581782
transform 1 0 28128 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_294
timestamp 1679581782
transform 1 0 28800 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_301
timestamp 1679581782
transform 1 0 29472 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_308
timestamp 1679581782
transform 1 0 30144 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_315
timestamp 1679581782
transform 1 0 30816 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_322
timestamp 1679581782
transform 1 0 31488 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_329
timestamp 1679581782
transform 1 0 32160 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_336
timestamp 1679581782
transform 1 0 32832 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_343
timestamp 1679581782
transform 1 0 33504 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_350
timestamp 1679581782
transform 1 0 34176 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_357
timestamp 1679581782
transform 1 0 34848 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_364
timestamp 1679581782
transform 1 0 35520 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_371
timestamp 1679581782
transform 1 0 36192 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_378
timestamp 1679581782
transform 1 0 36864 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_385
timestamp 1679581782
transform 1 0 37536 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_392
timestamp 1679581782
transform 1 0 38208 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_399
timestamp 1679581782
transform 1 0 38880 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_406
timestamp 1679581782
transform 1 0 39552 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_413
timestamp 1679581782
transform 1 0 40224 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_420
timestamp 1679581782
transform 1 0 40896 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_427
timestamp 1679581782
transform 1 0 41568 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_434
timestamp 1679581782
transform 1 0 42240 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_441
timestamp 1679581782
transform 1 0 42912 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_448
timestamp 1679581782
transform 1 0 43584 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_455
timestamp 1679581782
transform 1 0 44256 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_462
timestamp 1679581782
transform 1 0 44928 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_469
timestamp 1679581782
transform 1 0 45600 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_476
timestamp 1679581782
transform 1 0 46272 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_483
timestamp 1679581782
transform 1 0 46944 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_490
timestamp 1679581782
transform 1 0 47616 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_497
timestamp 1679581782
transform 1 0 48288 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_504
timestamp 1679581782
transform 1 0 48960 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_511
timestamp 1679581782
transform 1 0 49632 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_518
timestamp 1679581782
transform 1 0 50304 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_525
timestamp 1679581782
transform 1 0 50976 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_532
timestamp 1679581782
transform 1 0 51648 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_539
timestamp 1679581782
transform 1 0 52320 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_546
timestamp 1679581782
transform 1 0 52992 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_553
timestamp 1679581782
transform 1 0 53664 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_560
timestamp 1679581782
transform 1 0 54336 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_567
timestamp 1679581782
transform 1 0 55008 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_574
timestamp 1679581782
transform 1 0 55680 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_581
timestamp 1679581782
transform 1 0 56352 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_588
timestamp 1679581782
transform 1 0 57024 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_595
timestamp 1679581782
transform 1 0 57696 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_602
timestamp 1679581782
transform 1 0 58368 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_609
timestamp 1679581782
transform 1 0 59040 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_616
timestamp 1679581782
transform 1 0 59712 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_623
timestamp 1679581782
transform 1 0 60384 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_630
timestamp 1679581782
transform 1 0 61056 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_637
timestamp 1679581782
transform 1 0 61728 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_644
timestamp 1679581782
transform 1 0 62400 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_651
timestamp 1679581782
transform 1 0 63072 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_658
timestamp 1679581782
transform 1 0 63744 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_665
timestamp 1679581782
transform 1 0 64416 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_672
timestamp 1679581782
transform 1 0 65088 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_679
timestamp 1679581782
transform 1 0 65760 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_686
timestamp 1679581782
transform 1 0 66432 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_693
timestamp 1679581782
transform 1 0 67104 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_700
timestamp 1679581782
transform 1 0 67776 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_707
timestamp 1679581782
transform 1 0 68448 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_714
timestamp 1679581782
transform 1 0 69120 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_721
timestamp 1679581782
transform 1 0 69792 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_728
timestamp 1679581782
transform 1 0 70464 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_735
timestamp 1679581782
transform 1 0 71136 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_742
timestamp 1679581782
transform 1 0 71808 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_749
timestamp 1679581782
transform 1 0 72480 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_756
timestamp 1679581782
transform 1 0 73152 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_763
timestamp 1679581782
transform 1 0 73824 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_770
timestamp 1679581782
transform 1 0 74496 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_777
timestamp 1679581782
transform 1 0 75168 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_784
timestamp 1679581782
transform 1 0 75840 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_791
timestamp 1679581782
transform 1 0 76512 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_798
timestamp 1679581782
transform 1 0 77184 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_805
timestamp 1679581782
transform 1 0 77856 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_812
timestamp 1679581782
transform 1 0 78528 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_819
timestamp 1679581782
transform 1 0 79200 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_826
timestamp 1679581782
transform 1 0 79872 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_833
timestamp 1679581782
transform 1 0 80544 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_840
timestamp 1679581782
transform 1 0 81216 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_847
timestamp 1679581782
transform 1 0 81888 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_854
timestamp 1679581782
transform 1 0 82560 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_861
timestamp 1679581782
transform 1 0 83232 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_868
timestamp 1679581782
transform 1 0 83904 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_875
timestamp 1679581782
transform 1 0 84576 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_882
timestamp 1679581782
transform 1 0 85248 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_889
timestamp 1679581782
transform 1 0 85920 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_896
timestamp 1679581782
transform 1 0 86592 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_903
timestamp 1679581782
transform 1 0 87264 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_910
timestamp 1679581782
transform 1 0 87936 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_917
timestamp 1679581782
transform 1 0 88608 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_924
timestamp 1679581782
transform 1 0 89280 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_931
timestamp 1679581782
transform 1 0 89952 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_938
timestamp 1679581782
transform 1 0 90624 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_945
timestamp 1679581782
transform 1 0 91296 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_952
timestamp 1679581782
transform 1 0 91968 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_959
timestamp 1679581782
transform 1 0 92640 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_966
timestamp 1679581782
transform 1 0 93312 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_973
timestamp 1679581782
transform 1 0 93984 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_980
timestamp 1679581782
transform 1 0 94656 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_987
timestamp 1679581782
transform 1 0 95328 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_994
timestamp 1679581782
transform 1 0 96000 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_1001
timestamp 1679581782
transform 1 0 96672 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_1008
timestamp 1679581782
transform 1 0 97344 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_1015
timestamp 1679581782
transform 1 0 98016 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_1022
timestamp 1679581782
transform 1 0 98688 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_4
timestamp 1679581782
transform 1 0 960 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_11
timestamp 1679581782
transform 1 0 1632 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_18
timestamp 1679581782
transform 1 0 2304 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_25
timestamp 1679581782
transform 1 0 2976 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_32
timestamp 1679581782
transform 1 0 3648 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_39
timestamp 1679581782
transform 1 0 4320 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_46
timestamp 1679581782
transform 1 0 4992 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_4  FILLER_73_53
timestamp 1679577901
transform 1 0 5664 0 -1 56700
box -48 -56 432 834
use sg13g2_fill_2  FILLER_73_57
timestamp 1677580104
transform 1 0 6048 0 -1 56700
box -48 -56 240 834
use sg13g2_decap_8  FILLER_73_67
timestamp 1679581782
transform 1 0 7008 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_74
timestamp 1679581782
transform 1 0 7680 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_81
timestamp 1679581782
transform 1 0 8352 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_88
timestamp 1679581782
transform 1 0 9024 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_95
timestamp 1679581782
transform 1 0 9696 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_102
timestamp 1679581782
transform 1 0 10368 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_109
timestamp 1679581782
transform 1 0 11040 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_116
timestamp 1679581782
transform 1 0 11712 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_123
timestamp 1679581782
transform 1 0 12384 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_130
timestamp 1679581782
transform 1 0 13056 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_137
timestamp 1679581782
transform 1 0 13728 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_144
timestamp 1679581782
transform 1 0 14400 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_151
timestamp 1679581782
transform 1 0 15072 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_158
timestamp 1679581782
transform 1 0 15744 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_165
timestamp 1679581782
transform 1 0 16416 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_172
timestamp 1679581782
transform 1 0 17088 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_179
timestamp 1679581782
transform 1 0 17760 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_186
timestamp 1679581782
transform 1 0 18432 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_193
timestamp 1679581782
transform 1 0 19104 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_200
timestamp 1679581782
transform 1 0 19776 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_207
timestamp 1679581782
transform 1 0 20448 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_214
timestamp 1679581782
transform 1 0 21120 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_221
timestamp 1679581782
transform 1 0 21792 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_228
timestamp 1679581782
transform 1 0 22464 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_235
timestamp 1679581782
transform 1 0 23136 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_242
timestamp 1679581782
transform 1 0 23808 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_249
timestamp 1679581782
transform 1 0 24480 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_256
timestamp 1679581782
transform 1 0 25152 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_263
timestamp 1679581782
transform 1 0 25824 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_270
timestamp 1679581782
transform 1 0 26496 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_277
timestamp 1679581782
transform 1 0 27168 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_284
timestamp 1679581782
transform 1 0 27840 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_291
timestamp 1679581782
transform 1 0 28512 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_298
timestamp 1679581782
transform 1 0 29184 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_305
timestamp 1679581782
transform 1 0 29856 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_312
timestamp 1679581782
transform 1 0 30528 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_319
timestamp 1679581782
transform 1 0 31200 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_326
timestamp 1679581782
transform 1 0 31872 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_333
timestamp 1679581782
transform 1 0 32544 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_340
timestamp 1679581782
transform 1 0 33216 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_347
timestamp 1679581782
transform 1 0 33888 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_354
timestamp 1679581782
transform 1 0 34560 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_361
timestamp 1679581782
transform 1 0 35232 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_368
timestamp 1679581782
transform 1 0 35904 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_375
timestamp 1679581782
transform 1 0 36576 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_382
timestamp 1679581782
transform 1 0 37248 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_389
timestamp 1679581782
transform 1 0 37920 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_396
timestamp 1679581782
transform 1 0 38592 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_403
timestamp 1679581782
transform 1 0 39264 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_410
timestamp 1679581782
transform 1 0 39936 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_417
timestamp 1679581782
transform 1 0 40608 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_424
timestamp 1679581782
transform 1 0 41280 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_431
timestamp 1679581782
transform 1 0 41952 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_438
timestamp 1679581782
transform 1 0 42624 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_445
timestamp 1679581782
transform 1 0 43296 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_452
timestamp 1679581782
transform 1 0 43968 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_459
timestamp 1679581782
transform 1 0 44640 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_466
timestamp 1679581782
transform 1 0 45312 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_473
timestamp 1679581782
transform 1 0 45984 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_480
timestamp 1679581782
transform 1 0 46656 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_487
timestamp 1679581782
transform 1 0 47328 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_494
timestamp 1679581782
transform 1 0 48000 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_501
timestamp 1679581782
transform 1 0 48672 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_508
timestamp 1679581782
transform 1 0 49344 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_515
timestamp 1679581782
transform 1 0 50016 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_522
timestamp 1679581782
transform 1 0 50688 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_529
timestamp 1679581782
transform 1 0 51360 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_536
timestamp 1679581782
transform 1 0 52032 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_543
timestamp 1679581782
transform 1 0 52704 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_550
timestamp 1679581782
transform 1 0 53376 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_557
timestamp 1679581782
transform 1 0 54048 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_564
timestamp 1679581782
transform 1 0 54720 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_571
timestamp 1679581782
transform 1 0 55392 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_578
timestamp 1679581782
transform 1 0 56064 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_585
timestamp 1679581782
transform 1 0 56736 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_592
timestamp 1679581782
transform 1 0 57408 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_599
timestamp 1679581782
transform 1 0 58080 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_606
timestamp 1679581782
transform 1 0 58752 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_613
timestamp 1679581782
transform 1 0 59424 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_620
timestamp 1679581782
transform 1 0 60096 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_627
timestamp 1679581782
transform 1 0 60768 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_634
timestamp 1679581782
transform 1 0 61440 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_641
timestamp 1679581782
transform 1 0 62112 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_648
timestamp 1679581782
transform 1 0 62784 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_655
timestamp 1679581782
transform 1 0 63456 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_662
timestamp 1679581782
transform 1 0 64128 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_669
timestamp 1679581782
transform 1 0 64800 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_676
timestamp 1679581782
transform 1 0 65472 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_683
timestamp 1679581782
transform 1 0 66144 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_690
timestamp 1679581782
transform 1 0 66816 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_697
timestamp 1679581782
transform 1 0 67488 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_704
timestamp 1679581782
transform 1 0 68160 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_711
timestamp 1679581782
transform 1 0 68832 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_718
timestamp 1679581782
transform 1 0 69504 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_725
timestamp 1679581782
transform 1 0 70176 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_732
timestamp 1679581782
transform 1 0 70848 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_739
timestamp 1679581782
transform 1 0 71520 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_746
timestamp 1679581782
transform 1 0 72192 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_753
timestamp 1679581782
transform 1 0 72864 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_760
timestamp 1679581782
transform 1 0 73536 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_767
timestamp 1679581782
transform 1 0 74208 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_774
timestamp 1679581782
transform 1 0 74880 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_781
timestamp 1679581782
transform 1 0 75552 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_788
timestamp 1679581782
transform 1 0 76224 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_795
timestamp 1679581782
transform 1 0 76896 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_802
timestamp 1679581782
transform 1 0 77568 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_809
timestamp 1679581782
transform 1 0 78240 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_816
timestamp 1679581782
transform 1 0 78912 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_823
timestamp 1679581782
transform 1 0 79584 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_830
timestamp 1679581782
transform 1 0 80256 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_837
timestamp 1679581782
transform 1 0 80928 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_844
timestamp 1679581782
transform 1 0 81600 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_851
timestamp 1679581782
transform 1 0 82272 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_858
timestamp 1679581782
transform 1 0 82944 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_865
timestamp 1679581782
transform 1 0 83616 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_872
timestamp 1679581782
transform 1 0 84288 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_879
timestamp 1679581782
transform 1 0 84960 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_886
timestamp 1679581782
transform 1 0 85632 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_893
timestamp 1679581782
transform 1 0 86304 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_900
timestamp 1679581782
transform 1 0 86976 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_907
timestamp 1679581782
transform 1 0 87648 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_914
timestamp 1679581782
transform 1 0 88320 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_921
timestamp 1679581782
transform 1 0 88992 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_928
timestamp 1679581782
transform 1 0 89664 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_935
timestamp 1679581782
transform 1 0 90336 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_942
timestamp 1679581782
transform 1 0 91008 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_949
timestamp 1679581782
transform 1 0 91680 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_956
timestamp 1679581782
transform 1 0 92352 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_963
timestamp 1679581782
transform 1 0 93024 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_970
timestamp 1679581782
transform 1 0 93696 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_977
timestamp 1679581782
transform 1 0 94368 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_984
timestamp 1679581782
transform 1 0 95040 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_991
timestamp 1679581782
transform 1 0 95712 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_998
timestamp 1679581782
transform 1 0 96384 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_1005
timestamp 1679581782
transform 1 0 97056 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_1012
timestamp 1679581782
transform 1 0 97728 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_1019
timestamp 1679581782
transform 1 0 98400 0 -1 56700
box -48 -56 720 834
use sg13g2_fill_2  FILLER_73_1026
timestamp 1677580104
transform 1 0 99072 0 -1 56700
box -48 -56 240 834
use sg13g2_fill_1  FILLER_73_1028
timestamp 1677579658
transform 1 0 99264 0 -1 56700
box -48 -56 144 834
use sg13g2_decap_8  FILLER_74_0
timestamp 1679581782
transform 1 0 576 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_7
timestamp 1679581782
transform 1 0 1248 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_14
timestamp 1679581782
transform 1 0 1920 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_21
timestamp 1679581782
transform 1 0 2592 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_28
timestamp 1679581782
transform 1 0 3264 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_35
timestamp 1679581782
transform 1 0 3936 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_42
timestamp 1679581782
transform 1 0 4608 0 1 56700
box -48 -56 720 834
use sg13g2_decap_4  FILLER_74_49
timestamp 1679577901
transform 1 0 5280 0 1 56700
box -48 -56 432 834
use sg13g2_fill_1  FILLER_74_53
timestamp 1677579658
transform 1 0 5664 0 1 56700
box -48 -56 144 834
use sg13g2_decap_8  FILLER_74_71
timestamp 1679581782
transform 1 0 7392 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_78
timestamp 1679581782
transform 1 0 8064 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_85
timestamp 1679581782
transform 1 0 8736 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_92
timestamp 1679581782
transform 1 0 9408 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_99
timestamp 1679581782
transform 1 0 10080 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_106
timestamp 1679581782
transform 1 0 10752 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_113
timestamp 1679581782
transform 1 0 11424 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_120
timestamp 1679581782
transform 1 0 12096 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_127
timestamp 1679581782
transform 1 0 12768 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_134
timestamp 1679581782
transform 1 0 13440 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_141
timestamp 1679581782
transform 1 0 14112 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_148
timestamp 1679581782
transform 1 0 14784 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_155
timestamp 1679581782
transform 1 0 15456 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_162
timestamp 1679581782
transform 1 0 16128 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_169
timestamp 1679581782
transform 1 0 16800 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_176
timestamp 1679581782
transform 1 0 17472 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_183
timestamp 1679581782
transform 1 0 18144 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_190
timestamp 1679581782
transform 1 0 18816 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_197
timestamp 1679581782
transform 1 0 19488 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_204
timestamp 1679581782
transform 1 0 20160 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_211
timestamp 1679581782
transform 1 0 20832 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_218
timestamp 1679581782
transform 1 0 21504 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_225
timestamp 1679581782
transform 1 0 22176 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_232
timestamp 1679581782
transform 1 0 22848 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_239
timestamp 1679581782
transform 1 0 23520 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_246
timestamp 1679581782
transform 1 0 24192 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_253
timestamp 1679581782
transform 1 0 24864 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_260
timestamp 1679581782
transform 1 0 25536 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_267
timestamp 1679581782
transform 1 0 26208 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_274
timestamp 1679581782
transform 1 0 26880 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_281
timestamp 1679581782
transform 1 0 27552 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_288
timestamp 1679581782
transform 1 0 28224 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_295
timestamp 1679581782
transform 1 0 28896 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_302
timestamp 1679581782
transform 1 0 29568 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_309
timestamp 1679581782
transform 1 0 30240 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_316
timestamp 1679581782
transform 1 0 30912 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_323
timestamp 1679581782
transform 1 0 31584 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_330
timestamp 1679581782
transform 1 0 32256 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_337
timestamp 1679581782
transform 1 0 32928 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_344
timestamp 1679581782
transform 1 0 33600 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_351
timestamp 1679581782
transform 1 0 34272 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_358
timestamp 1679581782
transform 1 0 34944 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_365
timestamp 1679581782
transform 1 0 35616 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_372
timestamp 1679581782
transform 1 0 36288 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_379
timestamp 1679581782
transform 1 0 36960 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_386
timestamp 1679581782
transform 1 0 37632 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_393
timestamp 1679581782
transform 1 0 38304 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_400
timestamp 1679581782
transform 1 0 38976 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_407
timestamp 1679581782
transform 1 0 39648 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_414
timestamp 1679581782
transform 1 0 40320 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_421
timestamp 1679581782
transform 1 0 40992 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_428
timestamp 1679581782
transform 1 0 41664 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_435
timestamp 1679581782
transform 1 0 42336 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_442
timestamp 1679581782
transform 1 0 43008 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_449
timestamp 1679581782
transform 1 0 43680 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_456
timestamp 1679581782
transform 1 0 44352 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_463
timestamp 1679581782
transform 1 0 45024 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_470
timestamp 1679581782
transform 1 0 45696 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_477
timestamp 1679581782
transform 1 0 46368 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_484
timestamp 1679581782
transform 1 0 47040 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_491
timestamp 1679581782
transform 1 0 47712 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_498
timestamp 1679581782
transform 1 0 48384 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_505
timestamp 1679581782
transform 1 0 49056 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_512
timestamp 1679581782
transform 1 0 49728 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_519
timestamp 1679581782
transform 1 0 50400 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_526
timestamp 1679581782
transform 1 0 51072 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_533
timestamp 1679581782
transform 1 0 51744 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_540
timestamp 1679581782
transform 1 0 52416 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_547
timestamp 1679581782
transform 1 0 53088 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_554
timestamp 1679581782
transform 1 0 53760 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_561
timestamp 1679581782
transform 1 0 54432 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_568
timestamp 1679581782
transform 1 0 55104 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_575
timestamp 1679581782
transform 1 0 55776 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_582
timestamp 1679581782
transform 1 0 56448 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_589
timestamp 1679581782
transform 1 0 57120 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_596
timestamp 1679581782
transform 1 0 57792 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_603
timestamp 1679581782
transform 1 0 58464 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_610
timestamp 1679581782
transform 1 0 59136 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_617
timestamp 1679581782
transform 1 0 59808 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_624
timestamp 1679581782
transform 1 0 60480 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_631
timestamp 1679581782
transform 1 0 61152 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_638
timestamp 1679581782
transform 1 0 61824 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_645
timestamp 1679581782
transform 1 0 62496 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_652
timestamp 1679581782
transform 1 0 63168 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_659
timestamp 1679581782
transform 1 0 63840 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_666
timestamp 1679581782
transform 1 0 64512 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_673
timestamp 1679581782
transform 1 0 65184 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_680
timestamp 1679581782
transform 1 0 65856 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_687
timestamp 1679581782
transform 1 0 66528 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_694
timestamp 1679581782
transform 1 0 67200 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_701
timestamp 1679581782
transform 1 0 67872 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_708
timestamp 1679581782
transform 1 0 68544 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_715
timestamp 1679581782
transform 1 0 69216 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_722
timestamp 1679581782
transform 1 0 69888 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_729
timestamp 1679581782
transform 1 0 70560 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_736
timestamp 1679581782
transform 1 0 71232 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_743
timestamp 1679581782
transform 1 0 71904 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_750
timestamp 1679581782
transform 1 0 72576 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_757
timestamp 1679581782
transform 1 0 73248 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_764
timestamp 1679581782
transform 1 0 73920 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_771
timestamp 1679581782
transform 1 0 74592 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_778
timestamp 1679581782
transform 1 0 75264 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_785
timestamp 1679581782
transform 1 0 75936 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_792
timestamp 1679581782
transform 1 0 76608 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_799
timestamp 1679581782
transform 1 0 77280 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_806
timestamp 1679581782
transform 1 0 77952 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_813
timestamp 1679581782
transform 1 0 78624 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_820
timestamp 1679581782
transform 1 0 79296 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_827
timestamp 1679581782
transform 1 0 79968 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_834
timestamp 1679581782
transform 1 0 80640 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_841
timestamp 1679581782
transform 1 0 81312 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_848
timestamp 1679581782
transform 1 0 81984 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_855
timestamp 1679581782
transform 1 0 82656 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_862
timestamp 1679581782
transform 1 0 83328 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_869
timestamp 1679581782
transform 1 0 84000 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_876
timestamp 1679581782
transform 1 0 84672 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_883
timestamp 1679581782
transform 1 0 85344 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_890
timestamp 1679581782
transform 1 0 86016 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_897
timestamp 1679581782
transform 1 0 86688 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_904
timestamp 1679581782
transform 1 0 87360 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_911
timestamp 1679581782
transform 1 0 88032 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_918
timestamp 1679581782
transform 1 0 88704 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_925
timestamp 1679581782
transform 1 0 89376 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_932
timestamp 1679581782
transform 1 0 90048 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_939
timestamp 1679581782
transform 1 0 90720 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_946
timestamp 1679581782
transform 1 0 91392 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_953
timestamp 1679581782
transform 1 0 92064 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_960
timestamp 1679581782
transform 1 0 92736 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_967
timestamp 1679581782
transform 1 0 93408 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_974
timestamp 1679581782
transform 1 0 94080 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_981
timestamp 1679581782
transform 1 0 94752 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_988
timestamp 1679581782
transform 1 0 95424 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_995
timestamp 1679581782
transform 1 0 96096 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_1002
timestamp 1679581782
transform 1 0 96768 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_1009
timestamp 1679581782
transform 1 0 97440 0 1 56700
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_1016
timestamp 1679581782
transform 1 0 98112 0 1 56700
box -48 -56 720 834
use sg13g2_decap_4  FILLER_74_1023
timestamp 1679577901
transform 1 0 98784 0 1 56700
box -48 -56 432 834
use sg13g2_fill_2  FILLER_74_1027
timestamp 1677580104
transform 1 0 99168 0 1 56700
box -48 -56 240 834
use sg13g2_decap_8  FILLER_75_0
timestamp 1679581782
transform 1 0 576 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_7
timestamp 1679581782
transform 1 0 1248 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_14
timestamp 1679581782
transform 1 0 1920 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_21
timestamp 1679581782
transform 1 0 2592 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_28
timestamp 1679581782
transform 1 0 3264 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_35
timestamp 1679581782
transform 1 0 3936 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_42
timestamp 1679581782
transform 1 0 4608 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_49
timestamp 1679581782
transform 1 0 5280 0 -1 58212
box -48 -56 720 834
use sg13g2_fill_2  FILLER_75_56
timestamp 1677580104
transform 1 0 5952 0 -1 58212
box -48 -56 240 834
use sg13g2_fill_1  FILLER_75_58
timestamp 1677579658
transform 1 0 6144 0 -1 58212
box -48 -56 144 834
use sg13g2_decap_8  FILLER_75_63
timestamp 1679581782
transform 1 0 6624 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_70
timestamp 1679581782
transform 1 0 7296 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_77
timestamp 1679581782
transform 1 0 7968 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_84
timestamp 1679581782
transform 1 0 8640 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_91
timestamp 1679581782
transform 1 0 9312 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_98
timestamp 1679581782
transform 1 0 9984 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_105
timestamp 1679581782
transform 1 0 10656 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_112
timestamp 1679581782
transform 1 0 11328 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_119
timestamp 1679581782
transform 1 0 12000 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_126
timestamp 1679581782
transform 1 0 12672 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_133
timestamp 1679581782
transform 1 0 13344 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_140
timestamp 1679581782
transform 1 0 14016 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_147
timestamp 1679581782
transform 1 0 14688 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_154
timestamp 1679581782
transform 1 0 15360 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_161
timestamp 1679581782
transform 1 0 16032 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_168
timestamp 1679581782
transform 1 0 16704 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_175
timestamp 1679581782
transform 1 0 17376 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_182
timestamp 1679581782
transform 1 0 18048 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_189
timestamp 1679581782
transform 1 0 18720 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_196
timestamp 1679581782
transform 1 0 19392 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_203
timestamp 1679581782
transform 1 0 20064 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_210
timestamp 1679581782
transform 1 0 20736 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_217
timestamp 1679581782
transform 1 0 21408 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_224
timestamp 1679581782
transform 1 0 22080 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_231
timestamp 1679581782
transform 1 0 22752 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_238
timestamp 1679581782
transform 1 0 23424 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_245
timestamp 1679581782
transform 1 0 24096 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_252
timestamp 1679581782
transform 1 0 24768 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_259
timestamp 1679581782
transform 1 0 25440 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_266
timestamp 1679581782
transform 1 0 26112 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_273
timestamp 1679581782
transform 1 0 26784 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_280
timestamp 1679581782
transform 1 0 27456 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_287
timestamp 1679581782
transform 1 0 28128 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_294
timestamp 1679581782
transform 1 0 28800 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_301
timestamp 1679581782
transform 1 0 29472 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_308
timestamp 1679581782
transform 1 0 30144 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_315
timestamp 1679581782
transform 1 0 30816 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_322
timestamp 1679581782
transform 1 0 31488 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_329
timestamp 1679581782
transform 1 0 32160 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_336
timestamp 1679581782
transform 1 0 32832 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_343
timestamp 1679581782
transform 1 0 33504 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_350
timestamp 1679581782
transform 1 0 34176 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_357
timestamp 1679581782
transform 1 0 34848 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_364
timestamp 1679581782
transform 1 0 35520 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_371
timestamp 1679581782
transform 1 0 36192 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_378
timestamp 1679581782
transform 1 0 36864 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_385
timestamp 1679581782
transform 1 0 37536 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_392
timestamp 1679581782
transform 1 0 38208 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_399
timestamp 1679581782
transform 1 0 38880 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_406
timestamp 1679581782
transform 1 0 39552 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_413
timestamp 1679581782
transform 1 0 40224 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_420
timestamp 1679581782
transform 1 0 40896 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_427
timestamp 1679581782
transform 1 0 41568 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_434
timestamp 1679581782
transform 1 0 42240 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_441
timestamp 1679581782
transform 1 0 42912 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_448
timestamp 1679581782
transform 1 0 43584 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_455
timestamp 1679581782
transform 1 0 44256 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_462
timestamp 1679581782
transform 1 0 44928 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_469
timestamp 1679581782
transform 1 0 45600 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_476
timestamp 1679581782
transform 1 0 46272 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_483
timestamp 1679581782
transform 1 0 46944 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_490
timestamp 1679581782
transform 1 0 47616 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_497
timestamp 1679581782
transform 1 0 48288 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_504
timestamp 1679581782
transform 1 0 48960 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_511
timestamp 1679581782
transform 1 0 49632 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_518
timestamp 1679581782
transform 1 0 50304 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_525
timestamp 1679581782
transform 1 0 50976 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_532
timestamp 1679581782
transform 1 0 51648 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_539
timestamp 1679581782
transform 1 0 52320 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_546
timestamp 1679581782
transform 1 0 52992 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_553
timestamp 1679581782
transform 1 0 53664 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_560
timestamp 1679581782
transform 1 0 54336 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_567
timestamp 1679581782
transform 1 0 55008 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_574
timestamp 1679581782
transform 1 0 55680 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_581
timestamp 1679581782
transform 1 0 56352 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_588
timestamp 1679581782
transform 1 0 57024 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_595
timestamp 1679581782
transform 1 0 57696 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_602
timestamp 1679581782
transform 1 0 58368 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_609
timestamp 1679581782
transform 1 0 59040 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_616
timestamp 1679581782
transform 1 0 59712 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_623
timestamp 1679581782
transform 1 0 60384 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_630
timestamp 1679581782
transform 1 0 61056 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_637
timestamp 1679581782
transform 1 0 61728 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_644
timestamp 1679581782
transform 1 0 62400 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_651
timestamp 1679581782
transform 1 0 63072 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_658
timestamp 1679581782
transform 1 0 63744 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_665
timestamp 1679581782
transform 1 0 64416 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_672
timestamp 1679581782
transform 1 0 65088 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_679
timestamp 1679581782
transform 1 0 65760 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_686
timestamp 1679581782
transform 1 0 66432 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_693
timestamp 1679581782
transform 1 0 67104 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_700
timestamp 1679581782
transform 1 0 67776 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_707
timestamp 1679581782
transform 1 0 68448 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_714
timestamp 1679581782
transform 1 0 69120 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_721
timestamp 1679581782
transform 1 0 69792 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_728
timestamp 1679581782
transform 1 0 70464 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_735
timestamp 1679581782
transform 1 0 71136 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_742
timestamp 1679581782
transform 1 0 71808 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_749
timestamp 1679581782
transform 1 0 72480 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_756
timestamp 1679581782
transform 1 0 73152 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_763
timestamp 1679581782
transform 1 0 73824 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_770
timestamp 1679581782
transform 1 0 74496 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_777
timestamp 1679581782
transform 1 0 75168 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_784
timestamp 1679581782
transform 1 0 75840 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_791
timestamp 1679581782
transform 1 0 76512 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_798
timestamp 1679581782
transform 1 0 77184 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_805
timestamp 1679581782
transform 1 0 77856 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_812
timestamp 1679581782
transform 1 0 78528 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_819
timestamp 1679581782
transform 1 0 79200 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_826
timestamp 1679581782
transform 1 0 79872 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_833
timestamp 1679581782
transform 1 0 80544 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_840
timestamp 1679581782
transform 1 0 81216 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_847
timestamp 1679581782
transform 1 0 81888 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_854
timestamp 1679581782
transform 1 0 82560 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_861
timestamp 1679581782
transform 1 0 83232 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_868
timestamp 1679581782
transform 1 0 83904 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_875
timestamp 1679581782
transform 1 0 84576 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_882
timestamp 1679581782
transform 1 0 85248 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_889
timestamp 1679581782
transform 1 0 85920 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_896
timestamp 1679581782
transform 1 0 86592 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_903
timestamp 1679581782
transform 1 0 87264 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_910
timestamp 1679581782
transform 1 0 87936 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_917
timestamp 1679581782
transform 1 0 88608 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_924
timestamp 1679581782
transform 1 0 89280 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_931
timestamp 1679581782
transform 1 0 89952 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_938
timestamp 1679581782
transform 1 0 90624 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_945
timestamp 1679581782
transform 1 0 91296 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_952
timestamp 1679581782
transform 1 0 91968 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_959
timestamp 1679581782
transform 1 0 92640 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_966
timestamp 1679581782
transform 1 0 93312 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_973
timestamp 1679581782
transform 1 0 93984 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_980
timestamp 1679581782
transform 1 0 94656 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_987
timestamp 1679581782
transform 1 0 95328 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_994
timestamp 1679581782
transform 1 0 96000 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_1001
timestamp 1679581782
transform 1 0 96672 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_1008
timestamp 1679581782
transform 1 0 97344 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_1015
timestamp 1679581782
transform 1 0 98016 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_1022
timestamp 1679581782
transform 1 0 98688 0 -1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_4
timestamp 1679581782
transform 1 0 960 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_11
timestamp 1679581782
transform 1 0 1632 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_18
timestamp 1679581782
transform 1 0 2304 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_25
timestamp 1679581782
transform 1 0 2976 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_32
timestamp 1679581782
transform 1 0 3648 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_39
timestamp 1679581782
transform 1 0 4320 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_46
timestamp 1679581782
transform 1 0 4992 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_53
timestamp 1679581782
transform 1 0 5664 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_60
timestamp 1679581782
transform 1 0 6336 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_67
timestamp 1679581782
transform 1 0 7008 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_74
timestamp 1679581782
transform 1 0 7680 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_81
timestamp 1679581782
transform 1 0 8352 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_88
timestamp 1679581782
transform 1 0 9024 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_95
timestamp 1679581782
transform 1 0 9696 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_102
timestamp 1679581782
transform 1 0 10368 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_109
timestamp 1679581782
transform 1 0 11040 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_116
timestamp 1679581782
transform 1 0 11712 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_123
timestamp 1679581782
transform 1 0 12384 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_130
timestamp 1679581782
transform 1 0 13056 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_137
timestamp 1679581782
transform 1 0 13728 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_144
timestamp 1679581782
transform 1 0 14400 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_151
timestamp 1679581782
transform 1 0 15072 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_158
timestamp 1679581782
transform 1 0 15744 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_165
timestamp 1679581782
transform 1 0 16416 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_172
timestamp 1679581782
transform 1 0 17088 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_179
timestamp 1679581782
transform 1 0 17760 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_186
timestamp 1679581782
transform 1 0 18432 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_193
timestamp 1679581782
transform 1 0 19104 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_200
timestamp 1679581782
transform 1 0 19776 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_207
timestamp 1679581782
transform 1 0 20448 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_214
timestamp 1679581782
transform 1 0 21120 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_221
timestamp 1679581782
transform 1 0 21792 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_228
timestamp 1679581782
transform 1 0 22464 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_235
timestamp 1679581782
transform 1 0 23136 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_242
timestamp 1679581782
transform 1 0 23808 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_249
timestamp 1679581782
transform 1 0 24480 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_256
timestamp 1679581782
transform 1 0 25152 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_263
timestamp 1679581782
transform 1 0 25824 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_270
timestamp 1679581782
transform 1 0 26496 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_277
timestamp 1679581782
transform 1 0 27168 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_284
timestamp 1679581782
transform 1 0 27840 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_291
timestamp 1679581782
transform 1 0 28512 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_298
timestamp 1679581782
transform 1 0 29184 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_305
timestamp 1679581782
transform 1 0 29856 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_312
timestamp 1679581782
transform 1 0 30528 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_319
timestamp 1679581782
transform 1 0 31200 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_326
timestamp 1679581782
transform 1 0 31872 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_333
timestamp 1679581782
transform 1 0 32544 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_340
timestamp 1679581782
transform 1 0 33216 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_347
timestamp 1679581782
transform 1 0 33888 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_354
timestamp 1679581782
transform 1 0 34560 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_361
timestamp 1679581782
transform 1 0 35232 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_368
timestamp 1679581782
transform 1 0 35904 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_375
timestamp 1679581782
transform 1 0 36576 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_382
timestamp 1679581782
transform 1 0 37248 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_389
timestamp 1679581782
transform 1 0 37920 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_396
timestamp 1679581782
transform 1 0 38592 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_403
timestamp 1679581782
transform 1 0 39264 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_410
timestamp 1679581782
transform 1 0 39936 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_417
timestamp 1679581782
transform 1 0 40608 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_424
timestamp 1679581782
transform 1 0 41280 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_431
timestamp 1679581782
transform 1 0 41952 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_438
timestamp 1679581782
transform 1 0 42624 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_445
timestamp 1679581782
transform 1 0 43296 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_452
timestamp 1679581782
transform 1 0 43968 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_459
timestamp 1679581782
transform 1 0 44640 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_466
timestamp 1679581782
transform 1 0 45312 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_473
timestamp 1679581782
transform 1 0 45984 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_480
timestamp 1679581782
transform 1 0 46656 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_487
timestamp 1679581782
transform 1 0 47328 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_494
timestamp 1679581782
transform 1 0 48000 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_501
timestamp 1679581782
transform 1 0 48672 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_508
timestamp 1679581782
transform 1 0 49344 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_515
timestamp 1679581782
transform 1 0 50016 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_522
timestamp 1679581782
transform 1 0 50688 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_529
timestamp 1679581782
transform 1 0 51360 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_536
timestamp 1679581782
transform 1 0 52032 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_543
timestamp 1679581782
transform 1 0 52704 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_550
timestamp 1679581782
transform 1 0 53376 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_557
timestamp 1679581782
transform 1 0 54048 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_564
timestamp 1679581782
transform 1 0 54720 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_571
timestamp 1679581782
transform 1 0 55392 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_578
timestamp 1679581782
transform 1 0 56064 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_585
timestamp 1679581782
transform 1 0 56736 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_592
timestamp 1679581782
transform 1 0 57408 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_599
timestamp 1679581782
transform 1 0 58080 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_606
timestamp 1679581782
transform 1 0 58752 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_613
timestamp 1679581782
transform 1 0 59424 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_620
timestamp 1679581782
transform 1 0 60096 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_627
timestamp 1679581782
transform 1 0 60768 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_634
timestamp 1679581782
transform 1 0 61440 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_641
timestamp 1679581782
transform 1 0 62112 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_648
timestamp 1679581782
transform 1 0 62784 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_655
timestamp 1679581782
transform 1 0 63456 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_662
timestamp 1679581782
transform 1 0 64128 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_669
timestamp 1679581782
transform 1 0 64800 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_676
timestamp 1679581782
transform 1 0 65472 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_683
timestamp 1679581782
transform 1 0 66144 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_690
timestamp 1679581782
transform 1 0 66816 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_697
timestamp 1679581782
transform 1 0 67488 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_704
timestamp 1679581782
transform 1 0 68160 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_711
timestamp 1679581782
transform 1 0 68832 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_718
timestamp 1679581782
transform 1 0 69504 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_725
timestamp 1679581782
transform 1 0 70176 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_732
timestamp 1679581782
transform 1 0 70848 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_739
timestamp 1679581782
transform 1 0 71520 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_746
timestamp 1679581782
transform 1 0 72192 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_753
timestamp 1679581782
transform 1 0 72864 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_760
timestamp 1679581782
transform 1 0 73536 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_767
timestamp 1679581782
transform 1 0 74208 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_774
timestamp 1679581782
transform 1 0 74880 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_781
timestamp 1679581782
transform 1 0 75552 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_788
timestamp 1679581782
transform 1 0 76224 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_795
timestamp 1679581782
transform 1 0 76896 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_802
timestamp 1679581782
transform 1 0 77568 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_809
timestamp 1679581782
transform 1 0 78240 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_816
timestamp 1679581782
transform 1 0 78912 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_823
timestamp 1679581782
transform 1 0 79584 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_830
timestamp 1679581782
transform 1 0 80256 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_837
timestamp 1679581782
transform 1 0 80928 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_844
timestamp 1679581782
transform 1 0 81600 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_851
timestamp 1679581782
transform 1 0 82272 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_858
timestamp 1679581782
transform 1 0 82944 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_865
timestamp 1679581782
transform 1 0 83616 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_872
timestamp 1679581782
transform 1 0 84288 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_879
timestamp 1679581782
transform 1 0 84960 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_886
timestamp 1679581782
transform 1 0 85632 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_893
timestamp 1679581782
transform 1 0 86304 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_900
timestamp 1679581782
transform 1 0 86976 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_907
timestamp 1679581782
transform 1 0 87648 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_914
timestamp 1679581782
transform 1 0 88320 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_921
timestamp 1679581782
transform 1 0 88992 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_928
timestamp 1679581782
transform 1 0 89664 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_935
timestamp 1679581782
transform 1 0 90336 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_942
timestamp 1679581782
transform 1 0 91008 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_949
timestamp 1679581782
transform 1 0 91680 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_956
timestamp 1679581782
transform 1 0 92352 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_963
timestamp 1679581782
transform 1 0 93024 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_970
timestamp 1679581782
transform 1 0 93696 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_977
timestamp 1679581782
transform 1 0 94368 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_984
timestamp 1679581782
transform 1 0 95040 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_991
timestamp 1679581782
transform 1 0 95712 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_998
timestamp 1679581782
transform 1 0 96384 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_1005
timestamp 1679581782
transform 1 0 97056 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_1012
timestamp 1679581782
transform 1 0 97728 0 1 58212
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_1019
timestamp 1679581782
transform 1 0 98400 0 1 58212
box -48 -56 720 834
use sg13g2_fill_2  FILLER_76_1026
timestamp 1677580104
transform 1 0 99072 0 1 58212
box -48 -56 240 834
use sg13g2_fill_1  FILLER_76_1028
timestamp 1677579658
transform 1 0 99264 0 1 58212
box -48 -56 144 834
use sg13g2_decap_8  FILLER_77_0
timestamp 1679581782
transform 1 0 576 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_7
timestamp 1679581782
transform 1 0 1248 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_14
timestamp 1679581782
transform 1 0 1920 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_21
timestamp 1679581782
transform 1 0 2592 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_28
timestamp 1679581782
transform 1 0 3264 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_35
timestamp 1679581782
transform 1 0 3936 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_42
timestamp 1679581782
transform 1 0 4608 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_49
timestamp 1679581782
transform 1 0 5280 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_56
timestamp 1679581782
transform 1 0 5952 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_63
timestamp 1679581782
transform 1 0 6624 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_70
timestamp 1679581782
transform 1 0 7296 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_77
timestamp 1679581782
transform 1 0 7968 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_84
timestamp 1679581782
transform 1 0 8640 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_91
timestamp 1679581782
transform 1 0 9312 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_98
timestamp 1679581782
transform 1 0 9984 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_105
timestamp 1679581782
transform 1 0 10656 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_112
timestamp 1679581782
transform 1 0 11328 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_119
timestamp 1679581782
transform 1 0 12000 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_126
timestamp 1679581782
transform 1 0 12672 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_133
timestamp 1679581782
transform 1 0 13344 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_140
timestamp 1679581782
transform 1 0 14016 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_147
timestamp 1679581782
transform 1 0 14688 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_154
timestamp 1679581782
transform 1 0 15360 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_161
timestamp 1679581782
transform 1 0 16032 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_168
timestamp 1679581782
transform 1 0 16704 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_175
timestamp 1679581782
transform 1 0 17376 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_182
timestamp 1679581782
transform 1 0 18048 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_189
timestamp 1679581782
transform 1 0 18720 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_196
timestamp 1679581782
transform 1 0 19392 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_203
timestamp 1679581782
transform 1 0 20064 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_210
timestamp 1679581782
transform 1 0 20736 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_217
timestamp 1679581782
transform 1 0 21408 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_224
timestamp 1679581782
transform 1 0 22080 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_231
timestamp 1679581782
transform 1 0 22752 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_238
timestamp 1679581782
transform 1 0 23424 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_245
timestamp 1679581782
transform 1 0 24096 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_252
timestamp 1679581782
transform 1 0 24768 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_259
timestamp 1679581782
transform 1 0 25440 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_266
timestamp 1679581782
transform 1 0 26112 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_273
timestamp 1679581782
transform 1 0 26784 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_280
timestamp 1679581782
transform 1 0 27456 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_287
timestamp 1679581782
transform 1 0 28128 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_294
timestamp 1679581782
transform 1 0 28800 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_301
timestamp 1679581782
transform 1 0 29472 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_308
timestamp 1679581782
transform 1 0 30144 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_315
timestamp 1679581782
transform 1 0 30816 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_322
timestamp 1679581782
transform 1 0 31488 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_329
timestamp 1679581782
transform 1 0 32160 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_336
timestamp 1679581782
transform 1 0 32832 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_343
timestamp 1679581782
transform 1 0 33504 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_350
timestamp 1679581782
transform 1 0 34176 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_357
timestamp 1679581782
transform 1 0 34848 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_364
timestamp 1679581782
transform 1 0 35520 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_371
timestamp 1679581782
transform 1 0 36192 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_378
timestamp 1679581782
transform 1 0 36864 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_385
timestamp 1679581782
transform 1 0 37536 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_392
timestamp 1679581782
transform 1 0 38208 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_399
timestamp 1679581782
transform 1 0 38880 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_406
timestamp 1679581782
transform 1 0 39552 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_413
timestamp 1679581782
transform 1 0 40224 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_420
timestamp 1679581782
transform 1 0 40896 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_427
timestamp 1679581782
transform 1 0 41568 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_434
timestamp 1679581782
transform 1 0 42240 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_441
timestamp 1679581782
transform 1 0 42912 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_448
timestamp 1679581782
transform 1 0 43584 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_455
timestamp 1679581782
transform 1 0 44256 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_462
timestamp 1679581782
transform 1 0 44928 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_469
timestamp 1679581782
transform 1 0 45600 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_476
timestamp 1679581782
transform 1 0 46272 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_483
timestamp 1679581782
transform 1 0 46944 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_490
timestamp 1679581782
transform 1 0 47616 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_497
timestamp 1679581782
transform 1 0 48288 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_504
timestamp 1679581782
transform 1 0 48960 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_511
timestamp 1679581782
transform 1 0 49632 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_518
timestamp 1679581782
transform 1 0 50304 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_525
timestamp 1679581782
transform 1 0 50976 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_532
timestamp 1679581782
transform 1 0 51648 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_539
timestamp 1679581782
transform 1 0 52320 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_546
timestamp 1679581782
transform 1 0 52992 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_553
timestamp 1679581782
transform 1 0 53664 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_560
timestamp 1679581782
transform 1 0 54336 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_567
timestamp 1679581782
transform 1 0 55008 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_574
timestamp 1679581782
transform 1 0 55680 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_581
timestamp 1679581782
transform 1 0 56352 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_588
timestamp 1679581782
transform 1 0 57024 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_595
timestamp 1679581782
transform 1 0 57696 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_602
timestamp 1679581782
transform 1 0 58368 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_609
timestamp 1679581782
transform 1 0 59040 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_616
timestamp 1679581782
transform 1 0 59712 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_623
timestamp 1679581782
transform 1 0 60384 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_630
timestamp 1679581782
transform 1 0 61056 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_637
timestamp 1679581782
transform 1 0 61728 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_644
timestamp 1679581782
transform 1 0 62400 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_651
timestamp 1679581782
transform 1 0 63072 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_658
timestamp 1679581782
transform 1 0 63744 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_665
timestamp 1679581782
transform 1 0 64416 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_672
timestamp 1679581782
transform 1 0 65088 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_679
timestamp 1679581782
transform 1 0 65760 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_686
timestamp 1679581782
transform 1 0 66432 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_693
timestamp 1679581782
transform 1 0 67104 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_700
timestamp 1679581782
transform 1 0 67776 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_707
timestamp 1679581782
transform 1 0 68448 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_714
timestamp 1679581782
transform 1 0 69120 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_721
timestamp 1679581782
transform 1 0 69792 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_728
timestamp 1679581782
transform 1 0 70464 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_735
timestamp 1679581782
transform 1 0 71136 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_742
timestamp 1679581782
transform 1 0 71808 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_749
timestamp 1679581782
transform 1 0 72480 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_756
timestamp 1679581782
transform 1 0 73152 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_763
timestamp 1679581782
transform 1 0 73824 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_770
timestamp 1679581782
transform 1 0 74496 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_777
timestamp 1679581782
transform 1 0 75168 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_784
timestamp 1679581782
transform 1 0 75840 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_791
timestamp 1679581782
transform 1 0 76512 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_798
timestamp 1679581782
transform 1 0 77184 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_805
timestamp 1679581782
transform 1 0 77856 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_812
timestamp 1679581782
transform 1 0 78528 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_819
timestamp 1679581782
transform 1 0 79200 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_826
timestamp 1679581782
transform 1 0 79872 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_833
timestamp 1679581782
transform 1 0 80544 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_840
timestamp 1679581782
transform 1 0 81216 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_847
timestamp 1679581782
transform 1 0 81888 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_854
timestamp 1679581782
transform 1 0 82560 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_861
timestamp 1679581782
transform 1 0 83232 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_868
timestamp 1679581782
transform 1 0 83904 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_875
timestamp 1679581782
transform 1 0 84576 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_882
timestamp 1679581782
transform 1 0 85248 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_889
timestamp 1679581782
transform 1 0 85920 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_896
timestamp 1679581782
transform 1 0 86592 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_903
timestamp 1679581782
transform 1 0 87264 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_910
timestamp 1679581782
transform 1 0 87936 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_917
timestamp 1679581782
transform 1 0 88608 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_924
timestamp 1679581782
transform 1 0 89280 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_931
timestamp 1679581782
transform 1 0 89952 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_938
timestamp 1679581782
transform 1 0 90624 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_945
timestamp 1679581782
transform 1 0 91296 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_952
timestamp 1679581782
transform 1 0 91968 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_959
timestamp 1679581782
transform 1 0 92640 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_966
timestamp 1679581782
transform 1 0 93312 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_973
timestamp 1679581782
transform 1 0 93984 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_980
timestamp 1679581782
transform 1 0 94656 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_987
timestamp 1679581782
transform 1 0 95328 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_994
timestamp 1679581782
transform 1 0 96000 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_1001
timestamp 1679581782
transform 1 0 96672 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_1008
timestamp 1679581782
transform 1 0 97344 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_1015
timestamp 1679581782
transform 1 0 98016 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_1022
timestamp 1679581782
transform 1 0 98688 0 -1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_4
timestamp 1679581782
transform 1 0 960 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_11
timestamp 1679581782
transform 1 0 1632 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_18
timestamp 1679581782
transform 1 0 2304 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_25
timestamp 1679581782
transform 1 0 2976 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_32
timestamp 1679581782
transform 1 0 3648 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_39
timestamp 1679581782
transform 1 0 4320 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_46
timestamp 1679581782
transform 1 0 4992 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_53
timestamp 1679581782
transform 1 0 5664 0 1 59724
box -48 -56 720 834
use sg13g2_fill_1  FILLER_78_60
timestamp 1677579658
transform 1 0 6336 0 1 59724
box -48 -56 144 834
use sg13g2_decap_8  FILLER_78_69
timestamp 1679581782
transform 1 0 7200 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_76
timestamp 1679581782
transform 1 0 7872 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_83
timestamp 1679581782
transform 1 0 8544 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_90
timestamp 1679581782
transform 1 0 9216 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_97
timestamp 1679581782
transform 1 0 9888 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_104
timestamp 1679581782
transform 1 0 10560 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_111
timestamp 1679581782
transform 1 0 11232 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_118
timestamp 1679581782
transform 1 0 11904 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_125
timestamp 1679581782
transform 1 0 12576 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_132
timestamp 1679581782
transform 1 0 13248 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_139
timestamp 1679581782
transform 1 0 13920 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_146
timestamp 1679581782
transform 1 0 14592 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_153
timestamp 1679581782
transform 1 0 15264 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_160
timestamp 1679581782
transform 1 0 15936 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_167
timestamp 1679581782
transform 1 0 16608 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_174
timestamp 1679581782
transform 1 0 17280 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_181
timestamp 1679581782
transform 1 0 17952 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_188
timestamp 1679581782
transform 1 0 18624 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_195
timestamp 1679581782
transform 1 0 19296 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_202
timestamp 1679581782
transform 1 0 19968 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_209
timestamp 1679581782
transform 1 0 20640 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_216
timestamp 1679581782
transform 1 0 21312 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_223
timestamp 1679581782
transform 1 0 21984 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_230
timestamp 1679581782
transform 1 0 22656 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_237
timestamp 1679581782
transform 1 0 23328 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_244
timestamp 1679581782
transform 1 0 24000 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_251
timestamp 1679581782
transform 1 0 24672 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_258
timestamp 1679581782
transform 1 0 25344 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_265
timestamp 1679581782
transform 1 0 26016 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_272
timestamp 1679581782
transform 1 0 26688 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_279
timestamp 1679581782
transform 1 0 27360 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_286
timestamp 1679581782
transform 1 0 28032 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_293
timestamp 1679581782
transform 1 0 28704 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_300
timestamp 1679581782
transform 1 0 29376 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_307
timestamp 1679581782
transform 1 0 30048 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_314
timestamp 1679581782
transform 1 0 30720 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_321
timestamp 1679581782
transform 1 0 31392 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_328
timestamp 1679581782
transform 1 0 32064 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_335
timestamp 1679581782
transform 1 0 32736 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_342
timestamp 1679581782
transform 1 0 33408 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_349
timestamp 1679581782
transform 1 0 34080 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_356
timestamp 1679581782
transform 1 0 34752 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_363
timestamp 1679581782
transform 1 0 35424 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_370
timestamp 1679581782
transform 1 0 36096 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_377
timestamp 1679581782
transform 1 0 36768 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_384
timestamp 1679581782
transform 1 0 37440 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_391
timestamp 1679581782
transform 1 0 38112 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_398
timestamp 1679581782
transform 1 0 38784 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_405
timestamp 1679581782
transform 1 0 39456 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_412
timestamp 1679581782
transform 1 0 40128 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_419
timestamp 1679581782
transform 1 0 40800 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_426
timestamp 1679581782
transform 1 0 41472 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_433
timestamp 1679581782
transform 1 0 42144 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_440
timestamp 1679581782
transform 1 0 42816 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_447
timestamp 1679581782
transform 1 0 43488 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_454
timestamp 1679581782
transform 1 0 44160 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_461
timestamp 1679581782
transform 1 0 44832 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_468
timestamp 1679581782
transform 1 0 45504 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_475
timestamp 1679581782
transform 1 0 46176 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_482
timestamp 1679581782
transform 1 0 46848 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_489
timestamp 1679581782
transform 1 0 47520 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_496
timestamp 1679581782
transform 1 0 48192 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_503
timestamp 1679581782
transform 1 0 48864 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_510
timestamp 1679581782
transform 1 0 49536 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_517
timestamp 1679581782
transform 1 0 50208 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_524
timestamp 1679581782
transform 1 0 50880 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_531
timestamp 1679581782
transform 1 0 51552 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_538
timestamp 1679581782
transform 1 0 52224 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_545
timestamp 1679581782
transform 1 0 52896 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_552
timestamp 1679581782
transform 1 0 53568 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_559
timestamp 1679581782
transform 1 0 54240 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_566
timestamp 1679581782
transform 1 0 54912 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_573
timestamp 1679581782
transform 1 0 55584 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_580
timestamp 1679581782
transform 1 0 56256 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_587
timestamp 1679581782
transform 1 0 56928 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_594
timestamp 1679581782
transform 1 0 57600 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_601
timestamp 1679581782
transform 1 0 58272 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_608
timestamp 1679581782
transform 1 0 58944 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_615
timestamp 1679581782
transform 1 0 59616 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_622
timestamp 1679581782
transform 1 0 60288 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_629
timestamp 1679581782
transform 1 0 60960 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_636
timestamp 1679581782
transform 1 0 61632 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_643
timestamp 1679581782
transform 1 0 62304 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_650
timestamp 1679581782
transform 1 0 62976 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_657
timestamp 1679581782
transform 1 0 63648 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_664
timestamp 1679581782
transform 1 0 64320 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_671
timestamp 1679581782
transform 1 0 64992 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_678
timestamp 1679581782
transform 1 0 65664 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_685
timestamp 1679581782
transform 1 0 66336 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_692
timestamp 1679581782
transform 1 0 67008 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_699
timestamp 1679581782
transform 1 0 67680 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_706
timestamp 1679581782
transform 1 0 68352 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_713
timestamp 1679581782
transform 1 0 69024 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_720
timestamp 1679581782
transform 1 0 69696 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_727
timestamp 1679581782
transform 1 0 70368 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_734
timestamp 1679581782
transform 1 0 71040 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_741
timestamp 1679581782
transform 1 0 71712 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_748
timestamp 1679581782
transform 1 0 72384 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_755
timestamp 1679581782
transform 1 0 73056 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_762
timestamp 1679581782
transform 1 0 73728 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_769
timestamp 1679581782
transform 1 0 74400 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_776
timestamp 1679581782
transform 1 0 75072 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_783
timestamp 1679581782
transform 1 0 75744 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_790
timestamp 1679581782
transform 1 0 76416 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_797
timestamp 1679581782
transform 1 0 77088 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_804
timestamp 1679581782
transform 1 0 77760 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_811
timestamp 1679581782
transform 1 0 78432 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_818
timestamp 1679581782
transform 1 0 79104 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_825
timestamp 1679581782
transform 1 0 79776 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_832
timestamp 1679581782
transform 1 0 80448 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_839
timestamp 1679581782
transform 1 0 81120 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_846
timestamp 1679581782
transform 1 0 81792 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_853
timestamp 1679581782
transform 1 0 82464 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_860
timestamp 1679581782
transform 1 0 83136 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_867
timestamp 1679581782
transform 1 0 83808 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_874
timestamp 1679581782
transform 1 0 84480 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_881
timestamp 1679581782
transform 1 0 85152 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_888
timestamp 1679581782
transform 1 0 85824 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_895
timestamp 1679581782
transform 1 0 86496 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_902
timestamp 1679581782
transform 1 0 87168 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_909
timestamp 1679581782
transform 1 0 87840 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_916
timestamp 1679581782
transform 1 0 88512 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_923
timestamp 1679581782
transform 1 0 89184 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_930
timestamp 1679581782
transform 1 0 89856 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_937
timestamp 1679581782
transform 1 0 90528 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_944
timestamp 1679581782
transform 1 0 91200 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_951
timestamp 1679581782
transform 1 0 91872 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_958
timestamp 1679581782
transform 1 0 92544 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_965
timestamp 1679581782
transform 1 0 93216 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_972
timestamp 1679581782
transform 1 0 93888 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_979
timestamp 1679581782
transform 1 0 94560 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_986
timestamp 1679581782
transform 1 0 95232 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_993
timestamp 1679581782
transform 1 0 95904 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_1000
timestamp 1679581782
transform 1 0 96576 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_1007
timestamp 1679581782
transform 1 0 97248 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_1014
timestamp 1679581782
transform 1 0 97920 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_1021
timestamp 1679581782
transform 1 0 98592 0 1 59724
box -48 -56 720 834
use sg13g2_fill_1  FILLER_78_1028
timestamp 1677579658
transform 1 0 99264 0 1 59724
box -48 -56 144 834
use sg13g2_decap_8  FILLER_79_0
timestamp 1679581782
transform 1 0 576 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_7
timestamp 1679581782
transform 1 0 1248 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_14
timestamp 1679581782
transform 1 0 1920 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_21
timestamp 1679581782
transform 1 0 2592 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_28
timestamp 1679581782
transform 1 0 3264 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_35
timestamp 1679581782
transform 1 0 3936 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_42
timestamp 1679581782
transform 1 0 4608 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_49
timestamp 1679581782
transform 1 0 5280 0 -1 61236
box -48 -56 720 834
use sg13g2_fill_2  FILLER_79_56
timestamp 1677580104
transform 1 0 5952 0 -1 61236
box -48 -56 240 834
use sg13g2_fill_1  FILLER_79_58
timestamp 1677579658
transform 1 0 6144 0 -1 61236
box -48 -56 144 834
use sg13g2_decap_8  FILLER_79_67
timestamp 1679581782
transform 1 0 7008 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_74
timestamp 1679581782
transform 1 0 7680 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_81
timestamp 1679581782
transform 1 0 8352 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_88
timestamp 1679581782
transform 1 0 9024 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_95
timestamp 1679581782
transform 1 0 9696 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_102
timestamp 1679581782
transform 1 0 10368 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_109
timestamp 1679581782
transform 1 0 11040 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_116
timestamp 1679581782
transform 1 0 11712 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_123
timestamp 1679581782
transform 1 0 12384 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_130
timestamp 1679581782
transform 1 0 13056 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_137
timestamp 1679581782
transform 1 0 13728 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_144
timestamp 1679581782
transform 1 0 14400 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_151
timestamp 1679581782
transform 1 0 15072 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_158
timestamp 1679581782
transform 1 0 15744 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_165
timestamp 1679581782
transform 1 0 16416 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_172
timestamp 1679581782
transform 1 0 17088 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_179
timestamp 1679581782
transform 1 0 17760 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_186
timestamp 1679581782
transform 1 0 18432 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_193
timestamp 1679581782
transform 1 0 19104 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_200
timestamp 1679581782
transform 1 0 19776 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_207
timestamp 1679581782
transform 1 0 20448 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_214
timestamp 1679581782
transform 1 0 21120 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_221
timestamp 1679581782
transform 1 0 21792 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_228
timestamp 1679581782
transform 1 0 22464 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_235
timestamp 1679581782
transform 1 0 23136 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_242
timestamp 1679581782
transform 1 0 23808 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_249
timestamp 1679581782
transform 1 0 24480 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_256
timestamp 1679581782
transform 1 0 25152 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_263
timestamp 1679581782
transform 1 0 25824 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_270
timestamp 1679581782
transform 1 0 26496 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_277
timestamp 1679581782
transform 1 0 27168 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_284
timestamp 1679581782
transform 1 0 27840 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_291
timestamp 1679581782
transform 1 0 28512 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_298
timestamp 1679581782
transform 1 0 29184 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_305
timestamp 1679581782
transform 1 0 29856 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_312
timestamp 1679581782
transform 1 0 30528 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_319
timestamp 1679581782
transform 1 0 31200 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_326
timestamp 1679581782
transform 1 0 31872 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_333
timestamp 1679581782
transform 1 0 32544 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_340
timestamp 1679581782
transform 1 0 33216 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_347
timestamp 1679581782
transform 1 0 33888 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_354
timestamp 1679581782
transform 1 0 34560 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_361
timestamp 1679581782
transform 1 0 35232 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_368
timestamp 1679581782
transform 1 0 35904 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_375
timestamp 1679581782
transform 1 0 36576 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_382
timestamp 1679581782
transform 1 0 37248 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_389
timestamp 1679581782
transform 1 0 37920 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_396
timestamp 1679581782
transform 1 0 38592 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_403
timestamp 1679581782
transform 1 0 39264 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_410
timestamp 1679581782
transform 1 0 39936 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_417
timestamp 1679581782
transform 1 0 40608 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_424
timestamp 1679581782
transform 1 0 41280 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_431
timestamp 1679581782
transform 1 0 41952 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_438
timestamp 1679581782
transform 1 0 42624 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_445
timestamp 1679581782
transform 1 0 43296 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_452
timestamp 1679581782
transform 1 0 43968 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_459
timestamp 1679581782
transform 1 0 44640 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_466
timestamp 1679581782
transform 1 0 45312 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_473
timestamp 1679581782
transform 1 0 45984 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_480
timestamp 1679581782
transform 1 0 46656 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_487
timestamp 1679581782
transform 1 0 47328 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_494
timestamp 1679581782
transform 1 0 48000 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_501
timestamp 1679581782
transform 1 0 48672 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_508
timestamp 1679581782
transform 1 0 49344 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_515
timestamp 1679581782
transform 1 0 50016 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_522
timestamp 1679581782
transform 1 0 50688 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_529
timestamp 1679581782
transform 1 0 51360 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_536
timestamp 1679581782
transform 1 0 52032 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_543
timestamp 1679581782
transform 1 0 52704 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_550
timestamp 1679581782
transform 1 0 53376 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_557
timestamp 1679581782
transform 1 0 54048 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_564
timestamp 1679581782
transform 1 0 54720 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_571
timestamp 1679581782
transform 1 0 55392 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_578
timestamp 1679581782
transform 1 0 56064 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_585
timestamp 1679581782
transform 1 0 56736 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_592
timestamp 1679581782
transform 1 0 57408 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_599
timestamp 1679581782
transform 1 0 58080 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_606
timestamp 1679581782
transform 1 0 58752 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_613
timestamp 1679581782
transform 1 0 59424 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_620
timestamp 1679581782
transform 1 0 60096 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_627
timestamp 1679581782
transform 1 0 60768 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_634
timestamp 1679581782
transform 1 0 61440 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_641
timestamp 1679581782
transform 1 0 62112 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_648
timestamp 1679581782
transform 1 0 62784 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_655
timestamp 1679581782
transform 1 0 63456 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_662
timestamp 1679581782
transform 1 0 64128 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_669
timestamp 1679581782
transform 1 0 64800 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_676
timestamp 1679581782
transform 1 0 65472 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_683
timestamp 1679581782
transform 1 0 66144 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_690
timestamp 1679581782
transform 1 0 66816 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_697
timestamp 1679581782
transform 1 0 67488 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_704
timestamp 1679581782
transform 1 0 68160 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_711
timestamp 1679581782
transform 1 0 68832 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_718
timestamp 1679581782
transform 1 0 69504 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_725
timestamp 1679581782
transform 1 0 70176 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_732
timestamp 1679581782
transform 1 0 70848 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_739
timestamp 1679581782
transform 1 0 71520 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_746
timestamp 1679581782
transform 1 0 72192 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_753
timestamp 1679581782
transform 1 0 72864 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_760
timestamp 1679581782
transform 1 0 73536 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_767
timestamp 1679581782
transform 1 0 74208 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_774
timestamp 1679581782
transform 1 0 74880 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_781
timestamp 1679581782
transform 1 0 75552 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_788
timestamp 1679581782
transform 1 0 76224 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_795
timestamp 1679581782
transform 1 0 76896 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_802
timestamp 1679581782
transform 1 0 77568 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_809
timestamp 1679581782
transform 1 0 78240 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_816
timestamp 1679581782
transform 1 0 78912 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_823
timestamp 1679581782
transform 1 0 79584 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_830
timestamp 1679581782
transform 1 0 80256 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_837
timestamp 1679581782
transform 1 0 80928 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_844
timestamp 1679581782
transform 1 0 81600 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_851
timestamp 1679581782
transform 1 0 82272 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_858
timestamp 1679581782
transform 1 0 82944 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_865
timestamp 1679581782
transform 1 0 83616 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_872
timestamp 1679581782
transform 1 0 84288 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_879
timestamp 1679581782
transform 1 0 84960 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_886
timestamp 1679581782
transform 1 0 85632 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_893
timestamp 1679581782
transform 1 0 86304 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_900
timestamp 1679581782
transform 1 0 86976 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_907
timestamp 1679581782
transform 1 0 87648 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_914
timestamp 1679581782
transform 1 0 88320 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_921
timestamp 1679581782
transform 1 0 88992 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_928
timestamp 1679581782
transform 1 0 89664 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_935
timestamp 1679581782
transform 1 0 90336 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_942
timestamp 1679581782
transform 1 0 91008 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_949
timestamp 1679581782
transform 1 0 91680 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_956
timestamp 1679581782
transform 1 0 92352 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_963
timestamp 1679581782
transform 1 0 93024 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_970
timestamp 1679581782
transform 1 0 93696 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_977
timestamp 1679581782
transform 1 0 94368 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_984
timestamp 1679581782
transform 1 0 95040 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_991
timestamp 1679581782
transform 1 0 95712 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_998
timestamp 1679581782
transform 1 0 96384 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_1005
timestamp 1679581782
transform 1 0 97056 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_1012
timestamp 1679581782
transform 1 0 97728 0 -1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_1019
timestamp 1679581782
transform 1 0 98400 0 -1 61236
box -48 -56 720 834
use sg13g2_fill_2  FILLER_79_1026
timestamp 1677580104
transform 1 0 99072 0 -1 61236
box -48 -56 240 834
use sg13g2_fill_1  FILLER_79_1028
timestamp 1677579658
transform 1 0 99264 0 -1 61236
box -48 -56 144 834
use sg13g2_decap_8  FILLER_80_0
timestamp 1679581782
transform 1 0 576 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_7
timestamp 1679581782
transform 1 0 1248 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_14
timestamp 1679581782
transform 1 0 1920 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_21
timestamp 1679581782
transform 1 0 2592 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_28
timestamp 1679581782
transform 1 0 3264 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_35
timestamp 1679581782
transform 1 0 3936 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_42
timestamp 1679581782
transform 1 0 4608 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_49
timestamp 1679581782
transform 1 0 5280 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_56
timestamp 1679581782
transform 1 0 5952 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_63
timestamp 1679581782
transform 1 0 6624 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_70
timestamp 1679581782
transform 1 0 7296 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_77
timestamp 1679581782
transform 1 0 7968 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_84
timestamp 1679581782
transform 1 0 8640 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_91
timestamp 1679581782
transform 1 0 9312 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_98
timestamp 1679581782
transform 1 0 9984 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_105
timestamp 1679581782
transform 1 0 10656 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_112
timestamp 1679581782
transform 1 0 11328 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_119
timestamp 1679581782
transform 1 0 12000 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_126
timestamp 1679581782
transform 1 0 12672 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_133
timestamp 1679581782
transform 1 0 13344 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_140
timestamp 1679581782
transform 1 0 14016 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_147
timestamp 1679581782
transform 1 0 14688 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_154
timestamp 1679581782
transform 1 0 15360 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_161
timestamp 1679581782
transform 1 0 16032 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_168
timestamp 1679581782
transform 1 0 16704 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_175
timestamp 1679581782
transform 1 0 17376 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_182
timestamp 1679581782
transform 1 0 18048 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_189
timestamp 1679581782
transform 1 0 18720 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_196
timestamp 1679581782
transform 1 0 19392 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_203
timestamp 1679581782
transform 1 0 20064 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_210
timestamp 1679581782
transform 1 0 20736 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_217
timestamp 1679581782
transform 1 0 21408 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_224
timestamp 1679581782
transform 1 0 22080 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_231
timestamp 1679581782
transform 1 0 22752 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_238
timestamp 1679581782
transform 1 0 23424 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_245
timestamp 1679581782
transform 1 0 24096 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_252
timestamp 1679581782
transform 1 0 24768 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_259
timestamp 1679581782
transform 1 0 25440 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_266
timestamp 1679581782
transform 1 0 26112 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_273
timestamp 1679581782
transform 1 0 26784 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_280
timestamp 1679581782
transform 1 0 27456 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_287
timestamp 1679581782
transform 1 0 28128 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_294
timestamp 1679581782
transform 1 0 28800 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_301
timestamp 1679581782
transform 1 0 29472 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_308
timestamp 1679581782
transform 1 0 30144 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_315
timestamp 1679581782
transform 1 0 30816 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_322
timestamp 1679581782
transform 1 0 31488 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_329
timestamp 1679581782
transform 1 0 32160 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_336
timestamp 1679581782
transform 1 0 32832 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_343
timestamp 1679581782
transform 1 0 33504 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_350
timestamp 1679581782
transform 1 0 34176 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_357
timestamp 1679581782
transform 1 0 34848 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_364
timestamp 1679581782
transform 1 0 35520 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_371
timestamp 1679581782
transform 1 0 36192 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_378
timestamp 1679581782
transform 1 0 36864 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_385
timestamp 1679581782
transform 1 0 37536 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_392
timestamp 1679581782
transform 1 0 38208 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_399
timestamp 1679581782
transform 1 0 38880 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_406
timestamp 1679581782
transform 1 0 39552 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_413
timestamp 1679581782
transform 1 0 40224 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_420
timestamp 1679581782
transform 1 0 40896 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_427
timestamp 1679581782
transform 1 0 41568 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_434
timestamp 1679581782
transform 1 0 42240 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_441
timestamp 1679581782
transform 1 0 42912 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_448
timestamp 1679581782
transform 1 0 43584 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_455
timestamp 1679581782
transform 1 0 44256 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_462
timestamp 1679581782
transform 1 0 44928 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_469
timestamp 1679581782
transform 1 0 45600 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_476
timestamp 1679581782
transform 1 0 46272 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_483
timestamp 1679581782
transform 1 0 46944 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_490
timestamp 1679581782
transform 1 0 47616 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_497
timestamp 1679581782
transform 1 0 48288 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_504
timestamp 1679581782
transform 1 0 48960 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_511
timestamp 1679581782
transform 1 0 49632 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_518
timestamp 1679581782
transform 1 0 50304 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_525
timestamp 1679581782
transform 1 0 50976 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_532
timestamp 1679581782
transform 1 0 51648 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_539
timestamp 1679581782
transform 1 0 52320 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_546
timestamp 1679581782
transform 1 0 52992 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_553
timestamp 1679581782
transform 1 0 53664 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_560
timestamp 1679581782
transform 1 0 54336 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_567
timestamp 1679581782
transform 1 0 55008 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_574
timestamp 1679581782
transform 1 0 55680 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_581
timestamp 1679581782
transform 1 0 56352 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_588
timestamp 1679581782
transform 1 0 57024 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_595
timestamp 1679581782
transform 1 0 57696 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_602
timestamp 1679581782
transform 1 0 58368 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_609
timestamp 1679581782
transform 1 0 59040 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_616
timestamp 1679581782
transform 1 0 59712 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_623
timestamp 1679581782
transform 1 0 60384 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_630
timestamp 1679581782
transform 1 0 61056 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_637
timestamp 1679581782
transform 1 0 61728 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_644
timestamp 1679581782
transform 1 0 62400 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_651
timestamp 1679581782
transform 1 0 63072 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_658
timestamp 1679581782
transform 1 0 63744 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_665
timestamp 1679581782
transform 1 0 64416 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_672
timestamp 1679581782
transform 1 0 65088 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_679
timestamp 1679581782
transform 1 0 65760 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_686
timestamp 1679581782
transform 1 0 66432 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_693
timestamp 1679581782
transform 1 0 67104 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_700
timestamp 1679581782
transform 1 0 67776 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_707
timestamp 1679581782
transform 1 0 68448 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_714
timestamp 1679581782
transform 1 0 69120 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_721
timestamp 1679581782
transform 1 0 69792 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_728
timestamp 1679581782
transform 1 0 70464 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_735
timestamp 1679581782
transform 1 0 71136 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_742
timestamp 1679581782
transform 1 0 71808 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_749
timestamp 1679581782
transform 1 0 72480 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_756
timestamp 1679581782
transform 1 0 73152 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_763
timestamp 1679581782
transform 1 0 73824 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_770
timestamp 1679581782
transform 1 0 74496 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_777
timestamp 1679581782
transform 1 0 75168 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_784
timestamp 1679581782
transform 1 0 75840 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_791
timestamp 1679581782
transform 1 0 76512 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_798
timestamp 1679581782
transform 1 0 77184 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_805
timestamp 1679581782
transform 1 0 77856 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_812
timestamp 1679581782
transform 1 0 78528 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_819
timestamp 1679581782
transform 1 0 79200 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_826
timestamp 1679581782
transform 1 0 79872 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_833
timestamp 1679581782
transform 1 0 80544 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_840
timestamp 1679581782
transform 1 0 81216 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_847
timestamp 1679581782
transform 1 0 81888 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_854
timestamp 1679581782
transform 1 0 82560 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_861
timestamp 1679581782
transform 1 0 83232 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_868
timestamp 1679581782
transform 1 0 83904 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_875
timestamp 1679581782
transform 1 0 84576 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_882
timestamp 1679581782
transform 1 0 85248 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_889
timestamp 1679581782
transform 1 0 85920 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_896
timestamp 1679581782
transform 1 0 86592 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_903
timestamp 1679581782
transform 1 0 87264 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_910
timestamp 1679581782
transform 1 0 87936 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_917
timestamp 1679581782
transform 1 0 88608 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_924
timestamp 1679581782
transform 1 0 89280 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_931
timestamp 1679581782
transform 1 0 89952 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_938
timestamp 1679581782
transform 1 0 90624 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_945
timestamp 1679581782
transform 1 0 91296 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_952
timestamp 1679581782
transform 1 0 91968 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_959
timestamp 1679581782
transform 1 0 92640 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_966
timestamp 1679581782
transform 1 0 93312 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_973
timestamp 1679581782
transform 1 0 93984 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_980
timestamp 1679581782
transform 1 0 94656 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_987
timestamp 1679581782
transform 1 0 95328 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_994
timestamp 1679581782
transform 1 0 96000 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_1001
timestamp 1679581782
transform 1 0 96672 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_1008
timestamp 1679581782
transform 1 0 97344 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_1015
timestamp 1679581782
transform 1 0 98016 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_1022
timestamp 1679581782
transform 1 0 98688 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_4
timestamp 1679581782
transform 1 0 960 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_11
timestamp 1679581782
transform 1 0 1632 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_18
timestamp 1679581782
transform 1 0 2304 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_25
timestamp 1679581782
transform 1 0 2976 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_32
timestamp 1679581782
transform 1 0 3648 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_39
timestamp 1679581782
transform 1 0 4320 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_46
timestamp 1679581782
transform 1 0 4992 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_53
timestamp 1679581782
transform 1 0 5664 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_60
timestamp 1679581782
transform 1 0 6336 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_67
timestamp 1679581782
transform 1 0 7008 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_74
timestamp 1679581782
transform 1 0 7680 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_81
timestamp 1679581782
transform 1 0 8352 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_88
timestamp 1679581782
transform 1 0 9024 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_95
timestamp 1679581782
transform 1 0 9696 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_102
timestamp 1679581782
transform 1 0 10368 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_109
timestamp 1679581782
transform 1 0 11040 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_116
timestamp 1679581782
transform 1 0 11712 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_123
timestamp 1679581782
transform 1 0 12384 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_130
timestamp 1679581782
transform 1 0 13056 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_137
timestamp 1679581782
transform 1 0 13728 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_144
timestamp 1679581782
transform 1 0 14400 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_151
timestamp 1679581782
transform 1 0 15072 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_158
timestamp 1679581782
transform 1 0 15744 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_165
timestamp 1679581782
transform 1 0 16416 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_172
timestamp 1679581782
transform 1 0 17088 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_179
timestamp 1679581782
transform 1 0 17760 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_186
timestamp 1679581782
transform 1 0 18432 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_193
timestamp 1679581782
transform 1 0 19104 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_200
timestamp 1679581782
transform 1 0 19776 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_207
timestamp 1679581782
transform 1 0 20448 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_214
timestamp 1679581782
transform 1 0 21120 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_221
timestamp 1679581782
transform 1 0 21792 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_228
timestamp 1679581782
transform 1 0 22464 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_235
timestamp 1679581782
transform 1 0 23136 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_242
timestamp 1679581782
transform 1 0 23808 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_249
timestamp 1679581782
transform 1 0 24480 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_256
timestamp 1679581782
transform 1 0 25152 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_263
timestamp 1679581782
transform 1 0 25824 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_270
timestamp 1679581782
transform 1 0 26496 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_277
timestamp 1679581782
transform 1 0 27168 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_284
timestamp 1679581782
transform 1 0 27840 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_291
timestamp 1679581782
transform 1 0 28512 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_298
timestamp 1679581782
transform 1 0 29184 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_305
timestamp 1679581782
transform 1 0 29856 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_312
timestamp 1679581782
transform 1 0 30528 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_319
timestamp 1679581782
transform 1 0 31200 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_326
timestamp 1679581782
transform 1 0 31872 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_333
timestamp 1679581782
transform 1 0 32544 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_340
timestamp 1679581782
transform 1 0 33216 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_347
timestamp 1679581782
transform 1 0 33888 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_354
timestamp 1679581782
transform 1 0 34560 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_361
timestamp 1679581782
transform 1 0 35232 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_368
timestamp 1679581782
transform 1 0 35904 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_375
timestamp 1679581782
transform 1 0 36576 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_382
timestamp 1679581782
transform 1 0 37248 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_389
timestamp 1679581782
transform 1 0 37920 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_396
timestamp 1679581782
transform 1 0 38592 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_403
timestamp 1679581782
transform 1 0 39264 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_410
timestamp 1679581782
transform 1 0 39936 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_417
timestamp 1679581782
transform 1 0 40608 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_424
timestamp 1679581782
transform 1 0 41280 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_431
timestamp 1679581782
transform 1 0 41952 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_438
timestamp 1679581782
transform 1 0 42624 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_445
timestamp 1679581782
transform 1 0 43296 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_452
timestamp 1679581782
transform 1 0 43968 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_459
timestamp 1679581782
transform 1 0 44640 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_466
timestamp 1679581782
transform 1 0 45312 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_473
timestamp 1679581782
transform 1 0 45984 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_480
timestamp 1679581782
transform 1 0 46656 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_487
timestamp 1679581782
transform 1 0 47328 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_494
timestamp 1679581782
transform 1 0 48000 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_501
timestamp 1679581782
transform 1 0 48672 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_508
timestamp 1679581782
transform 1 0 49344 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_515
timestamp 1679581782
transform 1 0 50016 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_522
timestamp 1679581782
transform 1 0 50688 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_529
timestamp 1679581782
transform 1 0 51360 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_536
timestamp 1679581782
transform 1 0 52032 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_543
timestamp 1679581782
transform 1 0 52704 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_550
timestamp 1679581782
transform 1 0 53376 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_557
timestamp 1679581782
transform 1 0 54048 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_564
timestamp 1679581782
transform 1 0 54720 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_571
timestamp 1679581782
transform 1 0 55392 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_578
timestamp 1679581782
transform 1 0 56064 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_585
timestamp 1679581782
transform 1 0 56736 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_592
timestamp 1679581782
transform 1 0 57408 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_599
timestamp 1679581782
transform 1 0 58080 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_606
timestamp 1679581782
transform 1 0 58752 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_613
timestamp 1679581782
transform 1 0 59424 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_620
timestamp 1679581782
transform 1 0 60096 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_627
timestamp 1679581782
transform 1 0 60768 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_634
timestamp 1679581782
transform 1 0 61440 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_641
timestamp 1679581782
transform 1 0 62112 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_648
timestamp 1679581782
transform 1 0 62784 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_655
timestamp 1679581782
transform 1 0 63456 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_662
timestamp 1679581782
transform 1 0 64128 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_669
timestamp 1679581782
transform 1 0 64800 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_676
timestamp 1679581782
transform 1 0 65472 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_683
timestamp 1679581782
transform 1 0 66144 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_690
timestamp 1679581782
transform 1 0 66816 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_697
timestamp 1679581782
transform 1 0 67488 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_704
timestamp 1679581782
transform 1 0 68160 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_711
timestamp 1679581782
transform 1 0 68832 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_718
timestamp 1679581782
transform 1 0 69504 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_725
timestamp 1679581782
transform 1 0 70176 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_732
timestamp 1679581782
transform 1 0 70848 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_739
timestamp 1679581782
transform 1 0 71520 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_746
timestamp 1679581782
transform 1 0 72192 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_753
timestamp 1679581782
transform 1 0 72864 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_760
timestamp 1679581782
transform 1 0 73536 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_767
timestamp 1679581782
transform 1 0 74208 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_774
timestamp 1679581782
transform 1 0 74880 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_781
timestamp 1679581782
transform 1 0 75552 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_788
timestamp 1679581782
transform 1 0 76224 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_795
timestamp 1679581782
transform 1 0 76896 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_802
timestamp 1679581782
transform 1 0 77568 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_809
timestamp 1679581782
transform 1 0 78240 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_816
timestamp 1679581782
transform 1 0 78912 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_823
timestamp 1679581782
transform 1 0 79584 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_830
timestamp 1679581782
transform 1 0 80256 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_837
timestamp 1679581782
transform 1 0 80928 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_844
timestamp 1679581782
transform 1 0 81600 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_851
timestamp 1679581782
transform 1 0 82272 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_858
timestamp 1679581782
transform 1 0 82944 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_865
timestamp 1679581782
transform 1 0 83616 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_872
timestamp 1679581782
transform 1 0 84288 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_879
timestamp 1679581782
transform 1 0 84960 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_886
timestamp 1679581782
transform 1 0 85632 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_893
timestamp 1679581782
transform 1 0 86304 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_900
timestamp 1679581782
transform 1 0 86976 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_907
timestamp 1679581782
transform 1 0 87648 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_914
timestamp 1679581782
transform 1 0 88320 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_921
timestamp 1679581782
transform 1 0 88992 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_928
timestamp 1679581782
transform 1 0 89664 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_935
timestamp 1679581782
transform 1 0 90336 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_942
timestamp 1679581782
transform 1 0 91008 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_949
timestamp 1679581782
transform 1 0 91680 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_956
timestamp 1679581782
transform 1 0 92352 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_963
timestamp 1679581782
transform 1 0 93024 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_970
timestamp 1679581782
transform 1 0 93696 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_977
timestamp 1679581782
transform 1 0 94368 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_984
timestamp 1679581782
transform 1 0 95040 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_991
timestamp 1679581782
transform 1 0 95712 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_998
timestamp 1679581782
transform 1 0 96384 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_1005
timestamp 1679581782
transform 1 0 97056 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_1012
timestamp 1679581782
transform 1 0 97728 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_1019
timestamp 1679581782
transform 1 0 98400 0 -1 62748
box -48 -56 720 834
use sg13g2_fill_2  FILLER_81_1026
timestamp 1677580104
transform 1 0 99072 0 -1 62748
box -48 -56 240 834
use sg13g2_fill_1  FILLER_81_1028
timestamp 1677579658
transform 1 0 99264 0 -1 62748
box -48 -56 144 834
use sg13g2_decap_8  FILLER_82_0
timestamp 1679581782
transform 1 0 576 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_7
timestamp 1679581782
transform 1 0 1248 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_14
timestamp 1679581782
transform 1 0 1920 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_21
timestamp 1679581782
transform 1 0 2592 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_28
timestamp 1679581782
transform 1 0 3264 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_35
timestamp 1679581782
transform 1 0 3936 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_42
timestamp 1679581782
transform 1 0 4608 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_49
timestamp 1679581782
transform 1 0 5280 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_56
timestamp 1679581782
transform 1 0 5952 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_63
timestamp 1679581782
transform 1 0 6624 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_70
timestamp 1679581782
transform 1 0 7296 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_77
timestamp 1679581782
transform 1 0 7968 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_84
timestamp 1679581782
transform 1 0 8640 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_91
timestamp 1679581782
transform 1 0 9312 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_98
timestamp 1679581782
transform 1 0 9984 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_105
timestamp 1679581782
transform 1 0 10656 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_112
timestamp 1679581782
transform 1 0 11328 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_119
timestamp 1679581782
transform 1 0 12000 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_126
timestamp 1679581782
transform 1 0 12672 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_133
timestamp 1679581782
transform 1 0 13344 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_140
timestamp 1679581782
transform 1 0 14016 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_147
timestamp 1679581782
transform 1 0 14688 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_154
timestamp 1679581782
transform 1 0 15360 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_161
timestamp 1679581782
transform 1 0 16032 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_168
timestamp 1679581782
transform 1 0 16704 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_175
timestamp 1679581782
transform 1 0 17376 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_182
timestamp 1679581782
transform 1 0 18048 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_189
timestamp 1679581782
transform 1 0 18720 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_196
timestamp 1679581782
transform 1 0 19392 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_203
timestamp 1679581782
transform 1 0 20064 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_210
timestamp 1679581782
transform 1 0 20736 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_217
timestamp 1679581782
transform 1 0 21408 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_224
timestamp 1679581782
transform 1 0 22080 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_231
timestamp 1679581782
transform 1 0 22752 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_238
timestamp 1679581782
transform 1 0 23424 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_245
timestamp 1679581782
transform 1 0 24096 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_252
timestamp 1679581782
transform 1 0 24768 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_259
timestamp 1679581782
transform 1 0 25440 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_266
timestamp 1679581782
transform 1 0 26112 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_273
timestamp 1679581782
transform 1 0 26784 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_280
timestamp 1679581782
transform 1 0 27456 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_287
timestamp 1679581782
transform 1 0 28128 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_294
timestamp 1679581782
transform 1 0 28800 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_301
timestamp 1679581782
transform 1 0 29472 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_308
timestamp 1679581782
transform 1 0 30144 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_315
timestamp 1679581782
transform 1 0 30816 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_322
timestamp 1679581782
transform 1 0 31488 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_329
timestamp 1679581782
transform 1 0 32160 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_336
timestamp 1679581782
transform 1 0 32832 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_343
timestamp 1679581782
transform 1 0 33504 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_350
timestamp 1679581782
transform 1 0 34176 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_357
timestamp 1679581782
transform 1 0 34848 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_364
timestamp 1679581782
transform 1 0 35520 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_371
timestamp 1679581782
transform 1 0 36192 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_378
timestamp 1679581782
transform 1 0 36864 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_385
timestamp 1679581782
transform 1 0 37536 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_392
timestamp 1679581782
transform 1 0 38208 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_399
timestamp 1679581782
transform 1 0 38880 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_406
timestamp 1679581782
transform 1 0 39552 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_413
timestamp 1679581782
transform 1 0 40224 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_420
timestamp 1679581782
transform 1 0 40896 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_427
timestamp 1679581782
transform 1 0 41568 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_434
timestamp 1679581782
transform 1 0 42240 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_441
timestamp 1679581782
transform 1 0 42912 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_448
timestamp 1679581782
transform 1 0 43584 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_455
timestamp 1679581782
transform 1 0 44256 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_462
timestamp 1679581782
transform 1 0 44928 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_469
timestamp 1679581782
transform 1 0 45600 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_476
timestamp 1679581782
transform 1 0 46272 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_483
timestamp 1679581782
transform 1 0 46944 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_490
timestamp 1679581782
transform 1 0 47616 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_497
timestamp 1679581782
transform 1 0 48288 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_504
timestamp 1679581782
transform 1 0 48960 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_511
timestamp 1679581782
transform 1 0 49632 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_518
timestamp 1679581782
transform 1 0 50304 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_525
timestamp 1679581782
transform 1 0 50976 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_532
timestamp 1679581782
transform 1 0 51648 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_539
timestamp 1679581782
transform 1 0 52320 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_546
timestamp 1679581782
transform 1 0 52992 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_553
timestamp 1679581782
transform 1 0 53664 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_560
timestamp 1679581782
transform 1 0 54336 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_567
timestamp 1679581782
transform 1 0 55008 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_574
timestamp 1679581782
transform 1 0 55680 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_581
timestamp 1679581782
transform 1 0 56352 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_588
timestamp 1679581782
transform 1 0 57024 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_595
timestamp 1679581782
transform 1 0 57696 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_602
timestamp 1679581782
transform 1 0 58368 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_609
timestamp 1679581782
transform 1 0 59040 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_616
timestamp 1679581782
transform 1 0 59712 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_623
timestamp 1679581782
transform 1 0 60384 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_630
timestamp 1679581782
transform 1 0 61056 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_637
timestamp 1679581782
transform 1 0 61728 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_644
timestamp 1679581782
transform 1 0 62400 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_651
timestamp 1679581782
transform 1 0 63072 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_658
timestamp 1679581782
transform 1 0 63744 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_665
timestamp 1679581782
transform 1 0 64416 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_672
timestamp 1679581782
transform 1 0 65088 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_679
timestamp 1679581782
transform 1 0 65760 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_686
timestamp 1679581782
transform 1 0 66432 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_693
timestamp 1679581782
transform 1 0 67104 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_700
timestamp 1679581782
transform 1 0 67776 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_707
timestamp 1679581782
transform 1 0 68448 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_714
timestamp 1679581782
transform 1 0 69120 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_721
timestamp 1679581782
transform 1 0 69792 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_728
timestamp 1679581782
transform 1 0 70464 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_735
timestamp 1679581782
transform 1 0 71136 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_742
timestamp 1679581782
transform 1 0 71808 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_749
timestamp 1679581782
transform 1 0 72480 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_756
timestamp 1679581782
transform 1 0 73152 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_763
timestamp 1679581782
transform 1 0 73824 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_770
timestamp 1679581782
transform 1 0 74496 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_777
timestamp 1679581782
transform 1 0 75168 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_784
timestamp 1679581782
transform 1 0 75840 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_791
timestamp 1679581782
transform 1 0 76512 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_798
timestamp 1679581782
transform 1 0 77184 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_805
timestamp 1679581782
transform 1 0 77856 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_812
timestamp 1679581782
transform 1 0 78528 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_819
timestamp 1679581782
transform 1 0 79200 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_826
timestamp 1679581782
transform 1 0 79872 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_833
timestamp 1679581782
transform 1 0 80544 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_840
timestamp 1679581782
transform 1 0 81216 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_847
timestamp 1679581782
transform 1 0 81888 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_854
timestamp 1679581782
transform 1 0 82560 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_861
timestamp 1679581782
transform 1 0 83232 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_868
timestamp 1679581782
transform 1 0 83904 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_875
timestamp 1679581782
transform 1 0 84576 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_882
timestamp 1679581782
transform 1 0 85248 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_889
timestamp 1679581782
transform 1 0 85920 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_896
timestamp 1679581782
transform 1 0 86592 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_903
timestamp 1679581782
transform 1 0 87264 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_910
timestamp 1679581782
transform 1 0 87936 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_917
timestamp 1679581782
transform 1 0 88608 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_924
timestamp 1679581782
transform 1 0 89280 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_931
timestamp 1679581782
transform 1 0 89952 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_938
timestamp 1679581782
transform 1 0 90624 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_945
timestamp 1679581782
transform 1 0 91296 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_952
timestamp 1679581782
transform 1 0 91968 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_959
timestamp 1679581782
transform 1 0 92640 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_966
timestamp 1679581782
transform 1 0 93312 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_973
timestamp 1679581782
transform 1 0 93984 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_980
timestamp 1679581782
transform 1 0 94656 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_987
timestamp 1679581782
transform 1 0 95328 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_994
timestamp 1679581782
transform 1 0 96000 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_1001
timestamp 1679581782
transform 1 0 96672 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_1008
timestamp 1679581782
transform 1 0 97344 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_1015
timestamp 1679581782
transform 1 0 98016 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_1022
timestamp 1679581782
transform 1 0 98688 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_4
timestamp 1679581782
transform 1 0 960 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_11
timestamp 1679581782
transform 1 0 1632 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_18
timestamp 1679581782
transform 1 0 2304 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_25
timestamp 1679581782
transform 1 0 2976 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_32
timestamp 1679581782
transform 1 0 3648 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_39
timestamp 1679581782
transform 1 0 4320 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_46
timestamp 1679581782
transform 1 0 4992 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_53
timestamp 1679581782
transform 1 0 5664 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_60
timestamp 1679581782
transform 1 0 6336 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_67
timestamp 1679581782
transform 1 0 7008 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_74
timestamp 1679581782
transform 1 0 7680 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_81
timestamp 1679581782
transform 1 0 8352 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_88
timestamp 1679581782
transform 1 0 9024 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_95
timestamp 1679581782
transform 1 0 9696 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_102
timestamp 1679581782
transform 1 0 10368 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_109
timestamp 1679581782
transform 1 0 11040 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_116
timestamp 1679581782
transform 1 0 11712 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_123
timestamp 1679581782
transform 1 0 12384 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_130
timestamp 1679581782
transform 1 0 13056 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_137
timestamp 1679581782
transform 1 0 13728 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_144
timestamp 1679581782
transform 1 0 14400 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_151
timestamp 1679581782
transform 1 0 15072 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_158
timestamp 1679581782
transform 1 0 15744 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_165
timestamp 1679581782
transform 1 0 16416 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_172
timestamp 1679581782
transform 1 0 17088 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_179
timestamp 1679581782
transform 1 0 17760 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_186
timestamp 1679581782
transform 1 0 18432 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_193
timestamp 1679581782
transform 1 0 19104 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_200
timestamp 1679581782
transform 1 0 19776 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_207
timestamp 1679581782
transform 1 0 20448 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_214
timestamp 1679581782
transform 1 0 21120 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_221
timestamp 1679581782
transform 1 0 21792 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_228
timestamp 1679581782
transform 1 0 22464 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_235
timestamp 1679581782
transform 1 0 23136 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_242
timestamp 1679581782
transform 1 0 23808 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_249
timestamp 1679581782
transform 1 0 24480 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_256
timestamp 1679581782
transform 1 0 25152 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_263
timestamp 1679581782
transform 1 0 25824 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_270
timestamp 1679581782
transform 1 0 26496 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_277
timestamp 1679581782
transform 1 0 27168 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_284
timestamp 1679581782
transform 1 0 27840 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_291
timestamp 1679581782
transform 1 0 28512 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_298
timestamp 1679581782
transform 1 0 29184 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_305
timestamp 1679581782
transform 1 0 29856 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_312
timestamp 1679581782
transform 1 0 30528 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_319
timestamp 1679581782
transform 1 0 31200 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_326
timestamp 1679581782
transform 1 0 31872 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_333
timestamp 1679581782
transform 1 0 32544 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_340
timestamp 1679581782
transform 1 0 33216 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_347
timestamp 1679581782
transform 1 0 33888 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_354
timestamp 1679581782
transform 1 0 34560 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_361
timestamp 1679581782
transform 1 0 35232 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_368
timestamp 1679581782
transform 1 0 35904 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_375
timestamp 1679581782
transform 1 0 36576 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_382
timestamp 1679581782
transform 1 0 37248 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_389
timestamp 1679581782
transform 1 0 37920 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_396
timestamp 1679581782
transform 1 0 38592 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_403
timestamp 1679581782
transform 1 0 39264 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_410
timestamp 1679581782
transform 1 0 39936 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_417
timestamp 1679581782
transform 1 0 40608 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_424
timestamp 1679581782
transform 1 0 41280 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_431
timestamp 1679581782
transform 1 0 41952 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_438
timestamp 1679581782
transform 1 0 42624 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_445
timestamp 1679581782
transform 1 0 43296 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_452
timestamp 1679581782
transform 1 0 43968 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_459
timestamp 1679581782
transform 1 0 44640 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_466
timestamp 1679581782
transform 1 0 45312 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_473
timestamp 1679581782
transform 1 0 45984 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_480
timestamp 1679581782
transform 1 0 46656 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_487
timestamp 1679581782
transform 1 0 47328 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_494
timestamp 1679581782
transform 1 0 48000 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_501
timestamp 1679581782
transform 1 0 48672 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_508
timestamp 1679581782
transform 1 0 49344 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_515
timestamp 1679581782
transform 1 0 50016 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_522
timestamp 1679581782
transform 1 0 50688 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_529
timestamp 1679581782
transform 1 0 51360 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_536
timestamp 1679581782
transform 1 0 52032 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_543
timestamp 1679581782
transform 1 0 52704 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_550
timestamp 1679581782
transform 1 0 53376 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_557
timestamp 1679581782
transform 1 0 54048 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_564
timestamp 1679581782
transform 1 0 54720 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_571
timestamp 1679581782
transform 1 0 55392 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_578
timestamp 1679581782
transform 1 0 56064 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_585
timestamp 1679581782
transform 1 0 56736 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_592
timestamp 1679581782
transform 1 0 57408 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_599
timestamp 1679581782
transform 1 0 58080 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_606
timestamp 1679581782
transform 1 0 58752 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_613
timestamp 1679581782
transform 1 0 59424 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_620
timestamp 1679581782
transform 1 0 60096 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_627
timestamp 1679581782
transform 1 0 60768 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_634
timestamp 1679581782
transform 1 0 61440 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_641
timestamp 1679581782
transform 1 0 62112 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_648
timestamp 1679581782
transform 1 0 62784 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_655
timestamp 1679581782
transform 1 0 63456 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_662
timestamp 1679581782
transform 1 0 64128 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_669
timestamp 1679581782
transform 1 0 64800 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_676
timestamp 1679581782
transform 1 0 65472 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_683
timestamp 1679581782
transform 1 0 66144 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_690
timestamp 1679581782
transform 1 0 66816 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_697
timestamp 1679581782
transform 1 0 67488 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_704
timestamp 1679581782
transform 1 0 68160 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_711
timestamp 1679581782
transform 1 0 68832 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_718
timestamp 1679581782
transform 1 0 69504 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_725
timestamp 1679581782
transform 1 0 70176 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_732
timestamp 1679581782
transform 1 0 70848 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_739
timestamp 1679581782
transform 1 0 71520 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_746
timestamp 1679581782
transform 1 0 72192 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_753
timestamp 1679581782
transform 1 0 72864 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_760
timestamp 1679581782
transform 1 0 73536 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_767
timestamp 1679581782
transform 1 0 74208 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_774
timestamp 1679581782
transform 1 0 74880 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_781
timestamp 1679581782
transform 1 0 75552 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_788
timestamp 1679581782
transform 1 0 76224 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_795
timestamp 1679581782
transform 1 0 76896 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_802
timestamp 1679581782
transform 1 0 77568 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_809
timestamp 1679581782
transform 1 0 78240 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_816
timestamp 1679581782
transform 1 0 78912 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_823
timestamp 1679581782
transform 1 0 79584 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_830
timestamp 1679581782
transform 1 0 80256 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_837
timestamp 1679581782
transform 1 0 80928 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_844
timestamp 1679581782
transform 1 0 81600 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_851
timestamp 1679581782
transform 1 0 82272 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_858
timestamp 1679581782
transform 1 0 82944 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_865
timestamp 1679581782
transform 1 0 83616 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_872
timestamp 1679581782
transform 1 0 84288 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_879
timestamp 1679581782
transform 1 0 84960 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_886
timestamp 1679581782
transform 1 0 85632 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_893
timestamp 1679581782
transform 1 0 86304 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_900
timestamp 1679581782
transform 1 0 86976 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_907
timestamp 1679581782
transform 1 0 87648 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_914
timestamp 1679581782
transform 1 0 88320 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_921
timestamp 1679581782
transform 1 0 88992 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_928
timestamp 1679581782
transform 1 0 89664 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_935
timestamp 1679581782
transform 1 0 90336 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_942
timestamp 1679581782
transform 1 0 91008 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_949
timestamp 1679581782
transform 1 0 91680 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_956
timestamp 1679581782
transform 1 0 92352 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_963
timestamp 1679581782
transform 1 0 93024 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_970
timestamp 1679581782
transform 1 0 93696 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_977
timestamp 1679581782
transform 1 0 94368 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_984
timestamp 1679581782
transform 1 0 95040 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_991
timestamp 1679581782
transform 1 0 95712 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_998
timestamp 1679581782
transform 1 0 96384 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_1005
timestamp 1679581782
transform 1 0 97056 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_1012
timestamp 1679581782
transform 1 0 97728 0 -1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_1019
timestamp 1679581782
transform 1 0 98400 0 -1 64260
box -48 -56 720 834
use sg13g2_fill_2  FILLER_83_1026
timestamp 1677580104
transform 1 0 99072 0 -1 64260
box -48 -56 240 834
use sg13g2_fill_1  FILLER_83_1028
timestamp 1677579658
transform 1 0 99264 0 -1 64260
box -48 -56 144 834
use sg13g2_decap_8  FILLER_84_0
timestamp 1679581782
transform 1 0 576 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_7
timestamp 1679581782
transform 1 0 1248 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_14
timestamp 1679581782
transform 1 0 1920 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_21
timestamp 1679581782
transform 1 0 2592 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_28
timestamp 1679581782
transform 1 0 3264 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_35
timestamp 1679581782
transform 1 0 3936 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_42
timestamp 1679581782
transform 1 0 4608 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_49
timestamp 1679581782
transform 1 0 5280 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_56
timestamp 1679581782
transform 1 0 5952 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_63
timestamp 1679581782
transform 1 0 6624 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_70
timestamp 1679581782
transform 1 0 7296 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_77
timestamp 1679581782
transform 1 0 7968 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_84
timestamp 1679581782
transform 1 0 8640 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_91
timestamp 1679581782
transform 1 0 9312 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_98
timestamp 1679581782
transform 1 0 9984 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_105
timestamp 1679581782
transform 1 0 10656 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_112
timestamp 1679581782
transform 1 0 11328 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_119
timestamp 1679581782
transform 1 0 12000 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_126
timestamp 1679581782
transform 1 0 12672 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_133
timestamp 1679581782
transform 1 0 13344 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_140
timestamp 1679581782
transform 1 0 14016 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_147
timestamp 1679581782
transform 1 0 14688 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_154
timestamp 1679581782
transform 1 0 15360 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_161
timestamp 1679581782
transform 1 0 16032 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_168
timestamp 1679581782
transform 1 0 16704 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_175
timestamp 1679581782
transform 1 0 17376 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_182
timestamp 1679581782
transform 1 0 18048 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_189
timestamp 1679581782
transform 1 0 18720 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_196
timestamp 1679581782
transform 1 0 19392 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_203
timestamp 1679581782
transform 1 0 20064 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_210
timestamp 1679581782
transform 1 0 20736 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_217
timestamp 1679581782
transform 1 0 21408 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_224
timestamp 1679581782
transform 1 0 22080 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_231
timestamp 1679581782
transform 1 0 22752 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_238
timestamp 1679581782
transform 1 0 23424 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_245
timestamp 1679581782
transform 1 0 24096 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_252
timestamp 1679581782
transform 1 0 24768 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_259
timestamp 1679581782
transform 1 0 25440 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_266
timestamp 1679581782
transform 1 0 26112 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_273
timestamp 1679581782
transform 1 0 26784 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_280
timestamp 1679581782
transform 1 0 27456 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_287
timestamp 1679581782
transform 1 0 28128 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_294
timestamp 1679581782
transform 1 0 28800 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_301
timestamp 1679581782
transform 1 0 29472 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_308
timestamp 1679581782
transform 1 0 30144 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_315
timestamp 1679581782
transform 1 0 30816 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_322
timestamp 1679581782
transform 1 0 31488 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_329
timestamp 1679581782
transform 1 0 32160 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_336
timestamp 1679581782
transform 1 0 32832 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_343
timestamp 1679581782
transform 1 0 33504 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_350
timestamp 1679581782
transform 1 0 34176 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_357
timestamp 1679581782
transform 1 0 34848 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_364
timestamp 1679581782
transform 1 0 35520 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_371
timestamp 1679581782
transform 1 0 36192 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_378
timestamp 1679581782
transform 1 0 36864 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_385
timestamp 1679581782
transform 1 0 37536 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_392
timestamp 1679581782
transform 1 0 38208 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_399
timestamp 1679581782
transform 1 0 38880 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_406
timestamp 1679581782
transform 1 0 39552 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_413
timestamp 1679581782
transform 1 0 40224 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_420
timestamp 1679581782
transform 1 0 40896 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_427
timestamp 1679581782
transform 1 0 41568 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_434
timestamp 1679581782
transform 1 0 42240 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_441
timestamp 1679581782
transform 1 0 42912 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_448
timestamp 1679581782
transform 1 0 43584 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_455
timestamp 1679581782
transform 1 0 44256 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_462
timestamp 1679581782
transform 1 0 44928 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_469
timestamp 1679581782
transform 1 0 45600 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_476
timestamp 1679581782
transform 1 0 46272 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_483
timestamp 1679581782
transform 1 0 46944 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_490
timestamp 1679581782
transform 1 0 47616 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_497
timestamp 1679581782
transform 1 0 48288 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_504
timestamp 1679581782
transform 1 0 48960 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_511
timestamp 1679581782
transform 1 0 49632 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_518
timestamp 1679581782
transform 1 0 50304 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_525
timestamp 1679581782
transform 1 0 50976 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_532
timestamp 1679581782
transform 1 0 51648 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_539
timestamp 1679581782
transform 1 0 52320 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_546
timestamp 1679581782
transform 1 0 52992 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_553
timestamp 1679581782
transform 1 0 53664 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_560
timestamp 1679581782
transform 1 0 54336 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_567
timestamp 1679581782
transform 1 0 55008 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_574
timestamp 1679581782
transform 1 0 55680 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_581
timestamp 1679581782
transform 1 0 56352 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_588
timestamp 1679581782
transform 1 0 57024 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_595
timestamp 1679581782
transform 1 0 57696 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_602
timestamp 1679581782
transform 1 0 58368 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_609
timestamp 1679581782
transform 1 0 59040 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_616
timestamp 1679581782
transform 1 0 59712 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_623
timestamp 1679581782
transform 1 0 60384 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_630
timestamp 1679581782
transform 1 0 61056 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_637
timestamp 1679581782
transform 1 0 61728 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_644
timestamp 1679581782
transform 1 0 62400 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_651
timestamp 1679581782
transform 1 0 63072 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_658
timestamp 1679581782
transform 1 0 63744 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_665
timestamp 1679581782
transform 1 0 64416 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_672
timestamp 1679581782
transform 1 0 65088 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_679
timestamp 1679581782
transform 1 0 65760 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_686
timestamp 1679581782
transform 1 0 66432 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_693
timestamp 1679581782
transform 1 0 67104 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_700
timestamp 1679581782
transform 1 0 67776 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_707
timestamp 1679581782
transform 1 0 68448 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_714
timestamp 1679581782
transform 1 0 69120 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_721
timestamp 1679581782
transform 1 0 69792 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_728
timestamp 1679581782
transform 1 0 70464 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_735
timestamp 1679581782
transform 1 0 71136 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_742
timestamp 1679581782
transform 1 0 71808 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_749
timestamp 1679581782
transform 1 0 72480 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_756
timestamp 1679581782
transform 1 0 73152 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_763
timestamp 1679581782
transform 1 0 73824 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_770
timestamp 1679581782
transform 1 0 74496 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_777
timestamp 1679581782
transform 1 0 75168 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_784
timestamp 1679581782
transform 1 0 75840 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_791
timestamp 1679581782
transform 1 0 76512 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_798
timestamp 1679581782
transform 1 0 77184 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_805
timestamp 1679581782
transform 1 0 77856 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_812
timestamp 1679581782
transform 1 0 78528 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_819
timestamp 1679581782
transform 1 0 79200 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_826
timestamp 1679581782
transform 1 0 79872 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_833
timestamp 1679581782
transform 1 0 80544 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_840
timestamp 1679581782
transform 1 0 81216 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_847
timestamp 1679581782
transform 1 0 81888 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_854
timestamp 1679581782
transform 1 0 82560 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_861
timestamp 1679581782
transform 1 0 83232 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_868
timestamp 1679581782
transform 1 0 83904 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_875
timestamp 1679581782
transform 1 0 84576 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_882
timestamp 1679581782
transform 1 0 85248 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_889
timestamp 1679581782
transform 1 0 85920 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_896
timestamp 1679581782
transform 1 0 86592 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_903
timestamp 1679581782
transform 1 0 87264 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_910
timestamp 1679581782
transform 1 0 87936 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_917
timestamp 1679581782
transform 1 0 88608 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_924
timestamp 1679581782
transform 1 0 89280 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_931
timestamp 1679581782
transform 1 0 89952 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_938
timestamp 1679581782
transform 1 0 90624 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_945
timestamp 1679581782
transform 1 0 91296 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_952
timestamp 1679581782
transform 1 0 91968 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_959
timestamp 1679581782
transform 1 0 92640 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_966
timestamp 1679581782
transform 1 0 93312 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_973
timestamp 1679581782
transform 1 0 93984 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_980
timestamp 1679581782
transform 1 0 94656 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_987
timestamp 1679581782
transform 1 0 95328 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_994
timestamp 1679581782
transform 1 0 96000 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_1001
timestamp 1679581782
transform 1 0 96672 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_1008
timestamp 1679581782
transform 1 0 97344 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_1015
timestamp 1679581782
transform 1 0 98016 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_1022
timestamp 1679581782
transform 1 0 98688 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_0
timestamp 1679581782
transform 1 0 576 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_7
timestamp 1679581782
transform 1 0 1248 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_14
timestamp 1679581782
transform 1 0 1920 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_21
timestamp 1679581782
transform 1 0 2592 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_28
timestamp 1679581782
transform 1 0 3264 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_35
timestamp 1679581782
transform 1 0 3936 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_42
timestamp 1679581782
transform 1 0 4608 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_49
timestamp 1679581782
transform 1 0 5280 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_56
timestamp 1679581782
transform 1 0 5952 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_63
timestamp 1679581782
transform 1 0 6624 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_70
timestamp 1679581782
transform 1 0 7296 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_77
timestamp 1679581782
transform 1 0 7968 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_84
timestamp 1679581782
transform 1 0 8640 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_91
timestamp 1679581782
transform 1 0 9312 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_98
timestamp 1679581782
transform 1 0 9984 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_105
timestamp 1679581782
transform 1 0 10656 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_112
timestamp 1679581782
transform 1 0 11328 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_119
timestamp 1679581782
transform 1 0 12000 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_126
timestamp 1679581782
transform 1 0 12672 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_133
timestamp 1679581782
transform 1 0 13344 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_140
timestamp 1679581782
transform 1 0 14016 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_147
timestamp 1679581782
transform 1 0 14688 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_154
timestamp 1679581782
transform 1 0 15360 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_161
timestamp 1679581782
transform 1 0 16032 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_168
timestamp 1679581782
transform 1 0 16704 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_175
timestamp 1679581782
transform 1 0 17376 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_182
timestamp 1679581782
transform 1 0 18048 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_189
timestamp 1679581782
transform 1 0 18720 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_196
timestamp 1679581782
transform 1 0 19392 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_203
timestamp 1679581782
transform 1 0 20064 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_210
timestamp 1679581782
transform 1 0 20736 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_217
timestamp 1679581782
transform 1 0 21408 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_224
timestamp 1679581782
transform 1 0 22080 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_231
timestamp 1679581782
transform 1 0 22752 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_238
timestamp 1679581782
transform 1 0 23424 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_245
timestamp 1679581782
transform 1 0 24096 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_252
timestamp 1679581782
transform 1 0 24768 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_259
timestamp 1679581782
transform 1 0 25440 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_266
timestamp 1679581782
transform 1 0 26112 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_273
timestamp 1679581782
transform 1 0 26784 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_280
timestamp 1679581782
transform 1 0 27456 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_287
timestamp 1679581782
transform 1 0 28128 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_294
timestamp 1679581782
transform 1 0 28800 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_301
timestamp 1679581782
transform 1 0 29472 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_308
timestamp 1679581782
transform 1 0 30144 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_315
timestamp 1679581782
transform 1 0 30816 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_322
timestamp 1679581782
transform 1 0 31488 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_329
timestamp 1679581782
transform 1 0 32160 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_336
timestamp 1679581782
transform 1 0 32832 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_343
timestamp 1679581782
transform 1 0 33504 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_350
timestamp 1679581782
transform 1 0 34176 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_357
timestamp 1679581782
transform 1 0 34848 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_364
timestamp 1679581782
transform 1 0 35520 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_371
timestamp 1679581782
transform 1 0 36192 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_378
timestamp 1679581782
transform 1 0 36864 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_385
timestamp 1679581782
transform 1 0 37536 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_392
timestamp 1679581782
transform 1 0 38208 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_399
timestamp 1679581782
transform 1 0 38880 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_406
timestamp 1679581782
transform 1 0 39552 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_413
timestamp 1679581782
transform 1 0 40224 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_420
timestamp 1679581782
transform 1 0 40896 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_427
timestamp 1679581782
transform 1 0 41568 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_434
timestamp 1679581782
transform 1 0 42240 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_441
timestamp 1679581782
transform 1 0 42912 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_448
timestamp 1679581782
transform 1 0 43584 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_455
timestamp 1679581782
transform 1 0 44256 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_462
timestamp 1679581782
transform 1 0 44928 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_469
timestamp 1679581782
transform 1 0 45600 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_476
timestamp 1679581782
transform 1 0 46272 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_483
timestamp 1679581782
transform 1 0 46944 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_490
timestamp 1679581782
transform 1 0 47616 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_497
timestamp 1679581782
transform 1 0 48288 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_504
timestamp 1679581782
transform 1 0 48960 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_511
timestamp 1679581782
transform 1 0 49632 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_518
timestamp 1679581782
transform 1 0 50304 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_525
timestamp 1679581782
transform 1 0 50976 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_532
timestamp 1679581782
transform 1 0 51648 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_539
timestamp 1679581782
transform 1 0 52320 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_546
timestamp 1679581782
transform 1 0 52992 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_553
timestamp 1679581782
transform 1 0 53664 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_560
timestamp 1679581782
transform 1 0 54336 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_567
timestamp 1679581782
transform 1 0 55008 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_574
timestamp 1679581782
transform 1 0 55680 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_581
timestamp 1679581782
transform 1 0 56352 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_588
timestamp 1679581782
transform 1 0 57024 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_595
timestamp 1679581782
transform 1 0 57696 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_602
timestamp 1679581782
transform 1 0 58368 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_609
timestamp 1679581782
transform 1 0 59040 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_616
timestamp 1679581782
transform 1 0 59712 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_623
timestamp 1679581782
transform 1 0 60384 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_630
timestamp 1679581782
transform 1 0 61056 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_637
timestamp 1679581782
transform 1 0 61728 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_644
timestamp 1679581782
transform 1 0 62400 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_651
timestamp 1679581782
transform 1 0 63072 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_658
timestamp 1679581782
transform 1 0 63744 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_665
timestamp 1679581782
transform 1 0 64416 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_672
timestamp 1679581782
transform 1 0 65088 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_679
timestamp 1679581782
transform 1 0 65760 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_686
timestamp 1679581782
transform 1 0 66432 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_693
timestamp 1679581782
transform 1 0 67104 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_700
timestamp 1679581782
transform 1 0 67776 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_707
timestamp 1679581782
transform 1 0 68448 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_714
timestamp 1679581782
transform 1 0 69120 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_721
timestamp 1679581782
transform 1 0 69792 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_728
timestamp 1679581782
transform 1 0 70464 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_735
timestamp 1679581782
transform 1 0 71136 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_742
timestamp 1679581782
transform 1 0 71808 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_749
timestamp 1679581782
transform 1 0 72480 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_756
timestamp 1679581782
transform 1 0 73152 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_763
timestamp 1679581782
transform 1 0 73824 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_770
timestamp 1679581782
transform 1 0 74496 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_777
timestamp 1679581782
transform 1 0 75168 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_784
timestamp 1679581782
transform 1 0 75840 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_791
timestamp 1679581782
transform 1 0 76512 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_798
timestamp 1679581782
transform 1 0 77184 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_805
timestamp 1679581782
transform 1 0 77856 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_812
timestamp 1679581782
transform 1 0 78528 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_819
timestamp 1679581782
transform 1 0 79200 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_826
timestamp 1679581782
transform 1 0 79872 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_833
timestamp 1679581782
transform 1 0 80544 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_840
timestamp 1679581782
transform 1 0 81216 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_847
timestamp 1679581782
transform 1 0 81888 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_854
timestamp 1679581782
transform 1 0 82560 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_861
timestamp 1679581782
transform 1 0 83232 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_868
timestamp 1679581782
transform 1 0 83904 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_875
timestamp 1679581782
transform 1 0 84576 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_882
timestamp 1679581782
transform 1 0 85248 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_889
timestamp 1679581782
transform 1 0 85920 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_896
timestamp 1679581782
transform 1 0 86592 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_903
timestamp 1679581782
transform 1 0 87264 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_910
timestamp 1679581782
transform 1 0 87936 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_917
timestamp 1679581782
transform 1 0 88608 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_924
timestamp 1679581782
transform 1 0 89280 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_931
timestamp 1679581782
transform 1 0 89952 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_938
timestamp 1679581782
transform 1 0 90624 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_945
timestamp 1679581782
transform 1 0 91296 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_952
timestamp 1679581782
transform 1 0 91968 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_959
timestamp 1679581782
transform 1 0 92640 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_966
timestamp 1679581782
transform 1 0 93312 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_973
timestamp 1679581782
transform 1 0 93984 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_980
timestamp 1679581782
transform 1 0 94656 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_987
timestamp 1679581782
transform 1 0 95328 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_994
timestamp 1679581782
transform 1 0 96000 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_1001
timestamp 1679581782
transform 1 0 96672 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_1008
timestamp 1679581782
transform 1 0 97344 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_1015
timestamp 1679581782
transform 1 0 98016 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_1022
timestamp 1679581782
transform 1 0 98688 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_4
timestamp 1679581782
transform 1 0 960 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_11
timestamp 1679581782
transform 1 0 1632 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_18
timestamp 1679581782
transform 1 0 2304 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_25
timestamp 1679581782
transform 1 0 2976 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_32
timestamp 1679581782
transform 1 0 3648 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_39
timestamp 1679581782
transform 1 0 4320 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_46
timestamp 1679581782
transform 1 0 4992 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_53
timestamp 1679581782
transform 1 0 5664 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_60
timestamp 1679581782
transform 1 0 6336 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_67
timestamp 1679581782
transform 1 0 7008 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_74
timestamp 1679581782
transform 1 0 7680 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_81
timestamp 1679581782
transform 1 0 8352 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_88
timestamp 1679581782
transform 1 0 9024 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_95
timestamp 1679581782
transform 1 0 9696 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_102
timestamp 1679581782
transform 1 0 10368 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_109
timestamp 1679581782
transform 1 0 11040 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_116
timestamp 1679581782
transform 1 0 11712 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_123
timestamp 1679581782
transform 1 0 12384 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_130
timestamp 1679581782
transform 1 0 13056 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_137
timestamp 1679581782
transform 1 0 13728 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_144
timestamp 1679581782
transform 1 0 14400 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_151
timestamp 1679581782
transform 1 0 15072 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_158
timestamp 1679581782
transform 1 0 15744 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_165
timestamp 1679581782
transform 1 0 16416 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_172
timestamp 1679581782
transform 1 0 17088 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_179
timestamp 1679581782
transform 1 0 17760 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_186
timestamp 1679581782
transform 1 0 18432 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_193
timestamp 1679581782
transform 1 0 19104 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_200
timestamp 1679581782
transform 1 0 19776 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_207
timestamp 1679581782
transform 1 0 20448 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_214
timestamp 1679581782
transform 1 0 21120 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_221
timestamp 1679581782
transform 1 0 21792 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_228
timestamp 1679581782
transform 1 0 22464 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_235
timestamp 1679581782
transform 1 0 23136 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_242
timestamp 1679581782
transform 1 0 23808 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_249
timestamp 1679581782
transform 1 0 24480 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_256
timestamp 1679581782
transform 1 0 25152 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_263
timestamp 1679581782
transform 1 0 25824 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_270
timestamp 1679581782
transform 1 0 26496 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_277
timestamp 1679581782
transform 1 0 27168 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_284
timestamp 1679581782
transform 1 0 27840 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_291
timestamp 1679581782
transform 1 0 28512 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_298
timestamp 1679581782
transform 1 0 29184 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_305
timestamp 1679581782
transform 1 0 29856 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_312
timestamp 1679581782
transform 1 0 30528 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_319
timestamp 1679581782
transform 1 0 31200 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_326
timestamp 1679581782
transform 1 0 31872 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_333
timestamp 1679581782
transform 1 0 32544 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_340
timestamp 1679581782
transform 1 0 33216 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_347
timestamp 1679581782
transform 1 0 33888 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_354
timestamp 1679581782
transform 1 0 34560 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_361
timestamp 1679581782
transform 1 0 35232 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_368
timestamp 1679581782
transform 1 0 35904 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_375
timestamp 1679581782
transform 1 0 36576 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_382
timestamp 1679581782
transform 1 0 37248 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_389
timestamp 1679581782
transform 1 0 37920 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_396
timestamp 1679581782
transform 1 0 38592 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_403
timestamp 1679581782
transform 1 0 39264 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_410
timestamp 1679581782
transform 1 0 39936 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_417
timestamp 1679581782
transform 1 0 40608 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_424
timestamp 1679581782
transform 1 0 41280 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_431
timestamp 1679581782
transform 1 0 41952 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_438
timestamp 1679581782
transform 1 0 42624 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_445
timestamp 1679581782
transform 1 0 43296 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_452
timestamp 1679581782
transform 1 0 43968 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_459
timestamp 1679581782
transform 1 0 44640 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_466
timestamp 1679581782
transform 1 0 45312 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_473
timestamp 1679581782
transform 1 0 45984 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_480
timestamp 1679581782
transform 1 0 46656 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_487
timestamp 1679581782
transform 1 0 47328 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_494
timestamp 1679581782
transform 1 0 48000 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_501
timestamp 1679581782
transform 1 0 48672 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_508
timestamp 1679581782
transform 1 0 49344 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_515
timestamp 1679581782
transform 1 0 50016 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_522
timestamp 1679581782
transform 1 0 50688 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_529
timestamp 1679581782
transform 1 0 51360 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_536
timestamp 1679581782
transform 1 0 52032 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_543
timestamp 1679581782
transform 1 0 52704 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_550
timestamp 1679581782
transform 1 0 53376 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_557
timestamp 1679581782
transform 1 0 54048 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_564
timestamp 1679581782
transform 1 0 54720 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_571
timestamp 1679581782
transform 1 0 55392 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_578
timestamp 1679581782
transform 1 0 56064 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_585
timestamp 1679581782
transform 1 0 56736 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_592
timestamp 1679581782
transform 1 0 57408 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_599
timestamp 1679581782
transform 1 0 58080 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_606
timestamp 1679581782
transform 1 0 58752 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_613
timestamp 1679581782
transform 1 0 59424 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_620
timestamp 1679581782
transform 1 0 60096 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_627
timestamp 1679581782
transform 1 0 60768 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_634
timestamp 1679581782
transform 1 0 61440 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_641
timestamp 1679581782
transform 1 0 62112 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_648
timestamp 1679581782
transform 1 0 62784 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_655
timestamp 1679581782
transform 1 0 63456 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_662
timestamp 1679581782
transform 1 0 64128 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_669
timestamp 1679581782
transform 1 0 64800 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_676
timestamp 1679581782
transform 1 0 65472 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_683
timestamp 1679581782
transform 1 0 66144 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_690
timestamp 1679581782
transform 1 0 66816 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_697
timestamp 1679581782
transform 1 0 67488 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_704
timestamp 1679581782
transform 1 0 68160 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_711
timestamp 1679581782
transform 1 0 68832 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_718
timestamp 1679581782
transform 1 0 69504 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_725
timestamp 1679581782
transform 1 0 70176 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_732
timestamp 1679581782
transform 1 0 70848 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_739
timestamp 1679581782
transform 1 0 71520 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_746
timestamp 1679581782
transform 1 0 72192 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_753
timestamp 1679581782
transform 1 0 72864 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_760
timestamp 1679581782
transform 1 0 73536 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_767
timestamp 1679581782
transform 1 0 74208 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_774
timestamp 1679581782
transform 1 0 74880 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_781
timestamp 1679581782
transform 1 0 75552 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_788
timestamp 1679581782
transform 1 0 76224 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_795
timestamp 1679581782
transform 1 0 76896 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_802
timestamp 1679581782
transform 1 0 77568 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_809
timestamp 1679581782
transform 1 0 78240 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_816
timestamp 1679581782
transform 1 0 78912 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_823
timestamp 1679581782
transform 1 0 79584 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_830
timestamp 1679581782
transform 1 0 80256 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_837
timestamp 1679581782
transform 1 0 80928 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_844
timestamp 1679581782
transform 1 0 81600 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_851
timestamp 1679581782
transform 1 0 82272 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_858
timestamp 1679581782
transform 1 0 82944 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_865
timestamp 1679581782
transform 1 0 83616 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_872
timestamp 1679581782
transform 1 0 84288 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_879
timestamp 1679581782
transform 1 0 84960 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_886
timestamp 1679581782
transform 1 0 85632 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_893
timestamp 1679581782
transform 1 0 86304 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_900
timestamp 1679581782
transform 1 0 86976 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_907
timestamp 1679581782
transform 1 0 87648 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_914
timestamp 1679581782
transform 1 0 88320 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_921
timestamp 1679581782
transform 1 0 88992 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_928
timestamp 1679581782
transform 1 0 89664 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_935
timestamp 1679581782
transform 1 0 90336 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_942
timestamp 1679581782
transform 1 0 91008 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_949
timestamp 1679581782
transform 1 0 91680 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_956
timestamp 1679581782
transform 1 0 92352 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_963
timestamp 1679581782
transform 1 0 93024 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_970
timestamp 1679581782
transform 1 0 93696 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_977
timestamp 1679581782
transform 1 0 94368 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_984
timestamp 1679581782
transform 1 0 95040 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_991
timestamp 1679581782
transform 1 0 95712 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_998
timestamp 1679581782
transform 1 0 96384 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_1005
timestamp 1679581782
transform 1 0 97056 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_1012
timestamp 1679581782
transform 1 0 97728 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_1019
timestamp 1679581782
transform 1 0 98400 0 1 65772
box -48 -56 720 834
use sg13g2_fill_2  FILLER_86_1026
timestamp 1677580104
transform 1 0 99072 0 1 65772
box -48 -56 240 834
use sg13g2_fill_1  FILLER_86_1028
timestamp 1677579658
transform 1 0 99264 0 1 65772
box -48 -56 144 834
use sg13g2_decap_8  FILLER_87_0
timestamp 1679581782
transform 1 0 576 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_7
timestamp 1679581782
transform 1 0 1248 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_14
timestamp 1679581782
transform 1 0 1920 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_21
timestamp 1679581782
transform 1 0 2592 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_28
timestamp 1679581782
transform 1 0 3264 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_35
timestamp 1679581782
transform 1 0 3936 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_42
timestamp 1679581782
transform 1 0 4608 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_49
timestamp 1679581782
transform 1 0 5280 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_56
timestamp 1679581782
transform 1 0 5952 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_63
timestamp 1679581782
transform 1 0 6624 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_70
timestamp 1679581782
transform 1 0 7296 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_77
timestamp 1679581782
transform 1 0 7968 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_84
timestamp 1679581782
transform 1 0 8640 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_91
timestamp 1679581782
transform 1 0 9312 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_98
timestamp 1679581782
transform 1 0 9984 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_105
timestamp 1679581782
transform 1 0 10656 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_112
timestamp 1679581782
transform 1 0 11328 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_119
timestamp 1679581782
transform 1 0 12000 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_126
timestamp 1679581782
transform 1 0 12672 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_133
timestamp 1679581782
transform 1 0 13344 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_140
timestamp 1679581782
transform 1 0 14016 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_147
timestamp 1679581782
transform 1 0 14688 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_154
timestamp 1679581782
transform 1 0 15360 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_161
timestamp 1679581782
transform 1 0 16032 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_168
timestamp 1679581782
transform 1 0 16704 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_175
timestamp 1679581782
transform 1 0 17376 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_182
timestamp 1679581782
transform 1 0 18048 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_189
timestamp 1679581782
transform 1 0 18720 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_196
timestamp 1679581782
transform 1 0 19392 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_203
timestamp 1679581782
transform 1 0 20064 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_210
timestamp 1679581782
transform 1 0 20736 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_217
timestamp 1679581782
transform 1 0 21408 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_224
timestamp 1679581782
transform 1 0 22080 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_231
timestamp 1679581782
transform 1 0 22752 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_238
timestamp 1679581782
transform 1 0 23424 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_245
timestamp 1679581782
transform 1 0 24096 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_252
timestamp 1679581782
transform 1 0 24768 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_259
timestamp 1679581782
transform 1 0 25440 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_266
timestamp 1679581782
transform 1 0 26112 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_273
timestamp 1679581782
transform 1 0 26784 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_280
timestamp 1679581782
transform 1 0 27456 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_287
timestamp 1679581782
transform 1 0 28128 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_294
timestamp 1679581782
transform 1 0 28800 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_301
timestamp 1679581782
transform 1 0 29472 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_308
timestamp 1679581782
transform 1 0 30144 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_315
timestamp 1679581782
transform 1 0 30816 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_322
timestamp 1679581782
transform 1 0 31488 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_329
timestamp 1679581782
transform 1 0 32160 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_336
timestamp 1679581782
transform 1 0 32832 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_343
timestamp 1679581782
transform 1 0 33504 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_350
timestamp 1679581782
transform 1 0 34176 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_357
timestamp 1679581782
transform 1 0 34848 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_364
timestamp 1679581782
transform 1 0 35520 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_371
timestamp 1679581782
transform 1 0 36192 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_378
timestamp 1679581782
transform 1 0 36864 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_385
timestamp 1679581782
transform 1 0 37536 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_392
timestamp 1679581782
transform 1 0 38208 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_399
timestamp 1679581782
transform 1 0 38880 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_406
timestamp 1679581782
transform 1 0 39552 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_413
timestamp 1679581782
transform 1 0 40224 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_420
timestamp 1679581782
transform 1 0 40896 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_427
timestamp 1679581782
transform 1 0 41568 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_434
timestamp 1679581782
transform 1 0 42240 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_441
timestamp 1679581782
transform 1 0 42912 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_448
timestamp 1679581782
transform 1 0 43584 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_455
timestamp 1679581782
transform 1 0 44256 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_462
timestamp 1679581782
transform 1 0 44928 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_469
timestamp 1679581782
transform 1 0 45600 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_476
timestamp 1679581782
transform 1 0 46272 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_483
timestamp 1679581782
transform 1 0 46944 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_490
timestamp 1679581782
transform 1 0 47616 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_497
timestamp 1679581782
transform 1 0 48288 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_504
timestamp 1679581782
transform 1 0 48960 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_511
timestamp 1679581782
transform 1 0 49632 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_518
timestamp 1679581782
transform 1 0 50304 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_525
timestamp 1679581782
transform 1 0 50976 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_532
timestamp 1679581782
transform 1 0 51648 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_539
timestamp 1679581782
transform 1 0 52320 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_546
timestamp 1679581782
transform 1 0 52992 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_553
timestamp 1679581782
transform 1 0 53664 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_560
timestamp 1679581782
transform 1 0 54336 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_567
timestamp 1679581782
transform 1 0 55008 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_574
timestamp 1679581782
transform 1 0 55680 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_581
timestamp 1679581782
transform 1 0 56352 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_588
timestamp 1679581782
transform 1 0 57024 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_595
timestamp 1679581782
transform 1 0 57696 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_602
timestamp 1679581782
transform 1 0 58368 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_609
timestamp 1679581782
transform 1 0 59040 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_616
timestamp 1679581782
transform 1 0 59712 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_623
timestamp 1679581782
transform 1 0 60384 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_630
timestamp 1679581782
transform 1 0 61056 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_637
timestamp 1679581782
transform 1 0 61728 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_644
timestamp 1679581782
transform 1 0 62400 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_651
timestamp 1679581782
transform 1 0 63072 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_658
timestamp 1679581782
transform 1 0 63744 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_665
timestamp 1679581782
transform 1 0 64416 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_672
timestamp 1679581782
transform 1 0 65088 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_679
timestamp 1679581782
transform 1 0 65760 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_686
timestamp 1679581782
transform 1 0 66432 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_693
timestamp 1679581782
transform 1 0 67104 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_700
timestamp 1679581782
transform 1 0 67776 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_707
timestamp 1679581782
transform 1 0 68448 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_714
timestamp 1679581782
transform 1 0 69120 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_721
timestamp 1679581782
transform 1 0 69792 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_728
timestamp 1679581782
transform 1 0 70464 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_735
timestamp 1679581782
transform 1 0 71136 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_742
timestamp 1679581782
transform 1 0 71808 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_749
timestamp 1679581782
transform 1 0 72480 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_756
timestamp 1679581782
transform 1 0 73152 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_763
timestamp 1679581782
transform 1 0 73824 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_770
timestamp 1679581782
transform 1 0 74496 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_777
timestamp 1679581782
transform 1 0 75168 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_784
timestamp 1679581782
transform 1 0 75840 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_791
timestamp 1679581782
transform 1 0 76512 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_798
timestamp 1679581782
transform 1 0 77184 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_805
timestamp 1679581782
transform 1 0 77856 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_812
timestamp 1679581782
transform 1 0 78528 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_819
timestamp 1679581782
transform 1 0 79200 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_826
timestamp 1679581782
transform 1 0 79872 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_833
timestamp 1679581782
transform 1 0 80544 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_840
timestamp 1679581782
transform 1 0 81216 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_847
timestamp 1679581782
transform 1 0 81888 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_854
timestamp 1679581782
transform 1 0 82560 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_861
timestamp 1679581782
transform 1 0 83232 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_868
timestamp 1679581782
transform 1 0 83904 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_875
timestamp 1679581782
transform 1 0 84576 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_882
timestamp 1679581782
transform 1 0 85248 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_889
timestamp 1679581782
transform 1 0 85920 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_896
timestamp 1679581782
transform 1 0 86592 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_903
timestamp 1679581782
transform 1 0 87264 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_910
timestamp 1679581782
transform 1 0 87936 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_917
timestamp 1679581782
transform 1 0 88608 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_924
timestamp 1679581782
transform 1 0 89280 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_931
timestamp 1679581782
transform 1 0 89952 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_938
timestamp 1679581782
transform 1 0 90624 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_945
timestamp 1679581782
transform 1 0 91296 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_952
timestamp 1679581782
transform 1 0 91968 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_959
timestamp 1679581782
transform 1 0 92640 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_966
timestamp 1679581782
transform 1 0 93312 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_973
timestamp 1679581782
transform 1 0 93984 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_980
timestamp 1679581782
transform 1 0 94656 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_987
timestamp 1679581782
transform 1 0 95328 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_994
timestamp 1679581782
transform 1 0 96000 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_1001
timestamp 1679581782
transform 1 0 96672 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_1008
timestamp 1679581782
transform 1 0 97344 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_1015
timestamp 1679581782
transform 1 0 98016 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_1022
timestamp 1679581782
transform 1 0 98688 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_4
timestamp 1679581782
transform 1 0 960 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_11
timestamp 1679581782
transform 1 0 1632 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_18
timestamp 1679581782
transform 1 0 2304 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_25
timestamp 1679581782
transform 1 0 2976 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_32
timestamp 1679581782
transform 1 0 3648 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_39
timestamp 1679581782
transform 1 0 4320 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_46
timestamp 1679581782
transform 1 0 4992 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_53
timestamp 1679581782
transform 1 0 5664 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_60
timestamp 1679581782
transform 1 0 6336 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_67
timestamp 1679581782
transform 1 0 7008 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_74
timestamp 1679581782
transform 1 0 7680 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_81
timestamp 1679581782
transform 1 0 8352 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_88
timestamp 1679581782
transform 1 0 9024 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_95
timestamp 1679581782
transform 1 0 9696 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_102
timestamp 1679581782
transform 1 0 10368 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_109
timestamp 1679581782
transform 1 0 11040 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_116
timestamp 1679581782
transform 1 0 11712 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_123
timestamp 1679581782
transform 1 0 12384 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_130
timestamp 1679581782
transform 1 0 13056 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_137
timestamp 1679581782
transform 1 0 13728 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_144
timestamp 1679581782
transform 1 0 14400 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_151
timestamp 1679581782
transform 1 0 15072 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_158
timestamp 1679581782
transform 1 0 15744 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_165
timestamp 1679581782
transform 1 0 16416 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_172
timestamp 1679581782
transform 1 0 17088 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_179
timestamp 1679581782
transform 1 0 17760 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_186
timestamp 1679581782
transform 1 0 18432 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_193
timestamp 1679581782
transform 1 0 19104 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_200
timestamp 1679581782
transform 1 0 19776 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_207
timestamp 1679581782
transform 1 0 20448 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_214
timestamp 1679581782
transform 1 0 21120 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_221
timestamp 1679581782
transform 1 0 21792 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_228
timestamp 1679581782
transform 1 0 22464 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_235
timestamp 1679581782
transform 1 0 23136 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_242
timestamp 1679581782
transform 1 0 23808 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_249
timestamp 1679581782
transform 1 0 24480 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_256
timestamp 1679581782
transform 1 0 25152 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_263
timestamp 1679581782
transform 1 0 25824 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_270
timestamp 1679581782
transform 1 0 26496 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_277
timestamp 1679581782
transform 1 0 27168 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_284
timestamp 1679581782
transform 1 0 27840 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_291
timestamp 1679581782
transform 1 0 28512 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_298
timestamp 1679581782
transform 1 0 29184 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_305
timestamp 1679581782
transform 1 0 29856 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_312
timestamp 1679581782
transform 1 0 30528 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_319
timestamp 1679581782
transform 1 0 31200 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_326
timestamp 1679581782
transform 1 0 31872 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_333
timestamp 1679581782
transform 1 0 32544 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_340
timestamp 1679581782
transform 1 0 33216 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_347
timestamp 1679581782
transform 1 0 33888 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_354
timestamp 1679581782
transform 1 0 34560 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_361
timestamp 1679581782
transform 1 0 35232 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_368
timestamp 1679581782
transform 1 0 35904 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_375
timestamp 1679581782
transform 1 0 36576 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_382
timestamp 1679581782
transform 1 0 37248 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_389
timestamp 1679581782
transform 1 0 37920 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_396
timestamp 1679581782
transform 1 0 38592 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_403
timestamp 1679581782
transform 1 0 39264 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_410
timestamp 1679581782
transform 1 0 39936 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_417
timestamp 1679581782
transform 1 0 40608 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_424
timestamp 1679581782
transform 1 0 41280 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_431
timestamp 1679581782
transform 1 0 41952 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_438
timestamp 1679581782
transform 1 0 42624 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_445
timestamp 1679581782
transform 1 0 43296 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_452
timestamp 1679581782
transform 1 0 43968 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_459
timestamp 1679581782
transform 1 0 44640 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_466
timestamp 1679581782
transform 1 0 45312 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_473
timestamp 1679581782
transform 1 0 45984 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_480
timestamp 1679581782
transform 1 0 46656 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_487
timestamp 1679581782
transform 1 0 47328 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_494
timestamp 1679581782
transform 1 0 48000 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_501
timestamp 1679581782
transform 1 0 48672 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_508
timestamp 1679581782
transform 1 0 49344 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_515
timestamp 1679581782
transform 1 0 50016 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_522
timestamp 1679581782
transform 1 0 50688 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_529
timestamp 1679581782
transform 1 0 51360 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_536
timestamp 1679581782
transform 1 0 52032 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_543
timestamp 1679581782
transform 1 0 52704 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_550
timestamp 1679581782
transform 1 0 53376 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_557
timestamp 1679581782
transform 1 0 54048 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_564
timestamp 1679581782
transform 1 0 54720 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_571
timestamp 1679581782
transform 1 0 55392 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_578
timestamp 1679581782
transform 1 0 56064 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_585
timestamp 1679581782
transform 1 0 56736 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_592
timestamp 1679581782
transform 1 0 57408 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_599
timestamp 1679581782
transform 1 0 58080 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_606
timestamp 1679581782
transform 1 0 58752 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_613
timestamp 1679581782
transform 1 0 59424 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_620
timestamp 1679581782
transform 1 0 60096 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_627
timestamp 1679581782
transform 1 0 60768 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_634
timestamp 1679581782
transform 1 0 61440 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_641
timestamp 1679581782
transform 1 0 62112 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_648
timestamp 1679581782
transform 1 0 62784 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_655
timestamp 1679581782
transform 1 0 63456 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_662
timestamp 1679581782
transform 1 0 64128 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_669
timestamp 1679581782
transform 1 0 64800 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_676
timestamp 1679581782
transform 1 0 65472 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_683
timestamp 1679581782
transform 1 0 66144 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_690
timestamp 1679581782
transform 1 0 66816 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_697
timestamp 1679581782
transform 1 0 67488 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_704
timestamp 1679581782
transform 1 0 68160 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_711
timestamp 1679581782
transform 1 0 68832 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_718
timestamp 1679581782
transform 1 0 69504 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_725
timestamp 1679581782
transform 1 0 70176 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_732
timestamp 1679581782
transform 1 0 70848 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_739
timestamp 1679581782
transform 1 0 71520 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_746
timestamp 1679581782
transform 1 0 72192 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_753
timestamp 1679581782
transform 1 0 72864 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_760
timestamp 1679581782
transform 1 0 73536 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_767
timestamp 1679581782
transform 1 0 74208 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_774
timestamp 1679581782
transform 1 0 74880 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_781
timestamp 1679581782
transform 1 0 75552 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_788
timestamp 1679581782
transform 1 0 76224 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_795
timestamp 1679581782
transform 1 0 76896 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_802
timestamp 1679581782
transform 1 0 77568 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_809
timestamp 1679581782
transform 1 0 78240 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_816
timestamp 1679581782
transform 1 0 78912 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_823
timestamp 1679581782
transform 1 0 79584 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_830
timestamp 1679581782
transform 1 0 80256 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_837
timestamp 1679581782
transform 1 0 80928 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_844
timestamp 1679581782
transform 1 0 81600 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_851
timestamp 1679581782
transform 1 0 82272 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_858
timestamp 1679581782
transform 1 0 82944 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_865
timestamp 1679581782
transform 1 0 83616 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_872
timestamp 1679581782
transform 1 0 84288 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_879
timestamp 1679581782
transform 1 0 84960 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_886
timestamp 1679581782
transform 1 0 85632 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_893
timestamp 1679581782
transform 1 0 86304 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_900
timestamp 1679581782
transform 1 0 86976 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_907
timestamp 1679581782
transform 1 0 87648 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_914
timestamp 1679581782
transform 1 0 88320 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_921
timestamp 1679581782
transform 1 0 88992 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_928
timestamp 1679581782
transform 1 0 89664 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_935
timestamp 1679581782
transform 1 0 90336 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_942
timestamp 1679581782
transform 1 0 91008 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_949
timestamp 1679581782
transform 1 0 91680 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_956
timestamp 1679581782
transform 1 0 92352 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_963
timestamp 1679581782
transform 1 0 93024 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_970
timestamp 1679581782
transform 1 0 93696 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_977
timestamp 1679581782
transform 1 0 94368 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_984
timestamp 1679581782
transform 1 0 95040 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_991
timestamp 1679581782
transform 1 0 95712 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_998
timestamp 1679581782
transform 1 0 96384 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_1005
timestamp 1679581782
transform 1 0 97056 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_1012
timestamp 1679581782
transform 1 0 97728 0 1 67284
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_1019
timestamp 1679581782
transform 1 0 98400 0 1 67284
box -48 -56 720 834
use sg13g2_fill_2  FILLER_88_1026
timestamp 1677580104
transform 1 0 99072 0 1 67284
box -48 -56 240 834
use sg13g2_fill_1  FILLER_88_1028
timestamp 1677579658
transform 1 0 99264 0 1 67284
box -48 -56 144 834
use sg13g2_decap_8  FILLER_89_0
timestamp 1679581782
transform 1 0 576 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_7
timestamp 1679581782
transform 1 0 1248 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_14
timestamp 1679581782
transform 1 0 1920 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_21
timestamp 1679581782
transform 1 0 2592 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_28
timestamp 1679581782
transform 1 0 3264 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_35
timestamp 1679581782
transform 1 0 3936 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_42
timestamp 1679581782
transform 1 0 4608 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_49
timestamp 1679581782
transform 1 0 5280 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_56
timestamp 1679581782
transform 1 0 5952 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_63
timestamp 1679581782
transform 1 0 6624 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_70
timestamp 1679581782
transform 1 0 7296 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_77
timestamp 1679581782
transform 1 0 7968 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_84
timestamp 1679581782
transform 1 0 8640 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_91
timestamp 1679581782
transform 1 0 9312 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_98
timestamp 1679581782
transform 1 0 9984 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_105
timestamp 1679581782
transform 1 0 10656 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_112
timestamp 1679581782
transform 1 0 11328 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_119
timestamp 1679581782
transform 1 0 12000 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_126
timestamp 1679581782
transform 1 0 12672 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_133
timestamp 1679581782
transform 1 0 13344 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_140
timestamp 1679581782
transform 1 0 14016 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_147
timestamp 1679581782
transform 1 0 14688 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_154
timestamp 1679581782
transform 1 0 15360 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_161
timestamp 1679581782
transform 1 0 16032 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_168
timestamp 1679581782
transform 1 0 16704 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_175
timestamp 1679581782
transform 1 0 17376 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_182
timestamp 1679581782
transform 1 0 18048 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_189
timestamp 1679581782
transform 1 0 18720 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_196
timestamp 1679581782
transform 1 0 19392 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_203
timestamp 1679581782
transform 1 0 20064 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_210
timestamp 1679581782
transform 1 0 20736 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_217
timestamp 1679581782
transform 1 0 21408 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_224
timestamp 1679581782
transform 1 0 22080 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_231
timestamp 1679581782
transform 1 0 22752 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_238
timestamp 1679581782
transform 1 0 23424 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_245
timestamp 1679581782
transform 1 0 24096 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_252
timestamp 1679581782
transform 1 0 24768 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_259
timestamp 1679581782
transform 1 0 25440 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_266
timestamp 1679581782
transform 1 0 26112 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_273
timestamp 1679581782
transform 1 0 26784 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_280
timestamp 1679581782
transform 1 0 27456 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_287
timestamp 1679581782
transform 1 0 28128 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_294
timestamp 1679581782
transform 1 0 28800 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_301
timestamp 1679581782
transform 1 0 29472 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_308
timestamp 1679581782
transform 1 0 30144 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_315
timestamp 1679581782
transform 1 0 30816 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_322
timestamp 1679581782
transform 1 0 31488 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_329
timestamp 1679581782
transform 1 0 32160 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_336
timestamp 1679581782
transform 1 0 32832 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_343
timestamp 1679581782
transform 1 0 33504 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_350
timestamp 1679581782
transform 1 0 34176 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_357
timestamp 1679581782
transform 1 0 34848 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_364
timestamp 1679581782
transform 1 0 35520 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_371
timestamp 1679581782
transform 1 0 36192 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_378
timestamp 1679581782
transform 1 0 36864 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_385
timestamp 1679581782
transform 1 0 37536 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_392
timestamp 1679581782
transform 1 0 38208 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_399
timestamp 1679581782
transform 1 0 38880 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_406
timestamp 1679581782
transform 1 0 39552 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_413
timestamp 1679581782
transform 1 0 40224 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_420
timestamp 1679581782
transform 1 0 40896 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_427
timestamp 1679581782
transform 1 0 41568 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_434
timestamp 1679581782
transform 1 0 42240 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_441
timestamp 1679581782
transform 1 0 42912 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_448
timestamp 1679581782
transform 1 0 43584 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_455
timestamp 1679581782
transform 1 0 44256 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_462
timestamp 1679581782
transform 1 0 44928 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_469
timestamp 1679581782
transform 1 0 45600 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_476
timestamp 1679581782
transform 1 0 46272 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_483
timestamp 1679581782
transform 1 0 46944 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_490
timestamp 1679581782
transform 1 0 47616 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_497
timestamp 1679581782
transform 1 0 48288 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_504
timestamp 1679581782
transform 1 0 48960 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_511
timestamp 1679581782
transform 1 0 49632 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_518
timestamp 1679581782
transform 1 0 50304 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_525
timestamp 1679581782
transform 1 0 50976 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_532
timestamp 1679581782
transform 1 0 51648 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_539
timestamp 1679581782
transform 1 0 52320 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_546
timestamp 1679581782
transform 1 0 52992 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_553
timestamp 1679581782
transform 1 0 53664 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_560
timestamp 1679581782
transform 1 0 54336 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_567
timestamp 1679581782
transform 1 0 55008 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_574
timestamp 1679581782
transform 1 0 55680 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_581
timestamp 1679581782
transform 1 0 56352 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_588
timestamp 1679581782
transform 1 0 57024 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_595
timestamp 1679581782
transform 1 0 57696 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_602
timestamp 1679581782
transform 1 0 58368 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_609
timestamp 1679581782
transform 1 0 59040 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_616
timestamp 1679581782
transform 1 0 59712 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_623
timestamp 1679581782
transform 1 0 60384 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_630
timestamp 1679581782
transform 1 0 61056 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_637
timestamp 1679581782
transform 1 0 61728 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_644
timestamp 1679581782
transform 1 0 62400 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_651
timestamp 1679581782
transform 1 0 63072 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_658
timestamp 1679581782
transform 1 0 63744 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_665
timestamp 1679581782
transform 1 0 64416 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_672
timestamp 1679581782
transform 1 0 65088 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_679
timestamp 1679581782
transform 1 0 65760 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_686
timestamp 1679581782
transform 1 0 66432 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_693
timestamp 1679581782
transform 1 0 67104 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_700
timestamp 1679581782
transform 1 0 67776 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_707
timestamp 1679581782
transform 1 0 68448 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_714
timestamp 1679581782
transform 1 0 69120 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_721
timestamp 1679581782
transform 1 0 69792 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_728
timestamp 1679581782
transform 1 0 70464 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_735
timestamp 1679581782
transform 1 0 71136 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_742
timestamp 1679581782
transform 1 0 71808 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_749
timestamp 1679581782
transform 1 0 72480 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_756
timestamp 1679581782
transform 1 0 73152 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_763
timestamp 1679581782
transform 1 0 73824 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_770
timestamp 1679581782
transform 1 0 74496 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_777
timestamp 1679581782
transform 1 0 75168 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_784
timestamp 1679581782
transform 1 0 75840 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_791
timestamp 1679581782
transform 1 0 76512 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_798
timestamp 1679581782
transform 1 0 77184 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_805
timestamp 1679581782
transform 1 0 77856 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_812
timestamp 1679581782
transform 1 0 78528 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_819
timestamp 1679581782
transform 1 0 79200 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_826
timestamp 1679581782
transform 1 0 79872 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_833
timestamp 1679581782
transform 1 0 80544 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_840
timestamp 1679581782
transform 1 0 81216 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_847
timestamp 1679581782
transform 1 0 81888 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_854
timestamp 1679581782
transform 1 0 82560 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_861
timestamp 1679581782
transform 1 0 83232 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_868
timestamp 1679581782
transform 1 0 83904 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_875
timestamp 1679581782
transform 1 0 84576 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_882
timestamp 1679581782
transform 1 0 85248 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_889
timestamp 1679581782
transform 1 0 85920 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_896
timestamp 1679581782
transform 1 0 86592 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_903
timestamp 1679581782
transform 1 0 87264 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_910
timestamp 1679581782
transform 1 0 87936 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_917
timestamp 1679581782
transform 1 0 88608 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_924
timestamp 1679581782
transform 1 0 89280 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_931
timestamp 1679581782
transform 1 0 89952 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_938
timestamp 1679581782
transform 1 0 90624 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_945
timestamp 1679581782
transform 1 0 91296 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_952
timestamp 1679581782
transform 1 0 91968 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_959
timestamp 1679581782
transform 1 0 92640 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_966
timestamp 1679581782
transform 1 0 93312 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_973
timestamp 1679581782
transform 1 0 93984 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_980
timestamp 1679581782
transform 1 0 94656 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_987
timestamp 1679581782
transform 1 0 95328 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_994
timestamp 1679581782
transform 1 0 96000 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_1001
timestamp 1679581782
transform 1 0 96672 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_1008
timestamp 1679581782
transform 1 0 97344 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_1015
timestamp 1679581782
transform 1 0 98016 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_1022
timestamp 1679581782
transform 1 0 98688 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_4
timestamp 1679581782
transform 1 0 960 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_11
timestamp 1679581782
transform 1 0 1632 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_18
timestamp 1679581782
transform 1 0 2304 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_25
timestamp 1679581782
transform 1 0 2976 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_32
timestamp 1679581782
transform 1 0 3648 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_39
timestamp 1679581782
transform 1 0 4320 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_46
timestamp 1679581782
transform 1 0 4992 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_53
timestamp 1679581782
transform 1 0 5664 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_60
timestamp 1679581782
transform 1 0 6336 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_67
timestamp 1679581782
transform 1 0 7008 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_74
timestamp 1679581782
transform 1 0 7680 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_81
timestamp 1679581782
transform 1 0 8352 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_88
timestamp 1679581782
transform 1 0 9024 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_95
timestamp 1679581782
transform 1 0 9696 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_102
timestamp 1679581782
transform 1 0 10368 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_109
timestamp 1679581782
transform 1 0 11040 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_116
timestamp 1679581782
transform 1 0 11712 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_123
timestamp 1679581782
transform 1 0 12384 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_130
timestamp 1679581782
transform 1 0 13056 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_137
timestamp 1679581782
transform 1 0 13728 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_144
timestamp 1679581782
transform 1 0 14400 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_151
timestamp 1679581782
transform 1 0 15072 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_158
timestamp 1679581782
transform 1 0 15744 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_165
timestamp 1679581782
transform 1 0 16416 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_172
timestamp 1679581782
transform 1 0 17088 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_179
timestamp 1679581782
transform 1 0 17760 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_186
timestamp 1679581782
transform 1 0 18432 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_193
timestamp 1679581782
transform 1 0 19104 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_200
timestamp 1679581782
transform 1 0 19776 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_207
timestamp 1679581782
transform 1 0 20448 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_214
timestamp 1679581782
transform 1 0 21120 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_221
timestamp 1679581782
transform 1 0 21792 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_228
timestamp 1679581782
transform 1 0 22464 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_235
timestamp 1679581782
transform 1 0 23136 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_242
timestamp 1679581782
transform 1 0 23808 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_249
timestamp 1679581782
transform 1 0 24480 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_256
timestamp 1679581782
transform 1 0 25152 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_263
timestamp 1679581782
transform 1 0 25824 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_270
timestamp 1679581782
transform 1 0 26496 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_277
timestamp 1679581782
transform 1 0 27168 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_284
timestamp 1679581782
transform 1 0 27840 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_291
timestamp 1679581782
transform 1 0 28512 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_298
timestamp 1679581782
transform 1 0 29184 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_305
timestamp 1679581782
transform 1 0 29856 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_312
timestamp 1679581782
transform 1 0 30528 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_319
timestamp 1679581782
transform 1 0 31200 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_326
timestamp 1679581782
transform 1 0 31872 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_333
timestamp 1679581782
transform 1 0 32544 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_340
timestamp 1679581782
transform 1 0 33216 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_347
timestamp 1679581782
transform 1 0 33888 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_354
timestamp 1679581782
transform 1 0 34560 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_361
timestamp 1679581782
transform 1 0 35232 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_368
timestamp 1679581782
transform 1 0 35904 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_375
timestamp 1679581782
transform 1 0 36576 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_382
timestamp 1679581782
transform 1 0 37248 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_389
timestamp 1679581782
transform 1 0 37920 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_396
timestamp 1679581782
transform 1 0 38592 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_403
timestamp 1679581782
transform 1 0 39264 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_410
timestamp 1679581782
transform 1 0 39936 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_417
timestamp 1679581782
transform 1 0 40608 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_424
timestamp 1679581782
transform 1 0 41280 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_431
timestamp 1679581782
transform 1 0 41952 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_438
timestamp 1679581782
transform 1 0 42624 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_445
timestamp 1679581782
transform 1 0 43296 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_452
timestamp 1679581782
transform 1 0 43968 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_459
timestamp 1679581782
transform 1 0 44640 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_466
timestamp 1679581782
transform 1 0 45312 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_473
timestamp 1679581782
transform 1 0 45984 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_480
timestamp 1679581782
transform 1 0 46656 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_487
timestamp 1679581782
transform 1 0 47328 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_494
timestamp 1679581782
transform 1 0 48000 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_501
timestamp 1679581782
transform 1 0 48672 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_508
timestamp 1679581782
transform 1 0 49344 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_515
timestamp 1679581782
transform 1 0 50016 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_522
timestamp 1679581782
transform 1 0 50688 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_529
timestamp 1679581782
transform 1 0 51360 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_536
timestamp 1679581782
transform 1 0 52032 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_543
timestamp 1679581782
transform 1 0 52704 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_550
timestamp 1679581782
transform 1 0 53376 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_557
timestamp 1679581782
transform 1 0 54048 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_564
timestamp 1679581782
transform 1 0 54720 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_571
timestamp 1679581782
transform 1 0 55392 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_578
timestamp 1679581782
transform 1 0 56064 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_585
timestamp 1679581782
transform 1 0 56736 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_592
timestamp 1679581782
transform 1 0 57408 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_599
timestamp 1679581782
transform 1 0 58080 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_606
timestamp 1679581782
transform 1 0 58752 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_613
timestamp 1679581782
transform 1 0 59424 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_620
timestamp 1679581782
transform 1 0 60096 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_627
timestamp 1679581782
transform 1 0 60768 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_634
timestamp 1679581782
transform 1 0 61440 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_641
timestamp 1679581782
transform 1 0 62112 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_648
timestamp 1679581782
transform 1 0 62784 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_655
timestamp 1679581782
transform 1 0 63456 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_662
timestamp 1679581782
transform 1 0 64128 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_669
timestamp 1679581782
transform 1 0 64800 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_676
timestamp 1679581782
transform 1 0 65472 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_683
timestamp 1679581782
transform 1 0 66144 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_690
timestamp 1679581782
transform 1 0 66816 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_697
timestamp 1679581782
transform 1 0 67488 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_704
timestamp 1679581782
transform 1 0 68160 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_711
timestamp 1679581782
transform 1 0 68832 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_718
timestamp 1679581782
transform 1 0 69504 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_725
timestamp 1679581782
transform 1 0 70176 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_732
timestamp 1679581782
transform 1 0 70848 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_739
timestamp 1679581782
transform 1 0 71520 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_746
timestamp 1679581782
transform 1 0 72192 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_753
timestamp 1679581782
transform 1 0 72864 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_760
timestamp 1679581782
transform 1 0 73536 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_767
timestamp 1679581782
transform 1 0 74208 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_774
timestamp 1679581782
transform 1 0 74880 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_781
timestamp 1679581782
transform 1 0 75552 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_788
timestamp 1679581782
transform 1 0 76224 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_795
timestamp 1679581782
transform 1 0 76896 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_802
timestamp 1679581782
transform 1 0 77568 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_809
timestamp 1679581782
transform 1 0 78240 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_816
timestamp 1679581782
transform 1 0 78912 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_823
timestamp 1679581782
transform 1 0 79584 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_830
timestamp 1679581782
transform 1 0 80256 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_837
timestamp 1679581782
transform 1 0 80928 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_844
timestamp 1679581782
transform 1 0 81600 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_851
timestamp 1679581782
transform 1 0 82272 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_858
timestamp 1679581782
transform 1 0 82944 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_865
timestamp 1679581782
transform 1 0 83616 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_872
timestamp 1679581782
transform 1 0 84288 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_879
timestamp 1679581782
transform 1 0 84960 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_886
timestamp 1679581782
transform 1 0 85632 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_893
timestamp 1679581782
transform 1 0 86304 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_900
timestamp 1679581782
transform 1 0 86976 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_907
timestamp 1679581782
transform 1 0 87648 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_914
timestamp 1679581782
transform 1 0 88320 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_921
timestamp 1679581782
transform 1 0 88992 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_928
timestamp 1679581782
transform 1 0 89664 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_935
timestamp 1679581782
transform 1 0 90336 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_942
timestamp 1679581782
transform 1 0 91008 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_949
timestamp 1679581782
transform 1 0 91680 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_956
timestamp 1679581782
transform 1 0 92352 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_963
timestamp 1679581782
transform 1 0 93024 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_970
timestamp 1679581782
transform 1 0 93696 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_977
timestamp 1679581782
transform 1 0 94368 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_984
timestamp 1679581782
transform 1 0 95040 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_991
timestamp 1679581782
transform 1 0 95712 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_998
timestamp 1679581782
transform 1 0 96384 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_1005
timestamp 1679581782
transform 1 0 97056 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_1012
timestamp 1679581782
transform 1 0 97728 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_1019
timestamp 1679581782
transform 1 0 98400 0 1 68796
box -48 -56 720 834
use sg13g2_fill_2  FILLER_90_1026
timestamp 1677580104
transform 1 0 99072 0 1 68796
box -48 -56 240 834
use sg13g2_fill_1  FILLER_90_1028
timestamp 1677579658
transform 1 0 99264 0 1 68796
box -48 -56 144 834
use sg13g2_decap_8  FILLER_91_0
timestamp 1679581782
transform 1 0 576 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_7
timestamp 1679581782
transform 1 0 1248 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_14
timestamp 1679581782
transform 1 0 1920 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_21
timestamp 1679581782
transform 1 0 2592 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_28
timestamp 1679581782
transform 1 0 3264 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_35
timestamp 1679581782
transform 1 0 3936 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_42
timestamp 1679581782
transform 1 0 4608 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_49
timestamp 1679581782
transform 1 0 5280 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_56
timestamp 1679581782
transform 1 0 5952 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_63
timestamp 1679581782
transform 1 0 6624 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_70
timestamp 1679581782
transform 1 0 7296 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_77
timestamp 1679581782
transform 1 0 7968 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_84
timestamp 1679581782
transform 1 0 8640 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_91
timestamp 1679581782
transform 1 0 9312 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_98
timestamp 1679581782
transform 1 0 9984 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_105
timestamp 1679581782
transform 1 0 10656 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_112
timestamp 1679581782
transform 1 0 11328 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_119
timestamp 1679581782
transform 1 0 12000 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_126
timestamp 1679581782
transform 1 0 12672 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_133
timestamp 1679581782
transform 1 0 13344 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_140
timestamp 1679581782
transform 1 0 14016 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_147
timestamp 1679581782
transform 1 0 14688 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_154
timestamp 1679581782
transform 1 0 15360 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_161
timestamp 1679581782
transform 1 0 16032 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_168
timestamp 1679581782
transform 1 0 16704 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_175
timestamp 1679581782
transform 1 0 17376 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_182
timestamp 1679581782
transform 1 0 18048 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_189
timestamp 1679581782
transform 1 0 18720 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_196
timestamp 1679581782
transform 1 0 19392 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_203
timestamp 1679581782
transform 1 0 20064 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_210
timestamp 1679581782
transform 1 0 20736 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_217
timestamp 1679581782
transform 1 0 21408 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_224
timestamp 1679581782
transform 1 0 22080 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_231
timestamp 1679581782
transform 1 0 22752 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_238
timestamp 1679581782
transform 1 0 23424 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_245
timestamp 1679581782
transform 1 0 24096 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_252
timestamp 1679581782
transform 1 0 24768 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_259
timestamp 1679581782
transform 1 0 25440 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_266
timestamp 1679581782
transform 1 0 26112 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_273
timestamp 1679581782
transform 1 0 26784 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_280
timestamp 1679581782
transform 1 0 27456 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_287
timestamp 1679581782
transform 1 0 28128 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_294
timestamp 1679581782
transform 1 0 28800 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_301
timestamp 1679581782
transform 1 0 29472 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_308
timestamp 1679581782
transform 1 0 30144 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_315
timestamp 1679581782
transform 1 0 30816 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_322
timestamp 1679581782
transform 1 0 31488 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_329
timestamp 1679581782
transform 1 0 32160 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_336
timestamp 1679581782
transform 1 0 32832 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_343
timestamp 1679581782
transform 1 0 33504 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_350
timestamp 1679581782
transform 1 0 34176 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_357
timestamp 1679581782
transform 1 0 34848 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_364
timestamp 1679581782
transform 1 0 35520 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_371
timestamp 1679581782
transform 1 0 36192 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_378
timestamp 1679581782
transform 1 0 36864 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_385
timestamp 1679581782
transform 1 0 37536 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_392
timestamp 1679581782
transform 1 0 38208 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_399
timestamp 1679581782
transform 1 0 38880 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_406
timestamp 1679581782
transform 1 0 39552 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_413
timestamp 1679581782
transform 1 0 40224 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_420
timestamp 1679581782
transform 1 0 40896 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_427
timestamp 1679581782
transform 1 0 41568 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_434
timestamp 1679581782
transform 1 0 42240 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_441
timestamp 1679581782
transform 1 0 42912 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_448
timestamp 1679581782
transform 1 0 43584 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_455
timestamp 1679581782
transform 1 0 44256 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_462
timestamp 1679581782
transform 1 0 44928 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_469
timestamp 1679581782
transform 1 0 45600 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_476
timestamp 1679581782
transform 1 0 46272 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_483
timestamp 1679581782
transform 1 0 46944 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_490
timestamp 1679581782
transform 1 0 47616 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_497
timestamp 1679581782
transform 1 0 48288 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_504
timestamp 1679581782
transform 1 0 48960 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_511
timestamp 1679581782
transform 1 0 49632 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_518
timestamp 1679581782
transform 1 0 50304 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_525
timestamp 1679581782
transform 1 0 50976 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_532
timestamp 1679581782
transform 1 0 51648 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_539
timestamp 1679581782
transform 1 0 52320 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_546
timestamp 1679581782
transform 1 0 52992 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_553
timestamp 1679581782
transform 1 0 53664 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_560
timestamp 1679581782
transform 1 0 54336 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_567
timestamp 1679581782
transform 1 0 55008 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_574
timestamp 1679581782
transform 1 0 55680 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_581
timestamp 1679581782
transform 1 0 56352 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_588
timestamp 1679581782
transform 1 0 57024 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_595
timestamp 1679581782
transform 1 0 57696 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_602
timestamp 1679581782
transform 1 0 58368 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_609
timestamp 1679581782
transform 1 0 59040 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_616
timestamp 1679581782
transform 1 0 59712 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_623
timestamp 1679581782
transform 1 0 60384 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_630
timestamp 1679581782
transform 1 0 61056 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_637
timestamp 1679581782
transform 1 0 61728 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_644
timestamp 1679581782
transform 1 0 62400 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_651
timestamp 1679581782
transform 1 0 63072 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_658
timestamp 1679581782
transform 1 0 63744 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_665
timestamp 1679581782
transform 1 0 64416 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_672
timestamp 1679581782
transform 1 0 65088 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_679
timestamp 1679581782
transform 1 0 65760 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_686
timestamp 1679581782
transform 1 0 66432 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_693
timestamp 1679581782
transform 1 0 67104 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_700
timestamp 1679581782
transform 1 0 67776 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_707
timestamp 1679581782
transform 1 0 68448 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_714
timestamp 1679581782
transform 1 0 69120 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_721
timestamp 1679581782
transform 1 0 69792 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_728
timestamp 1679581782
transform 1 0 70464 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_735
timestamp 1679581782
transform 1 0 71136 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_742
timestamp 1679581782
transform 1 0 71808 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_749
timestamp 1679581782
transform 1 0 72480 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_756
timestamp 1679581782
transform 1 0 73152 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_763
timestamp 1679581782
transform 1 0 73824 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_770
timestamp 1679581782
transform 1 0 74496 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_777
timestamp 1679581782
transform 1 0 75168 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_784
timestamp 1679581782
transform 1 0 75840 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_791
timestamp 1679581782
transform 1 0 76512 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_798
timestamp 1679581782
transform 1 0 77184 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_805
timestamp 1679581782
transform 1 0 77856 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_812
timestamp 1679581782
transform 1 0 78528 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_819
timestamp 1679581782
transform 1 0 79200 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_826
timestamp 1679581782
transform 1 0 79872 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_833
timestamp 1679581782
transform 1 0 80544 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_840
timestamp 1679581782
transform 1 0 81216 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_847
timestamp 1679581782
transform 1 0 81888 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_854
timestamp 1679581782
transform 1 0 82560 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_861
timestamp 1679581782
transform 1 0 83232 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_868
timestamp 1679581782
transform 1 0 83904 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_875
timestamp 1679581782
transform 1 0 84576 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_882
timestamp 1679581782
transform 1 0 85248 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_889
timestamp 1679581782
transform 1 0 85920 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_896
timestamp 1679581782
transform 1 0 86592 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_903
timestamp 1679581782
transform 1 0 87264 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_910
timestamp 1679581782
transform 1 0 87936 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_917
timestamp 1679581782
transform 1 0 88608 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_924
timestamp 1679581782
transform 1 0 89280 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_931
timestamp 1679581782
transform 1 0 89952 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_938
timestamp 1679581782
transform 1 0 90624 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_945
timestamp 1679581782
transform 1 0 91296 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_952
timestamp 1679581782
transform 1 0 91968 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_959
timestamp 1679581782
transform 1 0 92640 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_966
timestamp 1679581782
transform 1 0 93312 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_973
timestamp 1679581782
transform 1 0 93984 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_980
timestamp 1679581782
transform 1 0 94656 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_987
timestamp 1679581782
transform 1 0 95328 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_994
timestamp 1679581782
transform 1 0 96000 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_1001
timestamp 1679581782
transform 1 0 96672 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_1008
timestamp 1679581782
transform 1 0 97344 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_1015
timestamp 1679581782
transform 1 0 98016 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_1022
timestamp 1679581782
transform 1 0 98688 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_0
timestamp 1679581782
transform 1 0 576 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_7
timestamp 1679581782
transform 1 0 1248 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_14
timestamp 1679581782
transform 1 0 1920 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_21
timestamp 1679581782
transform 1 0 2592 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_28
timestamp 1679581782
transform 1 0 3264 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_35
timestamp 1679581782
transform 1 0 3936 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_42
timestamp 1679581782
transform 1 0 4608 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_49
timestamp 1679581782
transform 1 0 5280 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_56
timestamp 1679581782
transform 1 0 5952 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_63
timestamp 1679581782
transform 1 0 6624 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_70
timestamp 1679581782
transform 1 0 7296 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_77
timestamp 1679581782
transform 1 0 7968 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_84
timestamp 1679581782
transform 1 0 8640 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_91
timestamp 1679581782
transform 1 0 9312 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_98
timestamp 1679581782
transform 1 0 9984 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_105
timestamp 1679581782
transform 1 0 10656 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_112
timestamp 1679581782
transform 1 0 11328 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_119
timestamp 1679581782
transform 1 0 12000 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_126
timestamp 1679581782
transform 1 0 12672 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_133
timestamp 1679581782
transform 1 0 13344 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_140
timestamp 1679581782
transform 1 0 14016 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_147
timestamp 1679581782
transform 1 0 14688 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_154
timestamp 1679581782
transform 1 0 15360 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_161
timestamp 1679581782
transform 1 0 16032 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_168
timestamp 1679581782
transform 1 0 16704 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_175
timestamp 1679581782
transform 1 0 17376 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_182
timestamp 1679581782
transform 1 0 18048 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_189
timestamp 1679581782
transform 1 0 18720 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_196
timestamp 1679581782
transform 1 0 19392 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_203
timestamp 1679581782
transform 1 0 20064 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_210
timestamp 1679581782
transform 1 0 20736 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_217
timestamp 1679581782
transform 1 0 21408 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_224
timestamp 1679581782
transform 1 0 22080 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_231
timestamp 1679581782
transform 1 0 22752 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_238
timestamp 1679581782
transform 1 0 23424 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_245
timestamp 1679581782
transform 1 0 24096 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_252
timestamp 1679581782
transform 1 0 24768 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_259
timestamp 1679581782
transform 1 0 25440 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_266
timestamp 1679581782
transform 1 0 26112 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_273
timestamp 1679581782
transform 1 0 26784 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_280
timestamp 1679581782
transform 1 0 27456 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_287
timestamp 1679581782
transform 1 0 28128 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_294
timestamp 1679581782
transform 1 0 28800 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_301
timestamp 1679581782
transform 1 0 29472 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_308
timestamp 1679581782
transform 1 0 30144 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_315
timestamp 1679581782
transform 1 0 30816 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_322
timestamp 1679581782
transform 1 0 31488 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_329
timestamp 1679581782
transform 1 0 32160 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_336
timestamp 1679581782
transform 1 0 32832 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_343
timestamp 1679581782
transform 1 0 33504 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_350
timestamp 1679581782
transform 1 0 34176 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_357
timestamp 1679581782
transform 1 0 34848 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_364
timestamp 1679581782
transform 1 0 35520 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_371
timestamp 1679581782
transform 1 0 36192 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_378
timestamp 1679581782
transform 1 0 36864 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_385
timestamp 1679581782
transform 1 0 37536 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_392
timestamp 1679581782
transform 1 0 38208 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_399
timestamp 1679581782
transform 1 0 38880 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_406
timestamp 1679581782
transform 1 0 39552 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_413
timestamp 1679581782
transform 1 0 40224 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_420
timestamp 1679581782
transform 1 0 40896 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_427
timestamp 1679581782
transform 1 0 41568 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_434
timestamp 1679581782
transform 1 0 42240 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_441
timestamp 1679581782
transform 1 0 42912 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_448
timestamp 1679581782
transform 1 0 43584 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_455
timestamp 1679581782
transform 1 0 44256 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_462
timestamp 1679581782
transform 1 0 44928 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_469
timestamp 1679581782
transform 1 0 45600 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_476
timestamp 1679581782
transform 1 0 46272 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_483
timestamp 1679581782
transform 1 0 46944 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_490
timestamp 1679581782
transform 1 0 47616 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_497
timestamp 1679581782
transform 1 0 48288 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_504
timestamp 1679581782
transform 1 0 48960 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_511
timestamp 1679581782
transform 1 0 49632 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_518
timestamp 1679581782
transform 1 0 50304 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_525
timestamp 1679581782
transform 1 0 50976 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_532
timestamp 1679581782
transform 1 0 51648 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_539
timestamp 1679581782
transform 1 0 52320 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_546
timestamp 1679581782
transform 1 0 52992 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_553
timestamp 1679581782
transform 1 0 53664 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_560
timestamp 1679581782
transform 1 0 54336 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_567
timestamp 1679581782
transform 1 0 55008 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_574
timestamp 1679581782
transform 1 0 55680 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_581
timestamp 1679581782
transform 1 0 56352 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_588
timestamp 1679581782
transform 1 0 57024 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_595
timestamp 1679581782
transform 1 0 57696 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_602
timestamp 1679581782
transform 1 0 58368 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_609
timestamp 1679581782
transform 1 0 59040 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_616
timestamp 1679581782
transform 1 0 59712 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_623
timestamp 1679581782
transform 1 0 60384 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_630
timestamp 1679581782
transform 1 0 61056 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_637
timestamp 1679581782
transform 1 0 61728 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_644
timestamp 1679581782
transform 1 0 62400 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_651
timestamp 1679581782
transform 1 0 63072 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_658
timestamp 1679581782
transform 1 0 63744 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_665
timestamp 1679581782
transform 1 0 64416 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_672
timestamp 1679581782
transform 1 0 65088 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_679
timestamp 1679581782
transform 1 0 65760 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_686
timestamp 1679581782
transform 1 0 66432 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_693
timestamp 1679581782
transform 1 0 67104 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_700
timestamp 1679581782
transform 1 0 67776 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_707
timestamp 1679581782
transform 1 0 68448 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_714
timestamp 1679581782
transform 1 0 69120 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_721
timestamp 1679581782
transform 1 0 69792 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_728
timestamp 1679581782
transform 1 0 70464 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_735
timestamp 1679581782
transform 1 0 71136 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_742
timestamp 1679581782
transform 1 0 71808 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_749
timestamp 1679581782
transform 1 0 72480 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_756
timestamp 1679581782
transform 1 0 73152 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_763
timestamp 1679581782
transform 1 0 73824 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_770
timestamp 1679581782
transform 1 0 74496 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_777
timestamp 1679581782
transform 1 0 75168 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_784
timestamp 1679581782
transform 1 0 75840 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_791
timestamp 1679581782
transform 1 0 76512 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_798
timestamp 1679581782
transform 1 0 77184 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_805
timestamp 1679581782
transform 1 0 77856 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_812
timestamp 1679581782
transform 1 0 78528 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_819
timestamp 1679581782
transform 1 0 79200 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_826
timestamp 1679581782
transform 1 0 79872 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_833
timestamp 1679581782
transform 1 0 80544 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_840
timestamp 1679581782
transform 1 0 81216 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_847
timestamp 1679581782
transform 1 0 81888 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_854
timestamp 1679581782
transform 1 0 82560 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_861
timestamp 1679581782
transform 1 0 83232 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_868
timestamp 1679581782
transform 1 0 83904 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_875
timestamp 1679581782
transform 1 0 84576 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_882
timestamp 1679581782
transform 1 0 85248 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_889
timestamp 1679581782
transform 1 0 85920 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_896
timestamp 1679581782
transform 1 0 86592 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_903
timestamp 1679581782
transform 1 0 87264 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_910
timestamp 1679581782
transform 1 0 87936 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_917
timestamp 1679581782
transform 1 0 88608 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_924
timestamp 1679581782
transform 1 0 89280 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_931
timestamp 1679581782
transform 1 0 89952 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_938
timestamp 1679581782
transform 1 0 90624 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_945
timestamp 1679581782
transform 1 0 91296 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_952
timestamp 1679581782
transform 1 0 91968 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_959
timestamp 1679581782
transform 1 0 92640 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_966
timestamp 1679581782
transform 1 0 93312 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_973
timestamp 1679581782
transform 1 0 93984 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_980
timestamp 1679581782
transform 1 0 94656 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_987
timestamp 1679581782
transform 1 0 95328 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_994
timestamp 1679581782
transform 1 0 96000 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_1001
timestamp 1679581782
transform 1 0 96672 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_1008
timestamp 1679581782
transform 1 0 97344 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_1015
timestamp 1679581782
transform 1 0 98016 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_1022
timestamp 1679581782
transform 1 0 98688 0 1 70308
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_5
timestamp 1679581782
transform 1 0 1056 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_12
timestamp 1679581782
transform 1 0 1728 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_19
timestamp 1679581782
transform 1 0 2400 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_26
timestamp 1679581782
transform 1 0 3072 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_33
timestamp 1679581782
transform 1 0 3744 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_40
timestamp 1679581782
transform 1 0 4416 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_47
timestamp 1679581782
transform 1 0 5088 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_54
timestamp 1679581782
transform 1 0 5760 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_61
timestamp 1679581782
transform 1 0 6432 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_68
timestamp 1679581782
transform 1 0 7104 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_75
timestamp 1679581782
transform 1 0 7776 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_82
timestamp 1679581782
transform 1 0 8448 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_89
timestamp 1679581782
transform 1 0 9120 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_96
timestamp 1679581782
transform 1 0 9792 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_103
timestamp 1679581782
transform 1 0 10464 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_110
timestamp 1679581782
transform 1 0 11136 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_117
timestamp 1679581782
transform 1 0 11808 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_124
timestamp 1679581782
transform 1 0 12480 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_131
timestamp 1679581782
transform 1 0 13152 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_138
timestamp 1679581782
transform 1 0 13824 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_145
timestamp 1679581782
transform 1 0 14496 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_152
timestamp 1679581782
transform 1 0 15168 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_159
timestamp 1679581782
transform 1 0 15840 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_166
timestamp 1679581782
transform 1 0 16512 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_173
timestamp 1679581782
transform 1 0 17184 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_180
timestamp 1679581782
transform 1 0 17856 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_187
timestamp 1679581782
transform 1 0 18528 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_194
timestamp 1679581782
transform 1 0 19200 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_201
timestamp 1679581782
transform 1 0 19872 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_208
timestamp 1679581782
transform 1 0 20544 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_215
timestamp 1679581782
transform 1 0 21216 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_222
timestamp 1679581782
transform 1 0 21888 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_229
timestamp 1679581782
transform 1 0 22560 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_236
timestamp 1679581782
transform 1 0 23232 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_243
timestamp 1679581782
transform 1 0 23904 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_250
timestamp 1679581782
transform 1 0 24576 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_257
timestamp 1679581782
transform 1 0 25248 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_264
timestamp 1679581782
transform 1 0 25920 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_271
timestamp 1679581782
transform 1 0 26592 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_278
timestamp 1679581782
transform 1 0 27264 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_285
timestamp 1679581782
transform 1 0 27936 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_292
timestamp 1679581782
transform 1 0 28608 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_299
timestamp 1679581782
transform 1 0 29280 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_306
timestamp 1679581782
transform 1 0 29952 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_313
timestamp 1679581782
transform 1 0 30624 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_320
timestamp 1679581782
transform 1 0 31296 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_327
timestamp 1679581782
transform 1 0 31968 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_334
timestamp 1679581782
transform 1 0 32640 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_341
timestamp 1679581782
transform 1 0 33312 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_348
timestamp 1679581782
transform 1 0 33984 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_355
timestamp 1679581782
transform 1 0 34656 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_362
timestamp 1679581782
transform 1 0 35328 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_369
timestamp 1679581782
transform 1 0 36000 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_376
timestamp 1679581782
transform 1 0 36672 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_383
timestamp 1679581782
transform 1 0 37344 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_390
timestamp 1679581782
transform 1 0 38016 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_397
timestamp 1679581782
transform 1 0 38688 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_404
timestamp 1679581782
transform 1 0 39360 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_411
timestamp 1679581782
transform 1 0 40032 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_418
timestamp 1679581782
transform 1 0 40704 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_425
timestamp 1679581782
transform 1 0 41376 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_432
timestamp 1679581782
transform 1 0 42048 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_439
timestamp 1679581782
transform 1 0 42720 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_446
timestamp 1679581782
transform 1 0 43392 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_453
timestamp 1679581782
transform 1 0 44064 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_460
timestamp 1679581782
transform 1 0 44736 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_467
timestamp 1679581782
transform 1 0 45408 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_474
timestamp 1679581782
transform 1 0 46080 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_481
timestamp 1679581782
transform 1 0 46752 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_488
timestamp 1679581782
transform 1 0 47424 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_495
timestamp 1679581782
transform 1 0 48096 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_502
timestamp 1679581782
transform 1 0 48768 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_509
timestamp 1679581782
transform 1 0 49440 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_516
timestamp 1679581782
transform 1 0 50112 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_523
timestamp 1679581782
transform 1 0 50784 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_530
timestamp 1679581782
transform 1 0 51456 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_537
timestamp 1679581782
transform 1 0 52128 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_544
timestamp 1679581782
transform 1 0 52800 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_551
timestamp 1679581782
transform 1 0 53472 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_558
timestamp 1679581782
transform 1 0 54144 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_565
timestamp 1679581782
transform 1 0 54816 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_572
timestamp 1679581782
transform 1 0 55488 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_579
timestamp 1679581782
transform 1 0 56160 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_586
timestamp 1679581782
transform 1 0 56832 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_593
timestamp 1679581782
transform 1 0 57504 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_600
timestamp 1679581782
transform 1 0 58176 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_607
timestamp 1679581782
transform 1 0 58848 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_614
timestamp 1679581782
transform 1 0 59520 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_621
timestamp 1679581782
transform 1 0 60192 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_628
timestamp 1679581782
transform 1 0 60864 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_635
timestamp 1679581782
transform 1 0 61536 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_642
timestamp 1679581782
transform 1 0 62208 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_649
timestamp 1679581782
transform 1 0 62880 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_656
timestamp 1679581782
transform 1 0 63552 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_663
timestamp 1679581782
transform 1 0 64224 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_670
timestamp 1679581782
transform 1 0 64896 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_677
timestamp 1679581782
transform 1 0 65568 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_684
timestamp 1679581782
transform 1 0 66240 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_691
timestamp 1679581782
transform 1 0 66912 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_698
timestamp 1679581782
transform 1 0 67584 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_705
timestamp 1679581782
transform 1 0 68256 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_712
timestamp 1679581782
transform 1 0 68928 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_719
timestamp 1679581782
transform 1 0 69600 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_726
timestamp 1679581782
transform 1 0 70272 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_733
timestamp 1679581782
transform 1 0 70944 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_740
timestamp 1679581782
transform 1 0 71616 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_747
timestamp 1679581782
transform 1 0 72288 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_754
timestamp 1679581782
transform 1 0 72960 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_761
timestamp 1679581782
transform 1 0 73632 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_768
timestamp 1679581782
transform 1 0 74304 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_775
timestamp 1679581782
transform 1 0 74976 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_782
timestamp 1679581782
transform 1 0 75648 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_789
timestamp 1679581782
transform 1 0 76320 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_796
timestamp 1679581782
transform 1 0 76992 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_803
timestamp 1679581782
transform 1 0 77664 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_810
timestamp 1679581782
transform 1 0 78336 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_817
timestamp 1679581782
transform 1 0 79008 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_824
timestamp 1679581782
transform 1 0 79680 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_831
timestamp 1679581782
transform 1 0 80352 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_838
timestamp 1679581782
transform 1 0 81024 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_845
timestamp 1679581782
transform 1 0 81696 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_852
timestamp 1679581782
transform 1 0 82368 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_859
timestamp 1679581782
transform 1 0 83040 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_866
timestamp 1679581782
transform 1 0 83712 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_873
timestamp 1679581782
transform 1 0 84384 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_880
timestamp 1679581782
transform 1 0 85056 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_887
timestamp 1679581782
transform 1 0 85728 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_894
timestamp 1679581782
transform 1 0 86400 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_901
timestamp 1679581782
transform 1 0 87072 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_908
timestamp 1679581782
transform 1 0 87744 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_915
timestamp 1679581782
transform 1 0 88416 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_922
timestamp 1679581782
transform 1 0 89088 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_929
timestamp 1679581782
transform 1 0 89760 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_936
timestamp 1679581782
transform 1 0 90432 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_943
timestamp 1679581782
transform 1 0 91104 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_950
timestamp 1679581782
transform 1 0 91776 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_957
timestamp 1679581782
transform 1 0 92448 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_964
timestamp 1679581782
transform 1 0 93120 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_971
timestamp 1679581782
transform 1 0 93792 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_978
timestamp 1679581782
transform 1 0 94464 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_985
timestamp 1679581782
transform 1 0 95136 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_992
timestamp 1679581782
transform 1 0 95808 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_999
timestamp 1679581782
transform 1 0 96480 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_1006
timestamp 1679581782
transform 1 0 97152 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_1013
timestamp 1679581782
transform 1 0 97824 0 -1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_1020
timestamp 1679581782
transform 1 0 98496 0 -1 71820
box -48 -56 720 834
use sg13g2_fill_2  FILLER_93_1027
timestamp 1677580104
transform 1 0 99168 0 -1 71820
box -48 -56 240 834
use sg13g2_decap_8  FILLER_94_0
timestamp 1679581782
transform 1 0 576 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_7
timestamp 1679581782
transform 1 0 1248 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_14
timestamp 1679581782
transform 1 0 1920 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_21
timestamp 1679581782
transform 1 0 2592 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_28
timestamp 1679581782
transform 1 0 3264 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_35
timestamp 1679581782
transform 1 0 3936 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_42
timestamp 1679581782
transform 1 0 4608 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_49
timestamp 1679581782
transform 1 0 5280 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_56
timestamp 1679581782
transform 1 0 5952 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_63
timestamp 1679581782
transform 1 0 6624 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_70
timestamp 1679581782
transform 1 0 7296 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_77
timestamp 1679581782
transform 1 0 7968 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_84
timestamp 1679581782
transform 1 0 8640 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_91
timestamp 1679581782
transform 1 0 9312 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_98
timestamp 1679581782
transform 1 0 9984 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_105
timestamp 1679581782
transform 1 0 10656 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_112
timestamp 1679581782
transform 1 0 11328 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_119
timestamp 1679581782
transform 1 0 12000 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_126
timestamp 1679581782
transform 1 0 12672 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_133
timestamp 1679581782
transform 1 0 13344 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_140
timestamp 1679581782
transform 1 0 14016 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_147
timestamp 1679581782
transform 1 0 14688 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_154
timestamp 1679581782
transform 1 0 15360 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_161
timestamp 1679581782
transform 1 0 16032 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_168
timestamp 1679581782
transform 1 0 16704 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_175
timestamp 1679581782
transform 1 0 17376 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_182
timestamp 1679581782
transform 1 0 18048 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_189
timestamp 1679581782
transform 1 0 18720 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_196
timestamp 1679581782
transform 1 0 19392 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_203
timestamp 1679581782
transform 1 0 20064 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_210
timestamp 1679581782
transform 1 0 20736 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_217
timestamp 1679581782
transform 1 0 21408 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_224
timestamp 1679581782
transform 1 0 22080 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_231
timestamp 1679581782
transform 1 0 22752 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_238
timestamp 1679581782
transform 1 0 23424 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_245
timestamp 1679581782
transform 1 0 24096 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_252
timestamp 1679581782
transform 1 0 24768 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_259
timestamp 1679581782
transform 1 0 25440 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_266
timestamp 1679581782
transform 1 0 26112 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_273
timestamp 1679581782
transform 1 0 26784 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_280
timestamp 1679581782
transform 1 0 27456 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_287
timestamp 1679581782
transform 1 0 28128 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_294
timestamp 1679581782
transform 1 0 28800 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_301
timestamp 1679581782
transform 1 0 29472 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_308
timestamp 1679581782
transform 1 0 30144 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_315
timestamp 1679581782
transform 1 0 30816 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_322
timestamp 1679581782
transform 1 0 31488 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_329
timestamp 1679581782
transform 1 0 32160 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_336
timestamp 1679581782
transform 1 0 32832 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_343
timestamp 1679581782
transform 1 0 33504 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_350
timestamp 1679581782
transform 1 0 34176 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_357
timestamp 1679581782
transform 1 0 34848 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_364
timestamp 1679581782
transform 1 0 35520 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_371
timestamp 1679581782
transform 1 0 36192 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_378
timestamp 1679581782
transform 1 0 36864 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_385
timestamp 1679581782
transform 1 0 37536 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_392
timestamp 1679581782
transform 1 0 38208 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_399
timestamp 1679581782
transform 1 0 38880 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_406
timestamp 1679581782
transform 1 0 39552 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_413
timestamp 1679581782
transform 1 0 40224 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_420
timestamp 1679581782
transform 1 0 40896 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_427
timestamp 1679581782
transform 1 0 41568 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_434
timestamp 1679581782
transform 1 0 42240 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_441
timestamp 1679581782
transform 1 0 42912 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_448
timestamp 1679581782
transform 1 0 43584 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_455
timestamp 1679581782
transform 1 0 44256 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_462
timestamp 1679581782
transform 1 0 44928 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_469
timestamp 1679581782
transform 1 0 45600 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_476
timestamp 1679581782
transform 1 0 46272 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_483
timestamp 1679581782
transform 1 0 46944 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_490
timestamp 1679581782
transform 1 0 47616 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_497
timestamp 1679581782
transform 1 0 48288 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_504
timestamp 1679581782
transform 1 0 48960 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_511
timestamp 1679581782
transform 1 0 49632 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_518
timestamp 1679581782
transform 1 0 50304 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_525
timestamp 1679581782
transform 1 0 50976 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_532
timestamp 1679581782
transform 1 0 51648 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_539
timestamp 1679581782
transform 1 0 52320 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_546
timestamp 1679581782
transform 1 0 52992 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_553
timestamp 1679581782
transform 1 0 53664 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_560
timestamp 1679581782
transform 1 0 54336 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_567
timestamp 1679581782
transform 1 0 55008 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_574
timestamp 1679581782
transform 1 0 55680 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_581
timestamp 1679581782
transform 1 0 56352 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_588
timestamp 1679581782
transform 1 0 57024 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_595
timestamp 1679581782
transform 1 0 57696 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_602
timestamp 1679581782
transform 1 0 58368 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_609
timestamp 1679581782
transform 1 0 59040 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_616
timestamp 1679581782
transform 1 0 59712 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_623
timestamp 1679581782
transform 1 0 60384 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_630
timestamp 1679581782
transform 1 0 61056 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_637
timestamp 1679581782
transform 1 0 61728 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_644
timestamp 1679581782
transform 1 0 62400 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_651
timestamp 1679581782
transform 1 0 63072 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_658
timestamp 1679581782
transform 1 0 63744 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_665
timestamp 1679581782
transform 1 0 64416 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_672
timestamp 1679581782
transform 1 0 65088 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_679
timestamp 1679581782
transform 1 0 65760 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_686
timestamp 1679581782
transform 1 0 66432 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_693
timestamp 1679581782
transform 1 0 67104 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_700
timestamp 1679581782
transform 1 0 67776 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_707
timestamp 1679581782
transform 1 0 68448 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_714
timestamp 1679581782
transform 1 0 69120 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_721
timestamp 1679581782
transform 1 0 69792 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_728
timestamp 1679581782
transform 1 0 70464 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_735
timestamp 1679581782
transform 1 0 71136 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_742
timestamp 1679581782
transform 1 0 71808 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_749
timestamp 1679581782
transform 1 0 72480 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_756
timestamp 1679581782
transform 1 0 73152 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_763
timestamp 1679581782
transform 1 0 73824 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_770
timestamp 1679581782
transform 1 0 74496 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_777
timestamp 1679581782
transform 1 0 75168 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_784
timestamp 1679581782
transform 1 0 75840 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_791
timestamp 1679581782
transform 1 0 76512 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_798
timestamp 1679581782
transform 1 0 77184 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_805
timestamp 1679581782
transform 1 0 77856 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_812
timestamp 1679581782
transform 1 0 78528 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_819
timestamp 1679581782
transform 1 0 79200 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_826
timestamp 1679581782
transform 1 0 79872 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_833
timestamp 1679581782
transform 1 0 80544 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_840
timestamp 1679581782
transform 1 0 81216 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_847
timestamp 1679581782
transform 1 0 81888 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_854
timestamp 1679581782
transform 1 0 82560 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_861
timestamp 1679581782
transform 1 0 83232 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_868
timestamp 1679581782
transform 1 0 83904 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_875
timestamp 1679581782
transform 1 0 84576 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_882
timestamp 1679581782
transform 1 0 85248 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_889
timestamp 1679581782
transform 1 0 85920 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_896
timestamp 1679581782
transform 1 0 86592 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_903
timestamp 1679581782
transform 1 0 87264 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_910
timestamp 1679581782
transform 1 0 87936 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_917
timestamp 1679581782
transform 1 0 88608 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_924
timestamp 1679581782
transform 1 0 89280 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_931
timestamp 1679581782
transform 1 0 89952 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_938
timestamp 1679581782
transform 1 0 90624 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_945
timestamp 1679581782
transform 1 0 91296 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_952
timestamp 1679581782
transform 1 0 91968 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_959
timestamp 1679581782
transform 1 0 92640 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_966
timestamp 1679581782
transform 1 0 93312 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_973
timestamp 1679581782
transform 1 0 93984 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_980
timestamp 1679581782
transform 1 0 94656 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_987
timestamp 1679581782
transform 1 0 95328 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_994
timestamp 1679581782
transform 1 0 96000 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_1001
timestamp 1679581782
transform 1 0 96672 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_1008
timestamp 1679581782
transform 1 0 97344 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_1015
timestamp 1679581782
transform 1 0 98016 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_1022
timestamp 1679581782
transform 1 0 98688 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_4
timestamp 1679581782
transform 1 0 960 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_11
timestamp 1679581782
transform 1 0 1632 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_18
timestamp 1679581782
transform 1 0 2304 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_25
timestamp 1679581782
transform 1 0 2976 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_32
timestamp 1679581782
transform 1 0 3648 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_39
timestamp 1679581782
transform 1 0 4320 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_46
timestamp 1679581782
transform 1 0 4992 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_53
timestamp 1679581782
transform 1 0 5664 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_60
timestamp 1679581782
transform 1 0 6336 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_67
timestamp 1679581782
transform 1 0 7008 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_74
timestamp 1679581782
transform 1 0 7680 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_81
timestamp 1679581782
transform 1 0 8352 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_88
timestamp 1679581782
transform 1 0 9024 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_95
timestamp 1679581782
transform 1 0 9696 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_102
timestamp 1679581782
transform 1 0 10368 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_109
timestamp 1679581782
transform 1 0 11040 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_116
timestamp 1679581782
transform 1 0 11712 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_123
timestamp 1679581782
transform 1 0 12384 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_130
timestamp 1679581782
transform 1 0 13056 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_137
timestamp 1679581782
transform 1 0 13728 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_144
timestamp 1679581782
transform 1 0 14400 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_151
timestamp 1679581782
transform 1 0 15072 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_158
timestamp 1679581782
transform 1 0 15744 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_165
timestamp 1679581782
transform 1 0 16416 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_172
timestamp 1679581782
transform 1 0 17088 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_179
timestamp 1679581782
transform 1 0 17760 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_186
timestamp 1679581782
transform 1 0 18432 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_193
timestamp 1679581782
transform 1 0 19104 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_200
timestamp 1679581782
transform 1 0 19776 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_207
timestamp 1679581782
transform 1 0 20448 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_214
timestamp 1679581782
transform 1 0 21120 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_221
timestamp 1679581782
transform 1 0 21792 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_228
timestamp 1679581782
transform 1 0 22464 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_235
timestamp 1679581782
transform 1 0 23136 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_242
timestamp 1679581782
transform 1 0 23808 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_249
timestamp 1679581782
transform 1 0 24480 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_256
timestamp 1679581782
transform 1 0 25152 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_263
timestamp 1679581782
transform 1 0 25824 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_270
timestamp 1679581782
transform 1 0 26496 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_277
timestamp 1679581782
transform 1 0 27168 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_284
timestamp 1679581782
transform 1 0 27840 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_291
timestamp 1679581782
transform 1 0 28512 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_298
timestamp 1679581782
transform 1 0 29184 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_305
timestamp 1679581782
transform 1 0 29856 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_312
timestamp 1679581782
transform 1 0 30528 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_319
timestamp 1679581782
transform 1 0 31200 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_326
timestamp 1679581782
transform 1 0 31872 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_333
timestamp 1679581782
transform 1 0 32544 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_340
timestamp 1679581782
transform 1 0 33216 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_347
timestamp 1679581782
transform 1 0 33888 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_354
timestamp 1679581782
transform 1 0 34560 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_361
timestamp 1679581782
transform 1 0 35232 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_368
timestamp 1679581782
transform 1 0 35904 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_375
timestamp 1679581782
transform 1 0 36576 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_382
timestamp 1679581782
transform 1 0 37248 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_389
timestamp 1679581782
transform 1 0 37920 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_396
timestamp 1679581782
transform 1 0 38592 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_403
timestamp 1679581782
transform 1 0 39264 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_410
timestamp 1679581782
transform 1 0 39936 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_417
timestamp 1679581782
transform 1 0 40608 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_424
timestamp 1679581782
transform 1 0 41280 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_431
timestamp 1679581782
transform 1 0 41952 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_438
timestamp 1679581782
transform 1 0 42624 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_445
timestamp 1679581782
transform 1 0 43296 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_452
timestamp 1679581782
transform 1 0 43968 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_459
timestamp 1679581782
transform 1 0 44640 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_466
timestamp 1679581782
transform 1 0 45312 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_473
timestamp 1679581782
transform 1 0 45984 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_480
timestamp 1679581782
transform 1 0 46656 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_487
timestamp 1679581782
transform 1 0 47328 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_494
timestamp 1679581782
transform 1 0 48000 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_501
timestamp 1679581782
transform 1 0 48672 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_508
timestamp 1679581782
transform 1 0 49344 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_515
timestamp 1679581782
transform 1 0 50016 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_522
timestamp 1679581782
transform 1 0 50688 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_529
timestamp 1679581782
transform 1 0 51360 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_536
timestamp 1679581782
transform 1 0 52032 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_543
timestamp 1679581782
transform 1 0 52704 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_550
timestamp 1679581782
transform 1 0 53376 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_557
timestamp 1679581782
transform 1 0 54048 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_564
timestamp 1679581782
transform 1 0 54720 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_571
timestamp 1679581782
transform 1 0 55392 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_578
timestamp 1679581782
transform 1 0 56064 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_585
timestamp 1679581782
transform 1 0 56736 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_592
timestamp 1679581782
transform 1 0 57408 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_599
timestamp 1679581782
transform 1 0 58080 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_606
timestamp 1679581782
transform 1 0 58752 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_613
timestamp 1679581782
transform 1 0 59424 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_620
timestamp 1679581782
transform 1 0 60096 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_627
timestamp 1679581782
transform 1 0 60768 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_634
timestamp 1679581782
transform 1 0 61440 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_641
timestamp 1679581782
transform 1 0 62112 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_648
timestamp 1679581782
transform 1 0 62784 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_655
timestamp 1679581782
transform 1 0 63456 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_662
timestamp 1679581782
transform 1 0 64128 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_669
timestamp 1679581782
transform 1 0 64800 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_676
timestamp 1679581782
transform 1 0 65472 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_683
timestamp 1679581782
transform 1 0 66144 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_690
timestamp 1679581782
transform 1 0 66816 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_697
timestamp 1679581782
transform 1 0 67488 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_704
timestamp 1679581782
transform 1 0 68160 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_711
timestamp 1679581782
transform 1 0 68832 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_718
timestamp 1679581782
transform 1 0 69504 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_725
timestamp 1679581782
transform 1 0 70176 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_732
timestamp 1679581782
transform 1 0 70848 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_739
timestamp 1679581782
transform 1 0 71520 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_746
timestamp 1679581782
transform 1 0 72192 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_753
timestamp 1679581782
transform 1 0 72864 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_760
timestamp 1679581782
transform 1 0 73536 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_767
timestamp 1679581782
transform 1 0 74208 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_774
timestamp 1679581782
transform 1 0 74880 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_781
timestamp 1679581782
transform 1 0 75552 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_788
timestamp 1679581782
transform 1 0 76224 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_795
timestamp 1679581782
transform 1 0 76896 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_802
timestamp 1679581782
transform 1 0 77568 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_809
timestamp 1679581782
transform 1 0 78240 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_816
timestamp 1679581782
transform 1 0 78912 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_823
timestamp 1679581782
transform 1 0 79584 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_830
timestamp 1679581782
transform 1 0 80256 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_837
timestamp 1679581782
transform 1 0 80928 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_844
timestamp 1679581782
transform 1 0 81600 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_851
timestamp 1679581782
transform 1 0 82272 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_858
timestamp 1679581782
transform 1 0 82944 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_865
timestamp 1679581782
transform 1 0 83616 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_872
timestamp 1679581782
transform 1 0 84288 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_879
timestamp 1679581782
transform 1 0 84960 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_886
timestamp 1679581782
transform 1 0 85632 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_893
timestamp 1679581782
transform 1 0 86304 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_900
timestamp 1679581782
transform 1 0 86976 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_907
timestamp 1679581782
transform 1 0 87648 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_914
timestamp 1679581782
transform 1 0 88320 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_921
timestamp 1679581782
transform 1 0 88992 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_928
timestamp 1679581782
transform 1 0 89664 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_935
timestamp 1679581782
transform 1 0 90336 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_942
timestamp 1679581782
transform 1 0 91008 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_949
timestamp 1679581782
transform 1 0 91680 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_956
timestamp 1679581782
transform 1 0 92352 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_963
timestamp 1679581782
transform 1 0 93024 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_970
timestamp 1679581782
transform 1 0 93696 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_977
timestamp 1679581782
transform 1 0 94368 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_984
timestamp 1679581782
transform 1 0 95040 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_991
timestamp 1679581782
transform 1 0 95712 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_998
timestamp 1679581782
transform 1 0 96384 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_1005
timestamp 1679581782
transform 1 0 97056 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_1012
timestamp 1679581782
transform 1 0 97728 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_1019
timestamp 1679581782
transform 1 0 98400 0 -1 73332
box -48 -56 720 834
use sg13g2_fill_2  FILLER_95_1026
timestamp 1677580104
transform 1 0 99072 0 -1 73332
box -48 -56 240 834
use sg13g2_fill_1  FILLER_95_1028
timestamp 1677579658
transform 1 0 99264 0 -1 73332
box -48 -56 144 834
use sg13g2_decap_8  FILLER_96_0
timestamp 1679581782
transform 1 0 576 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_7
timestamp 1679581782
transform 1 0 1248 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_14
timestamp 1679581782
transform 1 0 1920 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_21
timestamp 1679581782
transform 1 0 2592 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_28
timestamp 1679581782
transform 1 0 3264 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_35
timestamp 1679581782
transform 1 0 3936 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_42
timestamp 1679581782
transform 1 0 4608 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_49
timestamp 1679581782
transform 1 0 5280 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_56
timestamp 1679581782
transform 1 0 5952 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_63
timestamp 1679581782
transform 1 0 6624 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_70
timestamp 1679581782
transform 1 0 7296 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_77
timestamp 1679581782
transform 1 0 7968 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_84
timestamp 1679581782
transform 1 0 8640 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_91
timestamp 1679581782
transform 1 0 9312 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_98
timestamp 1679581782
transform 1 0 9984 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_105
timestamp 1679581782
transform 1 0 10656 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_112
timestamp 1679581782
transform 1 0 11328 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_119
timestamp 1679581782
transform 1 0 12000 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_126
timestamp 1679581782
transform 1 0 12672 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_133
timestamp 1679581782
transform 1 0 13344 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_140
timestamp 1679581782
transform 1 0 14016 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_147
timestamp 1679581782
transform 1 0 14688 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_154
timestamp 1679581782
transform 1 0 15360 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_161
timestamp 1679581782
transform 1 0 16032 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_168
timestamp 1679581782
transform 1 0 16704 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_175
timestamp 1679581782
transform 1 0 17376 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_182
timestamp 1679581782
transform 1 0 18048 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_189
timestamp 1679581782
transform 1 0 18720 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_196
timestamp 1679581782
transform 1 0 19392 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_203
timestamp 1679581782
transform 1 0 20064 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_210
timestamp 1679581782
transform 1 0 20736 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_217
timestamp 1679581782
transform 1 0 21408 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_224
timestamp 1679581782
transform 1 0 22080 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_231
timestamp 1679581782
transform 1 0 22752 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_238
timestamp 1679581782
transform 1 0 23424 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_245
timestamp 1679581782
transform 1 0 24096 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_252
timestamp 1679581782
transform 1 0 24768 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_259
timestamp 1679581782
transform 1 0 25440 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_266
timestamp 1679581782
transform 1 0 26112 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_273
timestamp 1679581782
transform 1 0 26784 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_280
timestamp 1679581782
transform 1 0 27456 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_287
timestamp 1679581782
transform 1 0 28128 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_294
timestamp 1679581782
transform 1 0 28800 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_301
timestamp 1679581782
transform 1 0 29472 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_308
timestamp 1679581782
transform 1 0 30144 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_315
timestamp 1679581782
transform 1 0 30816 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_322
timestamp 1679581782
transform 1 0 31488 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_329
timestamp 1679581782
transform 1 0 32160 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_336
timestamp 1679581782
transform 1 0 32832 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_343
timestamp 1679581782
transform 1 0 33504 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_350
timestamp 1679581782
transform 1 0 34176 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_357
timestamp 1679581782
transform 1 0 34848 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_364
timestamp 1679581782
transform 1 0 35520 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_371
timestamp 1679581782
transform 1 0 36192 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_378
timestamp 1679581782
transform 1 0 36864 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_385
timestamp 1679581782
transform 1 0 37536 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_392
timestamp 1679581782
transform 1 0 38208 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_399
timestamp 1679581782
transform 1 0 38880 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_406
timestamp 1679581782
transform 1 0 39552 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_413
timestamp 1679581782
transform 1 0 40224 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_420
timestamp 1679581782
transform 1 0 40896 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_427
timestamp 1679581782
transform 1 0 41568 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_434
timestamp 1679581782
transform 1 0 42240 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_441
timestamp 1679581782
transform 1 0 42912 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_448
timestamp 1679581782
transform 1 0 43584 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_455
timestamp 1679581782
transform 1 0 44256 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_462
timestamp 1679581782
transform 1 0 44928 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_469
timestamp 1679581782
transform 1 0 45600 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_476
timestamp 1679581782
transform 1 0 46272 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_483
timestamp 1679581782
transform 1 0 46944 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_490
timestamp 1679581782
transform 1 0 47616 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_497
timestamp 1679581782
transform 1 0 48288 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_504
timestamp 1679581782
transform 1 0 48960 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_511
timestamp 1679581782
transform 1 0 49632 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_518
timestamp 1679581782
transform 1 0 50304 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_525
timestamp 1679581782
transform 1 0 50976 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_532
timestamp 1679581782
transform 1 0 51648 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_539
timestamp 1679581782
transform 1 0 52320 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_546
timestamp 1679581782
transform 1 0 52992 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_553
timestamp 1679581782
transform 1 0 53664 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_560
timestamp 1679581782
transform 1 0 54336 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_567
timestamp 1679581782
transform 1 0 55008 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_574
timestamp 1679581782
transform 1 0 55680 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_581
timestamp 1679581782
transform 1 0 56352 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_588
timestamp 1679581782
transform 1 0 57024 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_595
timestamp 1679581782
transform 1 0 57696 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_602
timestamp 1679581782
transform 1 0 58368 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_609
timestamp 1679581782
transform 1 0 59040 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_616
timestamp 1679581782
transform 1 0 59712 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_623
timestamp 1679581782
transform 1 0 60384 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_630
timestamp 1679581782
transform 1 0 61056 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_637
timestamp 1679581782
transform 1 0 61728 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_644
timestamp 1679581782
transform 1 0 62400 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_651
timestamp 1679581782
transform 1 0 63072 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_658
timestamp 1679581782
transform 1 0 63744 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_665
timestamp 1679581782
transform 1 0 64416 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_672
timestamp 1679581782
transform 1 0 65088 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_679
timestamp 1679581782
transform 1 0 65760 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_686
timestamp 1679581782
transform 1 0 66432 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_693
timestamp 1679581782
transform 1 0 67104 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_700
timestamp 1679581782
transform 1 0 67776 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_707
timestamp 1679581782
transform 1 0 68448 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_714
timestamp 1679581782
transform 1 0 69120 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_721
timestamp 1679581782
transform 1 0 69792 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_728
timestamp 1679581782
transform 1 0 70464 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_735
timestamp 1679581782
transform 1 0 71136 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_742
timestamp 1679581782
transform 1 0 71808 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_749
timestamp 1679581782
transform 1 0 72480 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_756
timestamp 1679581782
transform 1 0 73152 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_763
timestamp 1679581782
transform 1 0 73824 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_770
timestamp 1679581782
transform 1 0 74496 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_777
timestamp 1679581782
transform 1 0 75168 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_784
timestamp 1679581782
transform 1 0 75840 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_791
timestamp 1679581782
transform 1 0 76512 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_798
timestamp 1679581782
transform 1 0 77184 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_805
timestamp 1679581782
transform 1 0 77856 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_812
timestamp 1679581782
transform 1 0 78528 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_819
timestamp 1679581782
transform 1 0 79200 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_826
timestamp 1679581782
transform 1 0 79872 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_833
timestamp 1679581782
transform 1 0 80544 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_840
timestamp 1679581782
transform 1 0 81216 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_847
timestamp 1679581782
transform 1 0 81888 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_854
timestamp 1679581782
transform 1 0 82560 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_861
timestamp 1679581782
transform 1 0 83232 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_868
timestamp 1679581782
transform 1 0 83904 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_875
timestamp 1679581782
transform 1 0 84576 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_882
timestamp 1679581782
transform 1 0 85248 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_889
timestamp 1679581782
transform 1 0 85920 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_896
timestamp 1679581782
transform 1 0 86592 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_903
timestamp 1679581782
transform 1 0 87264 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_910
timestamp 1679581782
transform 1 0 87936 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_917
timestamp 1679581782
transform 1 0 88608 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_924
timestamp 1679581782
transform 1 0 89280 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_931
timestamp 1679581782
transform 1 0 89952 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_938
timestamp 1679581782
transform 1 0 90624 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_945
timestamp 1679581782
transform 1 0 91296 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_952
timestamp 1679581782
transform 1 0 91968 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_959
timestamp 1679581782
transform 1 0 92640 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_966
timestamp 1679581782
transform 1 0 93312 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_973
timestamp 1679581782
transform 1 0 93984 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_980
timestamp 1679581782
transform 1 0 94656 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_987
timestamp 1679581782
transform 1 0 95328 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_994
timestamp 1679581782
transform 1 0 96000 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_1001
timestamp 1679581782
transform 1 0 96672 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_1008
timestamp 1679581782
transform 1 0 97344 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_1015
timestamp 1679581782
transform 1 0 98016 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_1022
timestamp 1679581782
transform 1 0 98688 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_0
timestamp 1679581782
transform 1 0 576 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_7
timestamp 1679581782
transform 1 0 1248 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_14
timestamp 1679581782
transform 1 0 1920 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_21
timestamp 1679581782
transform 1 0 2592 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_28
timestamp 1679581782
transform 1 0 3264 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_35
timestamp 1679581782
transform 1 0 3936 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_42
timestamp 1679581782
transform 1 0 4608 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_49
timestamp 1679581782
transform 1 0 5280 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_56
timestamp 1679581782
transform 1 0 5952 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_63
timestamp 1679581782
transform 1 0 6624 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_70
timestamp 1679581782
transform 1 0 7296 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_77
timestamp 1679581782
transform 1 0 7968 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_84
timestamp 1679581782
transform 1 0 8640 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_91
timestamp 1679581782
transform 1 0 9312 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_98
timestamp 1679581782
transform 1 0 9984 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_105
timestamp 1679581782
transform 1 0 10656 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_112
timestamp 1679581782
transform 1 0 11328 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_119
timestamp 1679581782
transform 1 0 12000 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_126
timestamp 1679581782
transform 1 0 12672 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_133
timestamp 1679581782
transform 1 0 13344 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_140
timestamp 1679581782
transform 1 0 14016 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_147
timestamp 1679581782
transform 1 0 14688 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_154
timestamp 1679581782
transform 1 0 15360 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_161
timestamp 1679581782
transform 1 0 16032 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_168
timestamp 1679581782
transform 1 0 16704 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_175
timestamp 1679581782
transform 1 0 17376 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_182
timestamp 1679581782
transform 1 0 18048 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_189
timestamp 1679581782
transform 1 0 18720 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_196
timestamp 1679581782
transform 1 0 19392 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_203
timestamp 1679581782
transform 1 0 20064 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_210
timestamp 1679581782
transform 1 0 20736 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_217
timestamp 1679581782
transform 1 0 21408 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_224
timestamp 1679581782
transform 1 0 22080 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_231
timestamp 1679581782
transform 1 0 22752 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_238
timestamp 1679581782
transform 1 0 23424 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_245
timestamp 1679581782
transform 1 0 24096 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_252
timestamp 1679581782
transform 1 0 24768 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_259
timestamp 1679581782
transform 1 0 25440 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_266
timestamp 1679581782
transform 1 0 26112 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_273
timestamp 1679581782
transform 1 0 26784 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_280
timestamp 1679581782
transform 1 0 27456 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_287
timestamp 1679581782
transform 1 0 28128 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_294
timestamp 1679581782
transform 1 0 28800 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_301
timestamp 1679581782
transform 1 0 29472 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_308
timestamp 1679581782
transform 1 0 30144 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_315
timestamp 1679581782
transform 1 0 30816 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_322
timestamp 1679581782
transform 1 0 31488 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_329
timestamp 1679581782
transform 1 0 32160 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_336
timestamp 1679581782
transform 1 0 32832 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_343
timestamp 1679581782
transform 1 0 33504 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_350
timestamp 1679581782
transform 1 0 34176 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_357
timestamp 1679581782
transform 1 0 34848 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_364
timestamp 1679581782
transform 1 0 35520 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_371
timestamp 1679581782
transform 1 0 36192 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_378
timestamp 1679581782
transform 1 0 36864 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_385
timestamp 1679581782
transform 1 0 37536 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_392
timestamp 1679581782
transform 1 0 38208 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_399
timestamp 1679581782
transform 1 0 38880 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_406
timestamp 1679581782
transform 1 0 39552 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_413
timestamp 1679581782
transform 1 0 40224 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_420
timestamp 1679581782
transform 1 0 40896 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_427
timestamp 1679581782
transform 1 0 41568 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_434
timestamp 1679581782
transform 1 0 42240 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_441
timestamp 1679581782
transform 1 0 42912 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_448
timestamp 1679581782
transform 1 0 43584 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_455
timestamp 1679581782
transform 1 0 44256 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_462
timestamp 1679581782
transform 1 0 44928 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_469
timestamp 1679581782
transform 1 0 45600 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_476
timestamp 1679581782
transform 1 0 46272 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_483
timestamp 1679581782
transform 1 0 46944 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_490
timestamp 1679581782
transform 1 0 47616 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_497
timestamp 1679581782
transform 1 0 48288 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_504
timestamp 1679581782
transform 1 0 48960 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_511
timestamp 1679581782
transform 1 0 49632 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_518
timestamp 1679581782
transform 1 0 50304 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_525
timestamp 1679581782
transform 1 0 50976 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_532
timestamp 1679581782
transform 1 0 51648 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_539
timestamp 1679581782
transform 1 0 52320 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_546
timestamp 1679581782
transform 1 0 52992 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_553
timestamp 1679581782
transform 1 0 53664 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_560
timestamp 1679581782
transform 1 0 54336 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_567
timestamp 1679581782
transform 1 0 55008 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_574
timestamp 1679581782
transform 1 0 55680 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_581
timestamp 1679581782
transform 1 0 56352 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_588
timestamp 1679581782
transform 1 0 57024 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_595
timestamp 1679581782
transform 1 0 57696 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_602
timestamp 1679581782
transform 1 0 58368 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_609
timestamp 1679581782
transform 1 0 59040 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_616
timestamp 1679581782
transform 1 0 59712 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_623
timestamp 1679581782
transform 1 0 60384 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_630
timestamp 1679581782
transform 1 0 61056 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_637
timestamp 1679581782
transform 1 0 61728 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_644
timestamp 1679581782
transform 1 0 62400 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_651
timestamp 1679581782
transform 1 0 63072 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_658
timestamp 1679581782
transform 1 0 63744 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_665
timestamp 1679581782
transform 1 0 64416 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_672
timestamp 1679581782
transform 1 0 65088 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_679
timestamp 1679581782
transform 1 0 65760 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_686
timestamp 1679581782
transform 1 0 66432 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_693
timestamp 1679581782
transform 1 0 67104 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_700
timestamp 1679581782
transform 1 0 67776 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_707
timestamp 1679581782
transform 1 0 68448 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_714
timestamp 1679581782
transform 1 0 69120 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_721
timestamp 1679581782
transform 1 0 69792 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_728
timestamp 1679581782
transform 1 0 70464 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_735
timestamp 1679581782
transform 1 0 71136 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_742
timestamp 1679581782
transform 1 0 71808 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_749
timestamp 1679581782
transform 1 0 72480 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_756
timestamp 1679581782
transform 1 0 73152 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_763
timestamp 1679581782
transform 1 0 73824 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_770
timestamp 1679581782
transform 1 0 74496 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_777
timestamp 1679581782
transform 1 0 75168 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_784
timestamp 1679581782
transform 1 0 75840 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_791
timestamp 1679581782
transform 1 0 76512 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_798
timestamp 1679581782
transform 1 0 77184 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_805
timestamp 1679581782
transform 1 0 77856 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_812
timestamp 1679581782
transform 1 0 78528 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_819
timestamp 1679581782
transform 1 0 79200 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_826
timestamp 1679581782
transform 1 0 79872 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_833
timestamp 1679581782
transform 1 0 80544 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_840
timestamp 1679581782
transform 1 0 81216 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_847
timestamp 1679581782
transform 1 0 81888 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_854
timestamp 1679581782
transform 1 0 82560 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_861
timestamp 1679581782
transform 1 0 83232 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_868
timestamp 1679581782
transform 1 0 83904 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_875
timestamp 1679581782
transform 1 0 84576 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_882
timestamp 1679581782
transform 1 0 85248 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_889
timestamp 1679581782
transform 1 0 85920 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_896
timestamp 1679581782
transform 1 0 86592 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_903
timestamp 1679581782
transform 1 0 87264 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_910
timestamp 1679581782
transform 1 0 87936 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_917
timestamp 1679581782
transform 1 0 88608 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_924
timestamp 1679581782
transform 1 0 89280 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_931
timestamp 1679581782
transform 1 0 89952 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_938
timestamp 1679581782
transform 1 0 90624 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_945
timestamp 1679581782
transform 1 0 91296 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_952
timestamp 1679581782
transform 1 0 91968 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_959
timestamp 1679581782
transform 1 0 92640 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_966
timestamp 1679581782
transform 1 0 93312 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_973
timestamp 1679581782
transform 1 0 93984 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_980
timestamp 1679581782
transform 1 0 94656 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_987
timestamp 1679581782
transform 1 0 95328 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_994
timestamp 1679581782
transform 1 0 96000 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_1001
timestamp 1679581782
transform 1 0 96672 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_1008
timestamp 1679581782
transform 1 0 97344 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_1015
timestamp 1679581782
transform 1 0 98016 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_1022
timestamp 1679581782
transform 1 0 98688 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_4
timestamp 1679581782
transform 1 0 960 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_11
timestamp 1679581782
transform 1 0 1632 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_18
timestamp 1679581782
transform 1 0 2304 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_25
timestamp 1679581782
transform 1 0 2976 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_32
timestamp 1679581782
transform 1 0 3648 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_39
timestamp 1679581782
transform 1 0 4320 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_46
timestamp 1679581782
transform 1 0 4992 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_53
timestamp 1679581782
transform 1 0 5664 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_60
timestamp 1679581782
transform 1 0 6336 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_67
timestamp 1679581782
transform 1 0 7008 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_74
timestamp 1679581782
transform 1 0 7680 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_81
timestamp 1679581782
transform 1 0 8352 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_88
timestamp 1679581782
transform 1 0 9024 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_95
timestamp 1679581782
transform 1 0 9696 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_102
timestamp 1679581782
transform 1 0 10368 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_109
timestamp 1679581782
transform 1 0 11040 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_116
timestamp 1679581782
transform 1 0 11712 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_123
timestamp 1679581782
transform 1 0 12384 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_130
timestamp 1679581782
transform 1 0 13056 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_137
timestamp 1679581782
transform 1 0 13728 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_144
timestamp 1679581782
transform 1 0 14400 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_151
timestamp 1679581782
transform 1 0 15072 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_158
timestamp 1679581782
transform 1 0 15744 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_165
timestamp 1679581782
transform 1 0 16416 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_172
timestamp 1679581782
transform 1 0 17088 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_179
timestamp 1679581782
transform 1 0 17760 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_186
timestamp 1679581782
transform 1 0 18432 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_193
timestamp 1679581782
transform 1 0 19104 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_200
timestamp 1679581782
transform 1 0 19776 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_207
timestamp 1679581782
transform 1 0 20448 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_214
timestamp 1679581782
transform 1 0 21120 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_221
timestamp 1679581782
transform 1 0 21792 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_228
timestamp 1679581782
transform 1 0 22464 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_235
timestamp 1679581782
transform 1 0 23136 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_242
timestamp 1679581782
transform 1 0 23808 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_249
timestamp 1679581782
transform 1 0 24480 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_256
timestamp 1679581782
transform 1 0 25152 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_263
timestamp 1679581782
transform 1 0 25824 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_270
timestamp 1679581782
transform 1 0 26496 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_277
timestamp 1679581782
transform 1 0 27168 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_284
timestamp 1679581782
transform 1 0 27840 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_291
timestamp 1679581782
transform 1 0 28512 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_298
timestamp 1679581782
transform 1 0 29184 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_305
timestamp 1679581782
transform 1 0 29856 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_312
timestamp 1679581782
transform 1 0 30528 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_319
timestamp 1679581782
transform 1 0 31200 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_326
timestamp 1679581782
transform 1 0 31872 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_333
timestamp 1679581782
transform 1 0 32544 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_340
timestamp 1679581782
transform 1 0 33216 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_347
timestamp 1679581782
transform 1 0 33888 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_354
timestamp 1679581782
transform 1 0 34560 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_361
timestamp 1679581782
transform 1 0 35232 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_368
timestamp 1679581782
transform 1 0 35904 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_375
timestamp 1679581782
transform 1 0 36576 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_382
timestamp 1679581782
transform 1 0 37248 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_389
timestamp 1679581782
transform 1 0 37920 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_396
timestamp 1679581782
transform 1 0 38592 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_403
timestamp 1679581782
transform 1 0 39264 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_410
timestamp 1679581782
transform 1 0 39936 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_417
timestamp 1679581782
transform 1 0 40608 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_424
timestamp 1679581782
transform 1 0 41280 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_431
timestamp 1679581782
transform 1 0 41952 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_438
timestamp 1679581782
transform 1 0 42624 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_445
timestamp 1679581782
transform 1 0 43296 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_452
timestamp 1679581782
transform 1 0 43968 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_459
timestamp 1679581782
transform 1 0 44640 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_466
timestamp 1679581782
transform 1 0 45312 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_473
timestamp 1679581782
transform 1 0 45984 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_480
timestamp 1679581782
transform 1 0 46656 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_487
timestamp 1679581782
transform 1 0 47328 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_494
timestamp 1679581782
transform 1 0 48000 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_501
timestamp 1679581782
transform 1 0 48672 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_508
timestamp 1679581782
transform 1 0 49344 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_515
timestamp 1679581782
transform 1 0 50016 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_522
timestamp 1679581782
transform 1 0 50688 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_529
timestamp 1679581782
transform 1 0 51360 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_536
timestamp 1679581782
transform 1 0 52032 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_543
timestamp 1679581782
transform 1 0 52704 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_550
timestamp 1679581782
transform 1 0 53376 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_557
timestamp 1679581782
transform 1 0 54048 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_564
timestamp 1679581782
transform 1 0 54720 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_571
timestamp 1679581782
transform 1 0 55392 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_578
timestamp 1679581782
transform 1 0 56064 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_585
timestamp 1679581782
transform 1 0 56736 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_592
timestamp 1679581782
transform 1 0 57408 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_599
timestamp 1679581782
transform 1 0 58080 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_606
timestamp 1679581782
transform 1 0 58752 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_613
timestamp 1679581782
transform 1 0 59424 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_620
timestamp 1679581782
transform 1 0 60096 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_627
timestamp 1679581782
transform 1 0 60768 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_634
timestamp 1679581782
transform 1 0 61440 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_641
timestamp 1679581782
transform 1 0 62112 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_648
timestamp 1679581782
transform 1 0 62784 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_655
timestamp 1679581782
transform 1 0 63456 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_662
timestamp 1679581782
transform 1 0 64128 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_669
timestamp 1679581782
transform 1 0 64800 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_676
timestamp 1679581782
transform 1 0 65472 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_683
timestamp 1679581782
transform 1 0 66144 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_690
timestamp 1679581782
transform 1 0 66816 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_697
timestamp 1679581782
transform 1 0 67488 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_704
timestamp 1679581782
transform 1 0 68160 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_711
timestamp 1679581782
transform 1 0 68832 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_718
timestamp 1679581782
transform 1 0 69504 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_725
timestamp 1679581782
transform 1 0 70176 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_732
timestamp 1679581782
transform 1 0 70848 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_739
timestamp 1679581782
transform 1 0 71520 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_746
timestamp 1679581782
transform 1 0 72192 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_753
timestamp 1679581782
transform 1 0 72864 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_760
timestamp 1679581782
transform 1 0 73536 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_767
timestamp 1679581782
transform 1 0 74208 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_774
timestamp 1679581782
transform 1 0 74880 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_781
timestamp 1679581782
transform 1 0 75552 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_788
timestamp 1679581782
transform 1 0 76224 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_795
timestamp 1679581782
transform 1 0 76896 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_802
timestamp 1679581782
transform 1 0 77568 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_809
timestamp 1679581782
transform 1 0 78240 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_816
timestamp 1679581782
transform 1 0 78912 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_823
timestamp 1679581782
transform 1 0 79584 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_830
timestamp 1679581782
transform 1 0 80256 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_837
timestamp 1679581782
transform 1 0 80928 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_844
timestamp 1679581782
transform 1 0 81600 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_851
timestamp 1679581782
transform 1 0 82272 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_858
timestamp 1679581782
transform 1 0 82944 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_865
timestamp 1679581782
transform 1 0 83616 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_872
timestamp 1679581782
transform 1 0 84288 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_879
timestamp 1679581782
transform 1 0 84960 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_886
timestamp 1679581782
transform 1 0 85632 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_893
timestamp 1679581782
transform 1 0 86304 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_900
timestamp 1679581782
transform 1 0 86976 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_907
timestamp 1679581782
transform 1 0 87648 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_914
timestamp 1679581782
transform 1 0 88320 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_921
timestamp 1679581782
transform 1 0 88992 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_928
timestamp 1679581782
transform 1 0 89664 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_935
timestamp 1679581782
transform 1 0 90336 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_942
timestamp 1679581782
transform 1 0 91008 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_949
timestamp 1679581782
transform 1 0 91680 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_956
timestamp 1679581782
transform 1 0 92352 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_963
timestamp 1679581782
transform 1 0 93024 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_970
timestamp 1679581782
transform 1 0 93696 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_977
timestamp 1679581782
transform 1 0 94368 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_984
timestamp 1679581782
transform 1 0 95040 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_991
timestamp 1679581782
transform 1 0 95712 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_998
timestamp 1679581782
transform 1 0 96384 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_1005
timestamp 1679581782
transform 1 0 97056 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_1012
timestamp 1679581782
transform 1 0 97728 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_1019
timestamp 1679581782
transform 1 0 98400 0 1 74844
box -48 -56 720 834
use sg13g2_fill_2  FILLER_98_1026
timestamp 1677580104
transform 1 0 99072 0 1 74844
box -48 -56 240 834
use sg13g2_fill_1  FILLER_98_1028
timestamp 1677579658
transform 1 0 99264 0 1 74844
box -48 -56 144 834
use sg13g2_decap_8  FILLER_99_0
timestamp 1679581782
transform 1 0 576 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_7
timestamp 1679581782
transform 1 0 1248 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_14
timestamp 1679581782
transform 1 0 1920 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_21
timestamp 1679581782
transform 1 0 2592 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_28
timestamp 1679581782
transform 1 0 3264 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_35
timestamp 1679581782
transform 1 0 3936 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_42
timestamp 1679581782
transform 1 0 4608 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_49
timestamp 1679581782
transform 1 0 5280 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_56
timestamp 1679581782
transform 1 0 5952 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_63
timestamp 1679581782
transform 1 0 6624 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_70
timestamp 1679581782
transform 1 0 7296 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_77
timestamp 1679581782
transform 1 0 7968 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_84
timestamp 1679581782
transform 1 0 8640 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_91
timestamp 1679581782
transform 1 0 9312 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_98
timestamp 1679581782
transform 1 0 9984 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_105
timestamp 1679581782
transform 1 0 10656 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_112
timestamp 1679581782
transform 1 0 11328 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_119
timestamp 1679581782
transform 1 0 12000 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_126
timestamp 1679581782
transform 1 0 12672 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_133
timestamp 1679581782
transform 1 0 13344 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_140
timestamp 1679581782
transform 1 0 14016 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_147
timestamp 1679581782
transform 1 0 14688 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_154
timestamp 1679581782
transform 1 0 15360 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_161
timestamp 1679581782
transform 1 0 16032 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_168
timestamp 1679581782
transform 1 0 16704 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_175
timestamp 1679581782
transform 1 0 17376 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_182
timestamp 1679581782
transform 1 0 18048 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_189
timestamp 1679581782
transform 1 0 18720 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_196
timestamp 1679581782
transform 1 0 19392 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_203
timestamp 1679581782
transform 1 0 20064 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_210
timestamp 1679581782
transform 1 0 20736 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_217
timestamp 1679581782
transform 1 0 21408 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_224
timestamp 1679581782
transform 1 0 22080 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_231
timestamp 1679581782
transform 1 0 22752 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_238
timestamp 1679581782
transform 1 0 23424 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_245
timestamp 1679581782
transform 1 0 24096 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_252
timestamp 1679581782
transform 1 0 24768 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_259
timestamp 1679581782
transform 1 0 25440 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_266
timestamp 1679581782
transform 1 0 26112 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_273
timestamp 1679581782
transform 1 0 26784 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_280
timestamp 1679581782
transform 1 0 27456 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_287
timestamp 1679581782
transform 1 0 28128 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_294
timestamp 1679581782
transform 1 0 28800 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_301
timestamp 1679581782
transform 1 0 29472 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_308
timestamp 1679581782
transform 1 0 30144 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_315
timestamp 1679581782
transform 1 0 30816 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_322
timestamp 1679581782
transform 1 0 31488 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_329
timestamp 1679581782
transform 1 0 32160 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_336
timestamp 1679581782
transform 1 0 32832 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_343
timestamp 1679581782
transform 1 0 33504 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_350
timestamp 1679581782
transform 1 0 34176 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_357
timestamp 1679581782
transform 1 0 34848 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_364
timestamp 1679581782
transform 1 0 35520 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_371
timestamp 1679581782
transform 1 0 36192 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_378
timestamp 1679581782
transform 1 0 36864 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_385
timestamp 1679581782
transform 1 0 37536 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_392
timestamp 1679581782
transform 1 0 38208 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_399
timestamp 1679581782
transform 1 0 38880 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_406
timestamp 1679581782
transform 1 0 39552 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_413
timestamp 1679581782
transform 1 0 40224 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_420
timestamp 1679581782
transform 1 0 40896 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_427
timestamp 1679581782
transform 1 0 41568 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_434
timestamp 1679581782
transform 1 0 42240 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_441
timestamp 1679581782
transform 1 0 42912 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_448
timestamp 1679581782
transform 1 0 43584 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_455
timestamp 1679581782
transform 1 0 44256 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_462
timestamp 1679581782
transform 1 0 44928 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_469
timestamp 1679581782
transform 1 0 45600 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_476
timestamp 1679581782
transform 1 0 46272 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_483
timestamp 1679581782
transform 1 0 46944 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_490
timestamp 1679581782
transform 1 0 47616 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_497
timestamp 1679581782
transform 1 0 48288 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_504
timestamp 1679581782
transform 1 0 48960 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_511
timestamp 1679581782
transform 1 0 49632 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_518
timestamp 1679581782
transform 1 0 50304 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_525
timestamp 1679581782
transform 1 0 50976 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_532
timestamp 1679581782
transform 1 0 51648 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_539
timestamp 1679581782
transform 1 0 52320 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_546
timestamp 1679581782
transform 1 0 52992 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_553
timestamp 1679581782
transform 1 0 53664 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_560
timestamp 1679581782
transform 1 0 54336 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_567
timestamp 1679581782
transform 1 0 55008 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_574
timestamp 1679581782
transform 1 0 55680 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_581
timestamp 1679581782
transform 1 0 56352 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_588
timestamp 1679581782
transform 1 0 57024 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_595
timestamp 1679581782
transform 1 0 57696 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_602
timestamp 1679581782
transform 1 0 58368 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_609
timestamp 1679581782
transform 1 0 59040 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_616
timestamp 1679581782
transform 1 0 59712 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_623
timestamp 1679581782
transform 1 0 60384 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_630
timestamp 1679581782
transform 1 0 61056 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_637
timestamp 1679581782
transform 1 0 61728 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_644
timestamp 1679581782
transform 1 0 62400 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_651
timestamp 1679581782
transform 1 0 63072 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_658
timestamp 1679581782
transform 1 0 63744 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_665
timestamp 1679581782
transform 1 0 64416 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_672
timestamp 1679581782
transform 1 0 65088 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_679
timestamp 1679581782
transform 1 0 65760 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_686
timestamp 1679581782
transform 1 0 66432 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_693
timestamp 1679581782
transform 1 0 67104 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_700
timestamp 1679581782
transform 1 0 67776 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_707
timestamp 1679581782
transform 1 0 68448 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_714
timestamp 1679581782
transform 1 0 69120 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_721
timestamp 1679581782
transform 1 0 69792 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_728
timestamp 1679581782
transform 1 0 70464 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_735
timestamp 1679581782
transform 1 0 71136 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_742
timestamp 1679581782
transform 1 0 71808 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_749
timestamp 1679581782
transform 1 0 72480 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_756
timestamp 1679581782
transform 1 0 73152 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_763
timestamp 1679581782
transform 1 0 73824 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_770
timestamp 1679581782
transform 1 0 74496 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_777
timestamp 1679581782
transform 1 0 75168 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_784
timestamp 1679581782
transform 1 0 75840 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_791
timestamp 1679581782
transform 1 0 76512 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_798
timestamp 1679581782
transform 1 0 77184 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_805
timestamp 1679581782
transform 1 0 77856 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_812
timestamp 1679581782
transform 1 0 78528 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_819
timestamp 1679581782
transform 1 0 79200 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_826
timestamp 1679581782
transform 1 0 79872 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_833
timestamp 1679581782
transform 1 0 80544 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_840
timestamp 1679581782
transform 1 0 81216 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_847
timestamp 1679581782
transform 1 0 81888 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_854
timestamp 1679581782
transform 1 0 82560 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_861
timestamp 1679581782
transform 1 0 83232 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_868
timestamp 1679581782
transform 1 0 83904 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_875
timestamp 1679581782
transform 1 0 84576 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_882
timestamp 1679581782
transform 1 0 85248 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_889
timestamp 1679581782
transform 1 0 85920 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_896
timestamp 1679581782
transform 1 0 86592 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_903
timestamp 1679581782
transform 1 0 87264 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_910
timestamp 1679581782
transform 1 0 87936 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_917
timestamp 1679581782
transform 1 0 88608 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_924
timestamp 1679581782
transform 1 0 89280 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_931
timestamp 1679581782
transform 1 0 89952 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_938
timestamp 1679581782
transform 1 0 90624 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_945
timestamp 1679581782
transform 1 0 91296 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_952
timestamp 1679581782
transform 1 0 91968 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_959
timestamp 1679581782
transform 1 0 92640 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_966
timestamp 1679581782
transform 1 0 93312 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_973
timestamp 1679581782
transform 1 0 93984 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_980
timestamp 1679581782
transform 1 0 94656 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_987
timestamp 1679581782
transform 1 0 95328 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_994
timestamp 1679581782
transform 1 0 96000 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_1001
timestamp 1679581782
transform 1 0 96672 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_1008
timestamp 1679581782
transform 1 0 97344 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_1015
timestamp 1679581782
transform 1 0 98016 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_1022
timestamp 1679581782
transform 1 0 98688 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_0
timestamp 1679581782
transform 1 0 576 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_7
timestamp 1679581782
transform 1 0 1248 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_14
timestamp 1679581782
transform 1 0 1920 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_21
timestamp 1679581782
transform 1 0 2592 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_28
timestamp 1679581782
transform 1 0 3264 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_35
timestamp 1679581782
transform 1 0 3936 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_42
timestamp 1679581782
transform 1 0 4608 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_49
timestamp 1679581782
transform 1 0 5280 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_56
timestamp 1679581782
transform 1 0 5952 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_63
timestamp 1679581782
transform 1 0 6624 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_70
timestamp 1679581782
transform 1 0 7296 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_77
timestamp 1679581782
transform 1 0 7968 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_84
timestamp 1679581782
transform 1 0 8640 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_91
timestamp 1679581782
transform 1 0 9312 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_98
timestamp 1679581782
transform 1 0 9984 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_105
timestamp 1679581782
transform 1 0 10656 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_112
timestamp 1679581782
transform 1 0 11328 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_119
timestamp 1679581782
transform 1 0 12000 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_126
timestamp 1679581782
transform 1 0 12672 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_133
timestamp 1679581782
transform 1 0 13344 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_140
timestamp 1679581782
transform 1 0 14016 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_147
timestamp 1679581782
transform 1 0 14688 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_154
timestamp 1679581782
transform 1 0 15360 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_161
timestamp 1679581782
transform 1 0 16032 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_168
timestamp 1679581782
transform 1 0 16704 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_175
timestamp 1679581782
transform 1 0 17376 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_182
timestamp 1679581782
transform 1 0 18048 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_189
timestamp 1679581782
transform 1 0 18720 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_196
timestamp 1679581782
transform 1 0 19392 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_203
timestamp 1679581782
transform 1 0 20064 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_210
timestamp 1679581782
transform 1 0 20736 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_217
timestamp 1679581782
transform 1 0 21408 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_224
timestamp 1679581782
transform 1 0 22080 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_231
timestamp 1679581782
transform 1 0 22752 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_238
timestamp 1679581782
transform 1 0 23424 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_245
timestamp 1679581782
transform 1 0 24096 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_252
timestamp 1679581782
transform 1 0 24768 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_259
timestamp 1679581782
transform 1 0 25440 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_266
timestamp 1679581782
transform 1 0 26112 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_273
timestamp 1679581782
transform 1 0 26784 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_280
timestamp 1679581782
transform 1 0 27456 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_287
timestamp 1679581782
transform 1 0 28128 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_294
timestamp 1679581782
transform 1 0 28800 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_301
timestamp 1679581782
transform 1 0 29472 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_308
timestamp 1679581782
transform 1 0 30144 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_315
timestamp 1679581782
transform 1 0 30816 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_322
timestamp 1679581782
transform 1 0 31488 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_329
timestamp 1679581782
transform 1 0 32160 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_336
timestamp 1679581782
transform 1 0 32832 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_343
timestamp 1679581782
transform 1 0 33504 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_350
timestamp 1679581782
transform 1 0 34176 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_357
timestamp 1679581782
transform 1 0 34848 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_364
timestamp 1679581782
transform 1 0 35520 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_371
timestamp 1679581782
transform 1 0 36192 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_378
timestamp 1679581782
transform 1 0 36864 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_385
timestamp 1679581782
transform 1 0 37536 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_392
timestamp 1679581782
transform 1 0 38208 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_399
timestamp 1679581782
transform 1 0 38880 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_406
timestamp 1679581782
transform 1 0 39552 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_413
timestamp 1679581782
transform 1 0 40224 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_420
timestamp 1679581782
transform 1 0 40896 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_427
timestamp 1679581782
transform 1 0 41568 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_434
timestamp 1679581782
transform 1 0 42240 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_441
timestamp 1679581782
transform 1 0 42912 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_448
timestamp 1679581782
transform 1 0 43584 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_455
timestamp 1679581782
transform 1 0 44256 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_462
timestamp 1679581782
transform 1 0 44928 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_469
timestamp 1679581782
transform 1 0 45600 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_476
timestamp 1679581782
transform 1 0 46272 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_483
timestamp 1679581782
transform 1 0 46944 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_490
timestamp 1679581782
transform 1 0 47616 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_497
timestamp 1679581782
transform 1 0 48288 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_504
timestamp 1679581782
transform 1 0 48960 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_511
timestamp 1679581782
transform 1 0 49632 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_518
timestamp 1679581782
transform 1 0 50304 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_525
timestamp 1679581782
transform 1 0 50976 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_532
timestamp 1679581782
transform 1 0 51648 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_539
timestamp 1679581782
transform 1 0 52320 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_546
timestamp 1679581782
transform 1 0 52992 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_553
timestamp 1679581782
transform 1 0 53664 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_560
timestamp 1679581782
transform 1 0 54336 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_567
timestamp 1679581782
transform 1 0 55008 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_574
timestamp 1679581782
transform 1 0 55680 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_581
timestamp 1679581782
transform 1 0 56352 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_588
timestamp 1679581782
transform 1 0 57024 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_595
timestamp 1679581782
transform 1 0 57696 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_602
timestamp 1679581782
transform 1 0 58368 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_609
timestamp 1679581782
transform 1 0 59040 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_616
timestamp 1679581782
transform 1 0 59712 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_623
timestamp 1679581782
transform 1 0 60384 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_630
timestamp 1679581782
transform 1 0 61056 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_637
timestamp 1679581782
transform 1 0 61728 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_644
timestamp 1679581782
transform 1 0 62400 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_651
timestamp 1679581782
transform 1 0 63072 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_658
timestamp 1679581782
transform 1 0 63744 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_665
timestamp 1679581782
transform 1 0 64416 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_672
timestamp 1679581782
transform 1 0 65088 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_679
timestamp 1679581782
transform 1 0 65760 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_686
timestamp 1679581782
transform 1 0 66432 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_693
timestamp 1679581782
transform 1 0 67104 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_700
timestamp 1679581782
transform 1 0 67776 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_707
timestamp 1679581782
transform 1 0 68448 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_714
timestamp 1679581782
transform 1 0 69120 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_721
timestamp 1679581782
transform 1 0 69792 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_728
timestamp 1679581782
transform 1 0 70464 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_735
timestamp 1679581782
transform 1 0 71136 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_742
timestamp 1679581782
transform 1 0 71808 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_749
timestamp 1679581782
transform 1 0 72480 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_756
timestamp 1679581782
transform 1 0 73152 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_763
timestamp 1679581782
transform 1 0 73824 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_770
timestamp 1679581782
transform 1 0 74496 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_777
timestamp 1679581782
transform 1 0 75168 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_784
timestamp 1679581782
transform 1 0 75840 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_791
timestamp 1679581782
transform 1 0 76512 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_798
timestamp 1679581782
transform 1 0 77184 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_805
timestamp 1679581782
transform 1 0 77856 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_812
timestamp 1679581782
transform 1 0 78528 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_819
timestamp 1679581782
transform 1 0 79200 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_826
timestamp 1679581782
transform 1 0 79872 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_833
timestamp 1679581782
transform 1 0 80544 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_840
timestamp 1679581782
transform 1 0 81216 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_847
timestamp 1679581782
transform 1 0 81888 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_854
timestamp 1679581782
transform 1 0 82560 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_861
timestamp 1679581782
transform 1 0 83232 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_868
timestamp 1679581782
transform 1 0 83904 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_875
timestamp 1679581782
transform 1 0 84576 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_882
timestamp 1679581782
transform 1 0 85248 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_889
timestamp 1679581782
transform 1 0 85920 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_896
timestamp 1679581782
transform 1 0 86592 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_903
timestamp 1679581782
transform 1 0 87264 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_910
timestamp 1679581782
transform 1 0 87936 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_917
timestamp 1679581782
transform 1 0 88608 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_924
timestamp 1679581782
transform 1 0 89280 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_931
timestamp 1679581782
transform 1 0 89952 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_938
timestamp 1679581782
transform 1 0 90624 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_945
timestamp 1679581782
transform 1 0 91296 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_952
timestamp 1679581782
transform 1 0 91968 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_959
timestamp 1679581782
transform 1 0 92640 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_966
timestamp 1679581782
transform 1 0 93312 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_973
timestamp 1679581782
transform 1 0 93984 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_980
timestamp 1679581782
transform 1 0 94656 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_987
timestamp 1679581782
transform 1 0 95328 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_994
timestamp 1679581782
transform 1 0 96000 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_1001
timestamp 1679581782
transform 1 0 96672 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_1008
timestamp 1679581782
transform 1 0 97344 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_1015
timestamp 1679581782
transform 1 0 98016 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_1022
timestamp 1679581782
transform 1 0 98688 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_0
timestamp 1679581782
transform 1 0 576 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_7
timestamp 1679581782
transform 1 0 1248 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_14
timestamp 1679581782
transform 1 0 1920 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_21
timestamp 1679581782
transform 1 0 2592 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_28
timestamp 1679581782
transform 1 0 3264 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_35
timestamp 1679581782
transform 1 0 3936 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_42
timestamp 1679581782
transform 1 0 4608 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_49
timestamp 1679581782
transform 1 0 5280 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_56
timestamp 1679581782
transform 1 0 5952 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_63
timestamp 1679581782
transform 1 0 6624 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_70
timestamp 1679581782
transform 1 0 7296 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_77
timestamp 1679581782
transform 1 0 7968 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_84
timestamp 1679581782
transform 1 0 8640 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_91
timestamp 1679581782
transform 1 0 9312 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_98
timestamp 1679581782
transform 1 0 9984 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_105
timestamp 1679581782
transform 1 0 10656 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_112
timestamp 1679581782
transform 1 0 11328 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_119
timestamp 1679581782
transform 1 0 12000 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_126
timestamp 1679581782
transform 1 0 12672 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_133
timestamp 1679581782
transform 1 0 13344 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_140
timestamp 1679581782
transform 1 0 14016 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_147
timestamp 1679581782
transform 1 0 14688 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_154
timestamp 1679581782
transform 1 0 15360 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_161
timestamp 1679581782
transform 1 0 16032 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_168
timestamp 1679581782
transform 1 0 16704 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_175
timestamp 1679581782
transform 1 0 17376 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_182
timestamp 1679581782
transform 1 0 18048 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_189
timestamp 1679581782
transform 1 0 18720 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_196
timestamp 1679581782
transform 1 0 19392 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_203
timestamp 1679581782
transform 1 0 20064 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_210
timestamp 1679581782
transform 1 0 20736 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_217
timestamp 1679581782
transform 1 0 21408 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_224
timestamp 1679581782
transform 1 0 22080 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_231
timestamp 1679581782
transform 1 0 22752 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_238
timestamp 1679581782
transform 1 0 23424 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_245
timestamp 1679581782
transform 1 0 24096 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_252
timestamp 1679581782
transform 1 0 24768 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_259
timestamp 1679581782
transform 1 0 25440 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_266
timestamp 1679581782
transform 1 0 26112 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_273
timestamp 1679581782
transform 1 0 26784 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_280
timestamp 1679581782
transform 1 0 27456 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_287
timestamp 1679581782
transform 1 0 28128 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_294
timestamp 1679581782
transform 1 0 28800 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_301
timestamp 1679581782
transform 1 0 29472 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_308
timestamp 1679581782
transform 1 0 30144 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_315
timestamp 1679581782
transform 1 0 30816 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_322
timestamp 1679581782
transform 1 0 31488 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_329
timestamp 1679581782
transform 1 0 32160 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_336
timestamp 1679581782
transform 1 0 32832 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_343
timestamp 1679581782
transform 1 0 33504 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_350
timestamp 1679581782
transform 1 0 34176 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_357
timestamp 1679581782
transform 1 0 34848 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_364
timestamp 1679581782
transform 1 0 35520 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_371
timestamp 1679581782
transform 1 0 36192 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_378
timestamp 1679581782
transform 1 0 36864 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_385
timestamp 1679581782
transform 1 0 37536 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_392
timestamp 1679581782
transform 1 0 38208 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_399
timestamp 1679581782
transform 1 0 38880 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_406
timestamp 1679581782
transform 1 0 39552 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_413
timestamp 1679581782
transform 1 0 40224 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_420
timestamp 1679581782
transform 1 0 40896 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_427
timestamp 1679581782
transform 1 0 41568 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_434
timestamp 1679581782
transform 1 0 42240 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_441
timestamp 1679581782
transform 1 0 42912 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_448
timestamp 1679581782
transform 1 0 43584 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_455
timestamp 1679581782
transform 1 0 44256 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_462
timestamp 1679581782
transform 1 0 44928 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_469
timestamp 1679581782
transform 1 0 45600 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_476
timestamp 1679581782
transform 1 0 46272 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_483
timestamp 1679581782
transform 1 0 46944 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_490
timestamp 1679581782
transform 1 0 47616 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_497
timestamp 1679581782
transform 1 0 48288 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_504
timestamp 1679581782
transform 1 0 48960 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_511
timestamp 1679581782
transform 1 0 49632 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_518
timestamp 1679581782
transform 1 0 50304 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_525
timestamp 1679581782
transform 1 0 50976 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_532
timestamp 1679581782
transform 1 0 51648 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_539
timestamp 1679581782
transform 1 0 52320 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_546
timestamp 1679581782
transform 1 0 52992 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_553
timestamp 1679581782
transform 1 0 53664 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_560
timestamp 1679581782
transform 1 0 54336 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_567
timestamp 1679581782
transform 1 0 55008 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_574
timestamp 1679581782
transform 1 0 55680 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_581
timestamp 1679581782
transform 1 0 56352 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_588
timestamp 1679581782
transform 1 0 57024 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_595
timestamp 1679581782
transform 1 0 57696 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_602
timestamp 1679581782
transform 1 0 58368 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_609
timestamp 1679581782
transform 1 0 59040 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_616
timestamp 1679581782
transform 1 0 59712 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_623
timestamp 1679581782
transform 1 0 60384 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_630
timestamp 1679581782
transform 1 0 61056 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_637
timestamp 1679581782
transform 1 0 61728 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_644
timestamp 1679581782
transform 1 0 62400 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_651
timestamp 1679581782
transform 1 0 63072 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_658
timestamp 1679581782
transform 1 0 63744 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_665
timestamp 1679581782
transform 1 0 64416 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_672
timestamp 1679581782
transform 1 0 65088 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_679
timestamp 1679581782
transform 1 0 65760 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_686
timestamp 1679581782
transform 1 0 66432 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_693
timestamp 1679581782
transform 1 0 67104 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_700
timestamp 1679581782
transform 1 0 67776 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_707
timestamp 1679581782
transform 1 0 68448 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_714
timestamp 1679581782
transform 1 0 69120 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_721
timestamp 1679581782
transform 1 0 69792 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_728
timestamp 1679581782
transform 1 0 70464 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_735
timestamp 1679581782
transform 1 0 71136 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_742
timestamp 1679581782
transform 1 0 71808 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_749
timestamp 1679581782
transform 1 0 72480 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_756
timestamp 1679581782
transform 1 0 73152 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_763
timestamp 1679581782
transform 1 0 73824 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_770
timestamp 1679581782
transform 1 0 74496 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_777
timestamp 1679581782
transform 1 0 75168 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_784
timestamp 1679581782
transform 1 0 75840 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_791
timestamp 1679581782
transform 1 0 76512 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_798
timestamp 1679581782
transform 1 0 77184 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_805
timestamp 1679581782
transform 1 0 77856 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_812
timestamp 1679581782
transform 1 0 78528 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_819
timestamp 1679581782
transform 1 0 79200 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_826
timestamp 1679581782
transform 1 0 79872 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_833
timestamp 1679581782
transform 1 0 80544 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_840
timestamp 1679581782
transform 1 0 81216 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_847
timestamp 1679581782
transform 1 0 81888 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_854
timestamp 1679581782
transform 1 0 82560 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_861
timestamp 1679581782
transform 1 0 83232 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_868
timestamp 1679581782
transform 1 0 83904 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_875
timestamp 1679581782
transform 1 0 84576 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_882
timestamp 1679581782
transform 1 0 85248 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_889
timestamp 1679581782
transform 1 0 85920 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_896
timestamp 1679581782
transform 1 0 86592 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_903
timestamp 1679581782
transform 1 0 87264 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_910
timestamp 1679581782
transform 1 0 87936 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_917
timestamp 1679581782
transform 1 0 88608 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_924
timestamp 1679581782
transform 1 0 89280 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_931
timestamp 1679581782
transform 1 0 89952 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_938
timestamp 1679581782
transform 1 0 90624 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_945
timestamp 1679581782
transform 1 0 91296 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_952
timestamp 1679581782
transform 1 0 91968 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_959
timestamp 1679581782
transform 1 0 92640 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_966
timestamp 1679581782
transform 1 0 93312 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_973
timestamp 1679581782
transform 1 0 93984 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_980
timestamp 1679581782
transform 1 0 94656 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_987
timestamp 1679581782
transform 1 0 95328 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_994
timestamp 1679581782
transform 1 0 96000 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_1001
timestamp 1679581782
transform 1 0 96672 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_1008
timestamp 1679581782
transform 1 0 97344 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_1015
timestamp 1679581782
transform 1 0 98016 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_1022
timestamp 1679581782
transform 1 0 98688 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_0
timestamp 1679581782
transform 1 0 576 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_7
timestamp 1679581782
transform 1 0 1248 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_14
timestamp 1679581782
transform 1 0 1920 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_21
timestamp 1679581782
transform 1 0 2592 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_28
timestamp 1679581782
transform 1 0 3264 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_35
timestamp 1679581782
transform 1 0 3936 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_42
timestamp 1679581782
transform 1 0 4608 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_49
timestamp 1679581782
transform 1 0 5280 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_56
timestamp 1679581782
transform 1 0 5952 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_63
timestamp 1679581782
transform 1 0 6624 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_70
timestamp 1679581782
transform 1 0 7296 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_77
timestamp 1679581782
transform 1 0 7968 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_84
timestamp 1679581782
transform 1 0 8640 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_91
timestamp 1679581782
transform 1 0 9312 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_98
timestamp 1679581782
transform 1 0 9984 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_105
timestamp 1679581782
transform 1 0 10656 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_112
timestamp 1679581782
transform 1 0 11328 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_119
timestamp 1679581782
transform 1 0 12000 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_126
timestamp 1679581782
transform 1 0 12672 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_133
timestamp 1679581782
transform 1 0 13344 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_140
timestamp 1679581782
transform 1 0 14016 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_147
timestamp 1679581782
transform 1 0 14688 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_154
timestamp 1679581782
transform 1 0 15360 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_161
timestamp 1679581782
transform 1 0 16032 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_168
timestamp 1679581782
transform 1 0 16704 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_175
timestamp 1679581782
transform 1 0 17376 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_182
timestamp 1679581782
transform 1 0 18048 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_189
timestamp 1679581782
transform 1 0 18720 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_196
timestamp 1679581782
transform 1 0 19392 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_203
timestamp 1679581782
transform 1 0 20064 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_210
timestamp 1679581782
transform 1 0 20736 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_217
timestamp 1679581782
transform 1 0 21408 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_224
timestamp 1679581782
transform 1 0 22080 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_231
timestamp 1679581782
transform 1 0 22752 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_238
timestamp 1679581782
transform 1 0 23424 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_245
timestamp 1679581782
transform 1 0 24096 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_252
timestamp 1679581782
transform 1 0 24768 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_259
timestamp 1679581782
transform 1 0 25440 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_266
timestamp 1679581782
transform 1 0 26112 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_273
timestamp 1679581782
transform 1 0 26784 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_280
timestamp 1679581782
transform 1 0 27456 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_287
timestamp 1679581782
transform 1 0 28128 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_294
timestamp 1679581782
transform 1 0 28800 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_301
timestamp 1679581782
transform 1 0 29472 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_308
timestamp 1679581782
transform 1 0 30144 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_315
timestamp 1679581782
transform 1 0 30816 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_322
timestamp 1679581782
transform 1 0 31488 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_329
timestamp 1679581782
transform 1 0 32160 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_336
timestamp 1679581782
transform 1 0 32832 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_343
timestamp 1679581782
transform 1 0 33504 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_350
timestamp 1679581782
transform 1 0 34176 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_357
timestamp 1679581782
transform 1 0 34848 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_364
timestamp 1679581782
transform 1 0 35520 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_371
timestamp 1679581782
transform 1 0 36192 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_378
timestamp 1679581782
transform 1 0 36864 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_385
timestamp 1679581782
transform 1 0 37536 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_392
timestamp 1679581782
transform 1 0 38208 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_399
timestamp 1679581782
transform 1 0 38880 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_406
timestamp 1679581782
transform 1 0 39552 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_413
timestamp 1679581782
transform 1 0 40224 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_420
timestamp 1679581782
transform 1 0 40896 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_427
timestamp 1679581782
transform 1 0 41568 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_434
timestamp 1679581782
transform 1 0 42240 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_441
timestamp 1679581782
transform 1 0 42912 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_448
timestamp 1679581782
transform 1 0 43584 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_455
timestamp 1679581782
transform 1 0 44256 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_462
timestamp 1679581782
transform 1 0 44928 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_469
timestamp 1679581782
transform 1 0 45600 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_476
timestamp 1679581782
transform 1 0 46272 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_483
timestamp 1679581782
transform 1 0 46944 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_490
timestamp 1679581782
transform 1 0 47616 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_497
timestamp 1679581782
transform 1 0 48288 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_504
timestamp 1679581782
transform 1 0 48960 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_511
timestamp 1679581782
transform 1 0 49632 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_518
timestamp 1679581782
transform 1 0 50304 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_525
timestamp 1679581782
transform 1 0 50976 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_532
timestamp 1679581782
transform 1 0 51648 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_539
timestamp 1679581782
transform 1 0 52320 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_546
timestamp 1679581782
transform 1 0 52992 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_553
timestamp 1679581782
transform 1 0 53664 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_560
timestamp 1679581782
transform 1 0 54336 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_567
timestamp 1679581782
transform 1 0 55008 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_574
timestamp 1679581782
transform 1 0 55680 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_581
timestamp 1679581782
transform 1 0 56352 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_588
timestamp 1679581782
transform 1 0 57024 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_595
timestamp 1679581782
transform 1 0 57696 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_602
timestamp 1679581782
transform 1 0 58368 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_609
timestamp 1679581782
transform 1 0 59040 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_616
timestamp 1679581782
transform 1 0 59712 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_623
timestamp 1679581782
transform 1 0 60384 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_630
timestamp 1679581782
transform 1 0 61056 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_637
timestamp 1679581782
transform 1 0 61728 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_644
timestamp 1679581782
transform 1 0 62400 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_651
timestamp 1679581782
transform 1 0 63072 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_658
timestamp 1679581782
transform 1 0 63744 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_665
timestamp 1679581782
transform 1 0 64416 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_672
timestamp 1679581782
transform 1 0 65088 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_679
timestamp 1679581782
transform 1 0 65760 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_686
timestamp 1679581782
transform 1 0 66432 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_693
timestamp 1679581782
transform 1 0 67104 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_700
timestamp 1679581782
transform 1 0 67776 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_707
timestamp 1679581782
transform 1 0 68448 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_714
timestamp 1679581782
transform 1 0 69120 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_721
timestamp 1679581782
transform 1 0 69792 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_728
timestamp 1679581782
transform 1 0 70464 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_735
timestamp 1679581782
transform 1 0 71136 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_742
timestamp 1679581782
transform 1 0 71808 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_749
timestamp 1679581782
transform 1 0 72480 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_756
timestamp 1679581782
transform 1 0 73152 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_763
timestamp 1679581782
transform 1 0 73824 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_770
timestamp 1679581782
transform 1 0 74496 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_777
timestamp 1679581782
transform 1 0 75168 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_784
timestamp 1679581782
transform 1 0 75840 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_791
timestamp 1679581782
transform 1 0 76512 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_798
timestamp 1679581782
transform 1 0 77184 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_805
timestamp 1679581782
transform 1 0 77856 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_812
timestamp 1679581782
transform 1 0 78528 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_819
timestamp 1679581782
transform 1 0 79200 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_826
timestamp 1679581782
transform 1 0 79872 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_833
timestamp 1679581782
transform 1 0 80544 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_840
timestamp 1679581782
transform 1 0 81216 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_847
timestamp 1679581782
transform 1 0 81888 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_854
timestamp 1679581782
transform 1 0 82560 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_861
timestamp 1679581782
transform 1 0 83232 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_868
timestamp 1679581782
transform 1 0 83904 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_875
timestamp 1679581782
transform 1 0 84576 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_882
timestamp 1679581782
transform 1 0 85248 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_889
timestamp 1679581782
transform 1 0 85920 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_896
timestamp 1679581782
transform 1 0 86592 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_903
timestamp 1679581782
transform 1 0 87264 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_910
timestamp 1679581782
transform 1 0 87936 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_917
timestamp 1679581782
transform 1 0 88608 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_924
timestamp 1679581782
transform 1 0 89280 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_931
timestamp 1679581782
transform 1 0 89952 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_938
timestamp 1679581782
transform 1 0 90624 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_945
timestamp 1679581782
transform 1 0 91296 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_952
timestamp 1679581782
transform 1 0 91968 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_959
timestamp 1679581782
transform 1 0 92640 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_966
timestamp 1679581782
transform 1 0 93312 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_973
timestamp 1679581782
transform 1 0 93984 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_980
timestamp 1679581782
transform 1 0 94656 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_987
timestamp 1679581782
transform 1 0 95328 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_994
timestamp 1679581782
transform 1 0 96000 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_1001
timestamp 1679581782
transform 1 0 96672 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_1008
timestamp 1679581782
transform 1 0 97344 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_1015
timestamp 1679581782
transform 1 0 98016 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_1022
timestamp 1679581782
transform 1 0 98688 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_0
timestamp 1679581782
transform 1 0 576 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_7
timestamp 1679581782
transform 1 0 1248 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_14
timestamp 1679581782
transform 1 0 1920 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_21
timestamp 1679581782
transform 1 0 2592 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_28
timestamp 1679581782
transform 1 0 3264 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_35
timestamp 1679581782
transform 1 0 3936 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_42
timestamp 1679581782
transform 1 0 4608 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_49
timestamp 1679581782
transform 1 0 5280 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_56
timestamp 1679581782
transform 1 0 5952 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_63
timestamp 1679581782
transform 1 0 6624 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_70
timestamp 1679581782
transform 1 0 7296 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_77
timestamp 1679581782
transform 1 0 7968 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_84
timestamp 1679581782
transform 1 0 8640 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_91
timestamp 1679581782
transform 1 0 9312 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_98
timestamp 1679581782
transform 1 0 9984 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_105
timestamp 1679581782
transform 1 0 10656 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_112
timestamp 1679581782
transform 1 0 11328 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_119
timestamp 1679581782
transform 1 0 12000 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_126
timestamp 1679581782
transform 1 0 12672 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_133
timestamp 1679581782
transform 1 0 13344 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_140
timestamp 1679581782
transform 1 0 14016 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_147
timestamp 1679581782
transform 1 0 14688 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_154
timestamp 1679581782
transform 1 0 15360 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_161
timestamp 1679581782
transform 1 0 16032 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_168
timestamp 1679581782
transform 1 0 16704 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_175
timestamp 1679581782
transform 1 0 17376 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_182
timestamp 1679581782
transform 1 0 18048 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_189
timestamp 1679581782
transform 1 0 18720 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_196
timestamp 1679581782
transform 1 0 19392 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_203
timestamp 1679581782
transform 1 0 20064 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_210
timestamp 1679581782
transform 1 0 20736 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_217
timestamp 1679581782
transform 1 0 21408 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_224
timestamp 1679581782
transform 1 0 22080 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_231
timestamp 1679581782
transform 1 0 22752 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_238
timestamp 1679581782
transform 1 0 23424 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_245
timestamp 1679581782
transform 1 0 24096 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_252
timestamp 1679581782
transform 1 0 24768 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_259
timestamp 1679581782
transform 1 0 25440 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_266
timestamp 1679581782
transform 1 0 26112 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_273
timestamp 1679581782
transform 1 0 26784 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_280
timestamp 1679581782
transform 1 0 27456 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_287
timestamp 1679581782
transform 1 0 28128 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_294
timestamp 1679581782
transform 1 0 28800 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_301
timestamp 1679581782
transform 1 0 29472 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_308
timestamp 1679581782
transform 1 0 30144 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_315
timestamp 1679581782
transform 1 0 30816 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_322
timestamp 1679581782
transform 1 0 31488 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_329
timestamp 1679581782
transform 1 0 32160 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_336
timestamp 1679581782
transform 1 0 32832 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_343
timestamp 1679581782
transform 1 0 33504 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_350
timestamp 1679581782
transform 1 0 34176 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_357
timestamp 1679581782
transform 1 0 34848 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_364
timestamp 1679581782
transform 1 0 35520 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_371
timestamp 1679581782
transform 1 0 36192 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_378
timestamp 1679581782
transform 1 0 36864 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_385
timestamp 1679581782
transform 1 0 37536 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_392
timestamp 1679581782
transform 1 0 38208 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_399
timestamp 1679581782
transform 1 0 38880 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_406
timestamp 1679581782
transform 1 0 39552 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_413
timestamp 1679581782
transform 1 0 40224 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_420
timestamp 1679581782
transform 1 0 40896 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_427
timestamp 1679581782
transform 1 0 41568 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_434
timestamp 1679581782
transform 1 0 42240 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_441
timestamp 1679581782
transform 1 0 42912 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_448
timestamp 1679581782
transform 1 0 43584 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_455
timestamp 1679581782
transform 1 0 44256 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_462
timestamp 1679581782
transform 1 0 44928 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_469
timestamp 1679581782
transform 1 0 45600 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_476
timestamp 1679581782
transform 1 0 46272 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_483
timestamp 1679581782
transform 1 0 46944 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_490
timestamp 1679581782
transform 1 0 47616 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_497
timestamp 1679581782
transform 1 0 48288 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_504
timestamp 1679581782
transform 1 0 48960 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_511
timestamp 1679581782
transform 1 0 49632 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_518
timestamp 1679581782
transform 1 0 50304 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_525
timestamp 1679581782
transform 1 0 50976 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_532
timestamp 1679581782
transform 1 0 51648 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_539
timestamp 1679581782
transform 1 0 52320 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_546
timestamp 1679581782
transform 1 0 52992 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_553
timestamp 1679581782
transform 1 0 53664 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_560
timestamp 1679581782
transform 1 0 54336 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_567
timestamp 1679581782
transform 1 0 55008 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_574
timestamp 1679581782
transform 1 0 55680 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_581
timestamp 1679581782
transform 1 0 56352 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_588
timestamp 1679581782
transform 1 0 57024 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_595
timestamp 1679581782
transform 1 0 57696 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_602
timestamp 1679581782
transform 1 0 58368 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_609
timestamp 1679581782
transform 1 0 59040 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_616
timestamp 1679581782
transform 1 0 59712 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_623
timestamp 1679581782
transform 1 0 60384 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_630
timestamp 1679581782
transform 1 0 61056 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_637
timestamp 1679581782
transform 1 0 61728 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_644
timestamp 1679581782
transform 1 0 62400 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_651
timestamp 1679581782
transform 1 0 63072 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_658
timestamp 1679581782
transform 1 0 63744 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_665
timestamp 1679581782
transform 1 0 64416 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_672
timestamp 1679581782
transform 1 0 65088 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_679
timestamp 1679581782
transform 1 0 65760 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_686
timestamp 1679581782
transform 1 0 66432 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_693
timestamp 1679581782
transform 1 0 67104 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_700
timestamp 1679581782
transform 1 0 67776 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_707
timestamp 1679581782
transform 1 0 68448 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_714
timestamp 1679581782
transform 1 0 69120 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_721
timestamp 1679581782
transform 1 0 69792 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_728
timestamp 1679581782
transform 1 0 70464 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_735
timestamp 1679581782
transform 1 0 71136 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_742
timestamp 1679581782
transform 1 0 71808 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_749
timestamp 1679581782
transform 1 0 72480 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_756
timestamp 1679581782
transform 1 0 73152 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_763
timestamp 1679581782
transform 1 0 73824 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_770
timestamp 1679581782
transform 1 0 74496 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_777
timestamp 1679581782
transform 1 0 75168 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_784
timestamp 1679581782
transform 1 0 75840 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_791
timestamp 1679581782
transform 1 0 76512 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_798
timestamp 1679581782
transform 1 0 77184 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_805
timestamp 1679581782
transform 1 0 77856 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_812
timestamp 1679581782
transform 1 0 78528 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_819
timestamp 1679581782
transform 1 0 79200 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_826
timestamp 1679581782
transform 1 0 79872 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_833
timestamp 1679581782
transform 1 0 80544 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_840
timestamp 1679581782
transform 1 0 81216 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_847
timestamp 1679581782
transform 1 0 81888 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_854
timestamp 1679581782
transform 1 0 82560 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_861
timestamp 1679581782
transform 1 0 83232 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_868
timestamp 1679581782
transform 1 0 83904 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_875
timestamp 1679581782
transform 1 0 84576 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_882
timestamp 1679581782
transform 1 0 85248 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_889
timestamp 1679581782
transform 1 0 85920 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_896
timestamp 1679581782
transform 1 0 86592 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_903
timestamp 1679581782
transform 1 0 87264 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_910
timestamp 1679581782
transform 1 0 87936 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_917
timestamp 1679581782
transform 1 0 88608 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_924
timestamp 1679581782
transform 1 0 89280 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_931
timestamp 1679581782
transform 1 0 89952 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_938
timestamp 1679581782
transform 1 0 90624 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_945
timestamp 1679581782
transform 1 0 91296 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_952
timestamp 1679581782
transform 1 0 91968 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_959
timestamp 1679581782
transform 1 0 92640 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_966
timestamp 1679581782
transform 1 0 93312 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_973
timestamp 1679581782
transform 1 0 93984 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_980
timestamp 1679581782
transform 1 0 94656 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_987
timestamp 1679581782
transform 1 0 95328 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_994
timestamp 1679581782
transform 1 0 96000 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_1001
timestamp 1679581782
transform 1 0 96672 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_1008
timestamp 1679581782
transform 1 0 97344 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_1015
timestamp 1679581782
transform 1 0 98016 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_1022
timestamp 1679581782
transform 1 0 98688 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_0
timestamp 1679581782
transform 1 0 576 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_7
timestamp 1679581782
transform 1 0 1248 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_14
timestamp 1679581782
transform 1 0 1920 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_21
timestamp 1679581782
transform 1 0 2592 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_28
timestamp 1679581782
transform 1 0 3264 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_35
timestamp 1679581782
transform 1 0 3936 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_42
timestamp 1679581782
transform 1 0 4608 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_49
timestamp 1679581782
transform 1 0 5280 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_56
timestamp 1679581782
transform 1 0 5952 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_63
timestamp 1679581782
transform 1 0 6624 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_70
timestamp 1679581782
transform 1 0 7296 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_77
timestamp 1679581782
transform 1 0 7968 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_84
timestamp 1679581782
transform 1 0 8640 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_91
timestamp 1679581782
transform 1 0 9312 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_98
timestamp 1679581782
transform 1 0 9984 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_105
timestamp 1679581782
transform 1 0 10656 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_112
timestamp 1679581782
transform 1 0 11328 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_119
timestamp 1679581782
transform 1 0 12000 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_126
timestamp 1679581782
transform 1 0 12672 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_133
timestamp 1679581782
transform 1 0 13344 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_140
timestamp 1679581782
transform 1 0 14016 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_147
timestamp 1679581782
transform 1 0 14688 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_154
timestamp 1679581782
transform 1 0 15360 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_161
timestamp 1679581782
transform 1 0 16032 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_168
timestamp 1679581782
transform 1 0 16704 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_175
timestamp 1679581782
transform 1 0 17376 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_182
timestamp 1679581782
transform 1 0 18048 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_189
timestamp 1679581782
transform 1 0 18720 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_196
timestamp 1679581782
transform 1 0 19392 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_203
timestamp 1679581782
transform 1 0 20064 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_210
timestamp 1679581782
transform 1 0 20736 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_217
timestamp 1679581782
transform 1 0 21408 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_224
timestamp 1679581782
transform 1 0 22080 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_231
timestamp 1679581782
transform 1 0 22752 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_238
timestamp 1679581782
transform 1 0 23424 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_245
timestamp 1679581782
transform 1 0 24096 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_252
timestamp 1679581782
transform 1 0 24768 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_259
timestamp 1679581782
transform 1 0 25440 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_266
timestamp 1679581782
transform 1 0 26112 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_273
timestamp 1679581782
transform 1 0 26784 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_280
timestamp 1679581782
transform 1 0 27456 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_287
timestamp 1679581782
transform 1 0 28128 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_294
timestamp 1679581782
transform 1 0 28800 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_301
timestamp 1679581782
transform 1 0 29472 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_308
timestamp 1679581782
transform 1 0 30144 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_315
timestamp 1679581782
transform 1 0 30816 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_322
timestamp 1679581782
transform 1 0 31488 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_329
timestamp 1679581782
transform 1 0 32160 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_336
timestamp 1679581782
transform 1 0 32832 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_343
timestamp 1679581782
transform 1 0 33504 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_350
timestamp 1679581782
transform 1 0 34176 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_357
timestamp 1679581782
transform 1 0 34848 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_364
timestamp 1679581782
transform 1 0 35520 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_371
timestamp 1679581782
transform 1 0 36192 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_378
timestamp 1679581782
transform 1 0 36864 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_385
timestamp 1679581782
transform 1 0 37536 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_392
timestamp 1679581782
transform 1 0 38208 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_399
timestamp 1679581782
transform 1 0 38880 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_406
timestamp 1679581782
transform 1 0 39552 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_413
timestamp 1679581782
transform 1 0 40224 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_420
timestamp 1679581782
transform 1 0 40896 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_427
timestamp 1679581782
transform 1 0 41568 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_434
timestamp 1679581782
transform 1 0 42240 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_441
timestamp 1679581782
transform 1 0 42912 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_448
timestamp 1679581782
transform 1 0 43584 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_455
timestamp 1679581782
transform 1 0 44256 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_462
timestamp 1679581782
transform 1 0 44928 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_469
timestamp 1679581782
transform 1 0 45600 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_476
timestamp 1679581782
transform 1 0 46272 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_483
timestamp 1679581782
transform 1 0 46944 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_490
timestamp 1679581782
transform 1 0 47616 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_497
timestamp 1679581782
transform 1 0 48288 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_504
timestamp 1679581782
transform 1 0 48960 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_511
timestamp 1679581782
transform 1 0 49632 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_518
timestamp 1679581782
transform 1 0 50304 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_525
timestamp 1679581782
transform 1 0 50976 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_532
timestamp 1679581782
transform 1 0 51648 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_539
timestamp 1679581782
transform 1 0 52320 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_546
timestamp 1679581782
transform 1 0 52992 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_553
timestamp 1679581782
transform 1 0 53664 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_560
timestamp 1679581782
transform 1 0 54336 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_567
timestamp 1679581782
transform 1 0 55008 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_574
timestamp 1679581782
transform 1 0 55680 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_581
timestamp 1679581782
transform 1 0 56352 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_588
timestamp 1679581782
transform 1 0 57024 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_595
timestamp 1679581782
transform 1 0 57696 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_602
timestamp 1679581782
transform 1 0 58368 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_609
timestamp 1679581782
transform 1 0 59040 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_616
timestamp 1679581782
transform 1 0 59712 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_623
timestamp 1679581782
transform 1 0 60384 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_630
timestamp 1679581782
transform 1 0 61056 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_637
timestamp 1679581782
transform 1 0 61728 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_644
timestamp 1679581782
transform 1 0 62400 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_651
timestamp 1679581782
transform 1 0 63072 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_658
timestamp 1679581782
transform 1 0 63744 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_665
timestamp 1679581782
transform 1 0 64416 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_672
timestamp 1679581782
transform 1 0 65088 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_679
timestamp 1679581782
transform 1 0 65760 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_686
timestamp 1679581782
transform 1 0 66432 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_693
timestamp 1679581782
transform 1 0 67104 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_700
timestamp 1679581782
transform 1 0 67776 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_707
timestamp 1679581782
transform 1 0 68448 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_714
timestamp 1679581782
transform 1 0 69120 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_721
timestamp 1679581782
transform 1 0 69792 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_728
timestamp 1679581782
transform 1 0 70464 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_735
timestamp 1679581782
transform 1 0 71136 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_742
timestamp 1679581782
transform 1 0 71808 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_749
timestamp 1679581782
transform 1 0 72480 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_756
timestamp 1679581782
transform 1 0 73152 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_763
timestamp 1679581782
transform 1 0 73824 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_770
timestamp 1679581782
transform 1 0 74496 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_777
timestamp 1679581782
transform 1 0 75168 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_784
timestamp 1679581782
transform 1 0 75840 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_791
timestamp 1679581782
transform 1 0 76512 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_798
timestamp 1679581782
transform 1 0 77184 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_805
timestamp 1679581782
transform 1 0 77856 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_812
timestamp 1679581782
transform 1 0 78528 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_819
timestamp 1679581782
transform 1 0 79200 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_826
timestamp 1679581782
transform 1 0 79872 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_833
timestamp 1679581782
transform 1 0 80544 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_840
timestamp 1679581782
transform 1 0 81216 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_847
timestamp 1679581782
transform 1 0 81888 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_854
timestamp 1679581782
transform 1 0 82560 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_861
timestamp 1679581782
transform 1 0 83232 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_868
timestamp 1679581782
transform 1 0 83904 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_875
timestamp 1679581782
transform 1 0 84576 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_882
timestamp 1679581782
transform 1 0 85248 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_889
timestamp 1679581782
transform 1 0 85920 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_896
timestamp 1679581782
transform 1 0 86592 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_903
timestamp 1679581782
transform 1 0 87264 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_910
timestamp 1679581782
transform 1 0 87936 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_917
timestamp 1679581782
transform 1 0 88608 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_924
timestamp 1679581782
transform 1 0 89280 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_931
timestamp 1679581782
transform 1 0 89952 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_938
timestamp 1679581782
transform 1 0 90624 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_945
timestamp 1679581782
transform 1 0 91296 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_952
timestamp 1679581782
transform 1 0 91968 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_959
timestamp 1679581782
transform 1 0 92640 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_966
timestamp 1679581782
transform 1 0 93312 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_973
timestamp 1679581782
transform 1 0 93984 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_980
timestamp 1679581782
transform 1 0 94656 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_987
timestamp 1679581782
transform 1 0 95328 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_994
timestamp 1679581782
transform 1 0 96000 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_1001
timestamp 1679581782
transform 1 0 96672 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_1008
timestamp 1679581782
transform 1 0 97344 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_1015
timestamp 1679581782
transform 1 0 98016 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_1022
timestamp 1679581782
transform 1 0 98688 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_0
timestamp 1679581782
transform 1 0 576 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_7
timestamp 1679581782
transform 1 0 1248 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_14
timestamp 1679581782
transform 1 0 1920 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_21
timestamp 1679581782
transform 1 0 2592 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_28
timestamp 1679581782
transform 1 0 3264 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_35
timestamp 1679581782
transform 1 0 3936 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_42
timestamp 1679581782
transform 1 0 4608 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_49
timestamp 1679581782
transform 1 0 5280 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_56
timestamp 1679581782
transform 1 0 5952 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_63
timestamp 1679581782
transform 1 0 6624 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_70
timestamp 1679581782
transform 1 0 7296 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_77
timestamp 1679581782
transform 1 0 7968 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_84
timestamp 1679581782
transform 1 0 8640 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_91
timestamp 1679581782
transform 1 0 9312 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_98
timestamp 1679581782
transform 1 0 9984 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_105
timestamp 1679581782
transform 1 0 10656 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_112
timestamp 1679581782
transform 1 0 11328 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_119
timestamp 1679581782
transform 1 0 12000 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_126
timestamp 1679581782
transform 1 0 12672 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_133
timestamp 1679581782
transform 1 0 13344 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_140
timestamp 1679581782
transform 1 0 14016 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_147
timestamp 1679581782
transform 1 0 14688 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_154
timestamp 1679581782
transform 1 0 15360 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_161
timestamp 1679581782
transform 1 0 16032 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_168
timestamp 1679581782
transform 1 0 16704 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_175
timestamp 1679581782
transform 1 0 17376 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_182
timestamp 1679581782
transform 1 0 18048 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_189
timestamp 1679581782
transform 1 0 18720 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_196
timestamp 1679581782
transform 1 0 19392 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_203
timestamp 1679581782
transform 1 0 20064 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_210
timestamp 1679581782
transform 1 0 20736 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_217
timestamp 1679581782
transform 1 0 21408 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_224
timestamp 1679581782
transform 1 0 22080 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_231
timestamp 1679581782
transform 1 0 22752 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_238
timestamp 1679581782
transform 1 0 23424 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_245
timestamp 1679581782
transform 1 0 24096 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_252
timestamp 1679581782
transform 1 0 24768 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_259
timestamp 1679581782
transform 1 0 25440 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_266
timestamp 1679581782
transform 1 0 26112 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_273
timestamp 1679581782
transform 1 0 26784 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_280
timestamp 1679581782
transform 1 0 27456 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_287
timestamp 1679581782
transform 1 0 28128 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_294
timestamp 1679581782
transform 1 0 28800 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_301
timestamp 1679581782
transform 1 0 29472 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_308
timestamp 1679581782
transform 1 0 30144 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_315
timestamp 1679581782
transform 1 0 30816 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_322
timestamp 1679581782
transform 1 0 31488 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_329
timestamp 1679581782
transform 1 0 32160 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_336
timestamp 1679581782
transform 1 0 32832 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_343
timestamp 1679581782
transform 1 0 33504 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_350
timestamp 1679581782
transform 1 0 34176 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_357
timestamp 1679581782
transform 1 0 34848 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_364
timestamp 1679581782
transform 1 0 35520 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_371
timestamp 1679581782
transform 1 0 36192 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_378
timestamp 1679581782
transform 1 0 36864 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_385
timestamp 1679581782
transform 1 0 37536 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_392
timestamp 1679581782
transform 1 0 38208 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_399
timestamp 1679581782
transform 1 0 38880 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_406
timestamp 1679581782
transform 1 0 39552 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_413
timestamp 1679581782
transform 1 0 40224 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_420
timestamp 1679581782
transform 1 0 40896 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_427
timestamp 1679581782
transform 1 0 41568 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_434
timestamp 1679581782
transform 1 0 42240 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_441
timestamp 1679581782
transform 1 0 42912 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_448
timestamp 1679581782
transform 1 0 43584 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_455
timestamp 1679581782
transform 1 0 44256 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_462
timestamp 1679581782
transform 1 0 44928 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_469
timestamp 1679581782
transform 1 0 45600 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_476
timestamp 1679581782
transform 1 0 46272 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_483
timestamp 1679581782
transform 1 0 46944 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_490
timestamp 1679581782
transform 1 0 47616 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_497
timestamp 1679581782
transform 1 0 48288 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_504
timestamp 1679581782
transform 1 0 48960 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_511
timestamp 1679581782
transform 1 0 49632 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_518
timestamp 1679581782
transform 1 0 50304 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_525
timestamp 1679581782
transform 1 0 50976 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_532
timestamp 1679581782
transform 1 0 51648 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_539
timestamp 1679581782
transform 1 0 52320 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_546
timestamp 1679581782
transform 1 0 52992 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_553
timestamp 1679581782
transform 1 0 53664 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_560
timestamp 1679581782
transform 1 0 54336 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_567
timestamp 1679581782
transform 1 0 55008 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_574
timestamp 1679581782
transform 1 0 55680 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_581
timestamp 1679581782
transform 1 0 56352 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_588
timestamp 1679581782
transform 1 0 57024 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_595
timestamp 1679581782
transform 1 0 57696 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_602
timestamp 1679581782
transform 1 0 58368 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_609
timestamp 1679581782
transform 1 0 59040 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_616
timestamp 1679581782
transform 1 0 59712 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_623
timestamp 1679581782
transform 1 0 60384 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_630
timestamp 1679581782
transform 1 0 61056 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_637
timestamp 1679581782
transform 1 0 61728 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_644
timestamp 1679581782
transform 1 0 62400 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_651
timestamp 1679581782
transform 1 0 63072 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_658
timestamp 1679581782
transform 1 0 63744 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_665
timestamp 1679581782
transform 1 0 64416 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_672
timestamp 1679581782
transform 1 0 65088 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_679
timestamp 1679581782
transform 1 0 65760 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_686
timestamp 1679581782
transform 1 0 66432 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_693
timestamp 1679581782
transform 1 0 67104 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_700
timestamp 1679581782
transform 1 0 67776 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_707
timestamp 1679581782
transform 1 0 68448 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_714
timestamp 1679581782
transform 1 0 69120 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_721
timestamp 1679581782
transform 1 0 69792 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_728
timestamp 1679581782
transform 1 0 70464 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_735
timestamp 1679581782
transform 1 0 71136 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_742
timestamp 1679581782
transform 1 0 71808 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_749
timestamp 1679581782
transform 1 0 72480 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_756
timestamp 1679581782
transform 1 0 73152 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_763
timestamp 1679581782
transform 1 0 73824 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_770
timestamp 1679581782
transform 1 0 74496 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_777
timestamp 1679581782
transform 1 0 75168 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_784
timestamp 1679581782
transform 1 0 75840 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_791
timestamp 1679581782
transform 1 0 76512 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_798
timestamp 1679581782
transform 1 0 77184 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_805
timestamp 1679581782
transform 1 0 77856 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_812
timestamp 1679581782
transform 1 0 78528 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_819
timestamp 1679581782
transform 1 0 79200 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_826
timestamp 1679581782
transform 1 0 79872 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_833
timestamp 1679581782
transform 1 0 80544 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_840
timestamp 1679581782
transform 1 0 81216 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_847
timestamp 1679581782
transform 1 0 81888 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_854
timestamp 1679581782
transform 1 0 82560 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_861
timestamp 1679581782
transform 1 0 83232 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_868
timestamp 1679581782
transform 1 0 83904 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_875
timestamp 1679581782
transform 1 0 84576 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_882
timestamp 1679581782
transform 1 0 85248 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_889
timestamp 1679581782
transform 1 0 85920 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_896
timestamp 1679581782
transform 1 0 86592 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_903
timestamp 1679581782
transform 1 0 87264 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_910
timestamp 1679581782
transform 1 0 87936 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_917
timestamp 1679581782
transform 1 0 88608 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_924
timestamp 1679581782
transform 1 0 89280 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_931
timestamp 1679581782
transform 1 0 89952 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_938
timestamp 1679581782
transform 1 0 90624 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_945
timestamp 1679581782
transform 1 0 91296 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_952
timestamp 1679581782
transform 1 0 91968 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_959
timestamp 1679581782
transform 1 0 92640 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_966
timestamp 1679581782
transform 1 0 93312 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_973
timestamp 1679581782
transform 1 0 93984 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_980
timestamp 1679581782
transform 1 0 94656 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_987
timestamp 1679581782
transform 1 0 95328 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_994
timestamp 1679581782
transform 1 0 96000 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_1001
timestamp 1679581782
transform 1 0 96672 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_1008
timestamp 1679581782
transform 1 0 97344 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_1015
timestamp 1679581782
transform 1 0 98016 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_1022
timestamp 1679581782
transform 1 0 98688 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_0
timestamp 1679581782
transform 1 0 576 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_7
timestamp 1679581782
transform 1 0 1248 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_14
timestamp 1679581782
transform 1 0 1920 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_21
timestamp 1679581782
transform 1 0 2592 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_28
timestamp 1679581782
transform 1 0 3264 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_35
timestamp 1679581782
transform 1 0 3936 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_42
timestamp 1679581782
transform 1 0 4608 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_49
timestamp 1679581782
transform 1 0 5280 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_56
timestamp 1679581782
transform 1 0 5952 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_63
timestamp 1679581782
transform 1 0 6624 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_70
timestamp 1679581782
transform 1 0 7296 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_77
timestamp 1679581782
transform 1 0 7968 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_84
timestamp 1679581782
transform 1 0 8640 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_91
timestamp 1679581782
transform 1 0 9312 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_98
timestamp 1679581782
transform 1 0 9984 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_105
timestamp 1679581782
transform 1 0 10656 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_112
timestamp 1679581782
transform 1 0 11328 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_119
timestamp 1679581782
transform 1 0 12000 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_126
timestamp 1679581782
transform 1 0 12672 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_133
timestamp 1679581782
transform 1 0 13344 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_140
timestamp 1679581782
transform 1 0 14016 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_147
timestamp 1679581782
transform 1 0 14688 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_154
timestamp 1679581782
transform 1 0 15360 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_161
timestamp 1679581782
transform 1 0 16032 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_168
timestamp 1679581782
transform 1 0 16704 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_175
timestamp 1679581782
transform 1 0 17376 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_182
timestamp 1679581782
transform 1 0 18048 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_189
timestamp 1679581782
transform 1 0 18720 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_196
timestamp 1679581782
transform 1 0 19392 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_203
timestamp 1679581782
transform 1 0 20064 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_210
timestamp 1679581782
transform 1 0 20736 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_217
timestamp 1679581782
transform 1 0 21408 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_224
timestamp 1679581782
transform 1 0 22080 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_231
timestamp 1679581782
transform 1 0 22752 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_238
timestamp 1679581782
transform 1 0 23424 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_245
timestamp 1679581782
transform 1 0 24096 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_252
timestamp 1679581782
transform 1 0 24768 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_259
timestamp 1679581782
transform 1 0 25440 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_266
timestamp 1679581782
transform 1 0 26112 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_273
timestamp 1679581782
transform 1 0 26784 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_280
timestamp 1679581782
transform 1 0 27456 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_287
timestamp 1679581782
transform 1 0 28128 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_294
timestamp 1679581782
transform 1 0 28800 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_301
timestamp 1679581782
transform 1 0 29472 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_308
timestamp 1679581782
transform 1 0 30144 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_315
timestamp 1679581782
transform 1 0 30816 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_322
timestamp 1679581782
transform 1 0 31488 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_329
timestamp 1679581782
transform 1 0 32160 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_336
timestamp 1679581782
transform 1 0 32832 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_343
timestamp 1679581782
transform 1 0 33504 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_350
timestamp 1679581782
transform 1 0 34176 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_357
timestamp 1679581782
transform 1 0 34848 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_364
timestamp 1679581782
transform 1 0 35520 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_371
timestamp 1679581782
transform 1 0 36192 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_378
timestamp 1679581782
transform 1 0 36864 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_385
timestamp 1679581782
transform 1 0 37536 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_392
timestamp 1679581782
transform 1 0 38208 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_399
timestamp 1679581782
transform 1 0 38880 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_406
timestamp 1679581782
transform 1 0 39552 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_413
timestamp 1679581782
transform 1 0 40224 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_420
timestamp 1679581782
transform 1 0 40896 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_427
timestamp 1679581782
transform 1 0 41568 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_434
timestamp 1679581782
transform 1 0 42240 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_441
timestamp 1679581782
transform 1 0 42912 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_448
timestamp 1679581782
transform 1 0 43584 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_455
timestamp 1679581782
transform 1 0 44256 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_462
timestamp 1679581782
transform 1 0 44928 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_469
timestamp 1679581782
transform 1 0 45600 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_476
timestamp 1679581782
transform 1 0 46272 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_483
timestamp 1679581782
transform 1 0 46944 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_490
timestamp 1679581782
transform 1 0 47616 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_497
timestamp 1679581782
transform 1 0 48288 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_504
timestamp 1679581782
transform 1 0 48960 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_511
timestamp 1679581782
transform 1 0 49632 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_518
timestamp 1679581782
transform 1 0 50304 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_525
timestamp 1679581782
transform 1 0 50976 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_532
timestamp 1679581782
transform 1 0 51648 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_539
timestamp 1679581782
transform 1 0 52320 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_546
timestamp 1679581782
transform 1 0 52992 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_553
timestamp 1679581782
transform 1 0 53664 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_560
timestamp 1679581782
transform 1 0 54336 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_567
timestamp 1679581782
transform 1 0 55008 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_574
timestamp 1679581782
transform 1 0 55680 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_581
timestamp 1679581782
transform 1 0 56352 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_588
timestamp 1679581782
transform 1 0 57024 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_595
timestamp 1679581782
transform 1 0 57696 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_602
timestamp 1679581782
transform 1 0 58368 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_609
timestamp 1679581782
transform 1 0 59040 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_616
timestamp 1679581782
transform 1 0 59712 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_623
timestamp 1679581782
transform 1 0 60384 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_630
timestamp 1679581782
transform 1 0 61056 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_637
timestamp 1679581782
transform 1 0 61728 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_644
timestamp 1679581782
transform 1 0 62400 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_651
timestamp 1679581782
transform 1 0 63072 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_658
timestamp 1679581782
transform 1 0 63744 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_665
timestamp 1679581782
transform 1 0 64416 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_672
timestamp 1679581782
transform 1 0 65088 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_679
timestamp 1679581782
transform 1 0 65760 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_686
timestamp 1679581782
transform 1 0 66432 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_693
timestamp 1679581782
transform 1 0 67104 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_700
timestamp 1679581782
transform 1 0 67776 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_707
timestamp 1679581782
transform 1 0 68448 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_714
timestamp 1679581782
transform 1 0 69120 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_721
timestamp 1679581782
transform 1 0 69792 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_728
timestamp 1679581782
transform 1 0 70464 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_735
timestamp 1679581782
transform 1 0 71136 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_742
timestamp 1679581782
transform 1 0 71808 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_749
timestamp 1679581782
transform 1 0 72480 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_756
timestamp 1679581782
transform 1 0 73152 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_763
timestamp 1679581782
transform 1 0 73824 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_770
timestamp 1679581782
transform 1 0 74496 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_777
timestamp 1679581782
transform 1 0 75168 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_784
timestamp 1679581782
transform 1 0 75840 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_791
timestamp 1679581782
transform 1 0 76512 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_798
timestamp 1679581782
transform 1 0 77184 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_805
timestamp 1679581782
transform 1 0 77856 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_812
timestamp 1679581782
transform 1 0 78528 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_819
timestamp 1679581782
transform 1 0 79200 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_826
timestamp 1679581782
transform 1 0 79872 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_833
timestamp 1679581782
transform 1 0 80544 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_840
timestamp 1679581782
transform 1 0 81216 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_847
timestamp 1679581782
transform 1 0 81888 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_854
timestamp 1679581782
transform 1 0 82560 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_861
timestamp 1679581782
transform 1 0 83232 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_868
timestamp 1679581782
transform 1 0 83904 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_875
timestamp 1679581782
transform 1 0 84576 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_882
timestamp 1679581782
transform 1 0 85248 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_889
timestamp 1679581782
transform 1 0 85920 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_896
timestamp 1679581782
transform 1 0 86592 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_903
timestamp 1679581782
transform 1 0 87264 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_910
timestamp 1679581782
transform 1 0 87936 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_917
timestamp 1679581782
transform 1 0 88608 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_924
timestamp 1679581782
transform 1 0 89280 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_931
timestamp 1679581782
transform 1 0 89952 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_938
timestamp 1679581782
transform 1 0 90624 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_945
timestamp 1679581782
transform 1 0 91296 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_952
timestamp 1679581782
transform 1 0 91968 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_959
timestamp 1679581782
transform 1 0 92640 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_966
timestamp 1679581782
transform 1 0 93312 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_973
timestamp 1679581782
transform 1 0 93984 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_980
timestamp 1679581782
transform 1 0 94656 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_987
timestamp 1679581782
transform 1 0 95328 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_994
timestamp 1679581782
transform 1 0 96000 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_1001
timestamp 1679581782
transform 1 0 96672 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_1008
timestamp 1679581782
transform 1 0 97344 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_1015
timestamp 1679581782
transform 1 0 98016 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_106_1022
timestamp 1679581782
transform 1 0 98688 0 1 80892
box -48 -56 720 834
use sg13g2_tielo  heichips25_example_large_25
timestamp 1680000637
transform -1 0 960 0 1 32508
box -48 -56 432 834
use sg13g2_tielo  heichips25_example_large_26
timestamp 1680000637
transform -1 0 960 0 1 34020
box -48 -56 432 834
use sg13g2_tielo  heichips25_example_large_27
timestamp 1680000637
transform -1 0 960 0 1 35532
box -48 -56 432 834
use sg13g2_tielo  heichips25_example_large_28
timestamp 1680000637
transform -1 0 960 0 -1 38556
box -48 -56 432 834
use sg13g2_tielo  heichips25_example_large_29
timestamp 1680000637
transform -1 0 960 0 -1 40068
box -48 -56 432 834
use sg13g2_tielo  heichips25_example_large_30
timestamp 1680000637
transform -1 0 960 0 1 41580
box -48 -56 432 834
use sg13g2_tielo  heichips25_example_large_31
timestamp 1680000637
transform -1 0 960 0 1 43092
box -48 -56 432 834
use sg13g2_tielo  heichips25_example_large_32
timestamp 1680000637
transform -1 0 960 0 -1 46116
box -48 -56 432 834
use sg13g2_tielo  heichips25_example_large_33
timestamp 1680000637
transform -1 0 960 0 1 17388
box -48 -56 432 834
use sg13g2_tielo  heichips25_example_large_34
timestamp 1680000637
transform -1 0 960 0 1 18900
box -48 -56 432 834
use sg13g2_tielo  heichips25_example_large_35
timestamp 1680000637
transform -1 0 960 0 -1 21924
box -48 -56 432 834
use sg13g2_tielo  heichips25_example_large_36
timestamp 1680000637
transform -1 0 960 0 -1 23436
box -48 -56 432 834
use sg13g2_tielo  heichips25_example_large_37
timestamp 1680000637
transform -1 0 960 0 1 24948
box -48 -56 432 834
use sg13g2_tielo  heichips25_example_large_38
timestamp 1680000637
transform -1 0 960 0 1 26460
box -48 -56 432 834
use sg13g2_tielo  heichips25_example_large_39
timestamp 1680000637
transform -1 0 960 0 -1 29484
box -48 -56 432 834
use sg13g2_tielo  heichips25_example_large_40
timestamp 1680000637
transform -1 0 960 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  input1
timestamp 1676381911
transform 1 0 576 0 -1 47628
box -48 -56 432 834
use sg13g2_buf_1  input2
timestamp 1676381911
transform 1 0 576 0 1 49140
box -48 -56 432 834
use sg13g2_buf_1  input3
timestamp 1676381911
transform 1 0 576 0 1 50652
box -48 -56 432 834
use sg13g2_buf_1  input4
timestamp 1676381911
transform 1 0 576 0 1 52164
box -48 -56 432 834
use sg13g2_buf_1  input5
timestamp 1676381911
transform 1 0 576 0 -1 55188
box -48 -56 432 834
use sg13g2_buf_1  input6
timestamp 1676381911
transform 1 0 576 0 -1 56700
box -48 -56 432 834
use sg13g2_buf_1  input7
timestamp 1676381911
transform 1 0 576 0 1 58212
box -48 -56 432 834
use sg13g2_buf_1  input8
timestamp 1676381911
transform 1 0 576 0 1 59724
box -48 -56 432 834
use sg13g2_buf_1  input9
timestamp 1676381911
transform 1 0 576 0 -1 62748
box -48 -56 432 834
use sg13g2_buf_1  input10
timestamp 1676381911
transform 1 0 576 0 -1 64260
box -48 -56 432 834
use sg13g2_buf_1  input11
timestamp 1676381911
transform 1 0 576 0 1 65772
box -48 -56 432 834
use sg13g2_buf_1  input12
timestamp 1676381911
transform 1 0 576 0 1 67284
box -48 -56 432 834
use sg13g2_buf_1  input13
timestamp 1676381911
transform 1 0 576 0 1 68796
box -48 -56 432 834
use sg13g2_buf_2  input14
timestamp 1676381867
transform -1 0 1056 0 -1 71820
box -48 -56 528 834
use sg13g2_buf_1  input15
timestamp 1676381911
transform 1 0 576 0 -1 73332
box -48 -56 432 834
use sg13g2_buf_1  input16
timestamp 1676381911
transform 1 0 576 0 1 74844
box -48 -56 432 834
use sg13g2_buf_1  output17
timestamp 1676381911
transform -1 0 960 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  output18
timestamp 1676381911
transform -1 0 960 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  output19
timestamp 1676381911
transform -1 0 960 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  output20
timestamp 1676381911
transform -1 0 960 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  output21
timestamp 1676381911
transform -1 0 960 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  output22
timestamp 1676381911
transform -1 0 960 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  output23
timestamp 1676381911
transform -1 0 960 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  output24
timestamp 1676381911
transform -1 0 960 0 1 15876
box -48 -56 432 834
<< labels >>
flabel metal6 s 4316 630 4756 81692 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 19436 630 19876 81692 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 34556 630 34996 81692 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 49676 630 50116 81692 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 64796 630 65236 81692 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 79916 630 80356 81692 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 95036 630 95476 81692 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 3076 712 3516 81774 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 18196 712 18636 81774 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 33316 712 33756 81774 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 48436 712 48876 81774 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 63556 712 63996 81774 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 78676 712 79116 81774 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 93796 712 94236 81774 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 78332 80 78412 0 FreeSans 320 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 0 76484 80 76564 0 FreeSans 320 0 0 0 ena
port 3 nsew signal input
flabel metal3 s 0 80180 80 80260 0 FreeSans 320 0 0 0 rst_n
port 4 nsew signal input
flabel metal3 s 0 46916 80 46996 0 FreeSans 320 0 0 0 ui_in[0]
port 5 nsew signal input
flabel metal3 s 0 48764 80 48844 0 FreeSans 320 0 0 0 ui_in[1]
port 6 nsew signal input
flabel metal3 s 0 50612 80 50692 0 FreeSans 320 0 0 0 ui_in[2]
port 7 nsew signal input
flabel metal3 s 0 52460 80 52540 0 FreeSans 320 0 0 0 ui_in[3]
port 8 nsew signal input
flabel metal3 s 0 54308 80 54388 0 FreeSans 320 0 0 0 ui_in[4]
port 9 nsew signal input
flabel metal3 s 0 56156 80 56236 0 FreeSans 320 0 0 0 ui_in[5]
port 10 nsew signal input
flabel metal3 s 0 58004 80 58084 0 FreeSans 320 0 0 0 ui_in[6]
port 11 nsew signal input
flabel metal3 s 0 59852 80 59932 0 FreeSans 320 0 0 0 ui_in[7]
port 12 nsew signal input
flabel metal3 s 0 61700 80 61780 0 FreeSans 320 0 0 0 uio_in[0]
port 13 nsew signal input
flabel metal3 s 0 63548 80 63628 0 FreeSans 320 0 0 0 uio_in[1]
port 14 nsew signal input
flabel metal3 s 0 65396 80 65476 0 FreeSans 320 0 0 0 uio_in[2]
port 15 nsew signal input
flabel metal3 s 0 67244 80 67324 0 FreeSans 320 0 0 0 uio_in[3]
port 16 nsew signal input
flabel metal3 s 0 69092 80 69172 0 FreeSans 320 0 0 0 uio_in[4]
port 17 nsew signal input
flabel metal3 s 0 70940 80 71020 0 FreeSans 320 0 0 0 uio_in[5]
port 18 nsew signal input
flabel metal3 s 0 72788 80 72868 0 FreeSans 320 0 0 0 uio_in[6]
port 19 nsew signal input
flabel metal3 s 0 74636 80 74716 0 FreeSans 320 0 0 0 uio_in[7]
port 20 nsew signal input
flabel metal3 s 0 32132 80 32212 0 FreeSans 320 0 0 0 uio_oe[0]
port 21 nsew signal output
flabel metal3 s 0 33980 80 34060 0 FreeSans 320 0 0 0 uio_oe[1]
port 22 nsew signal output
flabel metal3 s 0 35828 80 35908 0 FreeSans 320 0 0 0 uio_oe[2]
port 23 nsew signal output
flabel metal3 s 0 37676 80 37756 0 FreeSans 320 0 0 0 uio_oe[3]
port 24 nsew signal output
flabel metal3 s 0 39524 80 39604 0 FreeSans 320 0 0 0 uio_oe[4]
port 25 nsew signal output
flabel metal3 s 0 41372 80 41452 0 FreeSans 320 0 0 0 uio_oe[5]
port 26 nsew signal output
flabel metal3 s 0 43220 80 43300 0 FreeSans 320 0 0 0 uio_oe[6]
port 27 nsew signal output
flabel metal3 s 0 45068 80 45148 0 FreeSans 320 0 0 0 uio_oe[7]
port 28 nsew signal output
flabel metal3 s 0 17348 80 17428 0 FreeSans 320 0 0 0 uio_out[0]
port 29 nsew signal output
flabel metal3 s 0 19196 80 19276 0 FreeSans 320 0 0 0 uio_out[1]
port 30 nsew signal output
flabel metal3 s 0 21044 80 21124 0 FreeSans 320 0 0 0 uio_out[2]
port 31 nsew signal output
flabel metal3 s 0 22892 80 22972 0 FreeSans 320 0 0 0 uio_out[3]
port 32 nsew signal output
flabel metal3 s 0 24740 80 24820 0 FreeSans 320 0 0 0 uio_out[4]
port 33 nsew signal output
flabel metal3 s 0 26588 80 26668 0 FreeSans 320 0 0 0 uio_out[5]
port 34 nsew signal output
flabel metal3 s 0 28436 80 28516 0 FreeSans 320 0 0 0 uio_out[6]
port 35 nsew signal output
flabel metal3 s 0 30284 80 30364 0 FreeSans 320 0 0 0 uio_out[7]
port 36 nsew signal output
flabel metal3 s 0 2564 80 2644 0 FreeSans 320 0 0 0 uo_out[0]
port 37 nsew signal output
flabel metal3 s 0 4412 80 4492 0 FreeSans 320 0 0 0 uo_out[1]
port 38 nsew signal output
flabel metal3 s 0 6260 80 6340 0 FreeSans 320 0 0 0 uo_out[2]
port 39 nsew signal output
flabel metal3 s 0 8108 80 8188 0 FreeSans 320 0 0 0 uo_out[3]
port 40 nsew signal output
flabel metal3 s 0 9956 80 10036 0 FreeSans 320 0 0 0 uo_out[4]
port 41 nsew signal output
flabel metal3 s 0 11804 80 11884 0 FreeSans 320 0 0 0 uo_out[5]
port 42 nsew signal output
flabel metal3 s 0 13652 80 13732 0 FreeSans 320 0 0 0 uo_out[6]
port 43 nsew signal output
flabel metal3 s 0 15500 80 15580 0 FreeSans 320 0 0 0 uo_out[7]
port 44 nsew signal output
rlabel via1 49968 80892 49968 80892 0 VGND
rlabel metal1 49968 81648 49968 81648 0 VPWR
rlabel metal3 14544 46452 14544 46452 0 _00_
rlabel metal2 13728 46788 13728 46788 0 _01_
rlabel metal2 14112 47334 14112 47334 0 _02_
rlabel metal3 11856 47964 11856 47964 0 _03_
rlabel metal2 3840 47208 3840 47208 0 _04_
rlabel metal3 8448 47292 8448 47292 0 _05_
rlabel metal2 7008 47208 7008 47208 0 _06_
rlabel metal2 2880 46872 2880 46872 0 _07_
rlabel metal2 4032 47376 4032 47376 0 _08_
rlabel metal2 5856 47334 5856 47334 0 _09_
rlabel metal2 5952 47250 5952 47250 0 _10_
rlabel metal2 6336 47712 6336 47712 0 _11_
rlabel metal2 3936 47712 3936 47712 0 _12_
rlabel metal3 5040 52500 5040 52500 0 _13_
rlabel metal2 3264 51912 3264 51912 0 _14_
rlabel metal2 3936 51870 3936 51870 0 _15_
rlabel metal2 5424 51828 5424 51828 0 _16_
rlabel metal3 3744 51828 3744 51828 0 _17_
rlabel metal2 5856 52458 5856 52458 0 _18_
rlabel metal2 6240 51744 6240 51744 0 _19_
rlabel metal2 2880 51282 2880 51282 0 _20_
rlabel metal2 5760 52542 5760 52542 0 _21_
rlabel metal2 5664 52248 5664 52248 0 _22_
rlabel metal2 5664 54558 5664 54558 0 _23_
rlabel metal3 6432 57078 6432 57078 0 _24_
rlabel metal2 7104 57330 7104 57330 0 _25_
rlabel metal2 6720 56616 6720 56616 0 _26_
rlabel metal2 7296 58128 7296 58128 0 _27_
rlabel metal2 6912 60438 6912 60438 0 _28_
rlabel metal2 14592 45444 14592 45444 0 net1
rlabel metal3 13584 47292 13584 47292 0 net10
rlabel metal3 1008 65940 1008 65940 0 net11
rlabel metal2 2736 46620 2736 46620 0 net12
rlabel metal3 1056 68964 1056 68964 0 net13
rlabel metal2 1008 56196 1008 56196 0 net14
rlabel metal2 5856 57456 5856 57456 0 net15
rlabel metal2 816 75012 816 75012 0 net16
rlabel metal2 1008 2688 1008 2688 0 net17
rlabel metal3 7680 4872 7680 4872 0 net18
rlabel metal2 864 15120 864 15120 0 net19
rlabel metal2 13152 47502 13152 47502 0 net2
rlabel metal3 3264 8736 3264 8736 0 net20
rlabel metal3 3792 10248 3792 10248 0 net21
rlabel metal3 1392 12432 1392 12432 0 net22
rlabel metal2 960 13944 960 13944 0 net23
rlabel metal3 3984 16296 3984 16296 0 net24
rlabel metal3 366 32172 366 32172 0 net25
rlabel metal3 366 34020 366 34020 0 net26
rlabel metal3 366 35868 366 35868 0 net27
rlabel metal3 366 37716 366 37716 0 net28
rlabel metal3 366 39564 366 39564 0 net29
rlabel metal2 7872 47712 7872 47712 0 net3
rlabel metal3 366 41412 366 41412 0 net30
rlabel metal3 366 43260 366 43260 0 net31
rlabel metal3 366 45108 366 45108 0 net32
rlabel metal3 366 17388 366 17388 0 net33
rlabel metal3 366 19236 366 19236 0 net34
rlabel metal3 366 21084 366 21084 0 net35
rlabel metal3 366 22932 366 22932 0 net36
rlabel metal3 366 24780 366 24780 0 net37
rlabel metal3 366 26628 366 26628 0 net38
rlabel metal3 366 28476 366 28476 0 net39
rlabel metal2 2640 46452 2640 46452 0 net4
rlabel metal3 366 30324 366 30324 0 net40
rlabel metal2 2304 52164 2304 52164 0 net5
rlabel metal2 6048 52584 6048 52584 0 net6
rlabel metal2 6240 57078 6240 57078 0 net7
rlabel metal2 6624 60606 6624 60606 0 net8
rlabel metal2 14208 45360 14208 45360 0 net9
rlabel metal3 366 46956 366 46956 0 ui_in[0]
rlabel metal3 366 48804 366 48804 0 ui_in[1]
rlabel metal3 366 50652 366 50652 0 ui_in[2]
rlabel metal3 366 52500 366 52500 0 ui_in[3]
rlabel metal3 366 54348 366 54348 0 ui_in[4]
rlabel metal3 366 56196 366 56196 0 ui_in[5]
rlabel metal3 366 58044 366 58044 0 ui_in[6]
rlabel metal3 366 59892 366 59892 0 ui_in[7]
rlabel metal3 366 61740 366 61740 0 uio_in[0]
rlabel metal3 366 63588 366 63588 0 uio_in[1]
rlabel metal3 366 65436 366 65436 0 uio_in[2]
rlabel metal3 366 67284 366 67284 0 uio_in[3]
rlabel metal3 366 69132 366 69132 0 uio_in[4]
rlabel metal3 366 70980 366 70980 0 uio_in[5]
rlabel metal3 366 72828 366 72828 0 uio_in[6]
rlabel metal3 366 74676 366 74676 0 uio_in[7]
rlabel metal3 366 2604 366 2604 0 uo_out[0]
rlabel metal3 366 4452 366 4452 0 uo_out[1]
rlabel metal3 366 6300 366 6300 0 uo_out[2]
rlabel metal3 366 8148 366 8148 0 uo_out[3]
rlabel metal3 366 9996 366 9996 0 uo_out[4]
rlabel metal3 366 11844 366 11844 0 uo_out[5]
rlabel metal3 366 13692 366 13692 0 uo_out[6]
rlabel metal3 366 15540 366 15540 0 uo_out[7]
<< properties >>
string FIXED_BBOX 0 0 100000 83000
<< end >>
